//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 0 1 0 0 0 1 0 0 1 1 0 0 1 0 0 0 1 0 0 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 0 1 0 1 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:16 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n448, new_n451, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n551, new_n553, new_n554, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n575, new_n576, new_n577, new_n578, new_n581, new_n582, new_n583,
    new_n584, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n618, new_n621, new_n622, new_n624, new_n625, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1230, new_n1231, new_n1232;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  XNOR2_X1  g015(.A(KEYINPUT64), .B(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n447), .B(KEYINPUT65), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT1), .ZN(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT66), .ZN(G217));
  NAND4_X1  g027(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n455), .A2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n457), .A2(G567), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n464), .A2(G2104), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n465), .B1(new_n466), .B2(KEYINPUT67), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  OR3_X1    g044(.A1(new_n469), .A2(KEYINPUT67), .A3(KEYINPUT3), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n467), .A2(new_n468), .A3(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n472), .A2(KEYINPUT68), .A3(G137), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n469), .A2(KEYINPUT3), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n465), .A2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(G125), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n474), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n469), .A2(G2105), .ZN(new_n479));
  AOI22_X1  g054(.A1(new_n478), .A2(G2105), .B1(G101), .B2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT68), .ZN(new_n481));
  INV_X1    g056(.A(G137), .ZN(new_n482));
  OAI21_X1  g057(.A(new_n481), .B1(new_n471), .B2(new_n482), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n473), .A2(new_n480), .A3(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G160));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n468), .ZN(new_n487));
  INV_X1    g062(.A(G136), .ZN(new_n488));
  INV_X1    g063(.A(G124), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n467), .A2(G2105), .A3(new_n470), .ZN(new_n490));
  OAI221_X1 g065(.A(new_n487), .B1(new_n471), .B2(new_n488), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(G162));
  NOR2_X1   g067(.A1(new_n469), .A2(KEYINPUT3), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n493), .A2(new_n466), .ZN(new_n494));
  AND2_X1   g069(.A1(new_n468), .A2(G138), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  OR2_X1    g072(.A1(G102), .A2(G2105), .ZN(new_n498));
  INV_X1    g073(.A(G114), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n469), .B1(new_n499), .B2(G2105), .ZN(new_n500));
  AOI22_X1  g075(.A1(new_n496), .A2(new_n497), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n467), .A2(G126), .A3(G2105), .A4(new_n470), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n467), .A2(KEYINPUT4), .A3(new_n470), .A4(new_n495), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(G164));
  INV_X1    g080(.A(KEYINPUT5), .ZN(new_n506));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n506), .B1(new_n507), .B2(KEYINPUT69), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT69), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n509), .A2(KEYINPUT5), .A3(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n511), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n512));
  INV_X1    g087(.A(G651), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  XNOR2_X1  g089(.A(KEYINPUT6), .B(G651), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n511), .A2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(G88), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n515), .A2(G543), .ZN(new_n518));
  INV_X1    g093(.A(G50), .ZN(new_n519));
  OAI22_X1  g094(.A1(new_n516), .A2(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n514), .A2(new_n520), .ZN(G166));
  AND2_X1   g096(.A1(new_n511), .A2(new_n515), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G89), .ZN(new_n523));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n524), .B(KEYINPUT7), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n515), .A2(G51), .A3(G543), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT70), .ZN(new_n528));
  NAND2_X1  g103(.A1(G63), .A2(G651), .ZN(new_n529));
  INV_X1    g104(.A(new_n529), .ZN(new_n530));
  AOI21_X1  g105(.A(new_n528), .B1(new_n511), .B2(new_n530), .ZN(new_n531));
  AOI211_X1 g106(.A(KEYINPUT70), .B(new_n529), .C1(new_n508), .C2(new_n510), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n527), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(KEYINPUT71), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT71), .ZN(new_n535));
  OAI211_X1 g110(.A(new_n535), .B(new_n527), .C1(new_n531), .C2(new_n532), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n526), .B1(new_n534), .B2(new_n536), .ZN(G168));
  AOI22_X1  g112(.A1(new_n511), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n538), .A2(new_n513), .ZN(new_n539));
  INV_X1    g114(.A(G90), .ZN(new_n540));
  INV_X1    g115(.A(G52), .ZN(new_n541));
  OAI22_X1  g116(.A1(new_n516), .A2(new_n540), .B1(new_n518), .B2(new_n541), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n539), .A2(new_n542), .ZN(G171));
  AOI22_X1  g118(.A1(new_n511), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n544), .A2(new_n513), .ZN(new_n545));
  INV_X1    g120(.A(G81), .ZN(new_n546));
  INV_X1    g121(.A(G43), .ZN(new_n547));
  OAI22_X1  g122(.A1(new_n516), .A2(new_n546), .B1(new_n518), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  AND3_X1   g125(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G36), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n551), .A2(new_n554), .ZN(G188));
  INV_X1    g130(.A(KEYINPUT72), .ZN(new_n556));
  INV_X1    g131(.A(G91), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n556), .B1(new_n516), .B2(new_n557), .ZN(new_n558));
  NAND4_X1  g133(.A1(new_n511), .A2(KEYINPUT72), .A3(G91), .A4(new_n515), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n515), .A2(G53), .A3(G543), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT9), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT74), .ZN(new_n563));
  AND2_X1   g138(.A1(KEYINPUT73), .A2(G65), .ZN(new_n564));
  NOR2_X1   g139(.A1(KEYINPUT73), .A2(G65), .ZN(new_n565));
  NOR2_X1   g140(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n511), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(G78), .A2(G543), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n563), .B1(new_n569), .B2(G651), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n511), .A2(new_n566), .B1(G78), .B2(G543), .ZN(new_n571));
  NOR3_X1   g146(.A1(new_n571), .A2(KEYINPUT74), .A3(new_n513), .ZN(new_n572));
  OAI211_X1 g147(.A(new_n560), .B(new_n562), .C1(new_n570), .C2(new_n572), .ZN(G299));
  XNOR2_X1  g148(.A(G171), .B(KEYINPUT75), .ZN(G301));
  NOR2_X1   g149(.A1(G168), .A2(KEYINPUT76), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT76), .ZN(new_n576));
  AOI211_X1 g151(.A(new_n576), .B(new_n526), .C1(new_n534), .C2(new_n536), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(new_n578), .ZN(G286));
  INV_X1    g154(.A(G166), .ZN(G303));
  NAND2_X1  g155(.A1(new_n522), .A2(G87), .ZN(new_n581));
  OAI21_X1  g156(.A(G651), .B1(new_n511), .B2(G74), .ZN(new_n582));
  AND2_X1   g157(.A1(new_n515), .A2(G543), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n583), .A2(G49), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n581), .A2(new_n582), .A3(new_n584), .ZN(G288));
  NAND2_X1  g160(.A1(new_n583), .A2(G48), .ZN(new_n586));
  XNOR2_X1  g161(.A(new_n586), .B(KEYINPUT78), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n522), .A2(G86), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n511), .A2(G61), .ZN(new_n589));
  NAND2_X1  g164(.A1(G73), .A2(G543), .ZN(new_n590));
  AOI21_X1  g165(.A(new_n513), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT77), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n591), .A2(new_n592), .ZN(new_n595));
  OAI211_X1 g170(.A(new_n587), .B(new_n588), .C1(new_n594), .C2(new_n595), .ZN(G305));
  NAND2_X1  g171(.A1(new_n522), .A2(G85), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n583), .A2(G47), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n511), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n599));
  OAI211_X1 g174(.A(new_n597), .B(new_n598), .C1(new_n513), .C2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT79), .ZN(new_n601));
  XNOR2_X1  g176(.A(new_n600), .B(new_n601), .ZN(G290));
  INV_X1    g177(.A(KEYINPUT10), .ZN(new_n603));
  INV_X1    g178(.A(G92), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n516), .B2(new_n604), .ZN(new_n605));
  NAND4_X1  g180(.A1(new_n511), .A2(KEYINPUT10), .A3(G92), .A4(new_n515), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n511), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n608));
  OR2_X1    g183(.A1(new_n608), .A2(new_n513), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n583), .A2(G54), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n607), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(G868), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(KEYINPUT75), .ZN(new_n614));
  XNOR2_X1  g189(.A(G171), .B(new_n614), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n613), .B1(new_n615), .B2(new_n612), .ZN(G321));
  XOR2_X1   g191(.A(G321), .B(KEYINPUT80), .Z(G284));
  NAND2_X1  g192(.A1(G299), .A2(new_n612), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n618), .B1(new_n578), .B2(new_n612), .ZN(G280));
  XNOR2_X1  g194(.A(G280), .B(KEYINPUT81), .ZN(G297));
  AND3_X1   g195(.A1(new_n607), .A2(new_n609), .A3(new_n610), .ZN(new_n621));
  INV_X1    g196(.A(G559), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(new_n622), .B2(G860), .ZN(G148));
  NAND2_X1  g198(.A1(new_n621), .A2(new_n622), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n624), .A2(G868), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n625), .B1(G868), .B2(new_n549), .ZN(G323));
  XNOR2_X1  g201(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g202(.A1(new_n494), .A2(new_n479), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT12), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT13), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2100), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n472), .A2(G135), .ZN(new_n632));
  INV_X1    g207(.A(G123), .ZN(new_n633));
  NOR2_X1   g208(.A1(G99), .A2(G2105), .ZN(new_n634));
  OAI21_X1  g209(.A(G2104), .B1(new_n468), .B2(G111), .ZN(new_n635));
  OAI221_X1 g210(.A(new_n632), .B1(new_n633), .B2(new_n490), .C1(new_n634), .C2(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(G2096), .Z(new_n637));
  NAND2_X1  g212(.A1(new_n631), .A2(new_n637), .ZN(G156));
  XNOR2_X1  g213(.A(G1341), .B(G1348), .ZN(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2451), .B(G2454), .ZN(new_n641));
  INV_X1    g216(.A(KEYINPUT82), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT16), .ZN(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT15), .B(G2430), .ZN(new_n645));
  AND2_X1   g220(.A1(new_n645), .A2(G2435), .ZN(new_n646));
  NOR2_X1   g221(.A1(new_n645), .A2(G2435), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2427), .B(G2438), .ZN(new_n648));
  OR3_X1    g223(.A1(new_n646), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n648), .B1(new_n646), .B2(new_n647), .ZN(new_n650));
  NAND4_X1  g225(.A1(new_n644), .A2(KEYINPUT14), .A3(new_n649), .A4(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2443), .B(G2446), .ZN(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  INV_X1    g228(.A(KEYINPUT16), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n643), .B(new_n654), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n649), .A2(new_n650), .A3(KEYINPUT14), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n651), .A2(new_n653), .A3(new_n657), .ZN(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  AOI21_X1  g234(.A(new_n653), .B1(new_n651), .B2(new_n657), .ZN(new_n660));
  OAI21_X1  g235(.A(new_n640), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n651), .A2(new_n657), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n662), .A2(new_n652), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n663), .A2(new_n639), .A3(new_n658), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n661), .A2(new_n664), .A3(G14), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(G401));
  XOR2_X1   g241(.A(G2084), .B(G2090), .Z(new_n667));
  XNOR2_X1  g242(.A(G2067), .B(G2678), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  AND2_X1   g244(.A1(new_n669), .A2(KEYINPUT17), .ZN(new_n670));
  OR2_X1    g245(.A1(new_n667), .A2(new_n668), .ZN(new_n671));
  AOI21_X1  g246(.A(KEYINPUT18), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G2072), .B(G2078), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT83), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n674), .B1(KEYINPUT18), .B2(new_n669), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n672), .B(new_n675), .Z(new_n676));
  XNOR2_X1  g251(.A(G2096), .B(G2100), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n676), .B(new_n677), .Z(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(G227));
  XNOR2_X1  g254(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1971), .B(G1976), .ZN(new_n682));
  INV_X1    g257(.A(KEYINPUT19), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1956), .B(G2474), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1961), .B(G1966), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n687), .A2(KEYINPUT84), .ZN(new_n688));
  INV_X1    g263(.A(KEYINPUT84), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n689), .B1(new_n685), .B2(new_n686), .ZN(new_n690));
  NAND3_X1  g265(.A1(new_n684), .A2(new_n688), .A3(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n691), .A2(KEYINPUT85), .ZN(new_n692));
  INV_X1    g267(.A(KEYINPUT85), .ZN(new_n693));
  NAND4_X1  g268(.A1(new_n684), .A2(new_n688), .A3(new_n693), .A4(new_n690), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(KEYINPUT20), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  AND2_X1   g272(.A1(new_n685), .A2(new_n686), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n682), .B(KEYINPUT19), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n698), .B1(new_n699), .B2(new_n687), .ZN(new_n700));
  INV_X1    g275(.A(KEYINPUT86), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n700), .B(new_n702), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n692), .A2(KEYINPUT20), .A3(new_n694), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n697), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(G1991), .B(G1996), .ZN(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  XOR2_X1   g283(.A(G1981), .B(G1986), .Z(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  NAND4_X1  g285(.A1(new_n697), .A2(new_n703), .A3(new_n706), .A4(new_n704), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n708), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n710), .B1(new_n708), .B2(new_n711), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n681), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(new_n714), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n716), .A2(new_n680), .A3(new_n712), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(new_n718), .ZN(G229));
  INV_X1    g294(.A(G16), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n720), .A2(G23), .ZN(new_n721));
  INV_X1    g296(.A(G288), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n721), .B1(new_n722), .B2(new_n720), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(KEYINPUT33), .Z(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(G1976), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n720), .A2(G22), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G166), .B2(new_n720), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n727), .A2(G1971), .ZN(new_n728));
  AND2_X1   g303(.A1(new_n727), .A2(G1971), .ZN(new_n729));
  AND2_X1   g304(.A1(new_n720), .A2(G6), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(G305), .B2(G16), .ZN(new_n731));
  XOR2_X1   g306(.A(KEYINPUT32), .B(G1981), .Z(new_n732));
  AOI211_X1 g307(.A(new_n728), .B(new_n729), .C1(new_n731), .C2(new_n732), .ZN(new_n733));
  OR2_X1    g308(.A1(new_n731), .A2(new_n732), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  OAI21_X1  g310(.A(KEYINPUT93), .B1(new_n725), .B2(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(G1976), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n724), .B(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(KEYINPUT93), .ZN(new_n739));
  NAND4_X1  g314(.A1(new_n738), .A2(new_n733), .A3(new_n739), .A4(new_n734), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n736), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g316(.A(KEYINPUT92), .B(KEYINPUT34), .ZN(new_n742));
  INV_X1    g317(.A(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n720), .A2(G24), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n600), .B(KEYINPUT79), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n745), .B1(new_n746), .B2(new_n720), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT91), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(G1986), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n736), .A2(new_n740), .A3(new_n742), .ZN(new_n750));
  INV_X1    g325(.A(KEYINPUT88), .ZN(new_n751));
  OR2_X1    g326(.A1(G95), .A2(G2105), .ZN(new_n752));
  INV_X1    g327(.A(KEYINPUT89), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n469), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  OAI221_X1 g329(.A(new_n754), .B1(new_n753), .B2(new_n752), .C1(G107), .C2(new_n468), .ZN(new_n755));
  INV_X1    g330(.A(G131), .ZN(new_n756));
  INV_X1    g331(.A(G119), .ZN(new_n757));
  OAI221_X1 g332(.A(new_n755), .B1(new_n471), .B2(new_n756), .C1(new_n757), .C2(new_n490), .ZN(new_n758));
  XOR2_X1   g333(.A(KEYINPUT87), .B(G29), .Z(new_n759));
  NAND2_X1  g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(new_n759), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n761), .A2(G25), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n751), .B1(new_n760), .B2(new_n762), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(new_n751), .B2(new_n762), .ZN(new_n764));
  XNOR2_X1  g339(.A(KEYINPUT35), .B(G1991), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT90), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n764), .B(new_n766), .ZN(new_n767));
  AND2_X1   g342(.A1(new_n767), .A2(KEYINPUT94), .ZN(new_n768));
  NAND4_X1  g343(.A1(new_n744), .A2(new_n749), .A3(new_n750), .A4(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(KEYINPUT36), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  AND2_X1   g346(.A1(new_n750), .A2(new_n768), .ZN(new_n772));
  NAND4_X1  g347(.A1(new_n772), .A2(KEYINPUT36), .A3(new_n749), .A4(new_n744), .ZN(new_n773));
  INV_X1    g348(.A(KEYINPUT96), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(G29), .B2(G33), .ZN(new_n775));
  OR3_X1    g350(.A1(new_n774), .A2(G29), .A3(G33), .ZN(new_n776));
  NAND4_X1  g351(.A1(new_n467), .A2(G139), .A3(new_n468), .A4(new_n470), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n778));
  INV_X1    g353(.A(KEYINPUT25), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n777), .A2(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(KEYINPUT97), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g358(.A1(new_n777), .A2(KEYINPUT97), .A3(new_n780), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(G115), .A2(G2104), .ZN(new_n786));
  INV_X1    g361(.A(G127), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n786), .B1(new_n476), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n788), .A2(G2105), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n785), .A2(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(G29), .ZN(new_n791));
  OAI211_X1 g366(.A(new_n775), .B(new_n776), .C1(new_n790), .C2(new_n791), .ZN(new_n792));
  INV_X1    g367(.A(G2072), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n761), .A2(G35), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(G162), .B2(new_n761), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(KEYINPUT29), .Z(new_n797));
  INV_X1    g372(.A(G2090), .ZN(new_n798));
  AOI21_X1  g373(.A(KEYINPUT28), .B1(new_n761), .B2(G26), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n761), .A2(KEYINPUT28), .A3(G26), .ZN(new_n800));
  INV_X1    g375(.A(new_n800), .ZN(new_n801));
  OR2_X1    g376(.A1(G104), .A2(G2105), .ZN(new_n802));
  OAI211_X1 g377(.A(new_n802), .B(G2104), .C1(G116), .C2(new_n468), .ZN(new_n803));
  INV_X1    g378(.A(G140), .ZN(new_n804));
  INV_X1    g379(.A(G128), .ZN(new_n805));
  OAI221_X1 g380(.A(new_n803), .B1(new_n471), .B2(new_n804), .C1(new_n805), .C2(new_n490), .ZN(new_n806));
  INV_X1    g381(.A(KEYINPUT95), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  AOI211_X1 g383(.A(new_n799), .B(new_n801), .C1(new_n808), .C2(G29), .ZN(new_n809));
  INV_X1    g384(.A(G2067), .ZN(new_n810));
  OAI22_X1  g385(.A1(new_n797), .A2(new_n798), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  AOI211_X1 g386(.A(new_n794), .B(new_n811), .C1(new_n810), .C2(new_n809), .ZN(new_n812));
  NOR2_X1   g387(.A1(G16), .A2(G21), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n813), .B1(G168), .B2(G16), .ZN(new_n814));
  INV_X1    g389(.A(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(G1966), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n720), .A2(G4), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n818), .B1(new_n621), .B2(new_n720), .ZN(new_n819));
  INV_X1    g394(.A(G1348), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(G171), .A2(G16), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(G5), .B2(G16), .ZN(new_n823));
  INV_X1    g398(.A(G1961), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n823), .A2(new_n824), .ZN(new_n826));
  XOR2_X1   g401(.A(KEYINPUT30), .B(G28), .Z(new_n827));
  OAI22_X1  g402(.A1(new_n636), .A2(new_n761), .B1(G29), .B2(new_n827), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n821), .A2(new_n825), .A3(new_n829), .ZN(new_n830));
  XOR2_X1   g405(.A(KEYINPUT31), .B(G11), .Z(new_n831));
  NAND2_X1  g406(.A1(new_n720), .A2(G19), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n832), .B1(new_n549), .B2(new_n720), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n833), .A2(G1341), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n761), .A2(G27), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n835), .B1(G164), .B2(new_n761), .ZN(new_n836));
  OR2_X1    g411(.A1(new_n836), .A2(G2078), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n836), .A2(G2078), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n833), .A2(G1341), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n837), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  NOR4_X1   g415(.A1(new_n830), .A2(new_n831), .A3(new_n834), .A4(new_n840), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n812), .A2(new_n817), .A3(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(KEYINPUT98), .B(KEYINPUT24), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(G34), .ZN(new_n844));
  OAI22_X1  g419(.A1(new_n484), .A2(new_n791), .B1(new_n759), .B2(new_n844), .ZN(new_n845));
  XOR2_X1   g420(.A(new_n845), .B(KEYINPUT99), .Z(new_n846));
  INV_X1    g421(.A(G2084), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(G299), .ZN(new_n849));
  OAI21_X1  g424(.A(KEYINPUT23), .B1(new_n849), .B2(new_n720), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n720), .A2(G20), .ZN(new_n851));
  MUX2_X1   g426(.A(KEYINPUT23), .B(new_n850), .S(new_n851), .Z(new_n852));
  OR2_X1    g427(.A1(new_n852), .A2(G1956), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n846), .A2(new_n847), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n852), .A2(G1956), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n853), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  AND2_X1   g431(.A1(new_n792), .A2(new_n793), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n857), .B1(new_n797), .B2(new_n798), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n858), .B1(new_n816), .B2(new_n815), .ZN(new_n859));
  NOR4_X1   g434(.A1(new_n842), .A2(new_n848), .A3(new_n856), .A4(new_n859), .ZN(new_n860));
  NOR2_X1   g435(.A1(G29), .A2(G32), .ZN(new_n861));
  AND2_X1   g436(.A1(new_n467), .A2(new_n470), .ZN(new_n862));
  NAND4_X1  g437(.A1(new_n862), .A2(KEYINPUT100), .A3(G129), .A4(G2105), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT100), .ZN(new_n864));
  INV_X1    g439(.A(G129), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n864), .B1(new_n490), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n863), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g442(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n868));
  XOR2_X1   g443(.A(new_n868), .B(KEYINPUT26), .Z(new_n869));
  NAND2_X1  g444(.A1(new_n479), .A2(G105), .ZN(new_n870));
  INV_X1    g445(.A(G141), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n870), .B1(new_n471), .B2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n867), .A2(new_n869), .A3(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n861), .B1(new_n875), .B2(G29), .ZN(new_n876));
  XNOR2_X1  g451(.A(KEYINPUT27), .B(G1996), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n876), .B(new_n877), .ZN(new_n878));
  NAND4_X1  g453(.A1(new_n771), .A2(new_n773), .A3(new_n860), .A4(new_n878), .ZN(G150));
  INV_X1    g454(.A(G150), .ZN(G311));
  AOI22_X1  g455(.A1(new_n522), .A2(G93), .B1(new_n583), .B2(G55), .ZN(new_n881));
  AOI22_X1  g456(.A1(new_n511), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n881), .B1(new_n513), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n883), .A2(G860), .ZN(new_n884));
  XOR2_X1   g459(.A(new_n884), .B(KEYINPUT37), .Z(new_n885));
  OR2_X1    g460(.A1(new_n883), .A2(new_n549), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n883), .A2(new_n549), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(KEYINPUT39), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n621), .A2(G559), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(KEYINPUT38), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n889), .B(new_n891), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n885), .B1(new_n892), .B2(G860), .ZN(G145));
  AOI21_X1  g468(.A(new_n872), .B1(new_n863), .B2(new_n866), .ZN(new_n894));
  AOI22_X1  g469(.A1(new_n783), .A2(new_n784), .B1(G2105), .B2(new_n788), .ZN(new_n895));
  OAI211_X1 g470(.A(new_n869), .B(new_n894), .C1(new_n895), .C2(KEYINPUT101), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT101), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n790), .A2(new_n874), .A3(new_n897), .ZN(new_n898));
  AND3_X1   g473(.A1(new_n896), .A2(new_n898), .A3(new_n808), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n808), .B1(new_n896), .B2(new_n898), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n504), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n896), .A2(new_n898), .ZN(new_n902));
  INV_X1    g477(.A(new_n808), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n896), .A2(new_n898), .A3(new_n808), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n904), .A2(G164), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n901), .A2(new_n906), .ZN(new_n907));
  OR2_X1    g482(.A1(G106), .A2(G2105), .ZN(new_n908));
  OAI211_X1 g483(.A(new_n908), .B(G2104), .C1(G118), .C2(new_n468), .ZN(new_n909));
  INV_X1    g484(.A(G142), .ZN(new_n910));
  INV_X1    g485(.A(G130), .ZN(new_n911));
  OAI221_X1 g486(.A(new_n909), .B1(new_n471), .B2(new_n910), .C1(new_n911), .C2(new_n490), .ZN(new_n912));
  XOR2_X1   g487(.A(new_n912), .B(new_n629), .Z(new_n913));
  INV_X1    g488(.A(new_n758), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n913), .B(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT102), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n907), .A2(new_n917), .ZN(new_n918));
  XNOR2_X1  g493(.A(G162), .B(new_n484), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n919), .B(new_n636), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n901), .A2(new_n906), .A3(new_n916), .A4(new_n915), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n918), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(G37), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(new_n915), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n907), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n901), .A2(new_n906), .A3(new_n915), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n920), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  OR3_X1    g503(.A1(new_n924), .A2(KEYINPUT103), .A3(new_n928), .ZN(new_n929));
  OAI21_X1  g504(.A(KEYINPUT103), .B1(new_n924), .B2(new_n928), .ZN(new_n930));
  AND3_X1   g505(.A1(new_n929), .A2(KEYINPUT40), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(KEYINPUT40), .B1(new_n929), .B2(new_n930), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n931), .A2(new_n932), .ZN(G395));
  NAND2_X1  g508(.A1(new_n883), .A2(new_n612), .ZN(new_n934));
  XOR2_X1   g509(.A(new_n888), .B(new_n624), .Z(new_n935));
  NAND2_X1  g510(.A1(G299), .A2(new_n621), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n569), .A2(new_n563), .A3(G651), .ZN(new_n937));
  OAI21_X1  g512(.A(KEYINPUT74), .B1(new_n571), .B2(new_n513), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n611), .A2(new_n939), .A3(new_n560), .A4(new_n562), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n936), .A2(new_n940), .A3(KEYINPUT104), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT104), .ZN(new_n942));
  NAND3_X1  g517(.A1(G299), .A2(new_n621), .A3(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n935), .A2(new_n945), .ZN(new_n946));
  OR2_X1    g521(.A1(new_n946), .A2(KEYINPUT105), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(KEYINPUT105), .ZN(new_n948));
  AOI21_X1  g523(.A(KEYINPUT41), .B1(new_n936), .B2(new_n940), .ZN(new_n949));
  XNOR2_X1  g524(.A(KEYINPUT106), .B(KEYINPUT41), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n949), .B1(new_n944), .B2(new_n950), .ZN(new_n951));
  OAI211_X1 g526(.A(new_n947), .B(new_n948), .C1(new_n951), .C2(new_n935), .ZN(new_n952));
  NOR2_X1   g527(.A1(G303), .A2(new_n722), .ZN(new_n953));
  NOR2_X1   g528(.A1(G166), .A2(G288), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(G305), .ZN(new_n956));
  OR2_X1    g531(.A1(new_n591), .A2(new_n592), .ZN(new_n957));
  AOI22_X1  g532(.A1(new_n957), .A2(new_n593), .B1(G86), .B2(new_n522), .ZN(new_n958));
  OAI211_X1 g533(.A(new_n958), .B(new_n587), .C1(new_n953), .C2(new_n954), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n956), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(G290), .A2(KEYINPUT107), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT107), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n746), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n960), .A2(new_n964), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n956), .A2(new_n961), .A3(new_n963), .A4(new_n959), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  XOR2_X1   g542(.A(new_n967), .B(KEYINPUT42), .Z(new_n968));
  XNOR2_X1  g543(.A(new_n952), .B(new_n968), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n934), .B1(new_n969), .B2(new_n612), .ZN(G295));
  OAI21_X1  g545(.A(new_n934), .B1(new_n969), .B2(new_n612), .ZN(G331));
  INV_X1    g546(.A(KEYINPUT44), .ZN(new_n972));
  INV_X1    g547(.A(G171), .ZN(new_n973));
  INV_X1    g548(.A(new_n526), .ZN(new_n974));
  AND3_X1   g549(.A1(new_n509), .A2(KEYINPUT5), .A3(G543), .ZN(new_n975));
  AOI21_X1  g550(.A(KEYINPUT5), .B1(new_n509), .B2(G543), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n530), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(KEYINPUT70), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n511), .A2(new_n528), .A3(new_n530), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n535), .B1(new_n980), .B2(new_n527), .ZN(new_n981));
  INV_X1    g556(.A(new_n536), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n974), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(new_n576), .ZN(new_n984));
  NAND2_X1  g559(.A1(G168), .A2(KEYINPUT76), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n973), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n615), .A2(new_n983), .ZN(new_n987));
  NOR3_X1   g562(.A1(new_n986), .A2(new_n987), .A3(new_n888), .ZN(new_n988));
  INV_X1    g563(.A(new_n888), .ZN(new_n989));
  OAI21_X1  g564(.A(G171), .B1(new_n575), .B2(new_n577), .ZN(new_n990));
  NAND2_X1  g565(.A1(G301), .A2(G168), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n989), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n950), .B1(new_n988), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n936), .A2(new_n940), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n888), .B1(new_n986), .B2(new_n987), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n990), .A2(new_n989), .A3(new_n991), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n994), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  AOI22_X1  g572(.A1(new_n945), .A2(new_n993), .B1(new_n997), .B2(KEYINPUT41), .ZN(new_n998));
  INV_X1    g573(.A(new_n967), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n951), .B1(new_n988), .B2(new_n992), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n995), .A2(new_n944), .A3(new_n996), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n967), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT108), .ZN(new_n1003));
  OAI22_X1  g578(.A1(new_n998), .A2(new_n999), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n995), .A2(new_n996), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n944), .B1(new_n1005), .B2(new_n950), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT41), .ZN(new_n1007));
  AOI211_X1 g582(.A(new_n1007), .B(new_n994), .C1(new_n995), .C2(new_n996), .ZN(new_n1008));
  OAI211_X1 g583(.A(KEYINPUT108), .B(new_n967), .C1(new_n1006), .C2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1004), .A2(new_n923), .A3(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n972), .B1(new_n1010), .B2(KEYINPUT43), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1002), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT43), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1000), .A2(new_n967), .A3(new_n1001), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n1012), .A2(new_n1013), .A3(new_n923), .A4(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(KEYINPUT109), .ZN(new_n1016));
  OR2_X1    g591(.A1(new_n1015), .A2(KEYINPUT109), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1011), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1004), .A2(new_n1013), .A3(new_n923), .A4(new_n1009), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1012), .A2(new_n923), .A3(new_n1014), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(KEYINPUT43), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(new_n972), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1018), .A2(new_n1023), .ZN(G397));
  INV_X1    g599(.A(G1384), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n504), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT45), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n473), .A2(G40), .A3(new_n480), .A4(new_n483), .ZN(new_n1029));
  NOR3_X1   g604(.A1(new_n1028), .A2(G1996), .A3(new_n1029), .ZN(new_n1030));
  XOR2_X1   g605(.A(new_n1030), .B(KEYINPUT110), .Z(new_n1031));
  NOR2_X1   g606(.A1(new_n1031), .A2(new_n874), .ZN(new_n1032));
  XNOR2_X1  g607(.A(new_n808), .B(new_n810), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n874), .A2(G1996), .ZN(new_n1034));
  AOI211_X1 g609(.A(new_n1029), .B(new_n1028), .C1(new_n1033), .C2(new_n1034), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1036));
  XNOR2_X1  g611(.A(new_n758), .B(new_n765), .ZN(new_n1037));
  AND2_X1   g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  OR3_X1    g613(.A1(new_n1032), .A2(new_n1035), .A3(new_n1038), .ZN(new_n1039));
  XNOR2_X1  g614(.A(G290), .B(G1986), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1039), .B1(new_n1036), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT115), .ZN(new_n1042));
  NAND2_X1  g617(.A1(G303), .A2(G8), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT55), .ZN(new_n1044));
  AND3_X1   g619(.A1(new_n1043), .A2(KEYINPUT113), .A3(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(KEYINPUT113), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1046));
  NAND3_X1  g621(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1047), .ZN(new_n1048));
  NOR3_X1   g623(.A1(new_n1045), .A2(new_n1046), .A3(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT50), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n504), .A2(new_n1051), .A3(new_n1025), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(KEYINPUT111), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT111), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n504), .A2(new_n1054), .A3(new_n1051), .A4(new_n1025), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1053), .A2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1029), .B1(KEYINPUT50), .B2(new_n1026), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1056), .A2(new_n798), .A3(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1029), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n504), .A2(KEYINPUT45), .A3(new_n1025), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1028), .A2(new_n1059), .A3(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(G1971), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT112), .ZN(new_n1064));
  AND3_X1   g639(.A1(new_n1058), .A2(new_n1063), .A3(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1064), .B1(new_n1058), .B2(new_n1063), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1050), .B1(new_n1067), .B2(G8), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT114), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1026), .A2(new_n1029), .ZN(new_n1070));
  INV_X1    g645(.A(G8), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1069), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  OAI211_X1 g647(.A(KEYINPUT114), .B(G8), .C1(new_n1026), .C2(new_n1029), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n722), .A2(G1976), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(KEYINPUT52), .ZN(new_n1077));
  NAND2_X1  g652(.A1(G305), .A2(G1981), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT49), .ZN(new_n1079));
  INV_X1    g654(.A(G1981), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n958), .A2(new_n1080), .A3(new_n587), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1078), .A2(new_n1079), .A3(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1079), .B1(new_n1078), .B2(new_n1081), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1074), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g660(.A(KEYINPUT52), .B1(G288), .B2(new_n737), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1074), .A2(new_n1075), .A3(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1077), .A2(new_n1085), .A3(new_n1087), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1042), .B1(new_n1068), .B2(new_n1088), .ZN(new_n1089));
  AND3_X1   g664(.A1(new_n1077), .A2(new_n1085), .A3(new_n1087), .ZN(new_n1090));
  NOR3_X1   g665(.A1(new_n1065), .A2(new_n1066), .A3(new_n1071), .ZN(new_n1091));
  OAI211_X1 g666(.A(new_n1090), .B(KEYINPUT115), .C1(new_n1091), .C2(new_n1050), .ZN(new_n1092));
  NOR4_X1   g667(.A1(new_n1065), .A2(new_n1066), .A3(new_n1071), .A4(new_n1049), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT63), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1056), .A2(new_n847), .A3(new_n1057), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1061), .A2(new_n816), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1071), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(new_n578), .ZN(new_n1098));
  NOR3_X1   g673(.A1(new_n1093), .A2(new_n1094), .A3(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1089), .A2(new_n1092), .A3(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1026), .A2(KEYINPUT50), .ZN(new_n1101));
  AND3_X1   g676(.A1(new_n1101), .A2(new_n1059), .A3(new_n1052), .ZN(new_n1102));
  AOI22_X1  g677(.A1(new_n1102), .A2(new_n798), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1049), .B1(new_n1103), .B2(new_n1071), .ZN(new_n1104));
  AND4_X1   g679(.A1(new_n1104), .A2(new_n1077), .A3(new_n1085), .A4(new_n1087), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1091), .A2(new_n1050), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1094), .B1(new_n1107), .B2(new_n1098), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1100), .A2(new_n1108), .ZN(new_n1109));
  NOR2_X1   g684(.A1(G305), .A2(G1981), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1080), .B1(new_n958), .B2(new_n587), .ZN(new_n1111));
  OAI21_X1  g686(.A(KEYINPUT49), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1112), .A2(new_n1082), .ZN(new_n1113));
  AOI21_X1  g688(.A(G1976), .B1(new_n1113), .B2(new_n1074), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1110), .B1(new_n1114), .B2(new_n722), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1074), .ZN(new_n1116));
  OAI22_X1  g691(.A1(new_n1106), .A2(new_n1088), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(G2078), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1028), .A2(new_n1059), .A3(new_n1118), .A4(new_n1060), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT53), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT122), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(new_n824), .ZN(new_n1125));
  OR2_X1    g700(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1119), .A2(KEYINPUT122), .A3(new_n1120), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1123), .A2(new_n1125), .A3(new_n1126), .A4(new_n1127), .ZN(new_n1128));
  AND2_X1   g703(.A1(new_n1128), .A2(new_n615), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1131), .A2(G8), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n983), .A2(G8), .ZN(new_n1133));
  AND2_X1   g708(.A1(new_n1133), .A2(KEYINPUT120), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1134), .A2(KEYINPUT51), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1135), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1132), .A2(new_n1136), .A3(new_n1133), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1097), .A2(new_n983), .ZN(new_n1138));
  OAI211_X1 g713(.A(new_n1135), .B(G8), .C1(new_n1131), .C2(new_n983), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1137), .A2(new_n1138), .A3(new_n1139), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1130), .B1(new_n1140), .B2(KEYINPUT62), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT62), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1137), .A2(new_n1139), .A3(new_n1142), .A4(new_n1138), .ZN(new_n1143));
  AND3_X1   g718(.A1(new_n1143), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1117), .B1(new_n1141), .B2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1109), .A2(new_n1145), .ZN(new_n1146));
  AND3_X1   g721(.A1(new_n1123), .A2(new_n1125), .A3(new_n1127), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT124), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1147), .A2(new_n1148), .A3(G301), .A4(new_n1126), .ZN(new_n1149));
  OAI21_X1  g724(.A(KEYINPUT124), .B1(new_n1128), .B2(new_n615), .ZN(new_n1150));
  AND2_X1   g725(.A1(new_n1028), .A2(new_n1060), .ZN(new_n1151));
  OR2_X1    g726(.A1(new_n1059), .A2(KEYINPUT123), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1059), .A2(KEYINPUT123), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n1120), .A2(G2078), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1151), .A2(new_n1152), .A3(new_n1153), .A4(new_n1154), .ZN(new_n1155));
  NAND4_X1  g730(.A1(new_n1123), .A2(new_n1125), .A3(new_n1127), .A4(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1156), .A2(G171), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1149), .A2(new_n1150), .A3(KEYINPUT54), .A4(new_n1157), .ZN(new_n1158));
  XOR2_X1   g733(.A(KEYINPUT121), .B(KEYINPUT54), .Z(new_n1159));
  NOR2_X1   g734(.A1(new_n1156), .A2(new_n615), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1159), .B1(new_n1129), .B2(new_n1160), .ZN(new_n1161));
  NAND4_X1  g736(.A1(new_n1104), .A2(new_n1077), .A3(new_n1085), .A4(new_n1087), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1093), .A2(new_n1162), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n1158), .A2(new_n1161), .A3(new_n1163), .A4(new_n1140), .ZN(new_n1164));
  XOR2_X1   g739(.A(G299), .B(KEYINPUT57), .Z(new_n1165));
  XNOR2_X1  g740(.A(KEYINPUT56), .B(G2072), .ZN(new_n1166));
  NAND4_X1  g741(.A1(new_n1028), .A2(new_n1059), .A3(new_n1060), .A4(new_n1166), .ZN(new_n1167));
  OR2_X1    g742(.A1(new_n1167), .A2(KEYINPUT116), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1167), .A2(KEYINPUT116), .ZN(new_n1169));
  AND2_X1   g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1057), .A2(new_n1052), .ZN(new_n1171));
  INV_X1    g746(.A(G1956), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1165), .B1(new_n1170), .B2(new_n1173), .ZN(new_n1174));
  AOI22_X1  g749(.A1(new_n1124), .A2(new_n820), .B1(new_n810), .B2(new_n1070), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1175), .A2(KEYINPUT60), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1176), .A2(KEYINPUT119), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT119), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1175), .A2(new_n1178), .A3(KEYINPUT60), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1177), .A2(new_n621), .A3(new_n1179), .ZN(new_n1180));
  OR2_X1    g755(.A1(new_n1175), .A2(KEYINPUT60), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1176), .A2(KEYINPUT119), .A3(new_n611), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1180), .A2(new_n1181), .A3(new_n1182), .ZN(new_n1183));
  XNOR2_X1  g758(.A(KEYINPUT58), .B(G1341), .ZN(new_n1184));
  OAI22_X1  g759(.A1(new_n1061), .A2(G1996), .B1(new_n1070), .B2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1185), .A2(new_n549), .ZN(new_n1186));
  NOR2_X1   g761(.A1(KEYINPUT117), .A2(KEYINPUT59), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  XNOR2_X1  g763(.A(KEYINPUT117), .B(KEYINPUT59), .ZN(new_n1189));
  NAND4_X1  g764(.A1(new_n1168), .A2(new_n1173), .A3(new_n1165), .A4(new_n1169), .ZN(new_n1190));
  OAI221_X1 g765(.A(new_n1188), .B1(new_n1186), .B2(new_n1189), .C1(new_n1190), .C2(KEYINPUT61), .ZN(new_n1191));
  OR2_X1    g766(.A1(KEYINPUT118), .A2(KEYINPUT61), .ZN(new_n1192));
  AND2_X1   g767(.A1(new_n1190), .A2(new_n1192), .ZN(new_n1193));
  NOR2_X1   g768(.A1(new_n1191), .A2(new_n1193), .ZN(new_n1194));
  AOI21_X1  g769(.A(new_n1174), .B1(new_n1183), .B2(new_n1194), .ZN(new_n1195));
  INV_X1    g770(.A(new_n1175), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1190), .A2(new_n1196), .A3(new_n621), .ZN(new_n1197));
  AOI21_X1  g772(.A(new_n1164), .B1(new_n1195), .B2(new_n1197), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n1041), .B1(new_n1146), .B2(new_n1198), .ZN(new_n1199));
  INV_X1    g774(.A(KEYINPUT125), .ZN(new_n1200));
  NOR2_X1   g775(.A1(new_n1200), .A2(KEYINPUT46), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1033), .A2(new_n875), .ZN(new_n1202));
  AOI21_X1  g777(.A(new_n1201), .B1(new_n1202), .B2(new_n1036), .ZN(new_n1203));
  AND3_X1   g778(.A1(new_n1031), .A2(new_n1200), .A3(KEYINPUT46), .ZN(new_n1204));
  AOI21_X1  g779(.A(new_n1031), .B1(new_n1200), .B2(KEYINPUT46), .ZN(new_n1205));
  OAI21_X1  g780(.A(new_n1203), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1206), .A2(KEYINPUT126), .ZN(new_n1207));
  INV_X1    g782(.A(KEYINPUT126), .ZN(new_n1208));
  OAI211_X1 g783(.A(new_n1208), .B(new_n1203), .C1(new_n1204), .C2(new_n1205), .ZN(new_n1209));
  NAND3_X1  g784(.A1(new_n1207), .A2(KEYINPUT47), .A3(new_n1209), .ZN(new_n1210));
  NOR4_X1   g785(.A1(new_n1032), .A2(new_n1035), .A3(new_n758), .A4(new_n765), .ZN(new_n1211));
  NOR2_X1   g786(.A1(new_n808), .A2(G2067), .ZN(new_n1212));
  OAI21_X1  g787(.A(new_n1036), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1210), .A2(new_n1213), .ZN(new_n1214));
  NOR4_X1   g789(.A1(G290), .A2(new_n1028), .A3(G1986), .A4(new_n1029), .ZN(new_n1215));
  XNOR2_X1  g790(.A(new_n1215), .B(KEYINPUT48), .ZN(new_n1216));
  NOR2_X1   g791(.A1(new_n1039), .A2(new_n1216), .ZN(new_n1217));
  AOI21_X1  g792(.A(KEYINPUT47), .B1(new_n1207), .B2(new_n1209), .ZN(new_n1218));
  NOR3_X1   g793(.A1(new_n1214), .A2(new_n1217), .A3(new_n1218), .ZN(new_n1219));
  NAND2_X1  g794(.A1(new_n1199), .A2(new_n1219), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g795(.A1(new_n665), .A2(new_n678), .ZN(new_n1222));
  AOI211_X1 g796(.A(new_n462), .B(new_n1222), .C1(new_n717), .C2(new_n715), .ZN(new_n1223));
  OAI21_X1  g797(.A(new_n1223), .B1(new_n924), .B2(new_n928), .ZN(new_n1224));
  AOI211_X1 g798(.A(KEYINPUT127), .B(new_n1224), .C1(new_n1019), .C2(new_n1021), .ZN(new_n1225));
  INV_X1    g799(.A(KEYINPUT127), .ZN(new_n1226));
  INV_X1    g800(.A(new_n1224), .ZN(new_n1227));
  AOI21_X1  g801(.A(new_n1226), .B1(new_n1022), .B2(new_n1227), .ZN(new_n1228));
  NOR2_X1   g802(.A1(new_n1225), .A2(new_n1228), .ZN(G308));
  NAND2_X1  g803(.A1(new_n1022), .A2(new_n1227), .ZN(new_n1230));
  NAND2_X1  g804(.A1(new_n1230), .A2(KEYINPUT127), .ZN(new_n1231));
  NAND3_X1  g805(.A1(new_n1022), .A2(new_n1226), .A3(new_n1227), .ZN(new_n1232));
  NAND2_X1  g806(.A1(new_n1231), .A2(new_n1232), .ZN(G225));
endmodule


