//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 1 0 0 0 1 0 1 1 1 1 1 0 1 1 1 1 1 1 1 1 1 0 0 1 1 1 1 1 1 0 0 1 1 1 0 1 1 0 0 1 0 0 1 0 1 1 1 1 0 0 1 1 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:55 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n722, new_n723, new_n724, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n734, new_n735, new_n736,
    new_n737, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n761, new_n762, new_n763, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n900, new_n901, new_n902, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n931, new_n932, new_n933, new_n934, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995;
  NAND2_X1  g000(.A1(KEYINPUT2), .A2(G113), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  NOR2_X1   g002(.A1(KEYINPUT2), .A2(G113), .ZN(new_n189));
  OAI21_X1  g003(.A(KEYINPUT69), .B1(new_n188), .B2(new_n189), .ZN(new_n190));
  OR2_X1    g004(.A1(KEYINPUT2), .A2(G113), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT69), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n191), .A2(new_n192), .A3(new_n187), .ZN(new_n193));
  AND2_X1   g007(.A1(new_n190), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G116), .ZN(new_n195));
  INV_X1    g009(.A(G119), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(G116), .A2(G119), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT70), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n197), .A2(KEYINPUT70), .A3(new_n198), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  OAI21_X1  g017(.A(KEYINPUT71), .B1(new_n194), .B2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n190), .A2(new_n193), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT71), .ZN(new_n206));
  NAND4_X1  g020(.A1(new_n205), .A2(new_n206), .A3(new_n201), .A4(new_n202), .ZN(new_n207));
  INV_X1    g021(.A(new_n199), .ZN(new_n208));
  NOR3_X1   g022(.A1(new_n208), .A2(new_n189), .A3(new_n188), .ZN(new_n209));
  INV_X1    g023(.A(new_n209), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n204), .A2(new_n207), .A3(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G146), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n213), .A2(G143), .ZN(new_n214));
  OR2_X1    g028(.A1(KEYINPUT64), .A2(G143), .ZN(new_n215));
  NAND2_X1  g029(.A1(KEYINPUT64), .A2(G143), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n214), .B1(new_n217), .B2(new_n213), .ZN(new_n218));
  XNOR2_X1  g032(.A(KEYINPUT0), .B(G128), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(G143), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n221), .A2(G146), .ZN(new_n222));
  AND2_X1   g036(.A1(KEYINPUT64), .A2(G143), .ZN(new_n223));
  NOR2_X1   g037(.A1(KEYINPUT64), .A2(G143), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n222), .B1(new_n225), .B2(G146), .ZN(new_n226));
  NAND2_X1  g040(.A1(KEYINPUT0), .A2(G128), .ZN(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n220), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT11), .ZN(new_n230));
  INV_X1    g044(.A(G134), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n230), .B1(new_n231), .B2(G137), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(G137), .ZN(new_n233));
  INV_X1    g047(.A(G137), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n234), .A2(KEYINPUT11), .A3(G134), .ZN(new_n235));
  AND3_X1   g049(.A1(new_n232), .A2(new_n233), .A3(new_n235), .ZN(new_n236));
  XOR2_X1   g050(.A(KEYINPUT65), .B(G131), .Z(new_n237));
  AOI21_X1  g051(.A(KEYINPUT66), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n232), .A2(new_n233), .A3(new_n235), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT66), .ZN(new_n240));
  XNOR2_X1  g054(.A(KEYINPUT65), .B(G131), .ZN(new_n241));
  NOR3_X1   g055(.A1(new_n239), .A2(new_n240), .A3(new_n241), .ZN(new_n242));
  AND3_X1   g056(.A1(new_n239), .A2(KEYINPUT67), .A3(G131), .ZN(new_n243));
  AOI21_X1  g057(.A(KEYINPUT67), .B1(new_n239), .B2(G131), .ZN(new_n244));
  OAI22_X1  g058(.A1(new_n238), .A2(new_n242), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n229), .A2(new_n245), .ZN(new_n246));
  AND2_X1   g060(.A1(new_n235), .A2(new_n233), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n247), .A2(new_n237), .A3(KEYINPUT66), .A4(new_n232), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n240), .B1(new_n239), .B2(new_n241), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT1), .ZN(new_n251));
  OAI21_X1  g065(.A(G128), .B1(new_n222), .B2(new_n251), .ZN(new_n252));
  AOI21_X1  g066(.A(G146), .B1(new_n215), .B2(new_n216), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n252), .B1(new_n253), .B2(new_n214), .ZN(new_n254));
  INV_X1    g068(.A(new_n222), .ZN(new_n255));
  INV_X1    g069(.A(G128), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n256), .A2(KEYINPUT1), .ZN(new_n257));
  OAI211_X1 g071(.A(new_n255), .B(new_n257), .C1(new_n217), .C2(new_n213), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n254), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n233), .A2(KEYINPUT68), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n260), .B1(new_n231), .B2(G137), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n233), .A2(KEYINPUT68), .ZN(new_n262));
  OAI21_X1  g076(.A(G131), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n250), .A2(new_n259), .A3(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n212), .A2(new_n246), .A3(new_n264), .ZN(new_n265));
  OR2_X1    g079(.A1(KEYINPUT74), .A2(G237), .ZN(new_n266));
  NAND2_X1  g080(.A1(KEYINPUT74), .A2(G237), .ZN(new_n267));
  AOI21_X1  g081(.A(G953), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(G210), .ZN(new_n269));
  XNOR2_X1  g083(.A(KEYINPUT75), .B(KEYINPUT27), .ZN(new_n270));
  XNOR2_X1  g084(.A(new_n269), .B(new_n270), .ZN(new_n271));
  XNOR2_X1  g085(.A(KEYINPUT26), .B(G101), .ZN(new_n272));
  XNOR2_X1  g086(.A(new_n271), .B(new_n272), .ZN(new_n273));
  AND2_X1   g087(.A1(new_n265), .A2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT67), .ZN(new_n275));
  INV_X1    g089(.A(G131), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n275), .B1(new_n236), .B2(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n239), .A2(KEYINPUT67), .A3(G131), .ZN(new_n278));
  AOI22_X1  g092(.A1(new_n277), .A2(new_n278), .B1(new_n248), .B2(new_n249), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n226), .A2(new_n228), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n280), .B1(new_n218), .B2(new_n219), .ZN(new_n281));
  OAI211_X1 g095(.A(new_n264), .B(KEYINPUT30), .C1(new_n279), .C2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT72), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n246), .A2(KEYINPUT72), .A3(KEYINPUT30), .A4(new_n264), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT73), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n246), .A2(new_n264), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT30), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n212), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  AND3_X1   g104(.A1(new_n286), .A2(new_n287), .A3(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n287), .B1(new_n286), .B2(new_n290), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n274), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(KEYINPUT31), .ZN(new_n294));
  INV_X1    g108(.A(new_n273), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT28), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n288), .A2(new_n211), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n296), .B1(new_n297), .B2(new_n265), .ZN(new_n298));
  AND2_X1   g112(.A1(new_n265), .A2(new_n296), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n295), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT31), .ZN(new_n301));
  OAI211_X1 g115(.A(new_n301), .B(new_n274), .C1(new_n291), .C2(new_n292), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n294), .A2(new_n300), .A3(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(KEYINPUT76), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT76), .ZN(new_n305));
  NAND4_X1  g119(.A1(new_n294), .A2(new_n300), .A3(new_n305), .A4(new_n302), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  NOR2_X1   g121(.A1(G472), .A2(G902), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT32), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  OAI211_X1 g125(.A(new_n265), .B(new_n295), .C1(new_n291), .C2(new_n292), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n273), .B1(new_n298), .B2(new_n299), .ZN(new_n313));
  AOI21_X1  g127(.A(KEYINPUT29), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  OAI21_X1  g128(.A(KEYINPUT77), .B1(new_n298), .B2(new_n299), .ZN(new_n315));
  OR2_X1    g129(.A1(new_n299), .A2(KEYINPUT77), .ZN(new_n316));
  NAND4_X1  g130(.A1(new_n315), .A2(new_n316), .A3(KEYINPUT29), .A4(new_n273), .ZN(new_n317));
  INV_X1    g131(.A(G902), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  OAI21_X1  g133(.A(G472), .B1(new_n314), .B2(new_n319), .ZN(new_n320));
  XNOR2_X1  g134(.A(new_n320), .B(KEYINPUT78), .ZN(new_n321));
  INV_X1    g135(.A(new_n308), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n322), .B1(new_n304), .B2(new_n306), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(KEYINPUT32), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n311), .A2(new_n321), .A3(new_n324), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n196), .A2(G128), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(KEYINPUT23), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT79), .ZN(new_n328));
  AOI22_X1  g142(.A1(new_n328), .A2(KEYINPUT23), .B1(new_n196), .B2(G128), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n329), .B1(new_n328), .B2(KEYINPUT23), .ZN(new_n330));
  XNOR2_X1  g144(.A(new_n330), .B(KEYINPUT80), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n327), .B1(new_n331), .B2(new_n326), .ZN(new_n332));
  XOR2_X1   g146(.A(KEYINPUT83), .B(G110), .Z(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  XNOR2_X1  g148(.A(G119), .B(G128), .ZN(new_n335));
  XNOR2_X1  g149(.A(KEYINPUT24), .B(G110), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  OAI22_X1  g151(.A1(new_n332), .A2(new_n334), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT16), .ZN(new_n339));
  XNOR2_X1  g153(.A(KEYINPUT81), .B(G125), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(G140), .ZN(new_n341));
  OR2_X1    g155(.A1(G125), .A2(G140), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n339), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(G140), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n340), .A2(KEYINPUT82), .A3(new_n339), .A4(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT82), .ZN(new_n347));
  INV_X1    g161(.A(new_n340), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n339), .A2(new_n345), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n347), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n344), .A2(G146), .A3(new_n346), .A4(new_n350), .ZN(new_n351));
  XNOR2_X1  g165(.A(G125), .B(G140), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(new_n213), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n338), .A2(new_n351), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n332), .A2(G110), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n350), .A2(new_n346), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n213), .B1(new_n356), .B2(new_n343), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(new_n351), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n337), .A2(new_n335), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n355), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n354), .A2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(G953), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n362), .A2(G221), .A3(G234), .ZN(new_n363));
  XNOR2_X1  g177(.A(new_n363), .B(KEYINPUT22), .ZN(new_n364));
  XNOR2_X1  g178(.A(new_n364), .B(G137), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n361), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n354), .A2(new_n360), .A3(new_n365), .ZN(new_n368));
  AND2_X1   g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT25), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n369), .A2(new_n370), .A3(new_n318), .ZN(new_n371));
  INV_X1    g185(.A(G234), .ZN(new_n372));
  OAI21_X1  g186(.A(G217), .B1(new_n372), .B2(G902), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n367), .A2(new_n368), .A3(new_n318), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n373), .B1(new_n374), .B2(KEYINPUT25), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n371), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n373), .A2(new_n318), .ZN(new_n377));
  XOR2_X1   g191(.A(new_n377), .B(KEYINPUT84), .Z(new_n378));
  NAND2_X1  g192(.A1(new_n369), .A2(new_n378), .ZN(new_n379));
  AND2_X1   g193(.A1(new_n376), .A2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(G104), .ZN(new_n381));
  OAI21_X1  g195(.A(KEYINPUT3), .B1(new_n381), .B2(G107), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT3), .ZN(new_n383));
  INV_X1    g197(.A(G107), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n383), .A2(new_n384), .A3(G104), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n381), .A2(G107), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n382), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT4), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n387), .A2(new_n388), .A3(G101), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(KEYINPUT86), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT86), .ZN(new_n391));
  NAND4_X1  g205(.A1(new_n387), .A2(new_n391), .A3(new_n388), .A4(G101), .ZN(new_n392));
  INV_X1    g206(.A(G101), .ZN(new_n393));
  NAND4_X1  g207(.A1(new_n382), .A2(new_n385), .A3(new_n393), .A4(new_n386), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n388), .B1(new_n387), .B2(G101), .ZN(new_n395));
  AOI22_X1  g209(.A1(new_n390), .A2(new_n392), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n211), .A2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(G113), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n195), .A2(KEYINPUT5), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n398), .B1(new_n399), .B2(new_n196), .ZN(new_n400));
  INV_X1    g214(.A(new_n203), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT5), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n400), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n381), .A2(G107), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n384), .A2(G104), .ZN(new_n405));
  OAI21_X1  g219(.A(G101), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n394), .A2(new_n406), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n209), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n403), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n397), .A2(new_n409), .ZN(new_n410));
  XNOR2_X1  g224(.A(G110), .B(G122), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  AOI22_X1  g227(.A1(new_n211), .A2(new_n396), .B1(new_n403), .B2(new_n408), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(new_n411), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n413), .A2(KEYINPUT6), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n259), .A2(new_n348), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n417), .B1(new_n281), .B2(new_n348), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n362), .A2(G224), .ZN(new_n419));
  XNOR2_X1  g233(.A(new_n418), .B(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT6), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n410), .A2(new_n421), .A3(new_n412), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n416), .A2(new_n420), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(KEYINPUT92), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT92), .ZN(new_n425));
  NAND4_X1  g239(.A1(new_n416), .A2(new_n420), .A3(new_n425), .A4(new_n422), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n419), .A2(KEYINPUT7), .ZN(new_n428));
  XOR2_X1   g242(.A(new_n418), .B(new_n428), .Z(new_n429));
  XOR2_X1   g243(.A(new_n411), .B(KEYINPUT8), .Z(new_n430));
  NAND2_X1  g244(.A1(new_n403), .A2(new_n210), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(new_n407), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n400), .B1(new_n208), .B2(new_n402), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n408), .A2(new_n433), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n430), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n429), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g250(.A(G902), .B1(new_n436), .B2(new_n415), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n427), .A2(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(G210), .B1(G237), .B2(G902), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n427), .A2(new_n439), .A3(new_n437), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  XNOR2_X1  g257(.A(G110), .B(G140), .ZN(new_n444));
  XNOR2_X1  g258(.A(new_n444), .B(KEYINPUT85), .ZN(new_n445));
  AND2_X1   g259(.A1(new_n362), .A2(G227), .ZN(new_n446));
  XOR2_X1   g260(.A(new_n445), .B(new_n446), .Z(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n213), .B1(new_n223), .B2(new_n224), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n256), .B1(new_n449), .B2(KEYINPUT1), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n258), .B1(new_n450), .B2(new_n226), .ZN(new_n451));
  INV_X1    g265(.A(new_n407), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT10), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n259), .A2(KEYINPUT10), .A3(new_n452), .ZN(new_n456));
  AND2_X1   g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n396), .A2(new_n229), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n279), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  XNOR2_X1  g273(.A(new_n245), .B(KEYINPUT87), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n458), .A2(new_n455), .A3(new_n456), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n448), .B1(new_n459), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(KEYINPUT91), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT91), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n465), .B(new_n448), .C1(new_n459), .C2(new_n462), .ZN(new_n466));
  OR2_X1    g280(.A1(new_n460), .A2(new_n461), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n254), .A2(new_n407), .A3(new_n258), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT88), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n254), .A2(new_n407), .A3(KEYINPUT88), .A4(new_n258), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n470), .A2(new_n453), .A3(new_n471), .ZN(new_n472));
  NAND4_X1  g286(.A1(new_n472), .A2(KEYINPUT89), .A3(KEYINPUT12), .A4(new_n245), .ZN(new_n473));
  AOI22_X1  g287(.A1(new_n469), .A2(new_n468), .B1(new_n451), .B2(new_n452), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n279), .B1(new_n474), .B2(new_n471), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n473), .B1(new_n475), .B2(KEYINPUT12), .ZN(new_n476));
  AOI21_X1  g290(.A(KEYINPUT89), .B1(new_n475), .B2(KEYINPUT12), .ZN(new_n477));
  OAI211_X1 g291(.A(new_n467), .B(new_n447), .C1(new_n476), .C2(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n464), .A2(new_n466), .A3(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(G469), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n479), .A2(new_n480), .A3(new_n318), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n480), .A2(new_n318), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n467), .B1(new_n476), .B2(new_n477), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(KEYINPUT90), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT90), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n467), .B(new_n486), .C1(new_n476), .C2(new_n477), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n485), .A2(new_n487), .A3(new_n448), .ZN(new_n488));
  OR3_X1    g302(.A1(new_n459), .A2(new_n462), .A3(new_n448), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  OAI211_X1 g304(.A(new_n481), .B(new_n483), .C1(new_n490), .C2(new_n480), .ZN(new_n491));
  NAND2_X1  g305(.A1(G234), .A2(G237), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n492), .A2(G952), .A3(new_n362), .ZN(new_n493));
  XNOR2_X1  g307(.A(KEYINPUT21), .B(G898), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n492), .A2(G902), .A3(G953), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n493), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  OAI21_X1  g311(.A(G214), .B1(G237), .B2(G902), .ZN(new_n498));
  AND2_X1   g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  XNOR2_X1  g313(.A(KEYINPUT9), .B(G234), .ZN(new_n500));
  OAI21_X1  g314(.A(G221), .B1(new_n500), .B2(G902), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n443), .A2(new_n491), .A3(new_n499), .A4(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT93), .ZN(new_n503));
  XNOR2_X1  g317(.A(KEYINPUT74), .B(G237), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n504), .A2(G214), .A3(new_n362), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n503), .B1(new_n505), .B2(new_n221), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n268), .A2(KEYINPUT93), .A3(G143), .A4(G214), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n505), .A2(new_n225), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n506), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  AND2_X1   g323(.A1(KEYINPUT18), .A2(G131), .ZN(new_n510));
  AND2_X1   g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n341), .A2(new_n342), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n353), .B1(new_n512), .B2(new_n213), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n513), .B1(new_n509), .B2(new_n510), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n509), .A2(KEYINPUT17), .A3(new_n241), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n516), .A2(new_n357), .A3(new_n351), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT95), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n509), .A2(new_n241), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT17), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n506), .A2(new_n237), .A3(new_n507), .A4(new_n508), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n517), .B1(new_n518), .B2(new_n522), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n519), .A2(KEYINPUT95), .A3(new_n520), .A4(new_n521), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n515), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  XNOR2_X1  g339(.A(G113), .B(G122), .ZN(new_n526));
  XNOR2_X1  g340(.A(new_n526), .B(new_n381), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(KEYINPUT96), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n318), .B1(new_n525), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n522), .A2(new_n518), .ZN(new_n532));
  AND3_X1   g346(.A1(new_n516), .A2(new_n357), .A3(new_n351), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n532), .A2(new_n533), .A3(new_n524), .ZN(new_n534));
  INV_X1    g348(.A(new_n515), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n536), .A2(new_n529), .ZN(new_n537));
  OAI21_X1  g351(.A(G475), .B1(new_n531), .B2(new_n537), .ZN(new_n538));
  XOR2_X1   g352(.A(KEYINPUT94), .B(KEYINPUT19), .Z(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(new_n352), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT19), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n540), .B1(new_n512), .B2(new_n541), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n351), .B1(G146), .B2(new_n542), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n543), .B1(new_n519), .B2(new_n521), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n528), .B1(new_n511), .B2(new_n514), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n546), .B1(new_n536), .B2(new_n527), .ZN(new_n547));
  NOR2_X1   g361(.A1(G475), .A2(G902), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n547), .A2(KEYINPUT20), .A3(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(new_n546), .ZN(new_n550));
  OAI211_X1 g364(.A(new_n550), .B(new_n548), .C1(new_n525), .C2(new_n528), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT20), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n538), .A2(new_n549), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(KEYINPUT97), .ZN(new_n555));
  AOI21_X1  g369(.A(G902), .B1(new_n536), .B2(new_n529), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n525), .A2(new_n530), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  AOI22_X1  g372(.A1(new_n558), .A2(G475), .B1(new_n551), .B2(new_n552), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT97), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n559), .A2(new_n560), .A3(new_n549), .ZN(new_n561));
  XNOR2_X1  g375(.A(G116), .B(G122), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(new_n384), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT98), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n562), .A2(KEYINPUT98), .A3(new_n384), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT14), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n562), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n195), .A2(G122), .ZN(new_n570));
  OAI211_X1 g384(.A(new_n569), .B(G107), .C1(new_n568), .C2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n567), .A2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n225), .A2(G128), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n256), .A2(G143), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n576), .A2(G134), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n231), .B1(new_n574), .B2(new_n575), .ZN(new_n578));
  OAI211_X1 g392(.A(new_n573), .B(KEYINPUT99), .C1(new_n577), .C2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT99), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n577), .A2(new_n578), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n580), .B1(new_n581), .B2(new_n572), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n579), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n574), .A2(KEYINPUT13), .A3(new_n575), .ZN(new_n584));
  OAI211_X1 g398(.A(new_n584), .B(G134), .C1(KEYINPUT13), .C2(new_n574), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n562), .B(new_n384), .ZN(new_n586));
  OAI211_X1 g400(.A(new_n585), .B(new_n586), .C1(G134), .C2(new_n576), .ZN(new_n587));
  INV_X1    g401(.A(new_n500), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n588), .A2(G217), .A3(new_n362), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n583), .A2(new_n587), .A3(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n590), .B1(new_n583), .B2(new_n587), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n318), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  OAI21_X1  g408(.A(G478), .B1(KEYINPUT100), .B2(KEYINPUT15), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n595), .B1(KEYINPUT100), .B2(KEYINPUT15), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n583), .A2(new_n587), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(new_n589), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(new_n591), .ZN(new_n600));
  INV_X1    g414(.A(new_n596), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n600), .A2(new_n318), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n597), .A2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n555), .A2(new_n561), .A3(new_n604), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n502), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n325), .A2(new_n380), .A3(new_n606), .ZN(new_n607));
  XNOR2_X1  g421(.A(KEYINPUT101), .B(G101), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n607), .B(new_n608), .ZN(G3));
  INV_X1    g423(.A(G472), .ZN(new_n610));
  AOI21_X1  g424(.A(G902), .B1(new_n304), .B2(new_n306), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n309), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  AND2_X1   g426(.A1(new_n491), .A2(new_n501), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(new_n380), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT33), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n600), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n599), .A2(KEYINPUT33), .A3(new_n591), .ZN(new_n618));
  NAND4_X1  g432(.A1(new_n617), .A2(G478), .A3(new_n318), .A4(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(G478), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n594), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n623), .B1(new_n555), .B2(new_n561), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n441), .A2(KEYINPUT102), .A3(new_n442), .ZN(new_n625));
  INV_X1    g439(.A(new_n498), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n439), .B1(new_n427), .B2(new_n437), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT102), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n626), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  AND4_X1   g443(.A1(new_n497), .A2(new_n624), .A3(new_n625), .A4(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n615), .A2(new_n630), .ZN(new_n631));
  XOR2_X1   g445(.A(KEYINPUT34), .B(G104), .Z(new_n632));
  XNOR2_X1  g446(.A(new_n631), .B(new_n632), .ZN(G6));
  NAND4_X1  g447(.A1(new_n603), .A2(new_n538), .A3(new_n549), .A4(new_n553), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  NAND4_X1  g449(.A1(new_n625), .A2(new_n629), .A3(new_n497), .A4(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(KEYINPUT103), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(new_n615), .ZN(new_n638));
  XOR2_X1   g452(.A(KEYINPUT35), .B(G107), .Z(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G9));
  INV_X1    g454(.A(new_n612), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n366), .A2(KEYINPUT36), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n361), .B(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(new_n378), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n376), .A2(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  NOR3_X1   g460(.A1(new_n502), .A2(new_n605), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n641), .A2(new_n647), .ZN(new_n648));
  XOR2_X1   g462(.A(KEYINPUT37), .B(G110), .Z(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G12));
  INV_X1    g464(.A(KEYINPUT78), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n320), .B(new_n651), .ZN(new_n652));
  AOI21_X1  g466(.A(KEYINPUT32), .B1(new_n307), .B2(new_n308), .ZN(new_n653));
  AOI211_X1 g467(.A(new_n310), .B(new_n322), .C1(new_n304), .C2(new_n306), .ZN(new_n654));
  NOR3_X1   g468(.A1(new_n652), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n625), .A2(new_n629), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n491), .A2(new_n645), .A3(new_n501), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  AND3_X1   g472(.A1(new_n538), .A2(new_n549), .A3(new_n553), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT104), .ZN(new_n660));
  OR2_X1    g474(.A1(new_n496), .A2(G900), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(new_n493), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n659), .A2(new_n660), .A3(new_n603), .A4(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(new_n662), .ZN(new_n664));
  OAI21_X1  g478(.A(KEYINPUT104), .B1(new_n634), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n658), .A2(new_n667), .ZN(new_n668));
  OAI21_X1  g482(.A(KEYINPUT105), .B1(new_n655), .B2(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT105), .ZN(new_n670));
  NOR3_X1   g484(.A1(new_n666), .A2(new_n656), .A3(new_n657), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n325), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G128), .ZN(G30));
  XNOR2_X1  g488(.A(new_n443), .B(KEYINPUT38), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n555), .A2(new_n561), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(new_n603), .ZN(new_n678));
  NOR3_X1   g492(.A1(new_n676), .A2(new_n626), .A3(new_n678), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n653), .A2(new_n654), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n265), .B1(new_n291), .B2(new_n292), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(new_n273), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n297), .A2(new_n295), .A3(new_n265), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n682), .A2(new_n318), .A3(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(G472), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n680), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n679), .A2(new_n646), .A3(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n662), .B(KEYINPUT39), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n613), .A2(KEYINPUT106), .A3(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT106), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n491), .A2(new_n501), .ZN(new_n691));
  INV_X1    g505(.A(new_n688), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n690), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n689), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(KEYINPUT40), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n687), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(new_n225), .ZN(G45));
  AOI21_X1  g511(.A(new_n560), .B1(new_n559), .B2(new_n549), .ZN(new_n698));
  AND4_X1   g512(.A1(new_n560), .A2(new_n538), .A3(new_n549), .A4(new_n553), .ZN(new_n699));
  OAI211_X1 g513(.A(new_n622), .B(new_n662), .C1(new_n698), .C2(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT107), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n624), .A2(KEYINPUT107), .A3(new_n662), .ZN(new_n703));
  AND2_X1   g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n704), .A2(new_n325), .A3(new_n658), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G146), .ZN(G48));
  INV_X1    g520(.A(new_n380), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n707), .B1(new_n680), .B2(new_n321), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT108), .ZN(new_n709));
  AND3_X1   g523(.A1(new_n479), .A2(new_n480), .A3(new_n318), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n480), .B1(new_n479), .B2(new_n318), .ZN(new_n711));
  INV_X1    g525(.A(new_n501), .ZN(new_n712));
  NOR3_X1   g526(.A1(new_n710), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n708), .A2(new_n709), .A3(new_n630), .A4(new_n713), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n325), .A2(new_n630), .A3(new_n380), .A4(new_n713), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(KEYINPUT108), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(KEYINPUT41), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G113), .ZN(G15));
  NAND3_X1  g533(.A1(new_n708), .A2(new_n637), .A3(new_n713), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G116), .ZN(G18));
  NAND4_X1  g535(.A1(new_n713), .A2(new_n625), .A3(new_n497), .A4(new_n629), .ZN(new_n722));
  NOR3_X1   g536(.A1(new_n722), .A2(new_n605), .A3(new_n646), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(new_n325), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G119), .ZN(G21));
  AND2_X1   g539(.A1(new_n315), .A2(new_n316), .ZN(new_n726));
  OAI211_X1 g540(.A(new_n294), .B(new_n302), .C1(new_n273), .C2(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(new_n308), .ZN(new_n728));
  OAI211_X1 g542(.A(new_n728), .B(new_n380), .C1(new_n611), .C2(new_n610), .ZN(new_n729));
  INV_X1    g543(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n722), .A2(new_n678), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G122), .ZN(G24));
  OAI211_X1 g547(.A(new_n728), .B(new_n645), .C1(new_n611), .C2(new_n610), .ZN(new_n734));
  INV_X1    g548(.A(new_n713), .ZN(new_n735));
  NOR3_X1   g549(.A1(new_n734), .A2(new_n656), .A3(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(new_n704), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G125), .ZN(G27));
  NAND2_X1  g552(.A1(new_n325), .A2(new_n380), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT109), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n691), .A2(new_n740), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n443), .A2(new_n626), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n491), .A2(KEYINPUT109), .A3(new_n501), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n741), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n739), .A2(new_n744), .ZN(new_n745));
  AOI21_X1  g559(.A(KEYINPUT42), .B1(new_n745), .B2(new_n704), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n311), .A2(KEYINPUT110), .A3(new_n324), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT110), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n748), .B1(new_n653), .B2(new_n654), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n747), .A2(new_n749), .A3(new_n321), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(new_n380), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT111), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n750), .A2(KEYINPUT111), .A3(new_n380), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n702), .A2(new_n703), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT42), .ZN(new_n757));
  NOR3_X1   g571(.A1(new_n756), .A2(new_n744), .A3(new_n757), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n746), .B1(new_n755), .B2(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(new_n276), .ZN(G33));
  XOR2_X1   g574(.A(new_n666), .B(KEYINPUT112), .Z(new_n761));
  NOR3_X1   g575(.A1(new_n761), .A2(new_n739), .A3(new_n744), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(KEYINPUT113), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(new_n231), .ZN(G36));
  INV_X1    g578(.A(KEYINPUT45), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n480), .B1(new_n490), .B2(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n488), .A2(KEYINPUT45), .A3(new_n489), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n482), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n768), .A2(KEYINPUT46), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n769), .A2(KEYINPUT114), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n710), .B1(new_n768), .B2(KEYINPUT46), .ZN(new_n771));
  AND2_X1   g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  OR2_X1    g586(.A1(new_n769), .A2(KEYINPUT114), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n712), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  AND2_X1   g588(.A1(new_n774), .A2(new_n688), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n555), .A2(new_n561), .A3(new_n622), .ZN(new_n776));
  NAND2_X1  g590(.A1(KEYINPUT115), .A2(KEYINPUT43), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  XOR2_X1   g592(.A(KEYINPUT115), .B(KEYINPUT43), .Z(new_n779));
  OAI21_X1  g593(.A(new_n778), .B1(new_n776), .B2(new_n779), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n780), .A2(new_n612), .A3(new_n645), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT44), .ZN(new_n782));
  OR2_X1    g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(new_n742), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n784), .B1(new_n781), .B2(new_n782), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n775), .A2(new_n783), .A3(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G137), .ZN(G39));
  NAND2_X1  g601(.A1(KEYINPUT116), .A2(KEYINPUT47), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n774), .A2(new_n788), .ZN(new_n789));
  NOR4_X1   g603(.A1(new_n325), .A2(new_n756), .A3(new_n380), .A4(new_n784), .ZN(new_n790));
  XOR2_X1   g604(.A(KEYINPUT116), .B(KEYINPUT47), .Z(new_n791));
  OAI211_X1 g605(.A(new_n789), .B(new_n790), .C1(new_n774), .C2(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G140), .ZN(G42));
  NAND2_X1  g607(.A1(new_n677), .A2(new_n623), .ZN(new_n794));
  AND4_X1   g608(.A1(new_n605), .A2(new_n794), .A3(new_n443), .A4(new_n499), .ZN(new_n795));
  AOI22_X1  g609(.A1(new_n615), .A2(new_n795), .B1(new_n730), .B2(new_n731), .ZN(new_n796));
  AOI22_X1  g610(.A1(new_n723), .A2(new_n325), .B1(new_n641), .B2(new_n647), .ZN(new_n797));
  AND3_X1   g611(.A1(new_n796), .A2(new_n797), .A3(new_n607), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n728), .B1(new_n611), .B2(new_n610), .ZN(new_n799));
  NOR3_X1   g613(.A1(new_n756), .A2(new_n744), .A3(new_n799), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n691), .A2(new_n664), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n554), .A2(new_n603), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n801), .A2(new_n742), .A3(new_n802), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n655), .A2(new_n803), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n645), .B1(new_n800), .B2(new_n804), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n798), .A2(new_n717), .A3(new_n720), .A4(new_n805), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n759), .A2(new_n806), .A3(new_n762), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n613), .A2(new_n625), .A3(new_n629), .A4(new_n645), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n808), .B1(new_n680), .B2(new_n321), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n704), .B1(new_n809), .B2(new_n736), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n678), .A2(new_n656), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n686), .A2(new_n811), .A3(new_n646), .A4(new_n801), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n673), .A2(new_n810), .A3(KEYINPUT52), .A4(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT117), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n673), .A2(new_n810), .A3(new_n812), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT52), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n815), .A2(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n816), .A2(new_n814), .A3(new_n817), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n807), .A2(new_n821), .A3(KEYINPUT53), .ZN(new_n822));
  INV_X1    g636(.A(new_n754), .ZN(new_n823));
  AOI21_X1  g637(.A(KEYINPUT111), .B1(new_n750), .B2(new_n380), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n758), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(new_n746), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n762), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(new_n806), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n818), .A2(new_n813), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n827), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT53), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT54), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n822), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n834), .A2(KEYINPUT118), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT118), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n822), .A2(new_n832), .A3(new_n836), .A4(new_n833), .ZN(new_n837));
  AOI21_X1  g651(.A(KEYINPUT53), .B1(new_n807), .B2(new_n821), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n830), .A2(new_n831), .ZN(new_n839));
  OAI21_X1  g653(.A(KEYINPUT54), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n835), .A2(new_n837), .A3(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(new_n493), .ZN(new_n842));
  AND2_X1   g656(.A1(new_n780), .A2(new_n842), .ZN(new_n843));
  AND2_X1   g657(.A1(new_n843), .A2(new_n730), .ZN(new_n844));
  NOR3_X1   g658(.A1(new_n675), .A2(new_n498), .A3(new_n735), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  XOR2_X1   g660(.A(new_n846), .B(KEYINPUT50), .Z(new_n847));
  NOR2_X1   g661(.A1(new_n784), .A2(new_n735), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n843), .A2(new_n848), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n849), .A2(new_n734), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n848), .A2(new_n380), .A3(new_n842), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n686), .A2(new_n851), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n677), .A2(new_n622), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n850), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n847), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(KEYINPUT119), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT51), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n789), .B1(new_n774), .B2(new_n791), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n710), .A2(new_n711), .ZN(new_n859));
  INV_X1    g673(.A(new_n859), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n858), .B1(new_n501), .B2(new_n860), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n844), .A2(new_n742), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n857), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT119), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n847), .A2(new_n864), .A3(new_n854), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n856), .A2(new_n863), .A3(new_n865), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n861), .A2(new_n862), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n857), .B1(new_n867), .B2(new_n855), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n849), .B1(new_n753), .B2(new_n754), .ZN(new_n869));
  XOR2_X1   g683(.A(new_n869), .B(KEYINPUT48), .Z(new_n870));
  NAND2_X1  g684(.A1(new_n852), .A2(new_n624), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n871), .A2(G952), .A3(new_n362), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n656), .A2(new_n735), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n872), .B1(new_n873), .B2(new_n844), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n866), .A2(new_n868), .A3(new_n870), .A4(new_n874), .ZN(new_n875));
  OAI22_X1  g689(.A1(new_n841), .A2(new_n875), .B1(G952), .B2(G953), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n380), .A2(new_n498), .A3(new_n501), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n877), .B1(KEYINPUT49), .B2(new_n860), .ZN(new_n878));
  OAI211_X1 g692(.A(new_n676), .B(new_n878), .C1(KEYINPUT49), .C2(new_n860), .ZN(new_n879));
  OR3_X1    g693(.A1(new_n879), .A2(new_n686), .A3(new_n776), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n876), .A2(new_n880), .ZN(G75));
  AOI21_X1  g695(.A(new_n318), .B1(new_n822), .B2(new_n832), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(G210), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n416), .A2(new_n422), .ZN(new_n884));
  XNOR2_X1  g698(.A(new_n884), .B(new_n420), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n885), .B(KEYINPUT55), .ZN(new_n886));
  XOR2_X1   g700(.A(KEYINPUT120), .B(KEYINPUT56), .Z(new_n887));
  AND3_X1   g701(.A1(new_n883), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT56), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n886), .B1(new_n883), .B2(new_n889), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n362), .A2(G952), .ZN(new_n891));
  NOR3_X1   g705(.A1(new_n888), .A2(new_n890), .A3(new_n891), .ZN(G51));
  XNOR2_X1  g706(.A(new_n482), .B(KEYINPUT57), .ZN(new_n893));
  AND3_X1   g707(.A1(new_n822), .A2(new_n832), .A3(new_n833), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n833), .B1(new_n822), .B2(new_n832), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n893), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n896), .A2(new_n479), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n882), .A2(new_n767), .A3(new_n766), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n891), .B1(new_n897), .B2(new_n898), .ZN(G54));
  AND2_X1   g713(.A1(KEYINPUT58), .A2(G475), .ZN(new_n900));
  AND3_X1   g714(.A1(new_n882), .A2(new_n547), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n547), .B1(new_n882), .B2(new_n900), .ZN(new_n902));
  NOR3_X1   g716(.A1(new_n901), .A2(new_n902), .A3(new_n891), .ZN(G60));
  XNOR2_X1  g717(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n620), .A2(new_n318), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n904), .B(new_n905), .ZN(new_n906));
  AND3_X1   g720(.A1(new_n617), .A2(new_n618), .A3(new_n906), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n907), .B1(new_n894), .B2(new_n895), .ZN(new_n908));
  INV_X1    g722(.A(new_n891), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n841), .A2(new_n906), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n617), .A2(new_n618), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n910), .B1(new_n911), .B2(new_n912), .ZN(G63));
  NAND2_X1  g727(.A1(new_n822), .A2(new_n832), .ZN(new_n914));
  NAND2_X1  g728(.A1(G217), .A2(G902), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n915), .B(KEYINPUT60), .ZN(new_n916));
  INV_X1    g730(.A(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n914), .A2(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(new_n369), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n891), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n916), .B1(new_n822), .B2(new_n832), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n921), .A2(new_n643), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT122), .ZN(new_n923));
  OAI211_X1 g737(.A(new_n920), .B(new_n922), .C1(new_n923), .C2(KEYINPUT61), .ZN(new_n924));
  OAI211_X1 g738(.A(new_n923), .B(new_n909), .C1(new_n921), .C2(new_n369), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT61), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n909), .B1(new_n921), .B2(new_n369), .ZN(new_n927));
  AND3_X1   g741(.A1(new_n914), .A2(new_n643), .A3(new_n917), .ZN(new_n928));
  OAI211_X1 g742(.A(new_n925), .B(new_n926), .C1(new_n927), .C2(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n924), .A2(new_n929), .ZN(G66));
  AND3_X1   g744(.A1(new_n798), .A2(new_n717), .A3(new_n720), .ZN(new_n931));
  AND2_X1   g745(.A1(G224), .A2(G953), .ZN(new_n932));
  AOI22_X1  g746(.A1(new_n931), .A2(new_n362), .B1(new_n495), .B2(new_n932), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n884), .B1(G898), .B2(new_n362), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n933), .B(new_n934), .ZN(G69));
  INV_X1    g749(.A(KEYINPUT125), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT123), .ZN(new_n937));
  AND3_X1   g751(.A1(new_n325), .A2(new_n670), .A3(new_n671), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n670), .B1(new_n325), .B2(new_n671), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n705), .A2(new_n737), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n937), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n673), .A2(new_n810), .A3(KEYINPUT123), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n696), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT62), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n936), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  OR2_X1    g760(.A1(new_n687), .A2(new_n695), .ZN(new_n947));
  AND3_X1   g761(.A1(new_n673), .A2(KEYINPUT123), .A3(new_n810), .ZN(new_n948));
  AOI21_X1  g762(.A(KEYINPUT123), .B1(new_n673), .B2(new_n810), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n947), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n950), .A2(KEYINPUT125), .A3(KEYINPUT62), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n946), .A2(new_n951), .ZN(new_n952));
  OAI211_X1 g766(.A(new_n945), .B(new_n947), .C1(new_n948), .C2(new_n949), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT124), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n942), .A2(new_n943), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n956), .A2(KEYINPUT124), .A3(new_n945), .A4(new_n947), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n794), .A2(new_n605), .A3(new_n742), .ZN(new_n959));
  OR3_X1    g773(.A1(new_n739), .A2(new_n694), .A3(new_n959), .ZN(new_n960));
  AND3_X1   g774(.A1(new_n786), .A2(new_n792), .A3(new_n960), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n952), .A2(new_n958), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n962), .A2(new_n362), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n288), .A2(new_n289), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n286), .A2(new_n964), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n965), .B(new_n542), .ZN(new_n966));
  INV_X1    g780(.A(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n963), .A2(new_n967), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT127), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n362), .B1(G227), .B2(G900), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n967), .B1(G900), .B2(G953), .ZN(new_n971));
  INV_X1    g785(.A(new_n971), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n775), .A2(new_n755), .A3(new_n811), .ZN(new_n973));
  NAND4_X1  g787(.A1(new_n973), .A2(new_n956), .A3(new_n786), .A4(new_n792), .ZN(new_n974));
  OAI21_X1  g788(.A(KEYINPUT126), .B1(new_n759), .B2(new_n762), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT126), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n827), .A2(new_n976), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n974), .B1(new_n975), .B2(new_n977), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n972), .B1(new_n978), .B2(new_n362), .ZN(new_n979));
  INV_X1    g793(.A(new_n979), .ZN(new_n980));
  NAND4_X1  g794(.A1(new_n968), .A2(new_n969), .A3(new_n970), .A4(new_n980), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n970), .A2(new_n969), .ZN(new_n982));
  OR2_X1    g796(.A1(new_n970), .A2(new_n969), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n966), .B1(new_n962), .B2(new_n362), .ZN(new_n984));
  OAI211_X1 g798(.A(new_n982), .B(new_n983), .C1(new_n984), .C2(new_n979), .ZN(new_n985));
  AND2_X1   g799(.A1(new_n981), .A2(new_n985), .ZN(G72));
  NOR2_X1   g800(.A1(new_n838), .A2(new_n839), .ZN(new_n987));
  NAND2_X1  g801(.A1(G472), .A2(G902), .ZN(new_n988));
  XOR2_X1   g802(.A(new_n988), .B(KEYINPUT63), .Z(new_n989));
  NAND3_X1  g803(.A1(new_n682), .A2(new_n312), .A3(new_n989), .ZN(new_n990));
  INV_X1    g804(.A(new_n989), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n991), .B1(new_n978), .B2(new_n931), .ZN(new_n992));
  OAI221_X1 g806(.A(new_n909), .B1(new_n987), .B2(new_n990), .C1(new_n992), .C2(new_n312), .ZN(new_n993));
  NAND4_X1  g807(.A1(new_n952), .A2(new_n958), .A3(new_n931), .A4(new_n961), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n682), .B1(new_n994), .B2(new_n989), .ZN(new_n995));
  NOR2_X1   g809(.A1(new_n993), .A2(new_n995), .ZN(G57));
endmodule


