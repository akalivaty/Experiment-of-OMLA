

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U552 ( .A1(G651), .A2(n632), .ZN(n655) );
  XOR2_X1 U553 ( .A(n745), .B(KEYINPUT32), .Z(n516) );
  OR2_X1 U554 ( .A1(n706), .A2(n705), .ZN(n517) );
  INV_X1 U555 ( .A(n736), .ZN(n720) );
  INV_X1 U556 ( .A(KEYINPUT28), .ZN(n715) );
  AND2_X1 U557 ( .A1(n744), .A2(n743), .ZN(n745) );
  NOR2_X1 U558 ( .A1(n766), .A2(n765), .ZN(n798) );
  INV_X1 U559 ( .A(G651), .ZN(n548) );
  NOR2_X2 U560 ( .A1(n523), .A2(G2105), .ZN(n893) );
  XOR2_X1 U561 ( .A(KEYINPUT17), .B(n520), .Z(n892) );
  XOR2_X1 U562 ( .A(KEYINPUT77), .B(n587), .Z(n972) );
  NOR2_X1 U563 ( .A1(n527), .A2(n526), .ZN(G160) );
  INV_X1 U564 ( .A(G2104), .ZN(n523) );
  NAND2_X1 U565 ( .A1(n893), .A2(G101), .ZN(n518) );
  XNOR2_X1 U566 ( .A(n518), .B(KEYINPUT65), .ZN(n519) );
  XNOR2_X1 U567 ( .A(n519), .B(KEYINPUT23), .ZN(n522) );
  NOR2_X1 U568 ( .A1(G2104), .A2(G2105), .ZN(n520) );
  NAND2_X1 U569 ( .A1(G137), .A2(n892), .ZN(n521) );
  NAND2_X1 U570 ( .A1(n522), .A2(n521), .ZN(n527) );
  AND2_X1 U571 ( .A1(n523), .A2(G2105), .ZN(n888) );
  NAND2_X1 U572 ( .A1(G125), .A2(n888), .ZN(n525) );
  AND2_X1 U573 ( .A1(G2104), .A2(G2105), .ZN(n889) );
  NAND2_X1 U574 ( .A1(G113), .A2(n889), .ZN(n524) );
  NAND2_X1 U575 ( .A1(n525), .A2(n524), .ZN(n526) );
  XOR2_X1 U576 ( .A(G2446), .B(G2454), .Z(n529) );
  XNOR2_X1 U577 ( .A(KEYINPUT104), .B(G2430), .ZN(n528) );
  XNOR2_X1 U578 ( .A(n529), .B(n528), .ZN(n530) );
  XOR2_X1 U579 ( .A(n530), .B(G2443), .Z(n532) );
  XNOR2_X1 U580 ( .A(G1348), .B(G2438), .ZN(n531) );
  XNOR2_X1 U581 ( .A(n532), .B(n531), .ZN(n536) );
  XOR2_X1 U582 ( .A(G2435), .B(KEYINPUT103), .Z(n534) );
  XNOR2_X1 U583 ( .A(G1341), .B(G2427), .ZN(n533) );
  XNOR2_X1 U584 ( .A(n534), .B(n533), .ZN(n535) );
  XOR2_X1 U585 ( .A(n536), .B(n535), .Z(n538) );
  XNOR2_X1 U586 ( .A(G2451), .B(KEYINPUT105), .ZN(n537) );
  XNOR2_X1 U587 ( .A(n538), .B(n537), .ZN(n539) );
  AND2_X1 U588 ( .A1(n539), .A2(G14), .ZN(G401) );
  AND2_X1 U589 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U590 ( .A(G57), .ZN(G237) );
  INV_X1 U591 ( .A(G132), .ZN(G219) );
  INV_X1 U592 ( .A(G82), .ZN(G220) );
  NOR2_X1 U593 ( .A1(G543), .A2(n548), .ZN(n540) );
  XOR2_X1 U594 ( .A(n540), .B(KEYINPUT68), .Z(n541) );
  XNOR2_X2 U595 ( .A(KEYINPUT1), .B(n541), .ZN(n647) );
  NAND2_X1 U596 ( .A1(G63), .A2(n647), .ZN(n542) );
  XOR2_X1 U597 ( .A(KEYINPUT79), .B(n542), .Z(n544) );
  XOR2_X1 U598 ( .A(G543), .B(KEYINPUT0), .Z(n632) );
  NAND2_X1 U599 ( .A1(n655), .A2(G51), .ZN(n543) );
  NAND2_X1 U600 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U601 ( .A(KEYINPUT6), .B(n545), .ZN(n553) );
  NOR2_X1 U602 ( .A1(G651), .A2(G543), .ZN(n646) );
  NAND2_X1 U603 ( .A1(G89), .A2(n646), .ZN(n546) );
  XNOR2_X1 U604 ( .A(n546), .B(KEYINPUT78), .ZN(n547) );
  XNOR2_X1 U605 ( .A(n547), .B(KEYINPUT4), .ZN(n550) );
  NOR2_X1 U606 ( .A1(n632), .A2(n548), .ZN(n651) );
  NAND2_X1 U607 ( .A1(G76), .A2(n651), .ZN(n549) );
  NAND2_X1 U608 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U609 ( .A(n551), .B(KEYINPUT5), .Z(n552) );
  NOR2_X1 U610 ( .A1(n553), .A2(n552), .ZN(n554) );
  XOR2_X1 U611 ( .A(KEYINPUT7), .B(n554), .Z(n555) );
  XNOR2_X1 U612 ( .A(KEYINPUT80), .B(n555), .ZN(G168) );
  XOR2_X1 U613 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U614 ( .A1(G7), .A2(G661), .ZN(n556) );
  XOR2_X1 U615 ( .A(n556), .B(KEYINPUT10), .Z(n835) );
  NAND2_X1 U616 ( .A1(n835), .A2(G567), .ZN(n557) );
  XOR2_X1 U617 ( .A(KEYINPUT11), .B(n557), .Z(G234) );
  XOR2_X1 U618 ( .A(KEYINPUT14), .B(KEYINPUT74), .Z(n559) );
  NAND2_X1 U619 ( .A1(G56), .A2(n647), .ZN(n558) );
  XNOR2_X1 U620 ( .A(n559), .B(n558), .ZN(n560) );
  XOR2_X1 U621 ( .A(KEYINPUT73), .B(n560), .Z(n566) );
  NAND2_X1 U622 ( .A1(n646), .A2(G81), .ZN(n561) );
  XNOR2_X1 U623 ( .A(n561), .B(KEYINPUT12), .ZN(n563) );
  NAND2_X1 U624 ( .A1(G68), .A2(n651), .ZN(n562) );
  NAND2_X1 U625 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U626 ( .A(KEYINPUT13), .B(n564), .Z(n565) );
  NOR2_X1 U627 ( .A1(n566), .A2(n565), .ZN(n568) );
  NAND2_X1 U628 ( .A1(n655), .A2(G43), .ZN(n567) );
  NAND2_X1 U629 ( .A1(n568), .A2(n567), .ZN(n977) );
  XNOR2_X1 U630 ( .A(G860), .B(KEYINPUT75), .ZN(n599) );
  NOR2_X1 U631 ( .A1(n977), .A2(n599), .ZN(n569) );
  XOR2_X1 U632 ( .A(KEYINPUT76), .B(n569), .Z(G153) );
  NAND2_X1 U633 ( .A1(G52), .A2(n655), .ZN(n570) );
  XNOR2_X1 U634 ( .A(n570), .B(KEYINPUT70), .ZN(n573) );
  NAND2_X1 U635 ( .A1(n647), .A2(G64), .ZN(n571) );
  XOR2_X1 U636 ( .A(KEYINPUT69), .B(n571), .Z(n572) );
  NAND2_X1 U637 ( .A1(n573), .A2(n572), .ZN(n579) );
  NAND2_X1 U638 ( .A1(n651), .A2(G77), .ZN(n574) );
  XOR2_X1 U639 ( .A(KEYINPUT71), .B(n574), .Z(n576) );
  NAND2_X1 U640 ( .A1(n646), .A2(G90), .ZN(n575) );
  NAND2_X1 U641 ( .A1(n576), .A2(n575), .ZN(n577) );
  XOR2_X1 U642 ( .A(KEYINPUT9), .B(n577), .Z(n578) );
  NOR2_X1 U643 ( .A1(n579), .A2(n578), .ZN(G171) );
  INV_X1 U644 ( .A(G171), .ZN(G301) );
  NAND2_X1 U645 ( .A1(G868), .A2(G301), .ZN(n589) );
  NAND2_X1 U646 ( .A1(G92), .A2(n646), .ZN(n581) );
  NAND2_X1 U647 ( .A1(G66), .A2(n647), .ZN(n580) );
  NAND2_X1 U648 ( .A1(n581), .A2(n580), .ZN(n585) );
  NAND2_X1 U649 ( .A1(G79), .A2(n651), .ZN(n583) );
  NAND2_X1 U650 ( .A1(G54), .A2(n655), .ZN(n582) );
  NAND2_X1 U651 ( .A1(n583), .A2(n582), .ZN(n584) );
  NOR2_X1 U652 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U653 ( .A(n586), .B(KEYINPUT15), .Z(n587) );
  INV_X1 U654 ( .A(n972), .ZN(n706) );
  INV_X1 U655 ( .A(G868), .ZN(n666) );
  NAND2_X1 U656 ( .A1(n706), .A2(n666), .ZN(n588) );
  NAND2_X1 U657 ( .A1(n589), .A2(n588), .ZN(G284) );
  NAND2_X1 U658 ( .A1(G91), .A2(n646), .ZN(n591) );
  NAND2_X1 U659 ( .A1(G65), .A2(n647), .ZN(n590) );
  NAND2_X1 U660 ( .A1(n591), .A2(n590), .ZN(n594) );
  NAND2_X1 U661 ( .A1(n651), .A2(G78), .ZN(n592) );
  XOR2_X1 U662 ( .A(KEYINPUT72), .B(n592), .Z(n593) );
  NOR2_X1 U663 ( .A1(n594), .A2(n593), .ZN(n596) );
  NAND2_X1 U664 ( .A1(n655), .A2(G53), .ZN(n595) );
  NAND2_X1 U665 ( .A1(n596), .A2(n595), .ZN(G299) );
  NAND2_X1 U666 ( .A1(G868), .A2(G286), .ZN(n598) );
  NAND2_X1 U667 ( .A1(G299), .A2(n666), .ZN(n597) );
  NAND2_X1 U668 ( .A1(n598), .A2(n597), .ZN(G297) );
  NAND2_X1 U669 ( .A1(n599), .A2(G559), .ZN(n600) );
  NAND2_X1 U670 ( .A1(n600), .A2(n972), .ZN(n601) );
  XNOR2_X1 U671 ( .A(n601), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U672 ( .A1(n706), .A2(n666), .ZN(n602) );
  XNOR2_X1 U673 ( .A(n602), .B(KEYINPUT81), .ZN(n603) );
  NOR2_X1 U674 ( .A1(G559), .A2(n603), .ZN(n604) );
  XNOR2_X1 U675 ( .A(n604), .B(KEYINPUT82), .ZN(n606) );
  NOR2_X1 U676 ( .A1(n977), .A2(G868), .ZN(n605) );
  NOR2_X1 U677 ( .A1(n606), .A2(n605), .ZN(G282) );
  NAND2_X1 U678 ( .A1(n888), .A2(G123), .ZN(n607) );
  XNOR2_X1 U679 ( .A(n607), .B(KEYINPUT18), .ZN(n609) );
  NAND2_X1 U680 ( .A1(G111), .A2(n889), .ZN(n608) );
  NAND2_X1 U681 ( .A1(n609), .A2(n608), .ZN(n613) );
  NAND2_X1 U682 ( .A1(G135), .A2(n892), .ZN(n611) );
  NAND2_X1 U683 ( .A1(G99), .A2(n893), .ZN(n610) );
  NAND2_X1 U684 ( .A1(n611), .A2(n610), .ZN(n612) );
  NOR2_X1 U685 ( .A1(n613), .A2(n612), .ZN(n918) );
  XNOR2_X1 U686 ( .A(G2096), .B(n918), .ZN(n614) );
  INV_X1 U687 ( .A(G2100), .ZN(n840) );
  NAND2_X1 U688 ( .A1(n614), .A2(n840), .ZN(G156) );
  NAND2_X1 U689 ( .A1(G93), .A2(n646), .ZN(n616) );
  NAND2_X1 U690 ( .A1(G67), .A2(n647), .ZN(n615) );
  NAND2_X1 U691 ( .A1(n616), .A2(n615), .ZN(n620) );
  NAND2_X1 U692 ( .A1(G80), .A2(n651), .ZN(n618) );
  NAND2_X1 U693 ( .A1(G55), .A2(n655), .ZN(n617) );
  NAND2_X1 U694 ( .A1(n618), .A2(n617), .ZN(n619) );
  OR2_X1 U695 ( .A1(n620), .A2(n619), .ZN(n665) );
  NAND2_X1 U696 ( .A1(G559), .A2(n972), .ZN(n621) );
  XNOR2_X1 U697 ( .A(n977), .B(n621), .ZN(n663) );
  NOR2_X1 U698 ( .A1(G860), .A2(n663), .ZN(n622) );
  XOR2_X1 U699 ( .A(KEYINPUT83), .B(n622), .Z(n623) );
  XOR2_X1 U700 ( .A(n665), .B(n623), .Z(G145) );
  NAND2_X1 U701 ( .A1(n646), .A2(G85), .ZN(n624) );
  XNOR2_X1 U702 ( .A(KEYINPUT66), .B(n624), .ZN(n631) );
  NAND2_X1 U703 ( .A1(n655), .A2(G47), .ZN(n626) );
  NAND2_X1 U704 ( .A1(G60), .A2(n647), .ZN(n625) );
  NAND2_X1 U705 ( .A1(n626), .A2(n625), .ZN(n629) );
  NAND2_X1 U706 ( .A1(G72), .A2(n651), .ZN(n627) );
  XNOR2_X1 U707 ( .A(KEYINPUT67), .B(n627), .ZN(n628) );
  NOR2_X1 U708 ( .A1(n629), .A2(n628), .ZN(n630) );
  NAND2_X1 U709 ( .A1(n631), .A2(n630), .ZN(G290) );
  NAND2_X1 U710 ( .A1(G87), .A2(n632), .ZN(n634) );
  NAND2_X1 U711 ( .A1(G74), .A2(G651), .ZN(n633) );
  NAND2_X1 U712 ( .A1(n634), .A2(n633), .ZN(n635) );
  NOR2_X1 U713 ( .A1(n647), .A2(n635), .ZN(n637) );
  NAND2_X1 U714 ( .A1(n655), .A2(G49), .ZN(n636) );
  NAND2_X1 U715 ( .A1(n637), .A2(n636), .ZN(G288) );
  NAND2_X1 U716 ( .A1(G88), .A2(n646), .ZN(n639) );
  NAND2_X1 U717 ( .A1(G75), .A2(n651), .ZN(n638) );
  NAND2_X1 U718 ( .A1(n639), .A2(n638), .ZN(n640) );
  XOR2_X1 U719 ( .A(KEYINPUT86), .B(n640), .Z(n642) );
  NAND2_X1 U720 ( .A1(G62), .A2(n647), .ZN(n641) );
  NAND2_X1 U721 ( .A1(n642), .A2(n641), .ZN(n645) );
  NAND2_X1 U722 ( .A1(G50), .A2(n655), .ZN(n643) );
  XNOR2_X1 U723 ( .A(KEYINPUT85), .B(n643), .ZN(n644) );
  NOR2_X1 U724 ( .A1(n645), .A2(n644), .ZN(G166) );
  NAND2_X1 U725 ( .A1(G86), .A2(n646), .ZN(n649) );
  NAND2_X1 U726 ( .A1(G61), .A2(n647), .ZN(n648) );
  NAND2_X1 U727 ( .A1(n649), .A2(n648), .ZN(n650) );
  XNOR2_X1 U728 ( .A(KEYINPUT84), .B(n650), .ZN(n654) );
  NAND2_X1 U729 ( .A1(n651), .A2(G73), .ZN(n652) );
  XOR2_X1 U730 ( .A(KEYINPUT2), .B(n652), .Z(n653) );
  NOR2_X1 U731 ( .A1(n654), .A2(n653), .ZN(n657) );
  NAND2_X1 U732 ( .A1(n655), .A2(G48), .ZN(n656) );
  NAND2_X1 U733 ( .A1(n657), .A2(n656), .ZN(G305) );
  XNOR2_X1 U734 ( .A(KEYINPUT19), .B(G290), .ZN(n658) );
  XNOR2_X1 U735 ( .A(n658), .B(G288), .ZN(n659) );
  XNOR2_X1 U736 ( .A(n659), .B(n665), .ZN(n661) );
  XOR2_X1 U737 ( .A(G299), .B(G166), .Z(n660) );
  XNOR2_X1 U738 ( .A(n661), .B(n660), .ZN(n662) );
  XNOR2_X1 U739 ( .A(n662), .B(G305), .ZN(n905) );
  XOR2_X1 U740 ( .A(n663), .B(n905), .Z(n664) );
  NAND2_X1 U741 ( .A1(n664), .A2(G868), .ZN(n668) );
  NAND2_X1 U742 ( .A1(n666), .A2(n665), .ZN(n667) );
  NAND2_X1 U743 ( .A1(n668), .A2(n667), .ZN(G295) );
  NAND2_X1 U744 ( .A1(G2084), .A2(G2078), .ZN(n669) );
  XNOR2_X1 U745 ( .A(n669), .B(KEYINPUT20), .ZN(n670) );
  XNOR2_X1 U746 ( .A(KEYINPUT87), .B(n670), .ZN(n671) );
  NAND2_X1 U747 ( .A1(n671), .A2(G2090), .ZN(n672) );
  XNOR2_X1 U748 ( .A(KEYINPUT21), .B(n672), .ZN(n673) );
  NAND2_X1 U749 ( .A1(n673), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U750 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U751 ( .A1(G220), .A2(G219), .ZN(n674) );
  XOR2_X1 U752 ( .A(KEYINPUT22), .B(n674), .Z(n675) );
  NOR2_X1 U753 ( .A1(G218), .A2(n675), .ZN(n676) );
  NAND2_X1 U754 ( .A1(G96), .A2(n676), .ZN(n1022) );
  NAND2_X1 U755 ( .A1(n1022), .A2(G2106), .ZN(n680) );
  NAND2_X1 U756 ( .A1(G120), .A2(G108), .ZN(n677) );
  NOR2_X1 U757 ( .A1(G237), .A2(n677), .ZN(n678) );
  NAND2_X1 U758 ( .A1(G69), .A2(n678), .ZN(n1023) );
  NAND2_X1 U759 ( .A1(n1023), .A2(G567), .ZN(n679) );
  NAND2_X1 U760 ( .A1(n680), .A2(n679), .ZN(n839) );
  NAND2_X1 U761 ( .A1(G483), .A2(G661), .ZN(n681) );
  NOR2_X1 U762 ( .A1(n839), .A2(n681), .ZN(n838) );
  NAND2_X1 U763 ( .A1(n838), .A2(G36), .ZN(G176) );
  NAND2_X1 U764 ( .A1(G138), .A2(n892), .ZN(n683) );
  NAND2_X1 U765 ( .A1(G102), .A2(n893), .ZN(n682) );
  NAND2_X1 U766 ( .A1(n683), .A2(n682), .ZN(n687) );
  NAND2_X1 U767 ( .A1(G126), .A2(n888), .ZN(n685) );
  NAND2_X1 U768 ( .A1(G114), .A2(n889), .ZN(n684) );
  NAND2_X1 U769 ( .A1(n685), .A2(n684), .ZN(n686) );
  NOR2_X1 U770 ( .A1(n687), .A2(n686), .ZN(G164) );
  XOR2_X1 U771 ( .A(G166), .B(KEYINPUT88), .Z(G303) );
  INV_X1 U772 ( .A(G1348), .ZN(n688) );
  NOR2_X1 U773 ( .A1(n688), .A2(n972), .ZN(n691) );
  XNOR2_X1 U774 ( .A(KEYINPUT64), .B(KEYINPUT26), .ZN(n700) );
  INV_X1 U775 ( .A(G1341), .ZN(n689) );
  NAND2_X1 U776 ( .A1(n700), .A2(n689), .ZN(n690) );
  NOR2_X1 U777 ( .A1(n691), .A2(n690), .ZN(n693) );
  NOR2_X1 U778 ( .A1(G164), .A2(G1384), .ZN(n768) );
  NAND2_X1 U779 ( .A1(G160), .A2(G40), .ZN(n767) );
  XOR2_X1 U780 ( .A(KEYINPUT92), .B(n767), .Z(n692) );
  NAND2_X2 U781 ( .A1(n768), .A2(n692), .ZN(n736) );
  NOR2_X1 U782 ( .A1(n693), .A2(n720), .ZN(n694) );
  NOR2_X1 U783 ( .A1(n977), .A2(n694), .ZN(n699) );
  NAND2_X1 U784 ( .A1(G1996), .A2(n700), .ZN(n696) );
  NAND2_X1 U785 ( .A1(G2067), .A2(n706), .ZN(n695) );
  NAND2_X1 U786 ( .A1(n696), .A2(n695), .ZN(n697) );
  NAND2_X1 U787 ( .A1(n720), .A2(n697), .ZN(n698) );
  NAND2_X1 U788 ( .A1(n699), .A2(n698), .ZN(n702) );
  NOR2_X1 U789 ( .A1(G1996), .A2(n700), .ZN(n701) );
  NOR2_X1 U790 ( .A1(n702), .A2(n701), .ZN(n712) );
  NAND2_X1 U791 ( .A1(G1348), .A2(n736), .ZN(n704) );
  NAND2_X1 U792 ( .A1(G2067), .A2(n720), .ZN(n703) );
  NAND2_X1 U793 ( .A1(n704), .A2(n703), .ZN(n705) );
  NAND2_X1 U794 ( .A1(n720), .A2(G2072), .ZN(n707) );
  XNOR2_X1 U795 ( .A(n707), .B(KEYINPUT27), .ZN(n709) );
  AND2_X1 U796 ( .A1(G1956), .A2(n736), .ZN(n708) );
  NOR2_X1 U797 ( .A1(n709), .A2(n708), .ZN(n714) );
  INV_X1 U798 ( .A(G299), .ZN(n713) );
  NAND2_X1 U799 ( .A1(n714), .A2(n713), .ZN(n710) );
  NAND2_X1 U800 ( .A1(n517), .A2(n710), .ZN(n711) );
  OR2_X1 U801 ( .A1(n712), .A2(n711), .ZN(n718) );
  NOR2_X1 U802 ( .A1(n714), .A2(n713), .ZN(n716) );
  XNOR2_X1 U803 ( .A(n716), .B(n715), .ZN(n717) );
  NAND2_X1 U804 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U805 ( .A(n719), .B(KEYINPUT29), .ZN(n725) );
  NOR2_X1 U806 ( .A1(n720), .A2(G1961), .ZN(n721) );
  XNOR2_X1 U807 ( .A(n721), .B(KEYINPUT94), .ZN(n723) );
  XOR2_X1 U808 ( .A(G2078), .B(KEYINPUT25), .Z(n946) );
  NOR2_X1 U809 ( .A1(n736), .A2(n946), .ZN(n722) );
  NOR2_X1 U810 ( .A1(n723), .A2(n722), .ZN(n729) );
  NOR2_X1 U811 ( .A1(G301), .A2(n729), .ZN(n724) );
  NOR2_X1 U812 ( .A1(n725), .A2(n724), .ZN(n734) );
  NAND2_X1 U813 ( .A1(G8), .A2(n736), .ZN(n807) );
  NOR2_X1 U814 ( .A1(G1966), .A2(n807), .ZN(n750) );
  NOR2_X1 U815 ( .A1(G2084), .A2(n736), .ZN(n746) );
  NOR2_X1 U816 ( .A1(n750), .A2(n746), .ZN(n726) );
  NAND2_X1 U817 ( .A1(G8), .A2(n726), .ZN(n727) );
  XNOR2_X1 U818 ( .A(KEYINPUT30), .B(n727), .ZN(n728) );
  NOR2_X1 U819 ( .A1(G168), .A2(n728), .ZN(n731) );
  AND2_X1 U820 ( .A1(G301), .A2(n729), .ZN(n730) );
  NOR2_X1 U821 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U822 ( .A(n732), .B(KEYINPUT31), .ZN(n733) );
  NOR2_X1 U823 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U824 ( .A(n735), .B(KEYINPUT95), .ZN(n748) );
  NAND2_X1 U825 ( .A1(n748), .A2(G286), .ZN(n744) );
  INV_X1 U826 ( .A(G8), .ZN(n742) );
  NOR2_X1 U827 ( .A1(G1971), .A2(n807), .ZN(n738) );
  NOR2_X1 U828 ( .A1(G2090), .A2(n736), .ZN(n737) );
  NOR2_X1 U829 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U830 ( .A1(G303), .A2(n739), .ZN(n740) );
  XNOR2_X1 U831 ( .A(n740), .B(KEYINPUT96), .ZN(n741) );
  OR2_X1 U832 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U833 ( .A1(G8), .A2(n746), .ZN(n747) );
  NAND2_X1 U834 ( .A1(n748), .A2(n747), .ZN(n749) );
  NOR2_X1 U835 ( .A1(n750), .A2(n749), .ZN(n751) );
  NOR2_X2 U836 ( .A1(n516), .A2(n751), .ZN(n801) );
  NOR2_X1 U837 ( .A1(G1976), .A2(G288), .ZN(n971) );
  NOR2_X1 U838 ( .A1(G303), .A2(G1971), .ZN(n752) );
  XOR2_X1 U839 ( .A(n752), .B(KEYINPUT97), .Z(n753) );
  NOR2_X1 U840 ( .A1(n971), .A2(n753), .ZN(n754) );
  XOR2_X1 U841 ( .A(KEYINPUT98), .B(n754), .Z(n755) );
  NOR2_X1 U842 ( .A1(n801), .A2(n755), .ZN(n758) );
  NAND2_X1 U843 ( .A1(G1976), .A2(G288), .ZN(n968) );
  NOR2_X1 U844 ( .A1(KEYINPUT99), .A2(n807), .ZN(n756) );
  NAND2_X1 U845 ( .A1(n968), .A2(n756), .ZN(n757) );
  NOR2_X1 U846 ( .A1(n758), .A2(n757), .ZN(n759) );
  NOR2_X1 U847 ( .A1(n759), .A2(KEYINPUT33), .ZN(n766) );
  INV_X1 U848 ( .A(KEYINPUT99), .ZN(n761) );
  NAND2_X1 U849 ( .A1(n971), .A2(KEYINPUT33), .ZN(n760) );
  NAND2_X1 U850 ( .A1(n761), .A2(n760), .ZN(n763) );
  NAND2_X1 U851 ( .A1(n971), .A2(KEYINPUT99), .ZN(n762) );
  NAND2_X1 U852 ( .A1(n763), .A2(n762), .ZN(n764) );
  NOR2_X1 U853 ( .A1(n807), .A2(n764), .ZN(n765) );
  XOR2_X1 U854 ( .A(G1981), .B(G305), .Z(n983) );
  NOR2_X1 U855 ( .A1(n768), .A2(n767), .ZN(n828) );
  NAND2_X1 U856 ( .A1(G140), .A2(n892), .ZN(n770) );
  NAND2_X1 U857 ( .A1(G104), .A2(n893), .ZN(n769) );
  NAND2_X1 U858 ( .A1(n770), .A2(n769), .ZN(n771) );
  XNOR2_X1 U859 ( .A(KEYINPUT34), .B(n771), .ZN(n776) );
  NAND2_X1 U860 ( .A1(G128), .A2(n888), .ZN(n773) );
  NAND2_X1 U861 ( .A1(G116), .A2(n889), .ZN(n772) );
  NAND2_X1 U862 ( .A1(n773), .A2(n772), .ZN(n774) );
  XOR2_X1 U863 ( .A(KEYINPUT35), .B(n774), .Z(n775) );
  NOR2_X1 U864 ( .A1(n776), .A2(n775), .ZN(n777) );
  XOR2_X1 U865 ( .A(KEYINPUT36), .B(n777), .Z(n870) );
  XOR2_X1 U866 ( .A(G2067), .B(KEYINPUT37), .Z(n825) );
  AND2_X1 U867 ( .A1(n870), .A2(n825), .ZN(n920) );
  NAND2_X1 U868 ( .A1(n828), .A2(n920), .ZN(n778) );
  XOR2_X1 U869 ( .A(KEYINPUT89), .B(n778), .Z(n823) );
  NAND2_X1 U870 ( .A1(G131), .A2(n892), .ZN(n780) );
  NAND2_X1 U871 ( .A1(G95), .A2(n893), .ZN(n779) );
  NAND2_X1 U872 ( .A1(n780), .A2(n779), .ZN(n781) );
  XOR2_X1 U873 ( .A(KEYINPUT90), .B(n781), .Z(n785) );
  NAND2_X1 U874 ( .A1(G119), .A2(n888), .ZN(n783) );
  NAND2_X1 U875 ( .A1(G107), .A2(n889), .ZN(n782) );
  AND2_X1 U876 ( .A1(n783), .A2(n782), .ZN(n784) );
  NAND2_X1 U877 ( .A1(n785), .A2(n784), .ZN(n869) );
  AND2_X1 U878 ( .A1(n869), .A2(G1991), .ZN(n795) );
  NAND2_X1 U879 ( .A1(G105), .A2(n893), .ZN(n786) );
  XNOR2_X1 U880 ( .A(n786), .B(KEYINPUT38), .ZN(n793) );
  NAND2_X1 U881 ( .A1(G129), .A2(n888), .ZN(n788) );
  NAND2_X1 U882 ( .A1(G117), .A2(n889), .ZN(n787) );
  NAND2_X1 U883 ( .A1(n788), .A2(n787), .ZN(n791) );
  NAND2_X1 U884 ( .A1(G141), .A2(n892), .ZN(n789) );
  XNOR2_X1 U885 ( .A(KEYINPUT91), .B(n789), .ZN(n790) );
  NOR2_X1 U886 ( .A1(n791), .A2(n790), .ZN(n792) );
  NAND2_X1 U887 ( .A1(n793), .A2(n792), .ZN(n899) );
  AND2_X1 U888 ( .A1(n899), .A2(G1996), .ZN(n794) );
  NOR2_X1 U889 ( .A1(n795), .A2(n794), .ZN(n924) );
  INV_X1 U890 ( .A(n924), .ZN(n796) );
  NAND2_X1 U891 ( .A1(n796), .A2(n828), .ZN(n817) );
  AND2_X1 U892 ( .A1(n823), .A2(n817), .ZN(n812) );
  AND2_X1 U893 ( .A1(n983), .A2(n812), .ZN(n797) );
  NAND2_X1 U894 ( .A1(n798), .A2(n797), .ZN(n814) );
  NOR2_X1 U895 ( .A1(G303), .A2(G2090), .ZN(n799) );
  NAND2_X1 U896 ( .A1(G8), .A2(n799), .ZN(n800) );
  XNOR2_X1 U897 ( .A(n800), .B(KEYINPUT100), .ZN(n803) );
  INV_X1 U898 ( .A(n801), .ZN(n802) );
  NAND2_X1 U899 ( .A1(n803), .A2(n802), .ZN(n804) );
  NAND2_X1 U900 ( .A1(n804), .A2(n807), .ZN(n810) );
  NOR2_X1 U901 ( .A1(G1981), .A2(G305), .ZN(n805) );
  XOR2_X1 U902 ( .A(n805), .B(KEYINPUT24), .Z(n806) );
  NOR2_X1 U903 ( .A1(n807), .A2(n806), .ZN(n808) );
  XNOR2_X1 U904 ( .A(KEYINPUT93), .B(n808), .ZN(n809) );
  NAND2_X1 U905 ( .A1(n810), .A2(n809), .ZN(n811) );
  NAND2_X1 U906 ( .A1(n812), .A2(n811), .ZN(n813) );
  NAND2_X1 U907 ( .A1(n814), .A2(n813), .ZN(n816) );
  XNOR2_X1 U908 ( .A(G1986), .B(G290), .ZN(n974) );
  NAND2_X1 U909 ( .A1(n974), .A2(n828), .ZN(n815) );
  NAND2_X1 U910 ( .A1(n816), .A2(n815), .ZN(n831) );
  NOR2_X1 U911 ( .A1(G1996), .A2(n899), .ZN(n927) );
  INV_X1 U912 ( .A(n817), .ZN(n820) );
  NOR2_X1 U913 ( .A1(G1986), .A2(G290), .ZN(n818) );
  NOR2_X1 U914 ( .A1(G1991), .A2(n869), .ZN(n919) );
  NOR2_X1 U915 ( .A1(n818), .A2(n919), .ZN(n819) );
  NOR2_X1 U916 ( .A1(n820), .A2(n819), .ZN(n821) );
  NOR2_X1 U917 ( .A1(n927), .A2(n821), .ZN(n822) );
  XNOR2_X1 U918 ( .A(n822), .B(KEYINPUT39), .ZN(n824) );
  NAND2_X1 U919 ( .A1(n824), .A2(n823), .ZN(n827) );
  NOR2_X1 U920 ( .A1(n825), .A2(n870), .ZN(n826) );
  XNOR2_X1 U921 ( .A(n826), .B(KEYINPUT101), .ZN(n932) );
  NAND2_X1 U922 ( .A1(n827), .A2(n932), .ZN(n829) );
  NAND2_X1 U923 ( .A1(n829), .A2(n828), .ZN(n830) );
  NAND2_X1 U924 ( .A1(n831), .A2(n830), .ZN(n833) );
  XNOR2_X1 U925 ( .A(KEYINPUT102), .B(KEYINPUT40), .ZN(n832) );
  XNOR2_X1 U926 ( .A(n833), .B(n832), .ZN(G329) );
  NAND2_X1 U927 ( .A1(n835), .A2(G2106), .ZN(n834) );
  XNOR2_X1 U928 ( .A(n834), .B(KEYINPUT106), .ZN(G217) );
  INV_X1 U929 ( .A(n835), .ZN(G223) );
  AND2_X1 U930 ( .A1(G15), .A2(G2), .ZN(n836) );
  NAND2_X1 U931 ( .A1(G661), .A2(n836), .ZN(G259) );
  NAND2_X1 U932 ( .A1(G3), .A2(G1), .ZN(n837) );
  NAND2_X1 U933 ( .A1(n838), .A2(n837), .ZN(G188) );
  INV_X1 U934 ( .A(n839), .ZN(G319) );
  XNOR2_X1 U935 ( .A(G2078), .B(G2072), .ZN(n841) );
  XOR2_X1 U936 ( .A(n841), .B(n840), .Z(n851) );
  XOR2_X1 U937 ( .A(KEYINPUT108), .B(G2678), .Z(n843) );
  XNOR2_X1 U938 ( .A(KEYINPUT109), .B(KEYINPUT42), .ZN(n842) );
  XNOR2_X1 U939 ( .A(n843), .B(n842), .ZN(n847) );
  XOR2_X1 U940 ( .A(KEYINPUT107), .B(G2096), .Z(n845) );
  XNOR2_X1 U941 ( .A(G2090), .B(KEYINPUT43), .ZN(n844) );
  XNOR2_X1 U942 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U943 ( .A(n847), .B(n846), .Z(n849) );
  XNOR2_X1 U944 ( .A(G2067), .B(G2084), .ZN(n848) );
  XNOR2_X1 U945 ( .A(n849), .B(n848), .ZN(n850) );
  XNOR2_X1 U946 ( .A(n851), .B(n850), .ZN(G227) );
  XOR2_X1 U947 ( .A(G1971), .B(G1961), .Z(n853) );
  XNOR2_X1 U948 ( .A(G1986), .B(G1966), .ZN(n852) );
  XNOR2_X1 U949 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U950 ( .A(n854), .B(KEYINPUT41), .Z(n856) );
  XNOR2_X1 U951 ( .A(G1996), .B(G1956), .ZN(n855) );
  XNOR2_X1 U952 ( .A(n856), .B(n855), .ZN(n860) );
  XOR2_X1 U953 ( .A(G2474), .B(G1976), .Z(n858) );
  XNOR2_X1 U954 ( .A(G1991), .B(G1981), .ZN(n857) );
  XNOR2_X1 U955 ( .A(n858), .B(n857), .ZN(n859) );
  XNOR2_X1 U956 ( .A(n860), .B(n859), .ZN(G229) );
  NAND2_X1 U957 ( .A1(G124), .A2(n888), .ZN(n861) );
  XNOR2_X1 U958 ( .A(n861), .B(KEYINPUT110), .ZN(n862) );
  XNOR2_X1 U959 ( .A(n862), .B(KEYINPUT44), .ZN(n864) );
  NAND2_X1 U960 ( .A1(G112), .A2(n889), .ZN(n863) );
  NAND2_X1 U961 ( .A1(n864), .A2(n863), .ZN(n868) );
  NAND2_X1 U962 ( .A1(G136), .A2(n892), .ZN(n866) );
  NAND2_X1 U963 ( .A1(G100), .A2(n893), .ZN(n865) );
  NAND2_X1 U964 ( .A1(n866), .A2(n865), .ZN(n867) );
  NOR2_X1 U965 ( .A1(n868), .A2(n867), .ZN(G162) );
  XNOR2_X1 U966 ( .A(G162), .B(n869), .ZN(n872) );
  XNOR2_X1 U967 ( .A(G160), .B(n870), .ZN(n871) );
  XNOR2_X1 U968 ( .A(n872), .B(n871), .ZN(n876) );
  XOR2_X1 U969 ( .A(KEYINPUT114), .B(KEYINPUT111), .Z(n874) );
  XNOR2_X1 U970 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n873) );
  XNOR2_X1 U971 ( .A(n874), .B(n873), .ZN(n875) );
  XOR2_X1 U972 ( .A(n876), .B(n875), .Z(n887) );
  NAND2_X1 U973 ( .A1(G139), .A2(n892), .ZN(n878) );
  NAND2_X1 U974 ( .A1(G103), .A2(n893), .ZN(n877) );
  NAND2_X1 U975 ( .A1(n878), .A2(n877), .ZN(n884) );
  NAND2_X1 U976 ( .A1(G127), .A2(n888), .ZN(n880) );
  NAND2_X1 U977 ( .A1(G115), .A2(n889), .ZN(n879) );
  NAND2_X1 U978 ( .A1(n880), .A2(n879), .ZN(n881) );
  XOR2_X1 U979 ( .A(KEYINPUT47), .B(n881), .Z(n882) );
  XNOR2_X1 U980 ( .A(KEYINPUT112), .B(n882), .ZN(n883) );
  NOR2_X1 U981 ( .A1(n884), .A2(n883), .ZN(n885) );
  XOR2_X1 U982 ( .A(KEYINPUT113), .B(n885), .Z(n934) );
  XNOR2_X1 U983 ( .A(G164), .B(n934), .ZN(n886) );
  XNOR2_X1 U984 ( .A(n887), .B(n886), .ZN(n903) );
  NAND2_X1 U985 ( .A1(G130), .A2(n888), .ZN(n891) );
  NAND2_X1 U986 ( .A1(G118), .A2(n889), .ZN(n890) );
  NAND2_X1 U987 ( .A1(n891), .A2(n890), .ZN(n898) );
  NAND2_X1 U988 ( .A1(G142), .A2(n892), .ZN(n895) );
  NAND2_X1 U989 ( .A1(G106), .A2(n893), .ZN(n894) );
  NAND2_X1 U990 ( .A1(n895), .A2(n894), .ZN(n896) );
  XOR2_X1 U991 ( .A(n896), .B(KEYINPUT45), .Z(n897) );
  NOR2_X1 U992 ( .A1(n898), .A2(n897), .ZN(n900) );
  XNOR2_X1 U993 ( .A(n900), .B(n899), .ZN(n901) );
  XNOR2_X1 U994 ( .A(n918), .B(n901), .ZN(n902) );
  XNOR2_X1 U995 ( .A(n903), .B(n902), .ZN(n904) );
  NOR2_X1 U996 ( .A1(G37), .A2(n904), .ZN(G395) );
  XOR2_X1 U997 ( .A(n905), .B(n972), .Z(n906) );
  XNOR2_X1 U998 ( .A(n906), .B(n977), .ZN(n908) );
  XNOR2_X1 U999 ( .A(G286), .B(G301), .ZN(n907) );
  XNOR2_X1 U1000 ( .A(n908), .B(n907), .ZN(n909) );
  NOR2_X1 U1001 ( .A1(G37), .A2(n909), .ZN(n910) );
  XOR2_X1 U1002 ( .A(KEYINPUT115), .B(n910), .Z(G397) );
  NOR2_X1 U1003 ( .A1(G227), .A2(G229), .ZN(n911) );
  XOR2_X1 U1004 ( .A(KEYINPUT49), .B(n911), .Z(n912) );
  NAND2_X1 U1005 ( .A1(G319), .A2(n912), .ZN(n913) );
  NOR2_X1 U1006 ( .A1(G401), .A2(n913), .ZN(n914) );
  XNOR2_X1 U1007 ( .A(KEYINPUT116), .B(n914), .ZN(n916) );
  NOR2_X1 U1008 ( .A1(G395), .A2(G397), .ZN(n915) );
  NAND2_X1 U1009 ( .A1(n916), .A2(n915), .ZN(G225) );
  XNOR2_X1 U1010 ( .A(KEYINPUT117), .B(G225), .ZN(G308) );
  XOR2_X1 U1011 ( .A(G108), .B(KEYINPUT118), .Z(G238) );
  XOR2_X1 U1013 ( .A(G2084), .B(G160), .Z(n917) );
  NOR2_X1 U1014 ( .A1(n918), .A2(n917), .ZN(n922) );
  NOR2_X1 U1015 ( .A1(n920), .A2(n919), .ZN(n921) );
  NAND2_X1 U1016 ( .A1(n922), .A2(n921), .ZN(n923) );
  XNOR2_X1 U1017 ( .A(KEYINPUT119), .B(n923), .ZN(n925) );
  NAND2_X1 U1018 ( .A1(n925), .A2(n924), .ZN(n930) );
  XOR2_X1 U1019 ( .A(G2090), .B(G162), .Z(n926) );
  NOR2_X1 U1020 ( .A1(n927), .A2(n926), .ZN(n928) );
  XNOR2_X1 U1021 ( .A(n928), .B(KEYINPUT51), .ZN(n929) );
  NOR2_X1 U1022 ( .A1(n930), .A2(n929), .ZN(n931) );
  XNOR2_X1 U1023 ( .A(n931), .B(KEYINPUT120), .ZN(n933) );
  NAND2_X1 U1024 ( .A1(n933), .A2(n932), .ZN(n939) );
  XOR2_X1 U1025 ( .A(G2072), .B(n934), .Z(n936) );
  XOR2_X1 U1026 ( .A(G164), .B(G2078), .Z(n935) );
  NOR2_X1 U1027 ( .A1(n936), .A2(n935), .ZN(n937) );
  XOR2_X1 U1028 ( .A(KEYINPUT50), .B(n937), .Z(n938) );
  NOR2_X1 U1029 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1030 ( .A(KEYINPUT52), .B(n940), .ZN(n942) );
  INV_X1 U1031 ( .A(KEYINPUT55), .ZN(n941) );
  NAND2_X1 U1032 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1033 ( .A1(n943), .A2(G29), .ZN(n1020) );
  XNOR2_X1 U1034 ( .A(G2090), .B(G35), .ZN(n959) );
  XOR2_X1 U1035 ( .A(G1991), .B(G25), .Z(n944) );
  NAND2_X1 U1036 ( .A1(n944), .A2(G28), .ZN(n945) );
  XNOR2_X1 U1037 ( .A(n945), .B(KEYINPUT121), .ZN(n954) );
  XNOR2_X1 U1038 ( .A(n946), .B(G27), .ZN(n952) );
  XNOR2_X1 U1039 ( .A(G2072), .B(KEYINPUT122), .ZN(n947) );
  XNOR2_X1 U1040 ( .A(n947), .B(G33), .ZN(n949) );
  XNOR2_X1 U1041 ( .A(G26), .B(G2067), .ZN(n948) );
  NOR2_X1 U1042 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1043 ( .A(KEYINPUT123), .B(n950), .ZN(n951) );
  NOR2_X1 U1044 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1045 ( .A1(n954), .A2(n953), .ZN(n956) );
  XNOR2_X1 U1046 ( .A(G32), .B(G1996), .ZN(n955) );
  NOR2_X1 U1047 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1048 ( .A(KEYINPUT53), .B(n957), .ZN(n958) );
  NOR2_X1 U1049 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1050 ( .A(n960), .B(KEYINPUT124), .ZN(n963) );
  XOR2_X1 U1051 ( .A(G2084), .B(G34), .Z(n961) );
  XNOR2_X1 U1052 ( .A(KEYINPUT54), .B(n961), .ZN(n962) );
  NAND2_X1 U1053 ( .A1(n963), .A2(n962), .ZN(n964) );
  XOR2_X1 U1054 ( .A(KEYINPUT55), .B(n964), .Z(n966) );
  INV_X1 U1055 ( .A(G29), .ZN(n965) );
  NAND2_X1 U1056 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1057 ( .A1(G11), .A2(n967), .ZN(n1018) );
  INV_X1 U1058 ( .A(G16), .ZN(n1014) );
  XOR2_X1 U1059 ( .A(n1014), .B(KEYINPUT56), .Z(n991) );
  XOR2_X1 U1060 ( .A(G1956), .B(G299), .Z(n969) );
  NAND2_X1 U1061 ( .A1(n969), .A2(n968), .ZN(n970) );
  NOR2_X1 U1062 ( .A1(n971), .A2(n970), .ZN(n976) );
  XOR2_X1 U1063 ( .A(G1348), .B(n972), .Z(n973) );
  NOR2_X1 U1064 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1065 ( .A1(n976), .A2(n975), .ZN(n980) );
  XOR2_X1 U1066 ( .A(G1341), .B(n977), .Z(n978) );
  XNOR2_X1 U1067 ( .A(KEYINPUT125), .B(n978), .ZN(n979) );
  NOR2_X1 U1068 ( .A1(n980), .A2(n979), .ZN(n989) );
  XOR2_X1 U1069 ( .A(G303), .B(G1971), .Z(n982) );
  XOR2_X1 U1070 ( .A(G301), .B(G1961), .Z(n981) );
  NAND2_X1 U1071 ( .A1(n982), .A2(n981), .ZN(n987) );
  XNOR2_X1 U1072 ( .A(G1966), .B(G168), .ZN(n984) );
  NAND2_X1 U1073 ( .A1(n984), .A2(n983), .ZN(n985) );
  XOR2_X1 U1074 ( .A(KEYINPUT57), .B(n985), .Z(n986) );
  NOR2_X1 U1075 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1076 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1077 ( .A1(n991), .A2(n990), .ZN(n1016) );
  XNOR2_X1 U1078 ( .A(G1348), .B(KEYINPUT59), .ZN(n992) );
  XNOR2_X1 U1079 ( .A(n992), .B(G4), .ZN(n996) );
  XNOR2_X1 U1080 ( .A(G1956), .B(G20), .ZN(n994) );
  XNOR2_X1 U1081 ( .A(G1341), .B(G19), .ZN(n993) );
  NOR2_X1 U1082 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1083 ( .A1(n996), .A2(n995), .ZN(n999) );
  XNOR2_X1 U1084 ( .A(KEYINPUT126), .B(G1981), .ZN(n997) );
  XNOR2_X1 U1085 ( .A(G6), .B(n997), .ZN(n998) );
  NOR2_X1 U1086 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XNOR2_X1 U1087 ( .A(KEYINPUT60), .B(n1000), .ZN(n1004) );
  XNOR2_X1 U1088 ( .A(G1966), .B(G21), .ZN(n1002) );
  XNOR2_X1 U1089 ( .A(G1961), .B(G5), .ZN(n1001) );
  NOR2_X1 U1090 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1091 ( .A1(n1004), .A2(n1003), .ZN(n1011) );
  XNOR2_X1 U1092 ( .A(G1976), .B(G23), .ZN(n1006) );
  XNOR2_X1 U1093 ( .A(G1971), .B(G22), .ZN(n1005) );
  NOR2_X1 U1094 ( .A1(n1006), .A2(n1005), .ZN(n1008) );
  XOR2_X1 U1095 ( .A(G1986), .B(G24), .Z(n1007) );
  NAND2_X1 U1096 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1097 ( .A(KEYINPUT58), .B(n1009), .ZN(n1010) );
  NOR2_X1 U1098 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1099 ( .A(KEYINPUT61), .B(n1012), .ZN(n1013) );
  NAND2_X1 U1100 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1101 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NOR2_X1 U1102 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1103 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XOR2_X1 U1104 ( .A(KEYINPUT62), .B(n1021), .Z(G311) );
  XNOR2_X1 U1105 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1106 ( .A(G120), .ZN(G236) );
  INV_X1 U1107 ( .A(G96), .ZN(G221) );
  NOR2_X1 U1108 ( .A1(n1023), .A2(n1022), .ZN(G325) );
  INV_X1 U1109 ( .A(G325), .ZN(G261) );
  INV_X1 U1110 ( .A(G69), .ZN(G235) );
endmodule

