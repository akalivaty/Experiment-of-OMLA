//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 1 1 0 1 1 1 0 1 0 0 0 1 1 1 0 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 0 1 1 1 0 0 1 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:57 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n720, new_n721, new_n722, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n744, new_n745, new_n746, new_n747, new_n749, new_n750,
    new_n751, new_n752, new_n754, new_n755, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n788, new_n789,
    new_n791, new_n792, new_n793, new_n794, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n844, new_n845, new_n846, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n898, new_n899, new_n901, new_n902, new_n903,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n913, new_n914, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n958, new_n959, new_n960;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202));
  OAI21_X1  g001(.A(KEYINPUT66), .B1(G169gat), .B2(G176gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT68), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT26), .ZN(new_n206));
  OAI21_X1  g005(.A(KEYINPUT66), .B1(new_n206), .B2(KEYINPUT68), .ZN(new_n207));
  NOR2_X1   g006(.A1(G169gat), .A2(G176gat), .ZN(new_n208));
  AOI22_X1  g007(.A1(new_n205), .A2(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(G169gat), .A2(G176gat), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n202), .B1(new_n209), .B2(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(KEYINPUT27), .B(G183gat), .ZN(new_n213));
  INV_X1    g012(.A(G190gat), .ZN(new_n214));
  AOI21_X1  g013(.A(KEYINPUT28), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  AND2_X1   g014(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n216));
  NOR2_X1   g015(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n217));
  OAI211_X1 g016(.A(KEYINPUT28), .B(new_n214), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(new_n218), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n215), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g019(.A(KEYINPUT69), .B1(new_n212), .B2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n213), .A2(new_n214), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT28), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(new_n218), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT69), .ZN(new_n226));
  AND2_X1   g025(.A1(new_n207), .A2(new_n208), .ZN(new_n227));
  AOI21_X1  g026(.A(KEYINPUT26), .B1(new_n203), .B2(new_n204), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n210), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  NAND4_X1  g028(.A1(new_n225), .A2(new_n226), .A3(new_n202), .A4(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n221), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(G176gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(KEYINPUT65), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT65), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(G176gat), .ZN(new_n235));
  AOI21_X1  g034(.A(G169gat), .B1(new_n233), .B2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(new_n208), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n210), .A2(KEYINPUT23), .ZN(new_n238));
  AOI22_X1  g037(.A1(new_n236), .A2(KEYINPUT23), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT64), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n240), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT24), .ZN(new_n242));
  AOI21_X1  g041(.A(KEYINPUT64), .B1(new_n202), .B2(new_n242), .ZN(new_n243));
  NAND3_X1  g042(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  OAI221_X1 g044(.A(new_n241), .B1(G183gat), .B2(G190gat), .C1(new_n243), .C2(new_n245), .ZN(new_n246));
  AOI21_X1  g045(.A(KEYINPUT25), .B1(new_n239), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n202), .A2(new_n242), .ZN(new_n248));
  OAI211_X1 g047(.A(new_n248), .B(new_n244), .C1(G183gat), .C2(G190gat), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT66), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n208), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n251), .A2(KEYINPUT23), .A3(new_n203), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n238), .B1(G169gat), .B2(G176gat), .ZN(new_n253));
  NAND4_X1  g052(.A1(new_n249), .A2(new_n252), .A3(new_n253), .A4(KEYINPUT25), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT67), .ZN(new_n256));
  NOR3_X1   g055(.A1(new_n247), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT25), .ZN(new_n258));
  INV_X1    g057(.A(G169gat), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n234), .A2(G176gat), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n232), .A2(KEYINPUT65), .ZN(new_n261));
  OAI211_X1 g060(.A(KEYINPUT23), .B(new_n259), .C1(new_n260), .C2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(new_n253), .ZN(new_n263));
  OAI22_X1  g062(.A1(new_n244), .A2(KEYINPUT64), .B1(G183gat), .B2(G190gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n240), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n264), .B1(new_n244), .B2(new_n265), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n258), .B1(new_n263), .B2(new_n266), .ZN(new_n267));
  AOI21_X1  g066(.A(KEYINPUT67), .B1(new_n267), .B2(new_n254), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n231), .B1(new_n257), .B2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT1), .ZN(new_n270));
  XNOR2_X1  g069(.A(G127gat), .B(G134gat), .ZN(new_n271));
  INV_X1    g070(.A(G113gat), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n272), .A2(KEYINPUT70), .A3(G120gat), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n273), .B1(new_n272), .B2(G120gat), .ZN(new_n274));
  AOI21_X1  g073(.A(KEYINPUT70), .B1(new_n272), .B2(G120gat), .ZN(new_n275));
  OAI211_X1 g074(.A(new_n270), .B(new_n271), .C1(new_n274), .C2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n271), .ZN(new_n277));
  XNOR2_X1  g076(.A(G113gat), .B(G120gat), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n277), .B1(KEYINPUT1), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n276), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT71), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n276), .A2(new_n279), .A3(KEYINPUT71), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n269), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(G227gat), .ZN(new_n285));
  INV_X1    g084(.A(G233gat), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n256), .B1(new_n247), .B2(new_n255), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n267), .A2(KEYINPUT67), .A3(new_n254), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND4_X1  g089(.A1(new_n290), .A2(new_n281), .A3(new_n280), .A4(new_n231), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n284), .A2(new_n287), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(KEYINPUT32), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT33), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(KEYINPUT72), .B(G71gat), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n296), .B(G99gat), .ZN(new_n297));
  XNOR2_X1  g096(.A(G15gat), .B(G43gat), .ZN(new_n298));
  XOR2_X1   g097(.A(new_n297), .B(new_n298), .Z(new_n299));
  NAND3_X1  g098(.A1(new_n293), .A2(new_n295), .A3(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(new_n299), .ZN(new_n301));
  OAI211_X1 g100(.A(new_n292), .B(KEYINPUT32), .C1(new_n294), .C2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n287), .B1(new_n284), .B2(new_n291), .ZN(new_n304));
  AND2_X1   g103(.A1(new_n304), .A2(KEYINPUT34), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n304), .A2(KEYINPUT34), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n303), .A2(new_n307), .ZN(new_n308));
  OAI211_X1 g107(.A(new_n300), .B(new_n302), .C1(new_n306), .C2(new_n305), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(G228gat), .A2(G233gat), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT29), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT80), .ZN(new_n313));
  AND2_X1   g112(.A1(G155gat), .A2(G162gat), .ZN(new_n314));
  NOR2_X1   g113(.A1(G155gat), .A2(G162gat), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  AND2_X1   g115(.A1(KEYINPUT79), .A2(G141gat), .ZN(new_n317));
  NOR2_X1   g116(.A1(KEYINPUT79), .A2(G141gat), .ZN(new_n318));
  OAI21_X1  g117(.A(G148gat), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(G141gat), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n320), .A2(G148gat), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n316), .B1(new_n319), .B2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT2), .ZN(new_n324));
  OR2_X1    g123(.A1(new_n314), .A2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(G148gat), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n326), .A2(G141gat), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n324), .B1(new_n321), .B2(new_n327), .ZN(new_n328));
  AOI22_X1  g127(.A1(new_n323), .A2(new_n325), .B1(new_n316), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT3), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n313), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  OR2_X1    g130(.A1(new_n314), .A2(new_n315), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT79), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(new_n320), .ZN(new_n334));
  NAND2_X1  g133(.A1(KEYINPUT79), .A2(G141gat), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n326), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  OAI211_X1 g135(.A(new_n332), .B(new_n325), .C1(new_n336), .C2(new_n321), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n328), .A2(new_n316), .ZN(new_n338));
  NAND4_X1  g137(.A1(new_n337), .A2(new_n313), .A3(new_n330), .A4(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n312), .B1(new_n331), .B2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT85), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  XOR2_X1   g142(.A(G211gat), .B(G218gat), .Z(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n345), .A2(KEYINPUT75), .ZN(new_n346));
  OR2_X1    g145(.A1(KEYINPUT74), .A2(G204gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(KEYINPUT74), .A2(G204gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(G197gat), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT22), .ZN(new_n352));
  INV_X1    g151(.A(G211gat), .ZN(new_n353));
  INV_X1    g152(.A(G218gat), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n352), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n347), .A2(G197gat), .A3(new_n348), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n351), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  XNOR2_X1  g156(.A(new_n346), .B(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n337), .A2(new_n330), .A3(new_n338), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(KEYINPUT80), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(new_n339), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n362), .A2(KEYINPUT85), .A3(new_n312), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n343), .A2(new_n359), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n358), .A2(new_n312), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n329), .B1(new_n365), .B2(new_n330), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n311), .B1(new_n364), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n341), .A2(new_n359), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n357), .A2(new_n345), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n337), .A2(new_n338), .ZN(new_n371));
  NAND4_X1  g170(.A1(new_n351), .A2(new_n344), .A3(new_n355), .A4(new_n356), .ZN(new_n372));
  NAND4_X1  g171(.A1(new_n370), .A2(new_n371), .A3(new_n312), .A4(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n371), .A2(KEYINPUT3), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT84), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n373), .A2(KEYINPUT84), .A3(new_n374), .ZN(new_n378));
  NAND4_X1  g177(.A1(new_n369), .A2(new_n311), .A3(new_n377), .A4(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  OAI21_X1  g179(.A(G50gat), .B1(new_n368), .B2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(G50gat), .ZN(new_n382));
  AOI21_X1  g181(.A(KEYINPUT85), .B1(new_n362), .B2(new_n312), .ZN(new_n383));
  AOI211_X1 g182(.A(new_n342), .B(KEYINPUT29), .C1(new_n361), .C2(new_n339), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n366), .B1(new_n385), .B2(new_n359), .ZN(new_n386));
  OAI211_X1 g185(.A(new_n382), .B(new_n379), .C1(new_n386), .C2(new_n311), .ZN(new_n387));
  XNOR2_X1  g186(.A(G78gat), .B(G106gat), .ZN(new_n388));
  XNOR2_X1  g187(.A(new_n388), .B(G22gat), .ZN(new_n389));
  XOR2_X1   g188(.A(KEYINPUT83), .B(KEYINPUT31), .Z(new_n390));
  XOR2_X1   g189(.A(new_n389), .B(new_n390), .Z(new_n391));
  AND3_X1   g190(.A1(new_n381), .A2(new_n387), .A3(new_n391), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n391), .B1(new_n381), .B2(new_n387), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  OAI21_X1  g193(.A(KEYINPUT90), .B1(new_n310), .B2(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n362), .A2(new_n280), .A3(new_n374), .ZN(new_n396));
  NAND4_X1  g195(.A1(new_n337), .A2(new_n276), .A3(new_n338), .A4(new_n279), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(KEYINPUT4), .ZN(new_n398));
  XNOR2_X1  g197(.A(KEYINPUT81), .B(KEYINPUT4), .ZN(new_n399));
  OAI211_X1 g198(.A(new_n398), .B(KEYINPUT82), .C1(new_n397), .C2(new_n399), .ZN(new_n400));
  OR3_X1    g199(.A1(new_n397), .A2(KEYINPUT82), .A3(new_n399), .ZN(new_n401));
  NAND2_X1  g200(.A1(G225gat), .A2(G233gat), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n403), .A2(KEYINPUT5), .ZN(new_n404));
  AND4_X1   g203(.A1(new_n396), .A2(new_n400), .A3(new_n401), .A4(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(new_n397), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(KEYINPUT4), .ZN(new_n407));
  INV_X1    g206(.A(new_n399), .ZN(new_n408));
  AOI22_X1  g207(.A1(new_n361), .A2(new_n339), .B1(KEYINPUT3), .B2(new_n371), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n408), .B1(new_n409), .B2(new_n280), .ZN(new_n410));
  OAI211_X1 g209(.A(new_n402), .B(new_n407), .C1(new_n410), .C2(new_n406), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n371), .A2(new_n280), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(new_n397), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(new_n403), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(KEYINPUT5), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n405), .B1(new_n411), .B2(new_n416), .ZN(new_n417));
  XNOR2_X1  g216(.A(KEYINPUT0), .B(G57gat), .ZN(new_n418));
  XNOR2_X1  g217(.A(new_n418), .B(G85gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(G1gat), .B(G29gat), .ZN(new_n420));
  XOR2_X1   g219(.A(new_n419), .B(new_n420), .Z(new_n421));
  AOI21_X1  g220(.A(KEYINPUT6), .B1(new_n417), .B2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(new_n421), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n396), .A2(new_n399), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n403), .B1(new_n424), .B2(new_n397), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n415), .B1(new_n425), .B2(new_n407), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n423), .B1(new_n426), .B2(new_n405), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n422), .A2(new_n427), .ZN(new_n428));
  OAI211_X1 g227(.A(KEYINPUT6), .B(new_n423), .C1(new_n426), .C2(new_n405), .ZN(new_n429));
  NAND2_X1  g228(.A1(G226gat), .A2(G233gat), .ZN(new_n430));
  XOR2_X1   g229(.A(new_n430), .B(KEYINPUT76), .Z(new_n431));
  NAND2_X1  g230(.A1(new_n269), .A2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT77), .ZN(new_n433));
  INV_X1    g232(.A(new_n431), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n212), .A2(new_n220), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n435), .B1(new_n267), .B2(new_n254), .ZN(new_n436));
  OAI211_X1 g235(.A(new_n433), .B(new_n434), .C1(new_n436), .C2(KEYINPUT29), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n267), .A2(new_n254), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n225), .A2(new_n202), .A3(new_n229), .ZN(new_n439));
  AOI21_X1  g238(.A(KEYINPUT29), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  OAI21_X1  g239(.A(KEYINPUT77), .B1(new_n440), .B2(new_n431), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n432), .A2(new_n437), .A3(new_n441), .A4(new_n358), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n436), .A2(new_n431), .ZN(new_n443));
  AOI22_X1  g242(.A1(new_n288), .A2(new_n289), .B1(new_n221), .B2(new_n230), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n434), .A2(new_n312), .ZN(new_n445));
  OAI211_X1 g244(.A(new_n443), .B(new_n359), .C1(new_n444), .C2(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n442), .A2(new_n446), .ZN(new_n447));
  XOR2_X1   g246(.A(G8gat), .B(G36gat), .Z(new_n448));
  XNOR2_X1  g247(.A(new_n448), .B(G64gat), .ZN(new_n449));
  XNOR2_X1  g248(.A(new_n449), .B(G92gat), .ZN(new_n450));
  XNOR2_X1  g249(.A(new_n450), .B(KEYINPUT78), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n447), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n442), .A2(new_n446), .A3(new_n450), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n452), .A2(KEYINPUT30), .A3(new_n453), .ZN(new_n454));
  OR2_X1    g253(.A1(new_n453), .A2(KEYINPUT30), .ZN(new_n455));
  AOI22_X1  g254(.A1(new_n428), .A2(new_n429), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n381), .A2(new_n387), .ZN(new_n457));
  INV_X1    g256(.A(new_n391), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n381), .A2(new_n387), .A3(new_n391), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT90), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n461), .A2(new_n462), .A3(new_n308), .A4(new_n309), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n395), .A2(new_n456), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(KEYINPUT35), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n308), .A2(KEYINPUT73), .A3(new_n309), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT73), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n303), .A2(new_n467), .A3(new_n307), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT35), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n469), .A2(new_n470), .A3(new_n456), .A4(new_n461), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n465), .A2(new_n471), .ZN(new_n472));
  AOI21_X1  g271(.A(KEYINPUT36), .B1(new_n466), .B2(new_n468), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n456), .A2(new_n461), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT36), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n475), .B1(new_n308), .B2(new_n309), .ZN(new_n476));
  NOR3_X1   g275(.A1(new_n473), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT38), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n453), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n447), .A2(KEYINPUT37), .ZN(new_n480));
  XNOR2_X1  g279(.A(KEYINPUT89), .B(KEYINPUT37), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n480), .B1(new_n447), .B2(new_n481), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n479), .B1(new_n482), .B2(new_n450), .ZN(new_n483));
  OAI211_X1 g282(.A(new_n443), .B(new_n358), .C1(new_n444), .C2(new_n445), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n432), .A2(new_n437), .A3(new_n441), .ZN(new_n485));
  OAI211_X1 g284(.A(KEYINPUT37), .B(new_n484), .C1(new_n485), .C2(new_n358), .ZN(new_n486));
  AND2_X1   g285(.A1(new_n451), .A2(new_n478), .ZN(new_n487));
  OAI211_X1 g286(.A(new_n486), .B(new_n487), .C1(new_n447), .C2(new_n481), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n483), .A2(new_n429), .A3(new_n488), .A4(new_n428), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n454), .A2(new_n455), .ZN(new_n490));
  INV_X1    g289(.A(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n396), .A2(new_n400), .A3(new_n401), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(new_n403), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n421), .B1(new_n493), .B2(KEYINPUT39), .ZN(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n412), .A2(new_n402), .A3(new_n397), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n493), .A2(KEYINPUT39), .A3(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n495), .A2(KEYINPUT40), .A3(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT88), .ZN(new_n499));
  AND2_X1   g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n498), .A2(new_n499), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n491), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  XOR2_X1   g301(.A(KEYINPUT86), .B(KEYINPUT40), .Z(new_n503));
  INV_X1    g302(.A(new_n497), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n503), .B1(new_n504), .B2(new_n494), .ZN(new_n505));
  OR2_X1    g304(.A1(new_n505), .A2(KEYINPUT87), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(KEYINPUT87), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n506), .A2(new_n427), .A3(new_n507), .ZN(new_n508));
  OAI211_X1 g307(.A(new_n461), .B(new_n489), .C1(new_n502), .C2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n477), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n472), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(G232gat), .A2(G233gat), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n513), .A2(KEYINPUT41), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n514), .B(KEYINPUT98), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n515), .B(G218gat), .ZN(new_n516));
  INV_X1    g315(.A(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT99), .ZN(new_n518));
  INV_X1    g317(.A(G99gat), .ZN(new_n519));
  INV_X1    g318(.A(G106gat), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND3_X1  g320(.A1(KEYINPUT99), .A2(G99gat), .A3(G106gat), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n521), .A2(KEYINPUT8), .A3(new_n522), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n523), .B1(G85gat), .B2(G92gat), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n524), .B(KEYINPUT100), .ZN(new_n525));
  NAND2_X1  g324(.A1(G85gat), .A2(G92gat), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n526), .B(KEYINPUT7), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  XOR2_X1   g327(.A(G99gat), .B(G106gat), .Z(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT101), .ZN(new_n531));
  INV_X1    g330(.A(new_n529), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n525), .A2(new_n532), .A3(new_n527), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n530), .A2(new_n531), .A3(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n528), .A2(KEYINPUT101), .A3(new_n529), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  OR3_X1    g335(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n537));
  OAI21_X1  g336(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n538));
  AOI22_X1  g337(.A1(new_n537), .A2(new_n538), .B1(G29gat), .B2(G36gat), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT15), .ZN(new_n540));
  XOR2_X1   g339(.A(G43gat), .B(G50gat), .Z(new_n541));
  OR3_X1    g340(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  OR2_X1    g341(.A1(new_n541), .A2(new_n540), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n541), .A2(new_n540), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n543), .A2(new_n544), .A3(new_n539), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n536), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n513), .A2(KEYINPUT41), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n542), .A2(new_n545), .A3(KEYINPUT17), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT17), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n546), .A2(new_n550), .ZN(new_n551));
  NAND4_X1  g350(.A1(new_n534), .A2(new_n535), .A3(new_n549), .A4(new_n551), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n547), .A2(new_n548), .A3(new_n552), .ZN(new_n553));
  XNOR2_X1  g352(.A(G134gat), .B(G162gat), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n554), .B(new_n214), .ZN(new_n555));
  AND2_X1   g354(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n553), .A2(new_n555), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n517), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  OR2_X1    g357(.A1(new_n553), .A2(new_n555), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n553), .A2(new_n555), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n559), .A2(new_n516), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(G127gat), .B(G155gat), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n563), .B(G211gat), .ZN(new_n564));
  AOI21_X1  g363(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n565));
  OR2_X1    g364(.A1(new_n565), .A2(KEYINPUT94), .ZN(new_n566));
  XOR2_X1   g365(.A(G57gat), .B(G64gat), .Z(new_n567));
  XNOR2_X1  g366(.A(G71gat), .B(G78gat), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n565), .A2(KEYINPUT94), .ZN(new_n569));
  NAND4_X1  g368(.A1(new_n566), .A2(new_n567), .A3(new_n568), .A4(new_n569), .ZN(new_n570));
  XOR2_X1   g369(.A(G71gat), .B(G78gat), .Z(new_n571));
  INV_X1    g370(.A(KEYINPUT9), .ZN(new_n572));
  XNOR2_X1  g371(.A(G57gat), .B(G64gat), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n571), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n570), .A2(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n575), .B(KEYINPUT97), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(KEYINPUT21), .ZN(new_n577));
  XNOR2_X1  g376(.A(G15gat), .B(G22gat), .ZN(new_n578));
  INV_X1    g377(.A(G1gat), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(KEYINPUT16), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n581), .B1(G1gat), .B2(new_n578), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n582), .A2(G8gat), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n582), .A2(G8gat), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n577), .A2(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n587), .B(G183gat), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n588), .A2(KEYINPUT96), .ZN(new_n589));
  INV_X1    g388(.A(G183gat), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n587), .B(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT96), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(G231gat), .A2(G233gat), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  AND3_X1   g394(.A1(new_n589), .A2(new_n593), .A3(new_n595), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n595), .B1(new_n589), .B2(new_n593), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n564), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n589), .A2(new_n593), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(new_n594), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n589), .A2(new_n593), .A3(new_n595), .ZN(new_n601));
  INV_X1    g400(.A(new_n564), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n600), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  XOR2_X1   g402(.A(KEYINPUT95), .B(KEYINPUT21), .Z(new_n604));
  NAND2_X1  g403(.A1(new_n575), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n606));
  XOR2_X1   g405(.A(new_n605), .B(new_n606), .Z(new_n607));
  AND3_X1   g406(.A1(new_n598), .A2(new_n603), .A3(new_n607), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n607), .B1(new_n598), .B2(new_n603), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n562), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n610), .A2(KEYINPUT102), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT102), .ZN(new_n612));
  OAI211_X1 g411(.A(new_n612), .B(new_n562), .C1(new_n608), .C2(new_n609), .ZN(new_n613));
  AND3_X1   g412(.A1(new_n511), .A2(new_n611), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n586), .A2(KEYINPUT91), .ZN(new_n615));
  INV_X1    g414(.A(new_n585), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(new_n583), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT91), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND4_X1  g418(.A1(new_n615), .A2(new_n619), .A3(new_n549), .A4(new_n551), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n617), .A2(new_n546), .ZN(new_n621));
  NAND2_X1  g420(.A1(G229gat), .A2(G233gat), .ZN(new_n622));
  NAND4_X1  g421(.A1(new_n620), .A2(KEYINPUT18), .A3(new_n621), .A4(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n617), .B(new_n546), .ZN(new_n624));
  XOR2_X1   g423(.A(new_n622), .B(KEYINPUT13), .Z(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  AND2_X1   g425(.A1(new_n623), .A2(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(KEYINPUT11), .B(G169gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(G197gat), .ZN(new_n629));
  XOR2_X1   g428(.A(G113gat), .B(G141gat), .Z(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n631), .B(KEYINPUT12), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n620), .A2(new_n621), .A3(new_n622), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT18), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n627), .A2(new_n632), .A3(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT92), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n633), .A2(KEYINPUT92), .A3(new_n634), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n638), .A2(new_n627), .A3(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT93), .ZN(new_n641));
  INV_X1    g440(.A(new_n632), .ZN(new_n642));
  AND3_X1   g441(.A1(new_n640), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n641), .B1(new_n640), .B2(new_n642), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n636), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n534), .A2(new_n575), .A3(new_n535), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT10), .ZN(new_n648));
  NAND4_X1  g447(.A1(new_n530), .A2(new_n574), .A3(new_n570), .A4(new_n533), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n647), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n536), .A2(KEYINPUT10), .A3(new_n576), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(G230gat), .A2(G233gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(KEYINPUT104), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n647), .A2(new_n649), .ZN(new_n656));
  INV_X1    g455(.A(new_n653), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(G176gat), .B(G204gat), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(G148gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(KEYINPUT103), .ZN(new_n662));
  INV_X1    g461(.A(G120gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n662), .B(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n659), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n652), .A2(new_n653), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n667), .A2(new_n658), .A3(new_n664), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n646), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n614), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n428), .A2(new_n429), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g472(.A(KEYINPUT105), .B(G1gat), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n673), .B(new_n674), .ZN(G1324gat));
  NOR2_X1   g474(.A1(new_n671), .A2(new_n490), .ZN(new_n676));
  NAND2_X1  g475(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n677));
  OR2_X1    g476(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n676), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT42), .ZN(new_n680));
  OR2_X1    g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n679), .A2(new_n680), .ZN(new_n682));
  INV_X1    g481(.A(G8gat), .ZN(new_n683));
  OAI211_X1 g482(.A(new_n681), .B(new_n682), .C1(new_n683), .C2(new_n676), .ZN(G1325gat));
  INV_X1    g483(.A(new_n671), .ZN(new_n685));
  AOI21_X1  g484(.A(G15gat), .B1(new_n685), .B2(new_n469), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n473), .A2(new_n476), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n688), .A2(G15gat), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(KEYINPUT106), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n686), .B1(new_n685), .B2(new_n690), .ZN(G1326gat));
  NOR2_X1   g490(.A1(new_n671), .A2(new_n461), .ZN(new_n692));
  XOR2_X1   g491(.A(KEYINPUT43), .B(G22gat), .Z(new_n693));
  XNOR2_X1  g492(.A(new_n692), .B(new_n693), .ZN(G1327gat));
  INV_X1    g493(.A(new_n562), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n511), .A2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(new_n696), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n608), .A2(new_n609), .ZN(new_n698));
  AND2_X1   g497(.A1(new_n698), .A2(new_n670), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  NOR3_X1   g499(.A1(new_n700), .A2(G29gat), .A3(new_n672), .ZN(new_n701));
  XOR2_X1   g500(.A(new_n701), .B(KEYINPUT45), .Z(new_n702));
  AOI22_X1  g501(.A1(new_n465), .A2(new_n471), .B1(new_n477), .B2(new_n509), .ZN(new_n703));
  OAI21_X1  g502(.A(KEYINPUT44), .B1(new_n703), .B2(new_n562), .ZN(new_n704));
  AND3_X1   g503(.A1(new_n558), .A2(KEYINPUT107), .A3(new_n561), .ZN(new_n705));
  AOI21_X1  g504(.A(KEYINPUT107), .B1(new_n558), .B2(new_n561), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n707), .A2(KEYINPUT44), .ZN(new_n708));
  AOI211_X1 g507(.A(KEYINPUT35), .B(new_n394), .C1(new_n466), .C2(new_n468), .ZN(new_n709));
  AOI22_X1  g508(.A1(KEYINPUT35), .A2(new_n464), .B1(new_n709), .B2(new_n456), .ZN(new_n710));
  INV_X1    g509(.A(new_n474), .ZN(new_n711));
  AND3_X1   g510(.A1(new_n687), .A2(new_n711), .A3(new_n509), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n708), .B1(new_n710), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n704), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(new_n699), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n715), .A2(new_n672), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(KEYINPUT108), .ZN(new_n717));
  INV_X1    g516(.A(G29gat), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n702), .B1(new_n717), .B2(new_n718), .ZN(G1328gat));
  NOR3_X1   g518(.A1(new_n700), .A2(G36gat), .A3(new_n490), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(KEYINPUT46), .ZN(new_n721));
  OAI21_X1  g520(.A(G36gat), .B1(new_n715), .B2(new_n490), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(G1329gat));
  INV_X1    g522(.A(G43gat), .ZN(new_n724));
  INV_X1    g523(.A(new_n469), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n724), .B1(new_n700), .B2(new_n725), .ZN(new_n726));
  NAND4_X1  g525(.A1(new_n714), .A2(G43gat), .A3(new_n688), .A4(new_n699), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT109), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n728), .B(new_n729), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(KEYINPUT47), .ZN(G1330gat));
  NOR3_X1   g530(.A1(new_n715), .A2(new_n382), .A3(new_n461), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n700), .B(KEYINPUT110), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(new_n394), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n732), .B1(new_n734), .B2(new_n382), .ZN(new_n735));
  XOR2_X1   g534(.A(new_n735), .B(KEYINPUT48), .Z(G1331gat));
  INV_X1    g535(.A(new_n669), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n737), .A2(new_n645), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n614), .A2(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(new_n672), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g542(.A1(new_n739), .A2(new_n490), .ZN(new_n744));
  NOR2_X1   g543(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n745));
  AND2_X1   g544(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n744), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n747), .B1(new_n744), .B2(new_n745), .ZN(G1333gat));
  OAI21_X1  g547(.A(G71gat), .B1(new_n739), .B2(new_n687), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n740), .A2(new_n469), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n749), .B1(new_n750), .B2(G71gat), .ZN(new_n751));
  XNOR2_X1  g550(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n751), .B(new_n752), .ZN(G1334gat));
  NOR2_X1   g552(.A1(new_n739), .A2(new_n461), .ZN(new_n754));
  XNOR2_X1  g553(.A(KEYINPUT112), .B(G78gat), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n754), .B(new_n755), .ZN(G1335gat));
  NAND2_X1  g555(.A1(new_n698), .A2(new_n646), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n757), .A2(new_n737), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n714), .A2(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(G85gat), .ZN(new_n760));
  NOR3_X1   g559(.A1(new_n759), .A2(new_n760), .A3(new_n672), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT51), .ZN(new_n762));
  INV_X1    g561(.A(new_n757), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n697), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  OAI21_X1  g563(.A(KEYINPUT51), .B1(new_n696), .B2(new_n757), .ZN(new_n765));
  AND3_X1   g564(.A1(new_n764), .A2(new_n669), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(new_n741), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n761), .B1(new_n767), .B2(new_n760), .ZN(G1336gat));
  NOR2_X1   g567(.A1(new_n490), .A2(G92gat), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n764), .A2(new_n765), .A3(new_n669), .A4(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT52), .ZN(new_n771));
  INV_X1    g570(.A(G92gat), .ZN(new_n772));
  INV_X1    g571(.A(new_n758), .ZN(new_n773));
  AOI211_X1 g572(.A(new_n490), .B(new_n773), .C1(new_n704), .C2(new_n713), .ZN(new_n774));
  OAI211_X1 g573(.A(new_n770), .B(new_n771), .C1(new_n772), .C2(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT113), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n776), .B1(new_n774), .B2(new_n772), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n714), .A2(new_n491), .A3(new_n758), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n778), .A2(KEYINPUT113), .A3(G92gat), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n777), .A2(new_n770), .A3(new_n779), .ZN(new_n780));
  AND3_X1   g579(.A1(new_n780), .A2(KEYINPUT114), .A3(KEYINPUT52), .ZN(new_n781));
  AOI21_X1  g580(.A(KEYINPUT114), .B1(new_n780), .B2(KEYINPUT52), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n775), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(KEYINPUT115), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT115), .ZN(new_n785));
  OAI211_X1 g584(.A(new_n785), .B(new_n775), .C1(new_n781), .C2(new_n782), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n784), .A2(new_n786), .ZN(G1337gat));
  NAND3_X1  g586(.A1(new_n766), .A2(new_n519), .A3(new_n469), .ZN(new_n788));
  OAI21_X1  g587(.A(G99gat), .B1(new_n759), .B2(new_n687), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(G1338gat));
  OAI22_X1  g589(.A1(new_n759), .A2(new_n461), .B1(KEYINPUT116), .B2(G106gat), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n791), .B1(KEYINPUT116), .B2(G106gat), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n461), .A2(G106gat), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n792), .B1(new_n766), .B2(new_n793), .ZN(new_n794));
  XOR2_X1   g593(.A(new_n794), .B(KEYINPUT53), .Z(G1339gat));
  INV_X1    g594(.A(new_n698), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT55), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n652), .A2(new_n654), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT54), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n657), .B1(new_n650), .B2(new_n651), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n798), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n652), .A2(new_n799), .A3(new_n654), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(new_n665), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n797), .B1(new_n801), .B2(new_n803), .ZN(new_n804));
  OAI211_X1 g603(.A(new_n667), .B(KEYINPUT54), .C1(new_n654), .C2(new_n652), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n805), .A2(KEYINPUT55), .A3(new_n665), .A4(new_n802), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n804), .A2(new_n645), .A3(new_n806), .A4(new_n668), .ZN(new_n807));
  INV_X1    g606(.A(new_n636), .ZN(new_n808));
  AND2_X1   g607(.A1(new_n620), .A2(new_n621), .ZN(new_n809));
  OAI22_X1  g608(.A1(new_n809), .A2(new_n622), .B1(new_n624), .B2(new_n625), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n808), .B1(new_n631), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n669), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n807), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(KEYINPUT117), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT117), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n807), .A2(new_n815), .A3(new_n812), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n814), .A2(new_n707), .A3(new_n816), .ZN(new_n817));
  NAND4_X1  g616(.A1(new_n804), .A2(new_n806), .A3(new_n668), .A4(new_n811), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n707), .A2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n796), .B1(new_n817), .B2(new_n820), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n611), .A2(new_n737), .A3(new_n646), .A4(new_n613), .ZN(new_n822));
  INV_X1    g621(.A(new_n822), .ZN(new_n823));
  OR2_X1    g622(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  AND3_X1   g623(.A1(new_n824), .A2(new_n395), .A3(new_n463), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n491), .A2(new_n672), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(new_n827), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n828), .A2(new_n272), .A3(new_n645), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n725), .A2(new_n394), .ZN(new_n830));
  AND2_X1   g629(.A1(new_n824), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(new_n826), .ZN(new_n832));
  INV_X1    g631(.A(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(new_n645), .ZN(new_n834));
  AND3_X1   g633(.A1(new_n834), .A2(KEYINPUT118), .A3(G113gat), .ZN(new_n835));
  AOI21_X1  g634(.A(KEYINPUT118), .B1(new_n834), .B2(G113gat), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n829), .B1(new_n835), .B2(new_n836), .ZN(G1340gat));
  NAND3_X1  g636(.A1(new_n828), .A2(new_n663), .A3(new_n669), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n663), .B1(new_n833), .B2(new_n669), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(KEYINPUT119), .ZN(new_n840));
  INV_X1    g639(.A(new_n840), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n839), .A2(KEYINPUT119), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n838), .B1(new_n841), .B2(new_n842), .ZN(G1341gat));
  INV_X1    g642(.A(G127gat), .ZN(new_n844));
  NOR3_X1   g643(.A1(new_n832), .A2(new_n844), .A3(new_n698), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n828), .A2(new_n796), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n845), .B1(new_n846), .B2(new_n844), .ZN(G1342gat));
  NAND2_X1  g646(.A1(new_n695), .A2(new_n490), .ZN(new_n848));
  NOR3_X1   g647(.A1(new_n848), .A2(G134gat), .A3(new_n672), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n825), .A2(new_n849), .ZN(new_n850));
  XOR2_X1   g649(.A(new_n850), .B(KEYINPUT56), .Z(new_n851));
  OAI21_X1  g650(.A(G134gat), .B1(new_n832), .B2(new_n562), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(G1343gat));
  NOR2_X1   g652(.A1(new_n317), .A2(new_n318), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n687), .A2(new_n826), .ZN(new_n855));
  INV_X1    g654(.A(new_n855), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n394), .B1(new_n821), .B2(new_n823), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT57), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n695), .B1(new_n807), .B2(new_n812), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n698), .B1(new_n861), .B2(new_n819), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n858), .B1(new_n862), .B2(new_n822), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(new_n394), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(KEYINPUT120), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT120), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n863), .A2(new_n866), .A3(new_n394), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n856), .B1(new_n860), .B2(new_n868), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n854), .B1(new_n869), .B2(new_n646), .ZN(new_n870));
  INV_X1    g669(.A(new_n857), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(new_n856), .ZN(new_n872));
  INV_X1    g671(.A(new_n872), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n873), .A2(new_n320), .A3(new_n645), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n870), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g674(.A(new_n875), .B(KEYINPUT58), .ZN(G1344gat));
  INV_X1    g675(.A(KEYINPUT59), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n857), .A2(KEYINPUT57), .ZN(new_n878));
  INV_X1    g677(.A(new_n861), .ZN(new_n879));
  OR2_X1    g678(.A1(new_n818), .A2(new_n562), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n796), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  OAI211_X1 g680(.A(new_n858), .B(new_n394), .C1(new_n823), .C2(new_n881), .ZN(new_n882));
  NAND4_X1  g681(.A1(new_n878), .A2(new_n669), .A3(new_n856), .A4(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n877), .B1(new_n883), .B2(G148gat), .ZN(new_n884));
  AND3_X1   g683(.A1(new_n863), .A2(new_n866), .A3(new_n394), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n866), .B1(new_n863), .B2(new_n394), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n855), .B1(new_n887), .B2(new_n859), .ZN(new_n888));
  AOI21_X1  g687(.A(KEYINPUT59), .B1(new_n888), .B2(new_n669), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n884), .B1(new_n889), .B2(G148gat), .ZN(new_n890));
  NOR3_X1   g689(.A1(new_n872), .A2(G148gat), .A3(new_n737), .ZN(new_n891));
  OAI21_X1  g690(.A(KEYINPUT121), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT121), .ZN(new_n893));
  INV_X1    g692(.A(new_n891), .ZN(new_n894));
  AOI211_X1 g693(.A(KEYINPUT59), .B(new_n326), .C1(new_n888), .C2(new_n669), .ZN(new_n895));
  OAI211_X1 g694(.A(new_n893), .B(new_n894), .C1(new_n895), .C2(new_n884), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n892), .A2(new_n896), .ZN(G1345gat));
  AOI21_X1  g696(.A(G155gat), .B1(new_n873), .B2(new_n796), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n869), .A2(new_n698), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n898), .B1(new_n899), .B2(G155gat), .ZN(G1346gat));
  OAI21_X1  g699(.A(G162gat), .B1(new_n869), .B2(new_n707), .ZN(new_n901));
  NOR3_X1   g700(.A1(new_n848), .A2(G162gat), .A3(new_n672), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n871), .A2(new_n687), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n901), .A2(new_n903), .ZN(G1347gat));
  NOR2_X1   g703(.A1(new_n741), .A2(new_n490), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n825), .A2(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(new_n906), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n907), .A2(new_n259), .A3(new_n645), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n824), .A2(new_n830), .A3(new_n905), .ZN(new_n909));
  XNOR2_X1  g708(.A(new_n909), .B(KEYINPUT122), .ZN(new_n910));
  AND2_X1   g709(.A1(new_n910), .A2(new_n645), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n908), .B1(new_n911), .B2(new_n259), .ZN(G1348gat));
  AOI21_X1  g711(.A(G176gat), .B1(new_n907), .B2(new_n669), .ZN(new_n913));
  NOR3_X1   g712(.A1(new_n737), .A2(new_n260), .A3(new_n261), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n913), .B1(new_n910), .B2(new_n914), .ZN(G1349gat));
  NAND3_X1  g714(.A1(new_n831), .A2(KEYINPUT122), .A3(new_n905), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT122), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n909), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n916), .A2(new_n796), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n919), .A2(G183gat), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n907), .A2(new_n213), .A3(new_n796), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(KEYINPUT60), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT60), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n920), .A2(new_n924), .A3(new_n921), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n923), .A2(new_n925), .ZN(G1350gat));
  INV_X1    g725(.A(new_n707), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n907), .A2(new_n214), .A3(new_n927), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT61), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n910), .A2(new_n695), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n929), .B1(new_n930), .B2(G190gat), .ZN(new_n931));
  AOI211_X1 g730(.A(KEYINPUT61), .B(new_n214), .C1(new_n910), .C2(new_n695), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n928), .B1(new_n931), .B2(new_n932), .ZN(G1351gat));
  NAND2_X1  g732(.A1(new_n687), .A2(new_n905), .ZN(new_n934));
  OR2_X1    g733(.A1(new_n857), .A2(new_n934), .ZN(new_n935));
  XOR2_X1   g734(.A(new_n935), .B(KEYINPUT123), .Z(new_n936));
  XOR2_X1   g735(.A(KEYINPUT124), .B(G197gat), .Z(new_n937));
  INV_X1    g736(.A(new_n937), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n936), .A2(new_n645), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n878), .A2(new_n882), .ZN(new_n940));
  NOR3_X1   g739(.A1(new_n940), .A2(new_n646), .A3(new_n934), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n939), .B1(new_n941), .B2(new_n938), .ZN(G1352gat));
  NOR3_X1   g741(.A1(new_n935), .A2(G204gat), .A3(new_n737), .ZN(new_n943));
  XNOR2_X1  g742(.A(KEYINPUT125), .B(KEYINPUT62), .ZN(new_n944));
  XNOR2_X1  g743(.A(new_n943), .B(new_n944), .ZN(new_n945));
  INV_X1    g744(.A(G204gat), .ZN(new_n946));
  NOR3_X1   g745(.A1(new_n940), .A2(new_n737), .A3(new_n934), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n945), .B1(new_n946), .B2(new_n947), .ZN(G1353gat));
  NOR2_X1   g747(.A1(new_n940), .A2(new_n934), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n949), .A2(new_n796), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(G211gat), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n951), .A2(KEYINPUT126), .A3(KEYINPUT63), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n936), .A2(new_n353), .A3(new_n796), .ZN(new_n953));
  NAND2_X1  g752(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n954));
  OR2_X1    g753(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n955));
  NAND4_X1  g754(.A1(new_n950), .A2(G211gat), .A3(new_n954), .A4(new_n955), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n952), .A2(new_n953), .A3(new_n956), .ZN(G1354gat));
  AOI21_X1  g756(.A(G218gat), .B1(new_n936), .B2(new_n927), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n695), .A2(G218gat), .ZN(new_n959));
  XNOR2_X1  g758(.A(new_n959), .B(KEYINPUT127), .ZN(new_n960));
  AOI21_X1  g759(.A(new_n958), .B1(new_n949), .B2(new_n960), .ZN(G1355gat));
endmodule


