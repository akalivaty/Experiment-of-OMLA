//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 0 1 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 0 1 1 0 0 1 1 1 0 1 0 1 0 1 1 1 1 1 1 1 1 1 1 1 1 1 0 0 1 0 1 1 0 0 1 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n649, new_n650, new_n651, new_n652,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n684, new_n685, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n720, new_n721,
    new_n722, new_n724, new_n725, new_n726, new_n728, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n813,
    new_n814, new_n816, new_n817, new_n818, new_n819, new_n820, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n870, new_n871, new_n872, new_n874, new_n875,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n886, new_n887, new_n888, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n939,
    new_n940, new_n941, new_n942, new_n943;
  XNOR2_X1  g000(.A(G197gat), .B(G204gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT71), .B(KEYINPUT22), .ZN(new_n203));
  INV_X1    g002(.A(G211gat), .ZN(new_n204));
  INV_X1    g003(.A(G218gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n202), .B1(new_n203), .B2(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G211gat), .B(G218gat), .ZN(new_n208));
  XNOR2_X1  g007(.A(new_n207), .B(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT3), .ZN(new_n210));
  AND2_X1   g009(.A1(G155gat), .A2(G162gat), .ZN(new_n211));
  NOR2_X1   g010(.A1(G155gat), .A2(G162gat), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(G141gat), .B(G148gat), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n213), .B1(new_n214), .B2(KEYINPUT2), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT2), .ZN(new_n216));
  AND2_X1   g015(.A1(KEYINPUT73), .A2(G155gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(KEYINPUT73), .A2(G155gat), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n216), .B1(new_n219), .B2(G162gat), .ZN(new_n220));
  INV_X1    g019(.A(G141gat), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n221), .A2(G148gat), .ZN(new_n222));
  INV_X1    g021(.A(G148gat), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n223), .A2(G141gat), .ZN(new_n224));
  OAI22_X1  g023(.A1(new_n222), .A2(new_n224), .B1(new_n212), .B2(new_n211), .ZN(new_n225));
  OAI211_X1 g024(.A(new_n210), .B(new_n215), .C1(new_n220), .C2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT75), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  XNOR2_X1  g027(.A(KEYINPUT73), .B(G155gat), .ZN(new_n229));
  INV_X1    g028(.A(G162gat), .ZN(new_n230));
  OAI21_X1  g029(.A(KEYINPUT2), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n213), .A2(new_n214), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND4_X1  g032(.A1(new_n233), .A2(KEYINPUT75), .A3(new_n210), .A4(new_n215), .ZN(new_n234));
  AND2_X1   g033(.A1(new_n228), .A2(new_n234), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n209), .B1(new_n235), .B2(KEYINPUT29), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n210), .B1(new_n209), .B2(KEYINPUT29), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n215), .B1(new_n220), .B2(new_n225), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n236), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(G228gat), .A2(G233gat), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n241), .B(G22gat), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n240), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g042(.A(G78gat), .B(G106gat), .ZN(new_n244));
  XNOR2_X1  g043(.A(KEYINPUT31), .B(G50gat), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n246), .B(KEYINPUT78), .ZN(new_n247));
  OR2_X1    g046(.A1(new_n243), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n243), .A2(KEYINPUT78), .A3(new_n246), .ZN(new_n249));
  AND2_X1   g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(G225gat), .A2(G233gat), .ZN(new_n251));
  XOR2_X1   g050(.A(G127gat), .B(G134gat), .Z(new_n252));
  XNOR2_X1  g051(.A(G113gat), .B(G120gat), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n252), .B1(KEYINPUT1), .B2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(G120gat), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(G113gat), .ZN(new_n256));
  INV_X1    g055(.A(G113gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(G120gat), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  XNOR2_X1  g058(.A(G127gat), .B(G134gat), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT1), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n259), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n254), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n216), .B1(new_n222), .B2(new_n224), .ZN(new_n265));
  AOI22_X1  g064(.A1(new_n231), .A2(new_n232), .B1(new_n265), .B2(new_n213), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n264), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  OAI21_X1  g067(.A(KEYINPUT4), .B1(new_n238), .B2(new_n263), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT74), .ZN(new_n271));
  INV_X1    g070(.A(new_n262), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n260), .B1(new_n261), .B2(new_n259), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n271), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n254), .A2(KEYINPUT74), .A3(new_n262), .ZN(new_n275));
  OAI211_X1 g074(.A(new_n274), .B(new_n275), .C1(new_n210), .C2(new_n266), .ZN(new_n276));
  OAI211_X1 g075(.A(new_n251), .B(new_n270), .C1(new_n235), .C2(new_n276), .ZN(new_n277));
  XOR2_X1   g076(.A(KEYINPUT76), .B(KEYINPUT5), .Z(new_n278));
  NAND3_X1  g077(.A1(new_n274), .A2(new_n238), .A3(new_n275), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n264), .A2(new_n266), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(new_n251), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n278), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n277), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n228), .A2(new_n234), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n238), .A2(KEYINPUT3), .ZN(new_n286));
  NAND4_X1  g085(.A1(new_n285), .A2(new_n275), .A3(new_n274), .A4(new_n286), .ZN(new_n287));
  NAND4_X1  g086(.A1(new_n287), .A2(new_n251), .A3(new_n270), .A4(new_n278), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n284), .A2(new_n288), .ZN(new_n289));
  XNOR2_X1  g088(.A(G1gat), .B(G29gat), .ZN(new_n290));
  INV_X1    g089(.A(G85gat), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n290), .B(new_n291), .ZN(new_n292));
  XNOR2_X1  g091(.A(KEYINPUT0), .B(G57gat), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n292), .B(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  AND4_X1   g094(.A1(KEYINPUT77), .A2(new_n289), .A3(KEYINPUT6), .A4(new_n295), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n294), .B1(new_n284), .B2(new_n288), .ZN(new_n297));
  AOI21_X1  g096(.A(KEYINPUT77), .B1(new_n297), .B2(KEYINPUT6), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  AND2_X1   g098(.A1(new_n284), .A2(new_n288), .ZN(new_n300));
  AOI21_X1  g099(.A(KEYINPUT6), .B1(new_n300), .B2(new_n294), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n301), .B1(new_n294), .B2(new_n300), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n299), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT25), .ZN(new_n304));
  NAND2_X1  g103(.A1(G169gat), .A2(G176gat), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT24), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n306), .A2(G183gat), .A3(G190gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(G183gat), .A2(G190gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(KEYINPUT24), .ZN(new_n309));
  NOR2_X1   g108(.A1(G183gat), .A2(G190gat), .ZN(new_n310));
  OAI211_X1 g109(.A(new_n305), .B(new_n307), .C1(new_n309), .C2(new_n310), .ZN(new_n311));
  OAI21_X1  g110(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  NOR3_X1   g112(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n304), .B1(new_n311), .B2(new_n315), .ZN(new_n316));
  AND2_X1   g115(.A1(new_n307), .A2(new_n305), .ZN(new_n317));
  INV_X1    g116(.A(new_n310), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n318), .A2(KEYINPUT24), .A3(new_n308), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT23), .ZN(new_n320));
  INV_X1    g119(.A(G169gat), .ZN(new_n321));
  INV_X1    g120(.A(G176gat), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n320), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(new_n312), .ZN(new_n324));
  NAND4_X1  g123(.A1(new_n317), .A2(new_n319), .A3(KEYINPUT25), .A4(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n316), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(G190gat), .ZN(new_n327));
  AND2_X1   g126(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n328));
  NOR2_X1   g127(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n327), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(KEYINPUT65), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT65), .ZN(new_n332));
  OAI211_X1 g131(.A(new_n332), .B(new_n327), .C1(new_n328), .C2(new_n329), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n331), .A2(KEYINPUT28), .A3(new_n333), .ZN(new_n334));
  OAI21_X1  g133(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n335));
  AND2_X1   g134(.A1(new_n335), .A2(new_n305), .ZN(new_n336));
  OR3_X1    g135(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n337));
  AOI22_X1  g136(.A1(new_n336), .A2(new_n337), .B1(G183gat), .B2(G190gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n334), .A2(new_n338), .ZN(new_n339));
  AOI21_X1  g138(.A(KEYINPUT28), .B1(new_n331), .B2(new_n333), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n326), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(G226gat), .A2(G233gat), .ZN(new_n342));
  XNOR2_X1  g141(.A(new_n342), .B(KEYINPUT72), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n341), .A2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(new_n209), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT28), .ZN(new_n347));
  XNOR2_X1  g146(.A(KEYINPUT27), .B(G183gat), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n332), .B1(new_n348), .B2(new_n327), .ZN(new_n349));
  INV_X1    g148(.A(new_n333), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n347), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n351), .A2(new_n334), .A3(new_n338), .ZN(new_n352));
  AOI21_X1  g151(.A(KEYINPUT29), .B1(new_n352), .B2(new_n326), .ZN(new_n353));
  INV_X1    g152(.A(new_n342), .ZN(new_n354));
  OAI211_X1 g153(.A(new_n345), .B(new_n346), .C1(new_n353), .C2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT29), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n341), .A2(new_n356), .ZN(new_n357));
  AOI22_X1  g156(.A1(new_n357), .A2(new_n343), .B1(new_n341), .B2(new_n354), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n355), .B1(new_n358), .B2(new_n346), .ZN(new_n359));
  XNOR2_X1  g158(.A(G8gat), .B(G36gat), .ZN(new_n360));
  XNOR2_X1  g159(.A(G64gat), .B(G92gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n360), .B(new_n361), .ZN(new_n362));
  OR2_X1    g161(.A1(new_n359), .A2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT30), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n364), .B1(new_n359), .B2(new_n362), .ZN(new_n365));
  OR2_X1    g164(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n363), .A2(new_n365), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n250), .B1(new_n303), .B2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT80), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n289), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n284), .A2(new_n288), .A3(KEYINPUT80), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n371), .A2(new_n295), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(new_n301), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n359), .A2(new_n362), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT37), .ZN(new_n376));
  OAI211_X1 g175(.A(new_n376), .B(new_n355), .C1(new_n358), .C2(new_n346), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT38), .ZN(new_n378));
  AND3_X1   g177(.A1(new_n377), .A2(new_n378), .A3(new_n362), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n341), .A2(new_n354), .ZN(new_n380));
  OAI211_X1 g179(.A(new_n380), .B(new_n346), .C1(new_n353), .C2(new_n344), .ZN(new_n381));
  AOI22_X1  g180(.A1(new_n357), .A2(new_n342), .B1(new_n341), .B2(new_n344), .ZN(new_n382));
  OAI22_X1  g181(.A1(KEYINPUT81), .A2(new_n381), .B1(new_n382), .B2(new_n346), .ZN(new_n383));
  AND2_X1   g182(.A1(new_n381), .A2(KEYINPUT81), .ZN(new_n384));
  OAI21_X1  g183(.A(KEYINPUT37), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n375), .B1(new_n379), .B2(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n299), .A2(new_n374), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(KEYINPUT82), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT82), .ZN(new_n389));
  NAND4_X1  g188(.A1(new_n299), .A2(new_n374), .A3(new_n386), .A4(new_n389), .ZN(new_n390));
  AND2_X1   g189(.A1(new_n359), .A2(KEYINPUT37), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n377), .A2(new_n362), .ZN(new_n392));
  OAI21_X1  g191(.A(KEYINPUT38), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n388), .A2(new_n390), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n248), .A2(new_n249), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n251), .B1(new_n287), .B2(new_n270), .ZN(new_n396));
  OAI21_X1  g195(.A(KEYINPUT39), .B1(new_n281), .B2(new_n282), .ZN(new_n397));
  OR2_X1    g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT39), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n295), .B1(new_n396), .B2(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n398), .A2(KEYINPUT40), .A3(new_n400), .ZN(new_n401));
  AND4_X1   g200(.A1(new_n366), .A2(new_n401), .A3(new_n367), .A4(new_n373), .ZN(new_n402));
  AOI21_X1  g201(.A(KEYINPUT40), .B1(new_n398), .B2(new_n400), .ZN(new_n403));
  XNOR2_X1  g202(.A(new_n403), .B(KEYINPUT79), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n395), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n369), .B1(new_n394), .B2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT70), .ZN(new_n407));
  NAND2_X1  g206(.A1(G227gat), .A2(G233gat), .ZN(new_n408));
  XOR2_X1   g207(.A(new_n408), .B(KEYINPUT64), .Z(new_n409));
  OAI211_X1 g208(.A(new_n264), .B(new_n326), .C1(new_n339), .C2(new_n340), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n264), .B1(new_n352), .B2(new_n326), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n409), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(KEYINPUT32), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT33), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  XNOR2_X1  g215(.A(G15gat), .B(G99gat), .ZN(new_n417));
  INV_X1    g216(.A(G43gat), .ZN(new_n418));
  XNOR2_X1  g217(.A(new_n417), .B(new_n418), .ZN(new_n419));
  XNOR2_X1  g218(.A(KEYINPUT66), .B(G71gat), .ZN(new_n420));
  XOR2_X1   g219(.A(new_n419), .B(new_n420), .Z(new_n421));
  NAND3_X1  g220(.A1(new_n414), .A2(new_n416), .A3(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(new_n421), .ZN(new_n423));
  OAI211_X1 g222(.A(new_n413), .B(KEYINPUT32), .C1(new_n415), .C2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n341), .A2(new_n263), .ZN(new_n426));
  INV_X1    g225(.A(new_n409), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n426), .A2(new_n427), .A3(new_n410), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(KEYINPUT34), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT67), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n428), .A2(KEYINPUT67), .A3(KEYINPUT34), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT34), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n426), .A2(new_n433), .A3(new_n427), .A4(new_n410), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT68), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n411), .A2(new_n412), .ZN(new_n437));
  NAND4_X1  g236(.A1(new_n437), .A2(KEYINPUT68), .A3(new_n433), .A4(new_n427), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n431), .A2(new_n432), .A3(new_n436), .A4(new_n438), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n425), .A2(new_n439), .ZN(new_n440));
  AND3_X1   g239(.A1(new_n428), .A2(KEYINPUT67), .A3(KEYINPUT34), .ZN(new_n441));
  AOI21_X1  g240(.A(KEYINPUT67), .B1(new_n428), .B2(KEYINPUT34), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  XNOR2_X1  g242(.A(new_n434), .B(KEYINPUT68), .ZN(new_n444));
  AOI22_X1  g243(.A1(new_n443), .A2(new_n444), .B1(new_n422), .B2(new_n424), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n440), .A2(new_n445), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n407), .B1(new_n446), .B2(KEYINPUT36), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT36), .ZN(new_n448));
  OAI211_X1 g247(.A(KEYINPUT70), .B(new_n448), .C1(new_n440), .C2(new_n445), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT69), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n427), .B1(new_n426), .B2(new_n410), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n421), .B1(new_n451), .B2(KEYINPUT33), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT32), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n424), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n450), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(new_n439), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n425), .A2(new_n439), .A3(new_n450), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n459), .A2(KEYINPUT36), .A3(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n447), .A2(new_n449), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n406), .A2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n368), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n464), .A2(KEYINPUT35), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n299), .A2(new_n374), .ZN(new_n466));
  NAND4_X1  g265(.A1(new_n465), .A2(new_n446), .A3(new_n250), .A4(new_n466), .ZN(new_n467));
  AND2_X1   g266(.A1(new_n459), .A2(new_n460), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(new_n250), .ZN(new_n469));
  INV_X1    g268(.A(new_n303), .ZN(new_n470));
  NOR3_X1   g269(.A1(new_n469), .A2(new_n470), .A3(new_n464), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT35), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n467), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n463), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(G229gat), .A2(G233gat), .ZN(new_n475));
  XNOR2_X1  g274(.A(G15gat), .B(G22gat), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT16), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n476), .B1(new_n477), .B2(G1gat), .ZN(new_n478));
  NAND2_X1  g277(.A1(KEYINPUT86), .A2(G8gat), .ZN(new_n479));
  OAI211_X1 g278(.A(new_n478), .B(new_n479), .C1(G1gat), .C2(new_n476), .ZN(new_n480));
  NOR2_X1   g279(.A1(KEYINPUT86), .A2(G8gat), .ZN(new_n481));
  XOR2_X1   g280(.A(new_n480), .B(new_n481), .Z(new_n482));
  INV_X1    g281(.A(KEYINPUT14), .ZN(new_n483));
  XOR2_X1   g282(.A(KEYINPUT84), .B(G36gat), .Z(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(G29gat), .ZN(new_n485));
  OR2_X1    g284(.A1(G29gat), .A2(G36gat), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n483), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  AND2_X1   g286(.A1(new_n486), .A2(new_n483), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(G50gat), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n418), .A2(new_n490), .ZN(new_n491));
  NOR2_X1   g290(.A1(G43gat), .A2(G50gat), .ZN(new_n492));
  OAI21_X1  g291(.A(KEYINPUT15), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  XOR2_X1   g292(.A(KEYINPUT85), .B(G43gat), .Z(new_n494));
  NOR2_X1   g293(.A1(new_n494), .A2(G50gat), .ZN(new_n495));
  OR2_X1    g294(.A1(new_n491), .A2(KEYINPUT15), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n493), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n489), .A2(new_n497), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n493), .B1(new_n487), .B2(new_n488), .ZN(new_n499));
  AND2_X1   g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT17), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT87), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n482), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n482), .A2(new_n503), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n500), .B1(new_n505), .B2(new_n501), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n475), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT18), .ZN(new_n508));
  OR2_X1    g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  XNOR2_X1  g308(.A(new_n500), .B(new_n482), .ZN(new_n510));
  XOR2_X1   g309(.A(new_n475), .B(KEYINPUT13), .Z(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AND2_X1   g311(.A1(new_n509), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n507), .A2(new_n508), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT88), .ZN(new_n515));
  XNOR2_X1  g314(.A(G113gat), .B(G141gat), .ZN(new_n516));
  INV_X1    g315(.A(G197gat), .ZN(new_n517));
  XNOR2_X1  g316(.A(new_n516), .B(new_n517), .ZN(new_n518));
  XNOR2_X1  g317(.A(KEYINPUT11), .B(G169gat), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n518), .B(new_n519), .ZN(new_n520));
  XOR2_X1   g319(.A(KEYINPUT83), .B(KEYINPUT12), .Z(new_n521));
  XNOR2_X1  g320(.A(new_n520), .B(new_n521), .ZN(new_n522));
  OAI211_X1 g321(.A(new_n513), .B(new_n514), .C1(new_n515), .C2(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n509), .A2(new_n515), .A3(new_n512), .ZN(new_n524));
  INV_X1    g323(.A(new_n522), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n509), .A2(new_n512), .ZN(new_n526));
  INV_X1    g325(.A(new_n514), .ZN(new_n527));
  OAI211_X1 g326(.A(new_n524), .B(new_n525), .C1(new_n526), .C2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n523), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n474), .A2(new_n529), .ZN(new_n530));
  XOR2_X1   g329(.A(new_n530), .B(KEYINPUT89), .Z(new_n531));
  NAND3_X1  g330(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n532));
  NAND2_X1  g331(.A1(G99gat), .A2(G106gat), .ZN(new_n533));
  INV_X1    g332(.A(G92gat), .ZN(new_n534));
  AOI22_X1  g333(.A1(KEYINPUT8), .A2(new_n533), .B1(new_n291), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(KEYINPUT94), .A2(KEYINPUT7), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n536), .B1(new_n291), .B2(new_n534), .ZN(new_n537));
  NAND4_X1  g336(.A1(KEYINPUT94), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n535), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  XOR2_X1   g338(.A(G99gat), .B(G106gat), .Z(new_n540));
  OR2_X1    g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n539), .A2(new_n540), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT95), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n544), .B1(new_n502), .B2(new_n545), .ZN(new_n546));
  AOI21_X1  g345(.A(KEYINPUT17), .B1(new_n544), .B2(new_n545), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n500), .A2(new_n547), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n532), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  XOR2_X1   g348(.A(G190gat), .B(G218gat), .Z(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  AOI21_X1  g350(.A(KEYINPUT96), .B1(new_n549), .B2(new_n551), .ZN(new_n552));
  XNOR2_X1  g351(.A(G134gat), .B(G162gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n553), .B(KEYINPUT93), .ZN(new_n554));
  AOI21_X1  g353(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n554), .B(new_n555), .ZN(new_n556));
  OR3_X1    g355(.A1(new_n552), .A2(KEYINPUT97), .A3(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n549), .B(new_n550), .ZN(new_n558));
  OAI21_X1  g357(.A(KEYINPUT97), .B1(new_n552), .B2(new_n556), .ZN(new_n559));
  AND3_X1   g358(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n558), .B1(new_n557), .B2(new_n559), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(G71gat), .A2(G78gat), .ZN(new_n563));
  NOR2_X1   g362(.A1(G71gat), .A2(G78gat), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT90), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n563), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n566), .B1(new_n565), .B2(new_n564), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT9), .ZN(new_n568));
  XNOR2_X1  g367(.A(G57gat), .B(G64gat), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n567), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT91), .ZN(new_n571));
  OR2_X1    g370(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n564), .A2(KEYINPUT9), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n573), .A2(new_n563), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n569), .A2(new_n571), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n572), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  AND2_X1   g375(.A1(new_n570), .A2(new_n576), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n577), .A2(KEYINPUT21), .ZN(new_n578));
  XOR2_X1   g377(.A(G127gat), .B(G155gat), .Z(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n581));
  XNOR2_X1  g380(.A(G183gat), .B(G211gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n581), .B(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n580), .B(new_n583), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n482), .B1(KEYINPUT21), .B2(new_n577), .ZN(new_n585));
  NAND2_X1  g384(.A1(G231gat), .A2(G233gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n586), .B(KEYINPUT92), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n585), .B(new_n587), .ZN(new_n588));
  OR2_X1    g387(.A1(new_n584), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n584), .A2(new_n588), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n544), .A2(new_n577), .A3(KEYINPUT10), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n541), .A2(KEYINPUT98), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n593), .A2(new_n542), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT99), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n539), .A2(KEYINPUT98), .A3(new_n540), .ZN(new_n596));
  NAND4_X1  g395(.A1(new_n594), .A2(new_n595), .A3(new_n577), .A4(new_n596), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n544), .A2(new_n577), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n598), .A2(KEYINPUT99), .ZN(new_n599));
  AND3_X1   g398(.A1(new_n594), .A2(new_n577), .A3(new_n596), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n597), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n592), .B1(new_n601), .B2(KEYINPUT10), .ZN(new_n602));
  NAND2_X1  g401(.A1(G230gat), .A2(G233gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n603), .B(KEYINPUT101), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n601), .A2(G230gat), .A3(G233gat), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  XOR2_X1   g406(.A(G176gat), .B(G204gat), .Z(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(KEYINPUT100), .ZN(new_n609));
  XNOR2_X1  g408(.A(G120gat), .B(G148gat), .ZN(new_n610));
  XOR2_X1   g409(.A(new_n609), .B(new_n610), .Z(new_n611));
  NAND2_X1  g410(.A1(new_n607), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n602), .A2(new_n603), .ZN(new_n613));
  INV_X1    g412(.A(new_n611), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n613), .A2(new_n606), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n612), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n562), .A2(new_n591), .A3(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n531), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n621), .A2(new_n470), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n622), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g422(.A1(new_n620), .A2(new_n368), .ZN(new_n624));
  INV_X1    g423(.A(G8gat), .ZN(new_n625));
  OAI21_X1  g424(.A(KEYINPUT42), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  XOR2_X1   g425(.A(KEYINPUT16), .B(G8gat), .Z(new_n627));
  NAND2_X1  g426(.A1(new_n624), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n624), .A2(KEYINPUT42), .A3(new_n627), .ZN(new_n630));
  AND2_X1   g429(.A1(new_n630), .A2(KEYINPUT102), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n630), .A2(KEYINPUT102), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n629), .B1(new_n631), .B2(new_n632), .ZN(G1325gat));
  NAND2_X1  g432(.A1(new_n461), .A2(new_n449), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n425), .A2(new_n439), .ZN(new_n635));
  NAND4_X1  g434(.A1(new_n443), .A2(new_n444), .A3(new_n424), .A4(new_n422), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  AOI21_X1  g436(.A(KEYINPUT70), .B1(new_n637), .B2(new_n448), .ZN(new_n638));
  OAI21_X1  g437(.A(KEYINPUT103), .B1(new_n634), .B2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT103), .ZN(new_n640));
  NAND4_X1  g439(.A1(new_n447), .A2(new_n640), .A3(new_n449), .A4(new_n461), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n621), .A2(G15gat), .A3(new_n643), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n620), .A2(new_n637), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n644), .B1(new_n645), .B2(G15gat), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT104), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(G1326gat));
  OR3_X1    g447(.A1(new_n620), .A2(G22gat), .A3(new_n250), .ZN(new_n649));
  OAI21_X1  g448(.A(G22gat), .B1(new_n620), .B2(new_n250), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(KEYINPUT105), .B(KEYINPUT43), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n651), .B(new_n652), .ZN(G1327gat));
  INV_X1    g452(.A(new_n562), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n616), .A2(new_n591), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  XOR2_X1   g455(.A(new_n656), .B(KEYINPUT106), .Z(new_n657));
  AND2_X1   g456(.A1(new_n531), .A2(new_n657), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n303), .A2(G29gat), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n660), .A2(KEYINPUT107), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT107), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n658), .A2(new_n662), .A3(new_n659), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT45), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n661), .A2(KEYINPUT45), .A3(new_n663), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT108), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT109), .ZN(new_n669));
  AND3_X1   g468(.A1(new_n406), .A2(new_n669), .A3(new_n642), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n669), .B1(new_n406), .B2(new_n642), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n473), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT44), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n672), .A2(new_n673), .A3(new_n654), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n474), .A2(new_n654), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(KEYINPUT44), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n668), .B1(new_n674), .B2(new_n676), .ZN(new_n677));
  AOI21_X1  g476(.A(KEYINPUT108), .B1(new_n675), .B2(KEYINPUT44), .ZN(new_n678));
  OR2_X1    g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  AND2_X1   g478(.A1(new_n529), .A2(new_n655), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  OAI21_X1  g480(.A(G29gat), .B1(new_n681), .B2(new_n303), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n666), .A2(new_n667), .A3(new_n682), .ZN(G1328gat));
  INV_X1    g482(.A(new_n484), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n658), .A2(new_n464), .A3(new_n684), .ZN(new_n685));
  XOR2_X1   g484(.A(new_n685), .B(KEYINPUT46), .Z(new_n686));
  OAI21_X1  g485(.A(new_n484), .B1(new_n681), .B2(new_n368), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(G1329gat));
  NAND3_X1  g487(.A1(new_n531), .A2(new_n446), .A3(new_n657), .ZN(new_n689));
  INV_X1    g488(.A(new_n494), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT110), .ZN(new_n691));
  AOI22_X1  g490(.A1(new_n689), .A2(new_n690), .B1(new_n691), .B2(KEYINPUT47), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n643), .A2(new_n494), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n692), .B1(new_n681), .B2(new_n693), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n691), .A2(KEYINPUT47), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT111), .ZN(new_n696));
  INV_X1    g495(.A(new_n696), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n694), .B(new_n697), .ZN(G1330gat));
  OAI21_X1  g497(.A(G50gat), .B1(new_n681), .B2(new_n250), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n395), .A2(new_n490), .ZN(new_n700));
  XOR2_X1   g499(.A(new_n700), .B(KEYINPUT112), .Z(new_n701));
  NAND2_X1  g500(.A1(new_n658), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n699), .A2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT48), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n699), .A2(KEYINPUT48), .A3(new_n702), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(G1331gat));
  AND2_X1   g506(.A1(new_n523), .A2(new_n528), .ZN(new_n708));
  NAND4_X1  g507(.A1(new_n562), .A2(new_n708), .A3(new_n591), .A4(new_n616), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n394), .A2(new_n405), .ZN(new_n710));
  INV_X1    g509(.A(new_n369), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n642), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(KEYINPUT109), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n406), .A2(new_n669), .A3(new_n642), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n709), .B1(new_n715), .B2(new_n473), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n303), .B(KEYINPUT113), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g518(.A1(new_n716), .A2(new_n464), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n720), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n721));
  XOR2_X1   g520(.A(KEYINPUT49), .B(G64gat), .Z(new_n722));
  OAI21_X1  g521(.A(new_n721), .B1(new_n720), .B2(new_n722), .ZN(G1333gat));
  AOI21_X1  g522(.A(G71gat), .B1(new_n716), .B2(new_n446), .ZN(new_n724));
  AND2_X1   g523(.A1(new_n643), .A2(G71gat), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n724), .B1(new_n716), .B2(new_n725), .ZN(new_n726));
  XOR2_X1   g525(.A(new_n726), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g526(.A1(new_n716), .A2(new_n395), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g528(.A1(new_n529), .A2(new_n591), .A3(new_n617), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n679), .A2(new_n470), .A3(new_n730), .ZN(new_n731));
  AND2_X1   g530(.A1(new_n731), .A2(KEYINPUT114), .ZN(new_n732));
  OAI21_X1  g531(.A(G85gat), .B1(new_n731), .B2(KEYINPUT114), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n562), .B1(new_n715), .B2(new_n473), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n529), .A2(new_n591), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n734), .A2(KEYINPUT51), .A3(new_n735), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n672), .A2(new_n654), .A3(new_n735), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT51), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n736), .A2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(new_n740), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n470), .A2(new_n291), .A3(new_n616), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(KEYINPUT115), .ZN(new_n743));
  OAI22_X1  g542(.A1(new_n732), .A2(new_n733), .B1(new_n741), .B2(new_n743), .ZN(G1336gat));
  NAND3_X1  g543(.A1(new_n679), .A2(new_n464), .A3(new_n730), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(G92gat), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n740), .A2(new_n616), .ZN(new_n747));
  INV_X1    g546(.A(new_n747), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n748), .A2(new_n534), .A3(new_n464), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n746), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(KEYINPUT52), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT52), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n746), .A2(new_n752), .A3(new_n749), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n751), .A2(new_n753), .ZN(G1337gat));
  INV_X1    g553(.A(G99gat), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n748), .A2(new_n755), .A3(new_n446), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n679), .A2(new_n643), .A3(new_n730), .ZN(new_n757));
  INV_X1    g556(.A(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n756), .B1(new_n758), .B2(new_n755), .ZN(G1338gat));
  OAI211_X1 g558(.A(new_n395), .B(new_n730), .C1(new_n677), .C2(new_n678), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(G106gat), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT53), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n250), .A2(G106gat), .ZN(new_n763));
  AOI21_X1  g562(.A(KEYINPUT51), .B1(new_n734), .B2(new_n735), .ZN(new_n764));
  AND4_X1   g563(.A1(KEYINPUT51), .A2(new_n672), .A3(new_n654), .A4(new_n735), .ZN(new_n765));
  OAI211_X1 g564(.A(new_n616), .B(new_n763), .C1(new_n764), .C2(new_n765), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n761), .A2(new_n762), .A3(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(KEYINPUT116), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT116), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n740), .A2(new_n769), .A3(new_n616), .A4(new_n763), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n761), .A2(new_n768), .A3(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT117), .ZN(new_n772));
  AND3_X1   g571(.A1(new_n771), .A2(new_n772), .A3(KEYINPUT53), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n772), .B1(new_n771), .B2(KEYINPUT53), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n767), .B1(new_n773), .B2(new_n774), .ZN(G1339gat));
  INV_X1    g574(.A(KEYINPUT55), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n613), .A2(KEYINPUT54), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n602), .A2(new_n604), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n611), .B1(new_n605), .B2(KEYINPUT54), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n776), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(new_n780), .ZN(new_n782));
  OAI211_X1 g581(.A(new_n613), .B(KEYINPUT54), .C1(new_n604), .C2(new_n602), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n782), .A2(KEYINPUT55), .A3(new_n783), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n781), .A2(new_n784), .A3(new_n615), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT118), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND4_X1  g586(.A1(new_n781), .A2(new_n784), .A3(KEYINPUT118), .A4(new_n615), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n708), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n513), .A2(new_n514), .A3(new_n522), .ZN(new_n790));
  NOR3_X1   g589(.A1(new_n504), .A2(new_n475), .A3(new_n506), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n510), .A2(new_n511), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n520), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  AND2_X1   g592(.A1(new_n790), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(new_n616), .ZN(new_n795));
  INV_X1    g594(.A(new_n795), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n562), .B1(new_n789), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n787), .A2(new_n788), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n798), .A2(new_n654), .A3(new_n794), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n591), .B1(new_n797), .B2(new_n799), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n618), .A2(new_n529), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NOR3_X1   g601(.A1(new_n802), .A2(new_n637), .A3(new_n395), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n464), .A2(new_n303), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  OAI21_X1  g604(.A(G113gat), .B1(new_n805), .B2(new_n708), .ZN(new_n806));
  OR2_X1    g605(.A1(new_n800), .A2(new_n801), .ZN(new_n807));
  AND2_X1   g606(.A1(new_n807), .A2(new_n717), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n469), .A2(new_n464), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n529), .A2(new_n257), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n806), .B1(new_n810), .B2(new_n811), .ZN(G1340gat));
  OAI21_X1  g611(.A(G120gat), .B1(new_n805), .B2(new_n617), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n616), .A2(new_n255), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n813), .B1(new_n810), .B2(new_n814), .ZN(G1341gat));
  INV_X1    g614(.A(new_n810), .ZN(new_n816));
  AOI21_X1  g615(.A(G127gat), .B1(new_n816), .B2(new_n591), .ZN(new_n817));
  NAND4_X1  g616(.A1(new_n803), .A2(G127gat), .A3(new_n591), .A4(new_n804), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n818), .A2(KEYINPUT119), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n818), .A2(KEYINPUT119), .ZN(new_n820));
  NOR3_X1   g619(.A1(new_n817), .A2(new_n819), .A3(new_n820), .ZN(G1342gat));
  INV_X1    g620(.A(G134gat), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n816), .A2(new_n822), .A3(new_n654), .ZN(new_n823));
  OR2_X1    g622(.A1(new_n823), .A2(KEYINPUT56), .ZN(new_n824));
  OAI21_X1  g623(.A(G134gat), .B1(new_n805), .B2(new_n562), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n823), .A2(KEYINPUT56), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n824), .A2(new_n825), .A3(new_n826), .ZN(G1343gat));
  NAND2_X1  g626(.A1(new_n642), .A2(new_n804), .ZN(new_n828));
  INV_X1    g627(.A(new_n828), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n395), .B1(new_n800), .B2(new_n801), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n829), .B1(new_n830), .B2(KEYINPUT57), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT120), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n785), .A2(new_n832), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n781), .A2(new_n784), .A3(KEYINPUT120), .A4(new_n615), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n833), .A2(new_n529), .A3(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT121), .ZN(new_n836));
  AND3_X1   g635(.A1(new_n835), .A2(new_n836), .A3(new_n795), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n836), .B1(new_n835), .B2(new_n795), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n562), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n591), .B1(new_n839), .B2(new_n799), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n395), .B1(new_n840), .B2(new_n801), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n831), .B1(KEYINPUT57), .B2(new_n841), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n221), .B1(new_n842), .B2(new_n529), .ZN(new_n843));
  INV_X1    g642(.A(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT58), .ZN(new_n845));
  NOR3_X1   g644(.A1(new_n643), .A2(new_n464), .A3(new_n250), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n808), .A2(new_n846), .ZN(new_n847));
  NOR3_X1   g646(.A1(new_n847), .A2(G141gat), .A3(new_n708), .ZN(new_n848));
  INV_X1    g647(.A(new_n848), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n844), .A2(new_n845), .A3(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(KEYINPUT58), .B1(new_n843), .B2(new_n848), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(G1344gat));
  INV_X1    g651(.A(new_n847), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n853), .A2(new_n223), .A3(new_n616), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT59), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n250), .A2(KEYINPUT57), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT123), .ZN(new_n857));
  OR3_X1    g656(.A1(new_n562), .A2(new_n857), .A3(new_n785), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n857), .B1(new_n562), .B2(new_n785), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n858), .A2(new_n794), .A3(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n591), .B1(new_n839), .B2(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n856), .B1(new_n861), .B2(new_n801), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n830), .A2(KEYINPUT57), .ZN(new_n863));
  AND3_X1   g662(.A1(new_n862), .A2(new_n616), .A3(new_n863), .ZN(new_n864));
  XOR2_X1   g663(.A(new_n828), .B(KEYINPUT122), .Z(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n855), .B1(new_n866), .B2(G148gat), .ZN(new_n867));
  AOI211_X1 g666(.A(KEYINPUT59), .B(new_n223), .C1(new_n842), .C2(new_n616), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n854), .B1(new_n867), .B2(new_n868), .ZN(G1345gat));
  AOI21_X1  g668(.A(new_n219), .B1(new_n853), .B2(new_n591), .ZN(new_n870));
  INV_X1    g669(.A(new_n591), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n871), .A2(new_n229), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n870), .B1(new_n842), .B2(new_n872), .ZN(G1346gat));
  AOI21_X1  g672(.A(new_n230), .B1(new_n842), .B2(new_n654), .ZN(new_n874));
  NOR3_X1   g673(.A1(new_n847), .A2(G162gat), .A3(new_n562), .ZN(new_n875));
  OR2_X1    g674(.A1(new_n874), .A2(new_n875), .ZN(G1347gat));
  OR2_X1    g675(.A1(new_n717), .A2(new_n368), .ZN(new_n877));
  XNOR2_X1  g676(.A(new_n877), .B(KEYINPUT124), .ZN(new_n878));
  INV_X1    g677(.A(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n803), .A2(new_n879), .ZN(new_n880));
  OAI21_X1  g679(.A(G169gat), .B1(new_n880), .B2(new_n708), .ZN(new_n881));
  NOR3_X1   g680(.A1(new_n802), .A2(new_n470), .A3(new_n368), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n882), .A2(new_n468), .A3(new_n250), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n529), .A2(new_n321), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n881), .B1(new_n883), .B2(new_n884), .ZN(G1348gat));
  NOR3_X1   g684(.A1(new_n880), .A2(new_n322), .A3(new_n617), .ZN(new_n886));
  INV_X1    g685(.A(new_n883), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n887), .A2(new_n616), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n886), .B1(new_n888), .B2(new_n322), .ZN(G1349gat));
  NAND3_X1  g688(.A1(new_n887), .A2(new_n348), .A3(new_n591), .ZN(new_n890));
  OAI21_X1  g689(.A(G183gat), .B1(new_n880), .B2(new_n871), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(KEYINPUT60), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT60), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n890), .A2(new_n894), .A3(new_n891), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n893), .A2(new_n895), .ZN(G1350gat));
  NAND3_X1  g695(.A1(new_n887), .A2(new_n327), .A3(new_n654), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n803), .A2(new_n654), .A3(new_n879), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT61), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n898), .A2(new_n899), .A3(G190gat), .ZN(new_n900));
  INV_X1    g699(.A(new_n900), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n899), .B1(new_n898), .B2(G190gat), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n897), .B1(new_n901), .B2(new_n902), .ZN(G1351gat));
  NOR2_X1   g702(.A1(new_n643), .A2(new_n250), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n882), .A2(new_n904), .ZN(new_n905));
  INV_X1    g704(.A(new_n905), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n906), .A2(new_n517), .A3(new_n529), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n878), .A2(new_n643), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n862), .A2(new_n863), .A3(new_n908), .ZN(new_n909));
  OAI21_X1  g708(.A(G197gat), .B1(new_n909), .B2(new_n708), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n907), .A2(new_n910), .ZN(G1352gat));
  OR2_X1    g710(.A1(new_n617), .A2(G204gat), .ZN(new_n912));
  NOR3_X1   g711(.A1(new_n905), .A2(KEYINPUT62), .A3(new_n912), .ZN(new_n913));
  OAI21_X1  g712(.A(KEYINPUT62), .B1(new_n905), .B2(new_n912), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(KEYINPUT125), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT125), .ZN(new_n916));
  OAI211_X1 g715(.A(new_n916), .B(KEYINPUT62), .C1(new_n905), .C2(new_n912), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n913), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n864), .A2(new_n908), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n919), .A2(G204gat), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n918), .A2(new_n920), .ZN(G1353gat));
  NAND3_X1  g720(.A1(new_n906), .A2(new_n204), .A3(new_n591), .ZN(new_n922));
  NAND4_X1  g721(.A1(new_n862), .A2(new_n591), .A3(new_n863), .A4(new_n908), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT126), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n204), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n835), .A2(new_n795), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n926), .A2(KEYINPUT121), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n835), .A2(new_n836), .A3(new_n795), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n654), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  INV_X1    g728(.A(new_n860), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n871), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  INV_X1    g730(.A(new_n801), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  AOI22_X1  g732(.A1(new_n933), .A2(new_n856), .B1(KEYINPUT57), .B2(new_n830), .ZN(new_n934));
  NAND4_X1  g733(.A1(new_n934), .A2(KEYINPUT126), .A3(new_n591), .A4(new_n908), .ZN(new_n935));
  AND3_X1   g734(.A1(new_n925), .A2(KEYINPUT63), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g735(.A(KEYINPUT63), .B1(new_n925), .B2(new_n935), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n922), .B1(new_n936), .B2(new_n937), .ZN(G1354gat));
  AOI21_X1  g737(.A(KEYINPUT127), .B1(new_n934), .B2(new_n908), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT127), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n654), .B1(new_n909), .B2(new_n940), .ZN(new_n941));
  OAI21_X1  g740(.A(G218gat), .B1(new_n939), .B2(new_n941), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n906), .A2(new_n205), .A3(new_n654), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(G1355gat));
endmodule


