//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 1 0 1 0 1 0 1 1 1 0 0 1 0 1 0 1 1 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 0 0 0 0 1 1 1 0 1 1 0 0 1 1 1 0 0 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:25 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n768, new_n769, new_n770,
    new_n772, new_n773, new_n774, new_n776, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n860, new_n861, new_n863,
    new_n864, new_n866, new_n867, new_n868, new_n869, new_n870, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n921, new_n922, new_n923,
    new_n924, new_n926, new_n927, new_n928, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n954, new_n955, new_n956,
    new_n957, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n983, new_n984, new_n985, new_n986, new_n988,
    new_n989;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G50gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(KEYINPUT90), .B(KEYINPUT31), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n205), .B(KEYINPUT91), .ZN(new_n206));
  XNOR2_X1  g005(.A(G197gat), .B(G204gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(G211gat), .A2(G218gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT22), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n207), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(G211gat), .ZN(new_n212));
  INV_X1    g011(.A(G218gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n211), .A2(new_n208), .A3(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n208), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n216), .A2(new_n207), .A3(new_n210), .ZN(new_n217));
  AND2_X1   g016(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(KEYINPUT75), .ZN(new_n219));
  AOI21_X1  g018(.A(KEYINPUT75), .B1(new_n215), .B2(new_n217), .ZN(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n219), .A2(KEYINPUT76), .A3(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT76), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n215), .A2(new_n217), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT75), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n223), .B1(new_n226), .B2(new_n220), .ZN(new_n227));
  AND2_X1   g026(.A1(new_n222), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(G148gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(KEYINPUT83), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT83), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(G148gat), .ZN(new_n232));
  AND3_X1   g031(.A1(new_n230), .A2(new_n232), .A3(G141gat), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT82), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n234), .B1(new_n229), .B2(G141gat), .ZN(new_n235));
  INV_X1    g034(.A(G141gat), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n236), .A2(KEYINPUT82), .A3(G148gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  OAI21_X1  g037(.A(KEYINPUT84), .B1(new_n233), .B2(new_n238), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n230), .A2(new_n232), .A3(G141gat), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT84), .ZN(new_n241));
  NAND4_X1  g040(.A1(new_n240), .A2(new_n241), .A3(new_n235), .A4(new_n237), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n239), .A2(new_n242), .ZN(new_n243));
  NOR2_X1   g042(.A1(G155gat), .A2(G162gat), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT2), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(G155gat), .A2(G162gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT80), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n247), .B1(new_n244), .B2(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(KEYINPUT80), .A2(G155gat), .A3(G162gat), .ZN(new_n251));
  AOI21_X1  g050(.A(KEYINPUT81), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n236), .A2(G148gat), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n229), .A2(G141gat), .ZN(new_n254));
  AOI22_X1  g053(.A1(new_n253), .A2(new_n254), .B1(KEYINPUT2), .B2(new_n247), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n252), .A2(new_n255), .ZN(new_n256));
  AND3_X1   g055(.A1(new_n250), .A2(KEYINPUT81), .A3(new_n251), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  AOI22_X1  g057(.A1(new_n243), .A2(new_n248), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  XOR2_X1   g058(.A(KEYINPUT86), .B(KEYINPUT3), .Z(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  XOR2_X1   g060(.A(KEYINPUT77), .B(KEYINPUT29), .Z(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n228), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(G228gat), .A2(G233gat), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT3), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n266), .B1(new_n218), .B2(KEYINPUT29), .ZN(new_n267));
  INV_X1    g066(.A(new_n242), .ZN(new_n268));
  AND3_X1   g067(.A1(new_n236), .A2(KEYINPUT82), .A3(G148gat), .ZN(new_n269));
  AOI21_X1  g068(.A(KEYINPUT82), .B1(new_n236), .B2(G148gat), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n241), .B1(new_n271), .B2(new_n240), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n248), .B1(new_n268), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n256), .A2(new_n258), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n265), .B1(new_n267), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n264), .A2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(G22gat), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n265), .B(KEYINPUT92), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n226), .A2(new_n220), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n280), .B1(new_n261), .B2(new_n262), .ZN(new_n281));
  OR2_X1    g080(.A1(new_n215), .A2(KEYINPUT93), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT93), .ZN(new_n283));
  OAI211_X1 g082(.A(new_n282), .B(new_n262), .C1(new_n283), .C2(new_n224), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n259), .B1(new_n284), .B2(new_n260), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n279), .B1(new_n281), .B2(new_n285), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n277), .A2(new_n278), .A3(new_n286), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n278), .B1(new_n277), .B2(new_n286), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n287), .B1(new_n288), .B2(KEYINPUT94), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n277), .A2(new_n286), .ZN(new_n290));
  AND3_X1   g089(.A1(new_n290), .A2(KEYINPUT94), .A3(G22gat), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n206), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n290), .A2(G22gat), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT95), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n288), .A2(KEYINPUT95), .ZN(new_n296));
  NAND4_X1  g095(.A1(new_n295), .A2(new_n296), .A3(new_n205), .A4(new_n287), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n292), .A2(new_n297), .ZN(new_n298));
  XOR2_X1   g097(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n299));
  INV_X1    g098(.A(KEYINPUT23), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n300), .B1(G169gat), .B2(G176gat), .ZN(new_n301));
  NOR2_X1   g100(.A1(G169gat), .A2(G176gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(KEYINPUT23), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT65), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n304), .B1(G169gat), .B2(G176gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(G169gat), .A2(G176gat), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n306), .A2(KEYINPUT65), .ZN(new_n307));
  OAI211_X1 g106(.A(new_n301), .B(new_n303), .C1(new_n305), .C2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(G183gat), .A2(G190gat), .ZN(new_n309));
  OAI21_X1  g108(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n310));
  AND2_X1   g109(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n311));
  AOI22_X1  g110(.A1(new_n309), .A2(new_n310), .B1(new_n311), .B2(G190gat), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n299), .B1(new_n308), .B2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT66), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  OAI211_X1 g114(.A(KEYINPUT66), .B(new_n299), .C1(new_n308), .C2(new_n312), .ZN(new_n316));
  INV_X1    g115(.A(new_n302), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(KEYINPUT67), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT67), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n302), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n318), .A2(KEYINPUT23), .A3(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(new_n312), .ZN(new_n322));
  OR2_X1    g121(.A1(new_n305), .A2(new_n307), .ZN(new_n323));
  AND2_X1   g122(.A1(new_n301), .A2(KEYINPUT25), .ZN(new_n324));
  NAND4_X1  g123(.A1(new_n321), .A2(new_n322), .A3(new_n323), .A4(new_n324), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n315), .A2(new_n316), .A3(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(G127gat), .B(G134gat), .ZN(new_n327));
  AND2_X1   g126(.A1(G113gat), .A2(G120gat), .ZN(new_n328));
  NOR2_X1   g127(.A1(G113gat), .A2(G120gat), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT1), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n327), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  OR2_X1    g131(.A1(KEYINPUT71), .A2(KEYINPUT1), .ZN(new_n333));
  INV_X1    g132(.A(G134gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(G127gat), .ZN(new_n335));
  INV_X1    g134(.A(G127gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(G134gat), .ZN(new_n337));
  NAND2_X1  g136(.A1(KEYINPUT71), .A2(KEYINPUT1), .ZN(new_n338));
  NAND4_X1  g137(.A1(new_n333), .A2(new_n335), .A3(new_n337), .A4(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT70), .ZN(new_n340));
  NOR3_X1   g139(.A1(new_n328), .A2(new_n329), .A3(new_n340), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n330), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(new_n340), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n332), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT28), .ZN(new_n347));
  XNOR2_X1  g146(.A(KEYINPUT27), .B(G183gat), .ZN(new_n348));
  INV_X1    g147(.A(G190gat), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n347), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT69), .ZN(new_n352));
  INV_X1    g151(.A(G183gat), .ZN(new_n353));
  OAI21_X1  g152(.A(KEYINPUT27), .B1(new_n353), .B2(KEYINPUT68), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT68), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT27), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n355), .A2(new_n356), .A3(G183gat), .ZN(new_n357));
  NAND4_X1  g156(.A1(new_n354), .A2(new_n357), .A3(new_n347), .A4(new_n349), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n351), .A2(new_n352), .A3(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n358), .ZN(new_n360));
  OAI21_X1  g159(.A(KEYINPUT69), .B1(new_n360), .B2(new_n350), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n317), .A2(KEYINPUT26), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n318), .A2(new_n320), .ZN(new_n363));
  OAI211_X1 g162(.A(new_n323), .B(new_n362), .C1(new_n363), .C2(KEYINPUT26), .ZN(new_n364));
  NAND4_X1  g163(.A1(new_n359), .A2(new_n361), .A3(new_n364), .A4(new_n309), .ZN(new_n365));
  AND3_X1   g164(.A1(new_n326), .A2(new_n346), .A3(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n346), .B1(new_n326), .B2(new_n365), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(G227gat), .ZN(new_n369));
  INV_X1    g168(.A(G233gat), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n368), .A2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT34), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  OAI221_X1 g173(.A(new_n373), .B1(new_n369), .B2(new_n370), .C1(new_n366), .C2(new_n367), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT32), .ZN(new_n379));
  XNOR2_X1  g178(.A(G15gat), .B(G43gat), .ZN(new_n380));
  XNOR2_X1  g179(.A(G71gat), .B(G99gat), .ZN(new_n381));
  XNOR2_X1  g180(.A(new_n380), .B(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n379), .B1(new_n383), .B2(KEYINPUT33), .ZN(new_n384));
  AOI21_X1  g183(.A(KEYINPUT72), .B1(new_n368), .B2(new_n371), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n326), .A2(new_n365), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(new_n345), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n326), .A2(new_n346), .A3(new_n365), .ZN(new_n388));
  NAND4_X1  g187(.A1(new_n387), .A2(KEYINPUT72), .A3(new_n371), .A4(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n384), .B1(new_n385), .B2(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n387), .A2(new_n371), .A3(new_n388), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT72), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  AOI22_X1  g193(.A1(new_n394), .A2(new_n389), .B1(new_n379), .B2(KEYINPUT33), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n391), .B1(new_n395), .B2(new_n382), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n378), .A2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(new_n396), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(new_n377), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n298), .A2(new_n397), .A3(new_n399), .ZN(new_n400));
  XNOR2_X1  g199(.A(G1gat), .B(G29gat), .ZN(new_n401));
  XNOR2_X1  g200(.A(new_n401), .B(KEYINPUT0), .ZN(new_n402));
  XNOR2_X1  g201(.A(G57gat), .B(G85gat), .ZN(new_n403));
  XOR2_X1   g202(.A(new_n402), .B(new_n403), .Z(new_n404));
  INV_X1    g203(.A(KEYINPUT4), .ZN(new_n405));
  NAND4_X1  g204(.A1(new_n273), .A2(new_n405), .A3(new_n345), .A4(new_n274), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT87), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n259), .A2(KEYINPUT87), .A3(new_n405), .A4(new_n345), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n273), .A2(new_n345), .A3(new_n274), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(KEYINPUT4), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n408), .A2(new_n409), .A3(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n345), .B1(new_n259), .B2(new_n260), .ZN(new_n413));
  INV_X1    g212(.A(new_n248), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n414), .B1(new_n239), .B2(new_n242), .ZN(new_n415));
  NOR3_X1   g214(.A1(new_n257), .A2(new_n252), .A3(new_n255), .ZN(new_n416));
  OAI21_X1  g215(.A(KEYINPUT3), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT85), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  OAI211_X1 g218(.A(KEYINPUT85), .B(KEYINPUT3), .C1(new_n415), .C2(new_n416), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n413), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(G225gat), .A2(G233gat), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n412), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT5), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n275), .A2(new_n346), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(new_n410), .ZN(new_n426));
  INV_X1    g225(.A(new_n422), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n424), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n423), .A2(new_n428), .ZN(new_n429));
  AOI21_X1  g228(.A(KEYINPUT5), .B1(new_n411), .B2(new_n406), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n430), .A2(new_n421), .A3(new_n422), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n404), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  XOR2_X1   g231(.A(KEYINPUT88), .B(KEYINPUT6), .Z(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  AND2_X1   g234(.A1(new_n421), .A2(new_n422), .ZN(new_n436));
  AOI22_X1  g235(.A1(new_n436), .A2(new_n430), .B1(new_n423), .B2(new_n428), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n433), .B1(new_n437), .B2(new_n404), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n429), .A2(new_n431), .ZN(new_n439));
  INV_X1    g238(.A(new_n404), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n435), .B1(new_n438), .B2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  AND2_X1   g242(.A1(G226gat), .A2(G233gat), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n386), .A2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n444), .B1(new_n386), .B2(new_n262), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n228), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(KEYINPUT29), .B1(new_n326), .B2(new_n365), .ZN(new_n449));
  OAI211_X1 g248(.A(new_n445), .B(new_n280), .C1(new_n444), .C2(new_n449), .ZN(new_n450));
  XNOR2_X1  g249(.A(G8gat), .B(G36gat), .ZN(new_n451));
  XNOR2_X1  g250(.A(new_n451), .B(KEYINPUT78), .ZN(new_n452));
  XNOR2_X1  g251(.A(G64gat), .B(G92gat), .ZN(new_n453));
  XOR2_X1   g252(.A(new_n452), .B(new_n453), .Z(new_n454));
  INV_X1    g253(.A(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n448), .A2(new_n450), .A3(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(KEYINPUT30), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n448), .A2(new_n450), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(new_n454), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT30), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n456), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n458), .A2(new_n460), .A3(new_n462), .ZN(new_n463));
  OR2_X1    g262(.A1(new_n463), .A2(KEYINPUT35), .ZN(new_n464));
  NOR3_X1   g263(.A1(new_n400), .A2(new_n443), .A3(new_n464), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n434), .B1(new_n439), .B2(new_n440), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n437), .A2(new_n404), .ZN(new_n467));
  AOI21_X1  g266(.A(KEYINPUT89), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n468), .B1(KEYINPUT89), .B2(new_n442), .ZN(new_n469));
  INV_X1    g268(.A(new_n462), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n460), .B1(new_n461), .B2(new_n456), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT79), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n458), .A2(KEYINPUT79), .A3(new_n460), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n469), .A2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT73), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n394), .A2(new_n389), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n379), .A2(KEYINPUT33), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n382), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(new_n384), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n481), .B1(new_n394), .B2(new_n389), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n477), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  OAI211_X1 g282(.A(new_n391), .B(KEYINPUT73), .C1(new_n395), .C2(new_n382), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n483), .A2(new_n484), .A3(new_n378), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT74), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n377), .B1(new_n396), .B2(new_n477), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n488), .A2(KEYINPUT74), .A3(new_n484), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  AOI22_X1  g289(.A1(new_n292), .A2(new_n297), .B1(new_n398), .B2(new_n377), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n476), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n465), .B1(new_n492), .B2(KEYINPUT35), .ZN(new_n493));
  INV_X1    g292(.A(new_n459), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT37), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n455), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n496), .B1(new_n495), .B2(new_n494), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(KEYINPUT38), .ZN(new_n498));
  OR2_X1    g297(.A1(new_n446), .A2(new_n447), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n449), .A2(new_n444), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n446), .A2(new_n500), .ZN(new_n501));
  OAI22_X1  g300(.A1(new_n499), .A2(new_n228), .B1(new_n501), .B2(new_n280), .ZN(new_n502));
  AOI21_X1  g301(.A(KEYINPUT38), .B1(new_n502), .B2(KEYINPUT37), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n457), .B1(new_n503), .B2(new_n496), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n498), .A2(new_n443), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n411), .A2(new_n406), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n422), .B1(new_n421), .B2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT39), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  OAI21_X1  g308(.A(KEYINPUT39), .B1(new_n426), .B2(new_n427), .ZN(new_n510));
  OAI211_X1 g309(.A(new_n509), .B(new_n404), .C1(new_n507), .C2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT40), .ZN(new_n512));
  OR2_X1    g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(new_n432), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n511), .A2(new_n512), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n463), .A2(new_n513), .A3(new_n514), .A4(new_n515), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n505), .A2(new_n298), .A3(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(new_n298), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n519), .B1(new_n469), .B2(new_n475), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n399), .A2(KEYINPUT36), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n521), .B1(new_n487), .B2(new_n489), .ZN(new_n522));
  AOI21_X1  g321(.A(KEYINPUT36), .B1(new_n399), .B2(new_n397), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n520), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n518), .B1(new_n524), .B2(KEYINPUT96), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT96), .ZN(new_n526));
  OAI211_X1 g325(.A(new_n520), .B(new_n526), .C1(new_n522), .C2(new_n523), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n493), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  XNOR2_X1  g327(.A(G15gat), .B(G22gat), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT16), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n529), .B1(new_n530), .B2(G1gat), .ZN(new_n531));
  OAI211_X1 g330(.A(new_n531), .B(KEYINPUT101), .C1(G1gat), .C2(new_n529), .ZN(new_n532));
  OAI211_X1 g331(.A(new_n532), .B(G8gat), .C1(KEYINPUT101), .C2(new_n531), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n533), .B(KEYINPUT102), .ZN(new_n534));
  XOR2_X1   g333(.A(KEYINPUT103), .B(G8gat), .Z(new_n535));
  OAI211_X1 g334(.A(new_n531), .B(new_n535), .C1(G1gat), .C2(new_n529), .ZN(new_n536));
  AND2_X1   g335(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  OAI21_X1  g336(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  OR3_X1    g338(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n539), .B1(new_n540), .B2(KEYINPUT98), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n541), .B1(KEYINPUT98), .B2(new_n540), .ZN(new_n542));
  NAND2_X1  g341(.A1(G29gat), .A2(G36gat), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(G43gat), .B(G50gat), .ZN(new_n545));
  OR2_X1    g344(.A1(new_n545), .A2(KEYINPUT97), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(KEYINPUT97), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n546), .A2(KEYINPUT15), .A3(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n544), .A2(new_n549), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n545), .A2(KEYINPUT15), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n551), .B1(G29gat), .B2(G36gat), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n548), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n540), .A2(new_n538), .ZN(new_n554));
  XOR2_X1   g353(.A(new_n554), .B(KEYINPUT99), .Z(new_n555));
  OAI21_X1  g354(.A(new_n550), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(KEYINPUT17), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT17), .ZN(new_n559));
  AOI21_X1  g358(.A(KEYINPUT100), .B1(new_n556), .B2(new_n559), .ZN(new_n560));
  AND3_X1   g359(.A1(new_n556), .A2(KEYINPUT100), .A3(new_n559), .ZN(new_n561));
  OAI211_X1 g360(.A(new_n537), .B(new_n558), .C1(new_n560), .C2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(G229gat), .A2(G233gat), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n534), .A2(new_n536), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n564), .A2(new_n556), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n562), .A2(new_n563), .A3(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT18), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND4_X1  g367(.A1(new_n562), .A2(KEYINPUT18), .A3(new_n563), .A4(new_n565), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n537), .A2(new_n557), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n570), .A2(new_n565), .ZN(new_n571));
  XOR2_X1   g370(.A(new_n563), .B(KEYINPUT13), .Z(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n568), .A2(new_n569), .A3(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(G113gat), .B(G141gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n575), .B(G197gat), .ZN(new_n576));
  XOR2_X1   g375(.A(KEYINPUT11), .B(G169gat), .Z(new_n577));
  XNOR2_X1  g376(.A(new_n576), .B(new_n577), .ZN(new_n578));
  XOR2_X1   g377(.A(new_n578), .B(KEYINPUT12), .Z(new_n579));
  NAND2_X1  g378(.A1(new_n574), .A2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n579), .ZN(new_n581));
  NAND4_X1  g380(.A1(new_n568), .A2(new_n581), .A3(new_n569), .A4(new_n573), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n528), .A2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(G57gat), .ZN(new_n586));
  AND2_X1   g385(.A1(new_n586), .A2(G64gat), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT104), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n586), .A2(G64gat), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n587), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  OAI21_X1  g389(.A(KEYINPUT104), .B1(new_n586), .B2(G64gat), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(G71gat), .A2(G78gat), .ZN(new_n593));
  OR2_X1    g392(.A1(G71gat), .A2(G78gat), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT9), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n593), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n592), .A2(new_n596), .ZN(new_n597));
  OAI21_X1  g396(.A(KEYINPUT9), .B1(new_n587), .B2(new_n589), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n598), .A2(new_n593), .A3(new_n594), .ZN(new_n599));
  AND2_X1   g398(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n600), .A2(KEYINPUT21), .ZN(new_n601));
  NAND2_X1  g400(.A1(G231gat), .A2(G233gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(G127gat), .B(G155gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n604), .B(KEYINPUT105), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n603), .B(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(G183gat), .B(G211gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n564), .B1(KEYINPUT21), .B2(new_n600), .ZN(new_n609));
  XOR2_X1   g408(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  OR2_X1    g410(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n608), .A2(new_n611), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(G85gat), .A2(G92gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n616), .B(KEYINPUT7), .ZN(new_n617));
  NAND2_X1  g416(.A1(G99gat), .A2(G106gat), .ZN(new_n618));
  INV_X1    g417(.A(G85gat), .ZN(new_n619));
  INV_X1    g418(.A(G92gat), .ZN(new_n620));
  AOI22_X1  g419(.A1(KEYINPUT8), .A2(new_n618), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n617), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(G99gat), .B(G106gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n622), .B(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(KEYINPUT106), .ZN(new_n625));
  OAI211_X1 g424(.A(new_n625), .B(new_n558), .C1(new_n561), .C2(new_n560), .ZN(new_n626));
  AND2_X1   g425(.A1(G232gat), .A2(G233gat), .ZN(new_n627));
  AOI22_X1  g426(.A1(new_n556), .A2(new_n624), .B1(KEYINPUT41), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(G190gat), .B(G218gat), .ZN(new_n630));
  XOR2_X1   g429(.A(new_n630), .B(KEYINPUT107), .Z(new_n631));
  OR2_X1    g430(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n629), .A2(new_n631), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n627), .A2(KEYINPUT41), .ZN(new_n635));
  XNOR2_X1  g434(.A(G134gat), .B(G162gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n634), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n632), .A2(new_n637), .A3(new_n633), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n615), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(G120gat), .B(G148gat), .ZN(new_n644));
  XNOR2_X1  g443(.A(G176gat), .B(G204gat), .ZN(new_n645));
  XOR2_X1   g444(.A(new_n644), .B(new_n645), .Z(new_n646));
  NAND2_X1  g445(.A1(G230gat), .A2(G233gat), .ZN(new_n647));
  XOR2_X1   g446(.A(new_n622), .B(new_n623), .Z(new_n648));
  NAND2_X1  g447(.A1(new_n597), .A2(new_n599), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n600), .A2(new_n624), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n650), .A2(KEYINPUT108), .A3(new_n651), .ZN(new_n652));
  OR3_X1    g451(.A1(new_n600), .A2(new_n624), .A3(KEYINPUT108), .ZN(new_n653));
  AOI21_X1  g452(.A(KEYINPUT10), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  AND3_X1   g453(.A1(new_n600), .A2(new_n624), .A3(KEYINPUT10), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n647), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  OR2_X1    g455(.A1(new_n656), .A2(KEYINPUT110), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(KEYINPUT110), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n647), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n652), .A2(new_n660), .A3(new_n653), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n646), .B1(new_n659), .B2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT109), .ZN(new_n663));
  OR2_X1    g462(.A1(new_n656), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n656), .A2(new_n663), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n661), .A2(new_n646), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n662), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n643), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n585), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n469), .ZN(new_n674));
  OR2_X1    g473(.A1(new_n674), .A2(KEYINPUT111), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(KEYINPUT111), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n673), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n678), .B(G1gat), .ZN(G1324gat));
  INV_X1    g478(.A(KEYINPUT112), .ZN(new_n680));
  INV_X1    g479(.A(new_n463), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n672), .A2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(G8gat), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n680), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  OAI211_X1 g483(.A(KEYINPUT112), .B(G8gat), .C1(new_n672), .C2(new_n681), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT42), .ZN(new_n686));
  XOR2_X1   g485(.A(KEYINPUT16), .B(G8gat), .Z(new_n687));
  AND3_X1   g486(.A1(new_n682), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n686), .B1(new_n682), .B2(new_n687), .ZN(new_n689));
  OAI211_X1 g488(.A(new_n684), .B(new_n685), .C1(new_n688), .C2(new_n689), .ZN(G1325gat));
  NAND2_X1  g489(.A1(new_n399), .A2(new_n397), .ZN(new_n691));
  OR3_X1    g490(.A1(new_n672), .A2(G15gat), .A3(new_n691), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n522), .A2(new_n523), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  OAI21_X1  g493(.A(G15gat), .B1(new_n672), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n692), .A2(new_n695), .ZN(G1326gat));
  NOR2_X1   g495(.A1(new_n672), .A2(new_n298), .ZN(new_n697));
  XOR2_X1   g496(.A(KEYINPUT43), .B(G22gat), .Z(new_n698));
  XNOR2_X1  g497(.A(new_n697), .B(new_n698), .ZN(G1327gat));
  NAND2_X1  g498(.A1(new_n614), .A2(new_n669), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n700), .A2(new_n642), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n585), .A2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(new_n677), .ZN(new_n703));
  NOR3_X1   g502(.A1(new_n702), .A2(G29gat), .A3(new_n703), .ZN(new_n704));
  OR2_X1    g503(.A1(new_n704), .A2(KEYINPUT45), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n524), .A2(KEYINPUT96), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n706), .A2(new_n527), .A3(new_n517), .ZN(new_n707));
  AND4_X1   g506(.A1(KEYINPUT74), .A2(new_n483), .A3(new_n484), .A4(new_n378), .ZN(new_n708));
  AOI21_X1  g507(.A(KEYINPUT74), .B1(new_n488), .B2(new_n484), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n491), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT89), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n466), .A2(new_n467), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n711), .B1(new_n712), .B2(new_n435), .ZN(new_n713));
  OAI211_X1 g512(.A(new_n474), .B(new_n473), .C1(new_n713), .C2(new_n468), .ZN(new_n714));
  OAI21_X1  g513(.A(KEYINPUT35), .B1(new_n710), .B2(new_n714), .ZN(new_n715));
  OR3_X1    g514(.A1(new_n400), .A2(new_n443), .A3(new_n464), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n707), .A2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT44), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n642), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  OAI211_X1 g520(.A(new_n517), .B(new_n520), .C1(new_n522), .C2(new_n523), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n717), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(new_n641), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(new_n719), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n700), .A2(new_n584), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n721), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(G29gat), .B1(new_n727), .B2(new_n703), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n704), .A2(KEYINPUT45), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n705), .A2(new_n728), .A3(new_n729), .ZN(G1328gat));
  INV_X1    g529(.A(new_n702), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT113), .ZN(new_n732));
  AOI211_X1 g531(.A(G36gat), .B(new_n681), .C1(new_n732), .C2(KEYINPUT46), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n734), .B1(new_n732), .B2(KEYINPUT46), .ZN(new_n735));
  OAI21_X1  g534(.A(G36gat), .B1(new_n727), .B2(new_n681), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n732), .A2(KEYINPUT46), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n731), .A2(new_n737), .A3(new_n733), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n735), .A2(new_n736), .A3(new_n738), .ZN(G1329gat));
  NOR2_X1   g538(.A1(new_n691), .A2(G43gat), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n731), .A2(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(new_n720), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n642), .B1(new_n717), .B2(new_n722), .ZN(new_n743));
  OAI22_X1  g542(.A1(new_n528), .A2(new_n742), .B1(new_n743), .B2(KEYINPUT44), .ZN(new_n744));
  INV_X1    g543(.A(new_n726), .ZN(new_n745));
  NOR3_X1   g544(.A1(new_n744), .A2(new_n694), .A3(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT115), .ZN(new_n747));
  OAI21_X1  g546(.A(G43gat), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NOR3_X1   g547(.A1(new_n727), .A2(KEYINPUT115), .A3(new_n694), .ZN(new_n749));
  OAI211_X1 g548(.A(KEYINPUT47), .B(new_n741), .C1(new_n748), .C2(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(G43gat), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n741), .B1(new_n746), .B2(new_n751), .ZN(new_n752));
  XNOR2_X1  g551(.A(KEYINPUT114), .B(KEYINPUT47), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n750), .A2(new_n754), .ZN(G1330gat));
  NOR2_X1   g554(.A1(new_n727), .A2(new_n298), .ZN(new_n756));
  INV_X1    g555(.A(G50gat), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n519), .A2(new_n757), .ZN(new_n758));
  OAI22_X1  g557(.A1(new_n756), .A2(new_n757), .B1(new_n702), .B2(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT48), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  OAI221_X1 g560(.A(KEYINPUT48), .B1(new_n702), .B2(new_n758), .C1(new_n756), .C2(new_n757), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(G1331gat));
  NOR3_X1   g562(.A1(new_n643), .A2(new_n583), .A3(new_n669), .ZN(new_n764));
  AND2_X1   g563(.A1(new_n723), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(new_n677), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g566(.A1(new_n765), .A2(new_n463), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n768), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n769));
  XOR2_X1   g568(.A(KEYINPUT49), .B(G64gat), .Z(new_n770));
  OAI21_X1  g569(.A(new_n769), .B1(new_n768), .B2(new_n770), .ZN(G1333gat));
  NAND2_X1  g570(.A1(new_n765), .A2(new_n693), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n691), .A2(G71gat), .ZN(new_n773));
  AOI22_X1  g572(.A1(new_n772), .A2(G71gat), .B1(new_n765), .B2(new_n773), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n774), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g574(.A1(new_n765), .A2(new_n519), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g576(.A1(new_n615), .A2(new_n583), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n743), .A2(KEYINPUT51), .A3(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT117), .ZN(new_n780));
  OR2_X1    g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n743), .A2(new_n778), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT51), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n779), .A2(new_n780), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n781), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  NAND4_X1  g585(.A1(new_n786), .A2(new_n619), .A3(new_n670), .A4(new_n677), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n778), .A2(new_n670), .ZN(new_n788));
  OAI21_X1  g587(.A(KEYINPUT116), .B1(new_n744), .B2(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT116), .ZN(new_n790));
  INV_X1    g589(.A(new_n788), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n721), .A2(new_n725), .A3(new_n790), .A4(new_n791), .ZN(new_n792));
  AND3_X1   g591(.A1(new_n789), .A2(new_n677), .A3(new_n792), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n787), .B1(new_n619), .B2(new_n793), .ZN(G1336gat));
  NOR3_X1   g593(.A1(new_n669), .A2(G92gat), .A3(new_n681), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n786), .A2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT52), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n721), .A2(new_n725), .A3(new_n791), .ZN(new_n798));
  OAI21_X1  g597(.A(G92gat), .B1(new_n798), .B2(new_n681), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n796), .A2(new_n797), .A3(new_n799), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n789), .A2(new_n463), .A3(new_n792), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n784), .A2(new_n779), .ZN(new_n802));
  AOI22_X1  g601(.A1(new_n801), .A2(G92gat), .B1(new_n802), .B2(new_n795), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n800), .B1(new_n803), .B2(new_n797), .ZN(G1337gat));
  NAND3_X1  g603(.A1(new_n789), .A2(new_n693), .A3(new_n792), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT118), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n789), .A2(KEYINPUT118), .A3(new_n792), .A4(new_n693), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n807), .A2(G99gat), .A3(new_n808), .ZN(new_n809));
  NOR3_X1   g608(.A1(new_n669), .A2(new_n691), .A3(G99gat), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n786), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n809), .A2(new_n811), .ZN(G1338gat));
  NOR3_X1   g611(.A1(new_n669), .A2(new_n298), .A3(G106gat), .ZN(new_n813));
  XOR2_X1   g612(.A(new_n813), .B(KEYINPUT119), .Z(new_n814));
  NAND2_X1  g613(.A1(new_n786), .A2(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT53), .ZN(new_n816));
  OAI21_X1  g615(.A(G106gat), .B1(new_n798), .B2(new_n298), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n815), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n789), .A2(new_n519), .A3(new_n792), .ZN(new_n819));
  AOI22_X1  g618(.A1(new_n819), .A2(G106gat), .B1(new_n802), .B2(new_n814), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n818), .B1(new_n820), .B2(new_n816), .ZN(G1339gat));
  NOR3_X1   g620(.A1(new_n643), .A2(new_n583), .A3(new_n670), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT54), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n654), .A2(new_n655), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(new_n660), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n823), .B1(new_n825), .B2(KEYINPUT120), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT120), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n824), .A2(new_n827), .A3(new_n660), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n826), .A2(new_n664), .A3(new_n665), .A4(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(new_n646), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n657), .A2(new_n823), .A3(new_n658), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n829), .A2(KEYINPUT55), .A3(new_n830), .A4(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(new_n668), .ZN(new_n833));
  AND2_X1   g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n571), .A2(new_n572), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n563), .B1(new_n562), .B2(new_n565), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n578), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  AND2_X1   g636(.A1(new_n582), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n825), .A2(KEYINPUT120), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n839), .A2(KEYINPUT54), .A3(new_n828), .ZN(new_n840));
  OAI211_X1 g639(.A(new_n830), .B(new_n831), .C1(new_n840), .C2(new_n666), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT55), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n834), .A2(new_n641), .A3(new_n838), .A4(new_n843), .ZN(new_n844));
  AOI22_X1  g643(.A1(new_n842), .A2(new_n841), .B1(new_n580), .B2(new_n582), .ZN(new_n845));
  AOI22_X1  g644(.A1(new_n834), .A2(new_n845), .B1(new_n670), .B2(new_n838), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n844), .B1(new_n846), .B2(new_n641), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n822), .B1(new_n847), .B2(new_n614), .ZN(new_n848));
  NOR3_X1   g647(.A1(new_n848), .A2(new_n463), .A3(new_n703), .ZN(new_n849));
  INV_X1    g648(.A(new_n400), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(G113gat), .ZN(new_n852));
  NOR3_X1   g651(.A1(new_n851), .A2(new_n852), .A3(new_n584), .ZN(new_n853));
  INV_X1    g652(.A(new_n710), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n849), .A2(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(new_n583), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n853), .B1(new_n852), .B2(new_n857), .ZN(G1340gat));
  INV_X1    g657(.A(G120gat), .ZN(new_n859));
  NOR3_X1   g658(.A1(new_n851), .A2(new_n859), .A3(new_n669), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n856), .A2(new_n670), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n860), .B1(new_n859), .B2(new_n861), .ZN(G1341gat));
  OAI21_X1  g661(.A(G127gat), .B1(new_n851), .B2(new_n614), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n615), .A2(new_n336), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n863), .B1(new_n855), .B2(new_n864), .ZN(G1342gat));
  NOR2_X1   g664(.A1(new_n642), .A2(G134gat), .ZN(new_n866));
  INV_X1    g665(.A(new_n866), .ZN(new_n867));
  OR3_X1    g666(.A1(new_n855), .A2(KEYINPUT56), .A3(new_n867), .ZN(new_n868));
  OAI21_X1  g667(.A(G134gat), .B1(new_n851), .B2(new_n642), .ZN(new_n869));
  OAI21_X1  g668(.A(KEYINPUT56), .B1(new_n855), .B2(new_n867), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n868), .A2(new_n869), .A3(new_n870), .ZN(G1343gat));
  NAND4_X1  g670(.A1(new_n843), .A2(new_n583), .A3(new_n833), .A4(new_n832), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n670), .A2(new_n838), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n641), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n843), .A2(new_n641), .A3(new_n838), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n832), .A2(new_n833), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n614), .B1(new_n874), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n671), .A2(new_n584), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n693), .A2(new_n298), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n880), .A2(new_n677), .A3(new_n881), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT122), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NOR3_X1   g683(.A1(new_n584), .A2(G141gat), .A3(new_n463), .ZN(new_n885));
  NAND4_X1  g684(.A1(new_n880), .A2(KEYINPUT122), .A3(new_n677), .A4(new_n881), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n884), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  XNOR2_X1  g686(.A(new_n887), .B(KEYINPUT123), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n677), .A2(new_n694), .A3(new_n681), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n298), .B1(new_n878), .B2(new_n879), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT57), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n889), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n844), .B1(new_n874), .B2(KEYINPUT121), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT121), .ZN(new_n894));
  NOR3_X1   g693(.A1(new_n846), .A2(new_n894), .A3(new_n641), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n614), .B1(new_n893), .B2(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n298), .B1(new_n896), .B2(new_n879), .ZN(new_n897));
  OAI211_X1 g696(.A(new_n583), .B(new_n892), .C1(new_n897), .C2(new_n891), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(G141gat), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT58), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  INV_X1    g700(.A(new_n882), .ZN(new_n902));
  AOI22_X1  g701(.A1(new_n898), .A2(G141gat), .B1(new_n902), .B2(new_n885), .ZN(new_n903));
  OAI22_X1  g702(.A1(new_n888), .A2(new_n901), .B1(new_n900), .B2(new_n903), .ZN(G1344gat));
  AND2_X1   g703(.A1(new_n230), .A2(new_n232), .ZN(new_n905));
  AND2_X1   g704(.A1(new_n670), .A2(new_n905), .ZN(new_n906));
  NAND4_X1  g705(.A1(new_n884), .A2(new_n681), .A3(new_n886), .A4(new_n906), .ZN(new_n907));
  OR2_X1    g706(.A1(new_n905), .A2(KEYINPUT59), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n897), .A2(new_n891), .ZN(new_n909));
  INV_X1    g708(.A(new_n892), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n908), .B1(new_n911), .B2(new_n670), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT59), .ZN(new_n913));
  OAI21_X1  g712(.A(KEYINPUT57), .B1(new_n848), .B2(new_n298), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n890), .A2(new_n891), .ZN(new_n915));
  AND2_X1   g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  INV_X1    g715(.A(new_n889), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n916), .A2(new_n670), .A3(new_n917), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n913), .B1(new_n918), .B2(G148gat), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n907), .B1(new_n912), .B2(new_n919), .ZN(G1345gat));
  NAND2_X1  g719(.A1(new_n911), .A2(new_n615), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(G155gat), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n614), .A2(G155gat), .ZN(new_n923));
  NAND4_X1  g722(.A1(new_n884), .A2(new_n681), .A3(new_n886), .A4(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n922), .A2(new_n924), .ZN(G1346gat));
  INV_X1    g724(.A(G162gat), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n642), .A2(new_n926), .ZN(new_n927));
  NAND4_X1  g726(.A1(new_n884), .A2(new_n681), .A3(new_n641), .A4(new_n886), .ZN(new_n928));
  AOI22_X1  g727(.A1(new_n911), .A2(new_n927), .B1(new_n926), .B2(new_n928), .ZN(G1347gat));
  NOR3_X1   g728(.A1(new_n848), .A2(new_n681), .A3(new_n677), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n930), .A2(new_n850), .ZN(new_n931));
  INV_X1    g730(.A(G169gat), .ZN(new_n932));
  NOR3_X1   g731(.A1(new_n931), .A2(new_n932), .A3(new_n584), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n930), .A2(new_n583), .A3(new_n854), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n933), .B1(new_n932), .B2(new_n934), .ZN(G1348gat));
  INV_X1    g734(.A(G176gat), .ZN(new_n936));
  NAND4_X1  g735(.A1(new_n880), .A2(new_n854), .A3(new_n463), .A4(new_n703), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n936), .B1(new_n937), .B2(new_n669), .ZN(new_n938));
  XNOR2_X1  g737(.A(new_n938), .B(KEYINPUT124), .ZN(new_n939));
  NOR3_X1   g738(.A1(new_n931), .A2(new_n936), .A3(new_n669), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n939), .A2(new_n940), .ZN(G1349gat));
  OAI21_X1  g740(.A(G183gat), .B1(new_n931), .B2(new_n614), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT125), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n615), .A2(new_n348), .ZN(new_n944));
  INV_X1    g743(.A(new_n944), .ZN(new_n945));
  NAND4_X1  g744(.A1(new_n930), .A2(new_n943), .A3(new_n854), .A4(new_n945), .ZN(new_n946));
  OAI21_X1  g745(.A(KEYINPUT125), .B1(new_n937), .B2(new_n944), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n942), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n949), .A2(KEYINPUT60), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT60), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n942), .A2(new_n948), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n950), .A2(new_n952), .ZN(G1350gat));
  OAI21_X1  g752(.A(G190gat), .B1(new_n931), .B2(new_n642), .ZN(new_n954));
  AND2_X1   g753(.A1(new_n954), .A2(KEYINPUT61), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n954), .A2(KEYINPUT61), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n641), .A2(new_n349), .ZN(new_n957));
  OAI22_X1  g756(.A1(new_n955), .A2(new_n956), .B1(new_n937), .B2(new_n957), .ZN(G1351gat));
  NOR3_X1   g757(.A1(new_n677), .A2(new_n693), .A3(new_n681), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n916), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g759(.A(G197gat), .B1(new_n960), .B2(new_n584), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n848), .A2(new_n677), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n694), .A2(new_n519), .A3(new_n463), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT126), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  AND2_X1   g764(.A1(new_n962), .A2(new_n965), .ZN(new_n966));
  OR2_X1    g765(.A1(new_n963), .A2(new_n964), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  OR2_X1    g767(.A1(new_n584), .A2(G197gat), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n961), .B1(new_n968), .B2(new_n969), .ZN(G1352gat));
  INV_X1    g769(.A(KEYINPUT62), .ZN(new_n971));
  NOR2_X1   g770(.A1(new_n669), .A2(G204gat), .ZN(new_n972));
  NAND4_X1  g771(.A1(new_n966), .A2(new_n971), .A3(new_n967), .A4(new_n972), .ZN(new_n973));
  NAND4_X1  g772(.A1(new_n914), .A2(new_n915), .A3(new_n670), .A4(new_n959), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n974), .A2(G204gat), .ZN(new_n975));
  NAND4_X1  g774(.A1(new_n962), .A2(new_n967), .A3(new_n965), .A4(new_n972), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n976), .A2(KEYINPUT62), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n973), .A2(new_n975), .A3(new_n977), .ZN(new_n978));
  INV_X1    g777(.A(KEYINPUT127), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND4_X1  g779(.A1(new_n973), .A2(new_n975), .A3(KEYINPUT127), .A4(new_n977), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n980), .A2(new_n981), .ZN(G1353gat));
  NAND4_X1  g781(.A1(new_n914), .A2(new_n915), .A3(new_n615), .A4(new_n959), .ZN(new_n983));
  AND3_X1   g782(.A1(new_n983), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n984));
  AOI21_X1  g783(.A(KEYINPUT63), .B1(new_n983), .B2(G211gat), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n615), .A2(new_n212), .ZN(new_n986));
  OAI22_X1  g785(.A1(new_n984), .A2(new_n985), .B1(new_n968), .B2(new_n986), .ZN(G1354gat));
  OAI21_X1  g786(.A(G218gat), .B1(new_n960), .B2(new_n642), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n641), .A2(new_n213), .ZN(new_n989));
  OAI21_X1  g788(.A(new_n988), .B1(new_n968), .B2(new_n989), .ZN(G1355gat));
endmodule


