//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 0 1 1 1 1 0 1 1 0 1 0 1 1 0 0 0 1 0 0 1 0 1 1 1 0 1 1 0 0 1 1 1 0 1 0 1 1 1 1 0 0 0 1 1 1 1 0 1 0 1 1 0 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:52 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n632, new_n633, new_n634, new_n635, new_n637, new_n638,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n682,
    new_n683, new_n684, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n722, new_n723, new_n724, new_n725, new_n727, new_n728, new_n729,
    new_n731, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n742, new_n743, new_n744, new_n746, new_n747,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n787, new_n789, new_n791, new_n792, new_n793, new_n794,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n846,
    new_n847, new_n849, new_n850, new_n852, new_n853, new_n854, new_n855,
    new_n857, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n887, new_n888,
    new_n889, new_n890, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n910, new_n911;
  INV_X1    g000(.A(KEYINPUT30), .ZN(new_n202));
  XNOR2_X1  g001(.A(G8gat), .B(G36gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(G64gat), .B(G92gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT78), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT28), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(KEYINPUT65), .ZN(new_n208));
  INV_X1    g007(.A(G190gat), .ZN(new_n209));
  AND2_X1   g008(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n210));
  NOR2_X1   g009(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n211));
  OAI211_X1 g010(.A(new_n208), .B(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT65), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(KEYINPUT28), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(KEYINPUT27), .B(G183gat), .ZN(new_n216));
  NAND4_X1  g015(.A1(new_n216), .A2(new_n213), .A3(KEYINPUT28), .A4(new_n209), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  OAI21_X1  g017(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(G169gat), .A2(G176gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(KEYINPUT66), .ZN(new_n222));
  NOR3_X1   g021(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(KEYINPUT67), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT67), .ZN(new_n225));
  OR2_X1    g024(.A1(G169gat), .A2(G176gat), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n225), .B1(new_n226), .B2(KEYINPUT26), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT66), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n219), .A2(new_n228), .A3(new_n220), .ZN(new_n229));
  NAND4_X1  g028(.A1(new_n222), .A2(new_n224), .A3(new_n227), .A4(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(G183gat), .A2(G190gat), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n218), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT24), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  NOR2_X1   g033(.A1(G183gat), .A2(G190gat), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT64), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND3_X1  g036(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n238));
  OAI21_X1  g037(.A(KEYINPUT64), .B1(G183gat), .B2(G190gat), .ZN(new_n239));
  AND4_X1   g038(.A1(new_n234), .A2(new_n237), .A3(new_n238), .A4(new_n239), .ZN(new_n240));
  NOR2_X1   g039(.A1(G169gat), .A2(G176gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(KEYINPUT23), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT23), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n243), .B1(G169gat), .B2(G176gat), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n242), .A2(new_n220), .A3(new_n244), .ZN(new_n245));
  OAI21_X1  g044(.A(KEYINPUT25), .B1(new_n240), .B2(new_n245), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n245), .A2(KEYINPUT25), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n234), .A2(new_n238), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n247), .B1(new_n248), .B2(new_n235), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n232), .A2(new_n246), .A3(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(G226gat), .A2(G233gat), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n250), .A2(KEYINPUT75), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT75), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n232), .A2(new_n254), .A3(new_n246), .A4(new_n249), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n251), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n257), .A2(KEYINPUT29), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n252), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(G211gat), .ZN(new_n260));
  INV_X1    g059(.A(G218gat), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n260), .A2(new_n261), .A3(KEYINPUT22), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n262), .B1(new_n260), .B2(new_n261), .ZN(new_n263));
  XNOR2_X1  g062(.A(G197gat), .B(G204gat), .ZN(new_n264));
  AND2_X1   g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(KEYINPUT73), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT73), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n264), .A2(KEYINPUT22), .ZN(new_n268));
  XOR2_X1   g067(.A(G211gat), .B(G218gat), .Z(new_n269));
  AOI21_X1  g068(.A(new_n267), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n266), .B1(new_n265), .B2(new_n270), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n271), .B(KEYINPUT74), .ZN(new_n272));
  AOI21_X1  g071(.A(KEYINPUT76), .B1(new_n259), .B2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(new_n258), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n274), .B1(new_n253), .B2(new_n255), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT74), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n271), .B(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT76), .ZN(new_n278));
  NOR4_X1   g077(.A1(new_n275), .A2(new_n277), .A3(new_n278), .A4(new_n252), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n273), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n256), .A2(new_n257), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT29), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n250), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(new_n251), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(KEYINPUT77), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT77), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n283), .A2(new_n286), .A3(new_n251), .ZN(new_n287));
  NAND4_X1  g086(.A1(new_n281), .A2(new_n285), .A3(new_n277), .A4(new_n287), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n206), .B1(new_n280), .B2(new_n288), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n248), .A2(new_n235), .ZN(new_n290));
  NOR3_X1   g089(.A1(new_n290), .A2(KEYINPUT25), .A3(new_n245), .ZN(new_n291));
  INV_X1    g090(.A(new_n231), .ZN(new_n292));
  AND3_X1   g091(.A1(new_n219), .A2(new_n228), .A3(new_n220), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n228), .B1(new_n219), .B2(new_n220), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(new_n223), .B(new_n225), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n292), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n291), .B1(new_n297), .B2(new_n218), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n254), .B1(new_n298), .B2(new_n246), .ZN(new_n299));
  INV_X1    g098(.A(new_n255), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n258), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n252), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n301), .A2(new_n272), .A3(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(new_n278), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n259), .A2(KEYINPUT76), .A3(new_n272), .ZN(new_n305));
  NAND4_X1  g104(.A1(new_n304), .A2(new_n206), .A3(new_n288), .A4(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n205), .B1(new_n289), .B2(new_n307), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n304), .A2(new_n288), .A3(new_n305), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n309), .A2(new_n205), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n202), .B1(new_n308), .B2(new_n311), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n310), .A2(KEYINPUT30), .ZN(new_n313));
  OAI21_X1  g112(.A(KEYINPUT84), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n205), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n309), .A2(KEYINPUT78), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n315), .B1(new_n316), .B2(new_n306), .ZN(new_n317));
  OAI21_X1  g116(.A(KEYINPUT30), .B1(new_n317), .B2(new_n310), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT84), .ZN(new_n319));
  INV_X1    g118(.A(new_n313), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n318), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  XOR2_X1   g120(.A(G127gat), .B(G134gat), .Z(new_n322));
  OR2_X1    g121(.A1(KEYINPUT68), .A2(KEYINPUT1), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  XNOR2_X1  g123(.A(G113gat), .B(G120gat), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n325), .A2(KEYINPUT1), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  OAI211_X1 g126(.A(new_n322), .B(new_n323), .C1(KEYINPUT1), .C2(new_n325), .ZN(new_n328));
  AND2_X1   g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT4), .ZN(new_n330));
  XNOR2_X1  g129(.A(G155gat), .B(G162gat), .ZN(new_n331));
  INV_X1    g130(.A(G155gat), .ZN(new_n332));
  INV_X1    g131(.A(G162gat), .ZN(new_n333));
  OAI21_X1  g132(.A(KEYINPUT2), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(G148gat), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n335), .A2(KEYINPUT79), .A3(G141gat), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n331), .A2(new_n334), .A3(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(G141gat), .B(G148gat), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT79), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  OR2_X1    g140(.A1(new_n339), .A2(KEYINPUT2), .ZN(new_n342));
  XOR2_X1   g141(.A(G155gat), .B(G162gat), .Z(new_n343));
  AOI22_X1  g142(.A1(new_n338), .A2(new_n341), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n329), .A2(new_n330), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n327), .A2(new_n328), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n343), .B1(KEYINPUT2), .B2(new_n339), .ZN(new_n347));
  INV_X1    g146(.A(new_n341), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n347), .B1(new_n348), .B2(new_n337), .ZN(new_n349));
  OAI21_X1  g148(.A(KEYINPUT4), .B1(new_n346), .B2(new_n349), .ZN(new_n350));
  AOI22_X1  g149(.A1(new_n349), .A2(KEYINPUT3), .B1(new_n327), .B2(new_n328), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT3), .ZN(new_n352));
  OAI211_X1 g151(.A(new_n347), .B(new_n352), .C1(new_n348), .C2(new_n337), .ZN(new_n353));
  AOI22_X1  g152(.A1(new_n345), .A2(new_n350), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(G225gat), .A2(G233gat), .ZN(new_n355));
  OR2_X1    g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n355), .ZN(new_n357));
  XNOR2_X1  g156(.A(new_n346), .B(new_n349), .ZN(new_n358));
  OAI211_X1 g157(.A(new_n356), .B(KEYINPUT39), .C1(new_n357), .C2(new_n358), .ZN(new_n359));
  XOR2_X1   g158(.A(G57gat), .B(G85gat), .Z(new_n360));
  XNOR2_X1  g159(.A(G1gat), .B(G29gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n360), .B(new_n361), .ZN(new_n362));
  XNOR2_X1  g161(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n363));
  XNOR2_X1  g162(.A(new_n362), .B(new_n363), .ZN(new_n364));
  OAI211_X1 g163(.A(new_n359), .B(new_n364), .C1(KEYINPUT39), .C2(new_n356), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT40), .ZN(new_n366));
  OR2_X1    g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT5), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n349), .A2(KEYINPUT3), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n369), .A2(new_n346), .A3(new_n353), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n330), .B1(new_n329), .B2(new_n344), .ZN(new_n371));
  NOR3_X1   g170(.A1(new_n346), .A2(new_n349), .A3(KEYINPUT4), .ZN(new_n372));
  OAI211_X1 g171(.A(new_n355), .B(new_n370), .C1(new_n371), .C2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n358), .A2(new_n357), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n368), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  AOI21_X1  g174(.A(KEYINPUT5), .B1(new_n354), .B2(new_n355), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(new_n364), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n365), .A2(new_n366), .ZN(new_n380));
  AND3_X1   g179(.A1(new_n367), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n314), .A2(new_n321), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n353), .A2(new_n282), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n272), .A2(new_n383), .ZN(new_n384));
  AND2_X1   g183(.A1(new_n271), .A2(new_n282), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n349), .B1(new_n385), .B2(KEYINPUT3), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(G228gat), .A2(G233gat), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND4_X1  g188(.A1(new_n384), .A2(G228gat), .A3(G233gat), .A4(new_n386), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(G22gat), .ZN(new_n392));
  INV_X1    g191(.A(G22gat), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n389), .A2(new_n393), .A3(new_n390), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT83), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n392), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  XNOR2_X1  g195(.A(G78gat), .B(G106gat), .ZN(new_n397));
  XNOR2_X1  g196(.A(KEYINPUT31), .B(G50gat), .ZN(new_n398));
  XNOR2_X1  g197(.A(new_n397), .B(new_n398), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n399), .B(KEYINPUT82), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n389), .A2(KEYINPUT83), .A3(new_n393), .A4(new_n390), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n396), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n392), .A2(new_n394), .A3(new_n399), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n316), .A2(KEYINPUT37), .A3(new_n306), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT37), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n309), .A2(new_n407), .ZN(new_n408));
  AND2_X1   g207(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  OAI21_X1  g208(.A(KEYINPUT38), .B1(new_n409), .B2(new_n315), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n364), .B1(new_n375), .B2(new_n376), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT81), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT6), .ZN(new_n414));
  OAI211_X1 g213(.A(KEYINPUT81), .B(new_n364), .C1(new_n375), .C2(new_n376), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n413), .A2(new_n379), .A3(new_n414), .A4(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n377), .A2(KEYINPUT6), .A3(new_n378), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n277), .B1(new_n275), .B2(new_n252), .ZN(new_n419));
  AND3_X1   g218(.A1(new_n281), .A2(new_n285), .A3(new_n287), .ZN(new_n420));
  OAI211_X1 g219(.A(KEYINPUT37), .B(new_n419), .C1(new_n420), .C2(new_n277), .ZN(new_n421));
  AOI21_X1  g220(.A(KEYINPUT38), .B1(new_n408), .B2(new_n421), .ZN(new_n422));
  AOI211_X1 g221(.A(new_n310), .B(new_n418), .C1(new_n422), .C2(new_n205), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n405), .B1(new_n410), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n382), .A2(new_n424), .ZN(new_n425));
  OR3_X1    g224(.A1(new_n250), .A2(KEYINPUT69), .A3(new_n346), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n250), .A2(new_n346), .ZN(new_n427));
  OAI21_X1  g226(.A(KEYINPUT69), .B1(new_n250), .B2(new_n346), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n426), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(G227gat), .A2(G233gat), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(KEYINPUT33), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  XOR2_X1   g231(.A(G71gat), .B(G99gat), .Z(new_n433));
  XNOR2_X1  g232(.A(new_n433), .B(KEYINPUT70), .ZN(new_n434));
  XNOR2_X1  g233(.A(G15gat), .B(G43gat), .ZN(new_n435));
  XNOR2_X1  g234(.A(new_n434), .B(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n432), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n429), .A2(new_n431), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(KEYINPUT32), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  OAI211_X1 g240(.A(KEYINPUT32), .B(new_n439), .C1(new_n432), .C2(new_n437), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND4_X1  g242(.A1(new_n426), .A2(new_n430), .A3(new_n427), .A4(new_n428), .ZN(new_n444));
  XNOR2_X1  g243(.A(KEYINPUT71), .B(KEYINPUT34), .ZN(new_n445));
  XNOR2_X1  g244(.A(new_n444), .B(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n443), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n441), .A2(new_n446), .A3(new_n442), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(KEYINPUT72), .A2(KEYINPUT36), .ZN(new_n451));
  OR2_X1    g250(.A1(KEYINPUT72), .A2(KEYINPUT36), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n450), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n448), .A2(new_n449), .A3(KEYINPUT72), .A4(KEYINPUT36), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n318), .A2(new_n418), .A3(new_n320), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n455), .B1(new_n456), .B2(new_n405), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n425), .A2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT35), .ZN(new_n459));
  AND3_X1   g258(.A1(new_n404), .A2(new_n450), .A3(new_n418), .ZN(new_n460));
  INV_X1    g259(.A(new_n321), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n319), .B1(new_n318), .B2(new_n320), .ZN(new_n462));
  OAI211_X1 g261(.A(new_n459), .B(new_n460), .C1(new_n461), .C2(new_n462), .ZN(new_n463));
  AOI22_X1  g262(.A1(new_n402), .A2(new_n403), .B1(new_n448), .B2(new_n449), .ZN(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  OAI21_X1  g264(.A(KEYINPUT35), .B1(new_n465), .B2(new_n456), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n463), .A2(new_n466), .ZN(new_n467));
  AND2_X1   g266(.A1(new_n458), .A2(new_n467), .ZN(new_n468));
  XNOR2_X1  g267(.A(G15gat), .B(G22gat), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT16), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n469), .B1(new_n470), .B2(G1gat), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n471), .B1(G1gat), .B2(new_n469), .ZN(new_n472));
  INV_X1    g271(.A(G8gat), .ZN(new_n473));
  XNOR2_X1  g272(.A(new_n472), .B(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(G43gat), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(G50gat), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT89), .ZN(new_n477));
  XNOR2_X1  g276(.A(new_n476), .B(new_n477), .ZN(new_n478));
  XNOR2_X1  g277(.A(KEYINPUT88), .B(G43gat), .ZN(new_n479));
  INV_X1    g278(.A(G50gat), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(KEYINPUT15), .B1(new_n478), .B2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT86), .ZN(new_n483));
  OR2_X1    g282(.A1(new_n483), .A2(KEYINPUT14), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(KEYINPUT14), .ZN(new_n485));
  INV_X1    g284(.A(G29gat), .ZN(new_n486));
  INV_X1    g285(.A(G36gat), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n484), .A2(new_n485), .A3(new_n488), .ZN(new_n489));
  OR2_X1    g288(.A1(new_n488), .A2(new_n485), .ZN(new_n490));
  OAI21_X1  g289(.A(KEYINPUT87), .B1(new_n486), .B2(new_n487), .ZN(new_n491));
  OR3_X1    g290(.A1(new_n486), .A2(new_n487), .A3(KEYINPUT87), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n489), .A2(new_n490), .A3(new_n491), .A4(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n476), .A2(KEYINPUT15), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n494), .B1(G43gat), .B2(new_n480), .ZN(new_n495));
  NOR3_X1   g294(.A1(new_n482), .A2(new_n493), .A3(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT90), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n497), .B1(new_n493), .B2(new_n495), .ZN(new_n498));
  OR2_X1    g297(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n496), .A2(KEYINPUT90), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n474), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n499), .A2(new_n500), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(KEYINPUT91), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT17), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n503), .A2(KEYINPUT92), .A3(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT92), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n502), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(KEYINPUT17), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n506), .B1(new_n502), .B2(KEYINPUT91), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n505), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n501), .B1(new_n510), .B2(new_n474), .ZN(new_n511));
  NAND2_X1  g310(.A1(G229gat), .A2(G233gat), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT18), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(new_n474), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n502), .A2(new_n516), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n517), .A2(new_n501), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n512), .B(KEYINPUT13), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n511), .A2(KEYINPUT18), .A3(new_n512), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n515), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  XNOR2_X1  g322(.A(G113gat), .B(G141gat), .ZN(new_n524));
  INV_X1    g323(.A(G197gat), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n524), .B(new_n525), .ZN(new_n526));
  XNOR2_X1  g325(.A(KEYINPUT11), .B(G169gat), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n526), .B(new_n527), .ZN(new_n528));
  XOR2_X1   g327(.A(new_n528), .B(KEYINPUT12), .Z(new_n529));
  AND3_X1   g328(.A1(new_n523), .A2(KEYINPUT85), .A3(new_n529), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n529), .B1(new_n523), .B2(KEYINPUT85), .ZN(new_n531));
  OAI21_X1  g330(.A(KEYINPUT93), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(new_n529), .ZN(new_n533));
  AND3_X1   g332(.A1(new_n511), .A2(KEYINPUT18), .A3(new_n512), .ZN(new_n534));
  AOI21_X1  g333(.A(KEYINPUT18), .B1(new_n511), .B2(new_n512), .ZN(new_n535));
  NOR3_X1   g334(.A1(new_n534), .A2(new_n535), .A3(new_n520), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT85), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n533), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT93), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n523), .A2(KEYINPUT85), .A3(new_n529), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n532), .A2(new_n541), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n468), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(G232gat), .A2(G233gat), .ZN(new_n544));
  XOR2_X1   g343(.A(new_n544), .B(KEYINPUT96), .Z(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  OR2_X1    g345(.A1(new_n546), .A2(KEYINPUT41), .ZN(new_n547));
  XOR2_X1   g346(.A(G190gat), .B(G218gat), .Z(new_n548));
  INV_X1    g347(.A(KEYINPUT99), .ZN(new_n549));
  OR2_X1    g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n547), .B(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  XNOR2_X1  g351(.A(KEYINPUT97), .B(KEYINPUT7), .ZN(new_n553));
  NAND2_X1  g352(.A1(G85gat), .A2(G92gat), .ZN(new_n554));
  OR2_X1    g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(G99gat), .A2(G106gat), .ZN(new_n556));
  INV_X1    g355(.A(G85gat), .ZN(new_n557));
  INV_X1    g356(.A(G92gat), .ZN(new_n558));
  AOI22_X1  g357(.A1(KEYINPUT8), .A2(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n553), .A2(new_n554), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n555), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(G99gat), .B(G106gat), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n561), .B(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n510), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT98), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  AOI22_X1  g366(.A1(new_n502), .A2(new_n563), .B1(KEYINPUT41), .B2(new_n546), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n510), .A2(KEYINPUT98), .A3(new_n564), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n548), .A2(new_n549), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n552), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(G134gat), .B(G162gat), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n570), .A2(new_n552), .A3(new_n571), .ZN(new_n575));
  AND3_X1   g374(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n574), .B1(new_n573), .B2(new_n575), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  AND2_X1   g377(.A1(G71gat), .A2(G78gat), .ZN(new_n579));
  OR2_X1    g378(.A1(new_n579), .A2(KEYINPUT9), .ZN(new_n580));
  XOR2_X1   g379(.A(G57gat), .B(G64gat), .Z(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  XOR2_X1   g381(.A(G71gat), .B(G78gat), .Z(new_n583));
  OR2_X1    g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n582), .A2(new_n583), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  XOR2_X1   g385(.A(new_n586), .B(KEYINPUT94), .Z(new_n587));
  AOI21_X1  g386(.A(new_n516), .B1(new_n587), .B2(KEYINPUT21), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(KEYINPUT95), .ZN(new_n589));
  XOR2_X1   g388(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n590));
  XNOR2_X1  g389(.A(new_n589), .B(new_n590), .ZN(new_n591));
  AOI21_X1  g390(.A(KEYINPUT21), .B1(new_n584), .B2(new_n585), .ZN(new_n592));
  XNOR2_X1  g391(.A(G183gat), .B(G211gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n592), .B(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n591), .B(new_n594), .ZN(new_n595));
  XOR2_X1   g394(.A(G127gat), .B(G155gat), .Z(new_n596));
  NAND2_X1  g395(.A1(G231gat), .A2(G233gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n595), .B(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(G120gat), .B(G148gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(G176gat), .B(G204gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n563), .B(new_n586), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT10), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n587), .A2(KEYINPUT10), .A3(new_n563), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(G230gat), .A2(G233gat), .ZN(new_n608));
  XOR2_X1   g407(.A(new_n608), .B(KEYINPUT100), .Z(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(KEYINPUT101), .ZN(new_n610));
  AND2_X1   g409(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n609), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n603), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n602), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n609), .B1(new_n605), .B2(new_n606), .ZN(new_n615));
  NOR3_X1   g414(.A1(new_n615), .A2(new_n613), .A3(new_n602), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n614), .A2(new_n617), .ZN(new_n618));
  NOR3_X1   g417(.A1(new_n578), .A2(new_n599), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n543), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n620), .B(KEYINPUT102), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n621), .A2(new_n418), .ZN(new_n622));
  XNOR2_X1  g421(.A(KEYINPUT103), .B(G1gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n622), .B(new_n623), .ZN(G1324gat));
  NOR2_X1   g423(.A1(new_n461), .A2(new_n462), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n621), .A2(new_n626), .ZN(new_n627));
  XOR2_X1   g426(.A(KEYINPUT16), .B(G8gat), .Z(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(KEYINPUT42), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n630), .B1(new_n473), .B2(new_n627), .ZN(G1325gat));
  INV_X1    g430(.A(new_n621), .ZN(new_n632));
  AOI21_X1  g431(.A(G15gat), .B1(new_n632), .B2(new_n450), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n455), .A2(G15gat), .ZN(new_n634));
  XOR2_X1   g433(.A(new_n634), .B(KEYINPUT104), .Z(new_n635));
  AOI21_X1  g434(.A(new_n633), .B1(new_n632), .B2(new_n635), .ZN(G1326gat));
  NOR2_X1   g435(.A1(new_n621), .A2(new_n404), .ZN(new_n637));
  XOR2_X1   g436(.A(KEYINPUT43), .B(G22gat), .Z(new_n638));
  XNOR2_X1  g437(.A(new_n637), .B(new_n638), .ZN(G1327gat));
  INV_X1    g438(.A(new_n618), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n578), .A2(new_n599), .A3(new_n640), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n543), .B1(KEYINPUT105), .B2(new_n641), .ZN(new_n642));
  AND2_X1   g441(.A1(new_n641), .A2(KEYINPUT105), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n418), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n644), .A2(new_n486), .A3(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n646), .B(KEYINPUT45), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n599), .A2(new_n640), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n530), .A2(new_n531), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT44), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n578), .A2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT108), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT106), .ZN(new_n654));
  AND3_X1   g453(.A1(new_n425), .A2(new_n654), .A3(new_n457), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n654), .B1(new_n425), .B2(new_n457), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT107), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n467), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n463), .A2(KEYINPUT107), .A3(new_n466), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n653), .B1(new_n657), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n458), .A2(KEYINPUT106), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n425), .A2(new_n654), .A3(new_n457), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  AND3_X1   g464(.A1(new_n463), .A2(KEYINPUT107), .A3(new_n466), .ZN(new_n666));
  AOI21_X1  g465(.A(KEYINPUT107), .B1(new_n463), .B2(new_n466), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n665), .A2(new_n668), .A3(KEYINPUT108), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n652), .B1(new_n662), .B2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n578), .ZN(new_n671));
  OAI21_X1  g470(.A(KEYINPUT44), .B1(new_n468), .B2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n650), .B1(new_n670), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n674), .A2(KEYINPUT109), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT109), .ZN(new_n676));
  OAI211_X1 g475(.A(new_n676), .B(new_n650), .C1(new_n670), .C2(new_n673), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n418), .B1(new_n675), .B2(new_n677), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n647), .B1(new_n678), .B2(new_n486), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT110), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(G1328gat));
  NAND3_X1  g480(.A1(new_n644), .A2(new_n487), .A3(new_n625), .ZN(new_n682));
  XOR2_X1   g481(.A(new_n682), .B(KEYINPUT46), .Z(new_n683));
  AOI21_X1  g482(.A(new_n626), .B1(new_n675), .B2(new_n677), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n683), .B1(new_n684), .B2(new_n487), .ZN(G1329gat));
  OR2_X1    g484(.A1(new_n642), .A2(new_n643), .ZN(new_n686));
  INV_X1    g485(.A(new_n450), .ZN(new_n687));
  NOR3_X1   g486(.A1(new_n686), .A2(new_n687), .A3(new_n479), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n455), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n479), .B1(new_n674), .B2(new_n690), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n689), .A2(KEYINPUT47), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n675), .A2(new_n677), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(new_n455), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n688), .B1(new_n694), .B2(new_n479), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n692), .B1(new_n695), .B2(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g495(.A(KEYINPUT111), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n480), .B1(new_n644), .B2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n404), .B1(new_n644), .B2(new_n697), .ZN(new_n700));
  AOI21_X1  g499(.A(KEYINPUT48), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n404), .B1(new_n675), .B2(new_n677), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n701), .B1(new_n702), .B2(new_n480), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT112), .ZN(new_n704));
  INV_X1    g503(.A(new_n674), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n480), .B1(new_n705), .B2(new_n405), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n405), .B1(new_n686), .B2(KEYINPUT111), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n707), .A2(new_n698), .ZN(new_n708));
  OAI21_X1  g507(.A(KEYINPUT48), .B1(new_n706), .B2(new_n708), .ZN(new_n709));
  AND3_X1   g508(.A1(new_n703), .A2(new_n704), .A3(new_n709), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n704), .B1(new_n703), .B2(new_n709), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n710), .A2(new_n711), .ZN(G1331gat));
  INV_X1    g511(.A(new_n599), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n671), .A2(new_n649), .A3(new_n713), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n714), .A2(new_n640), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(KEYINPUT113), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n662), .A2(new_n669), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(new_n645), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g520(.A1(new_n718), .A2(new_n626), .ZN(new_n722));
  NOR2_X1   g521(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n723));
  AND2_X1   g522(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n722), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n725), .B1(new_n722), .B2(new_n723), .ZN(G1333gat));
  OAI21_X1  g525(.A(G71gat), .B1(new_n718), .B2(new_n690), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n719), .A2(new_n450), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n727), .B1(new_n728), .B2(G71gat), .ZN(new_n729));
  XOR2_X1   g528(.A(new_n729), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g529(.A1(new_n719), .A2(new_n405), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g531(.A1(new_n599), .A2(new_n649), .ZN(new_n733));
  INV_X1    g532(.A(new_n733), .ZN(new_n734));
  OAI211_X1 g533(.A(new_n618), .B(new_n734), .C1(new_n670), .C2(new_n673), .ZN(new_n735));
  NOR3_X1   g534(.A1(new_n735), .A2(new_n557), .A3(new_n418), .ZN(new_n736));
  OAI211_X1 g535(.A(new_n578), .B(new_n734), .C1(new_n657), .C2(new_n661), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(KEYINPUT51), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n738), .A2(new_n640), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(new_n645), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n736), .B1(new_n740), .B2(new_n557), .ZN(G1336gat));
  NOR3_X1   g540(.A1(new_n735), .A2(new_n558), .A3(new_n626), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n739), .A2(new_n625), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n742), .B1(new_n558), .B2(new_n743), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(KEYINPUT52), .ZN(G1337gat));
  XNOR2_X1  g544(.A(KEYINPUT114), .B(G99gat), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n687), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n739), .A2(new_n747), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n746), .B1(new_n735), .B2(new_n690), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(G1338gat));
  INV_X1    g549(.A(G106gat), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n739), .A2(new_n751), .A3(new_n405), .ZN(new_n752));
  OAI21_X1  g551(.A(G106gat), .B1(new_n735), .B2(new_n404), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(KEYINPUT53), .ZN(G1339gat));
  OR3_X1    g554(.A1(new_n607), .A2(KEYINPUT115), .A3(new_n610), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n607), .A2(new_n610), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n615), .A2(KEYINPUT115), .ZN(new_n758));
  OAI211_X1 g557(.A(new_n756), .B(KEYINPUT54), .C1(new_n757), .C2(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(new_n602), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT54), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n760), .B1(new_n611), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n759), .A2(new_n762), .ZN(new_n763));
  OR2_X1    g562(.A1(new_n763), .A2(KEYINPUT55), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(KEYINPUT55), .ZN(new_n765));
  AND2_X1   g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NOR3_X1   g565(.A1(new_n649), .A2(new_n616), .A3(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n518), .A2(new_n519), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n768), .B1(new_n511), .B2(new_n512), .ZN(new_n769));
  AOI22_X1  g568(.A1(new_n536), .A2(new_n533), .B1(new_n528), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(new_n618), .ZN(new_n771));
  INV_X1    g570(.A(new_n771), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n671), .B1(new_n767), .B2(new_n772), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n616), .B1(new_n764), .B2(new_n765), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n578), .A2(new_n774), .A3(new_n770), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n713), .B1(new_n773), .B2(new_n775), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n714), .A2(new_n618), .ZN(new_n777));
  OR2_X1    g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n778), .A2(new_n645), .A3(new_n626), .A4(new_n464), .ZN(new_n779));
  INV_X1    g578(.A(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(G113gat), .ZN(new_n781));
  INV_X1    g580(.A(new_n649), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n780), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  OR2_X1    g582(.A1(new_n779), .A2(new_n542), .ZN(new_n784));
  INV_X1    g583(.A(new_n784), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n783), .B1(new_n785), .B2(new_n781), .ZN(G1340gat));
  NAND2_X1  g585(.A1(new_n780), .A2(new_n618), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n787), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g587(.A1(new_n780), .A2(new_n713), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n789), .B(G127gat), .ZN(G1342gat));
  NAND2_X1  g589(.A1(new_n780), .A2(new_n578), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n791), .A2(G134gat), .ZN(new_n792));
  XNOR2_X1  g591(.A(new_n792), .B(KEYINPUT56), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n791), .A2(G134gat), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(G1343gat));
  OAI21_X1  g594(.A(new_n405), .B1(new_n776), .B2(new_n777), .ZN(new_n796));
  INV_X1    g595(.A(new_n796), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n455), .A2(new_n418), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT117), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  AOI21_X1  g600(.A(KEYINPUT117), .B1(new_n797), .B2(new_n798), .ZN(new_n802));
  NOR3_X1   g601(.A1(new_n801), .A2(new_n625), .A3(new_n802), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n542), .A2(G141gat), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n532), .A2(new_n541), .A3(new_n774), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(new_n771), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(new_n671), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(new_n775), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n777), .B1(new_n809), .B2(new_n599), .ZN(new_n810));
  OAI21_X1  g609(.A(KEYINPUT57), .B1(new_n810), .B2(new_n404), .ZN(new_n811));
  NOR3_X1   g610(.A1(new_n625), .A2(new_n418), .A3(new_n455), .ZN(new_n812));
  OAI211_X1 g611(.A(new_n811), .B(new_n812), .C1(KEYINPUT57), .C2(new_n796), .ZN(new_n813));
  OAI21_X1  g612(.A(G141gat), .B1(new_n813), .B2(new_n542), .ZN(new_n814));
  XOR2_X1   g613(.A(KEYINPUT118), .B(KEYINPUT58), .Z(new_n815));
  NAND3_X1  g614(.A1(new_n805), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n804), .A2(new_n626), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n799), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g617(.A(new_n818), .B(KEYINPUT116), .ZN(new_n819));
  OR2_X1    g618(.A1(new_n813), .A2(new_n649), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n819), .B1(new_n820), .B2(G141gat), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT58), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n816), .B1(new_n821), .B2(new_n822), .ZN(G1344gat));
  NAND3_X1  g622(.A1(new_n803), .A2(new_n335), .A3(new_n618), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT59), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT120), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n808), .A2(new_n826), .A3(new_n775), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n578), .B1(new_n806), .B2(new_n771), .ZN(new_n828));
  INV_X1    g627(.A(new_n775), .ZN(new_n829));
  OAI21_X1  g628(.A(KEYINPUT120), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n827), .A2(new_n599), .A3(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n619), .A2(new_n542), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT57), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n833), .A2(new_n834), .A3(new_n405), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n796), .A2(KEYINPUT57), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(new_n812), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(KEYINPUT119), .ZN(new_n839));
  OR2_X1    g638(.A1(new_n838), .A2(KEYINPUT119), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n837), .A2(new_n618), .A3(new_n839), .A4(new_n840), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n825), .B1(new_n841), .B2(G148gat), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n825), .B1(new_n813), .B2(new_n640), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n843), .A2(new_n335), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n824), .B1(new_n842), .B2(new_n844), .ZN(G1345gat));
  NOR3_X1   g644(.A1(new_n813), .A2(new_n332), .A3(new_n599), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n803), .A2(new_n713), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n846), .B1(new_n847), .B2(new_n332), .ZN(G1346gat));
  NOR3_X1   g647(.A1(new_n813), .A2(new_n333), .A3(new_n671), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n803), .A2(new_n578), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n849), .B1(new_n850), .B2(new_n333), .ZN(G1347gat));
  NOR2_X1   g650(.A1(new_n626), .A2(new_n645), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n778), .A2(new_n464), .A3(new_n852), .ZN(new_n853));
  OAI21_X1  g652(.A(G169gat), .B1(new_n853), .B2(new_n542), .ZN(new_n854));
  OR2_X1    g653(.A1(new_n853), .A2(G169gat), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n854), .B1(new_n855), .B2(new_n649), .ZN(G1348gat));
  NOR2_X1   g655(.A1(new_n853), .A2(new_n640), .ZN(new_n857));
  XOR2_X1   g656(.A(new_n857), .B(G176gat), .Z(G1349gat));
  INV_X1    g657(.A(KEYINPUT121), .ZN(new_n859));
  OR2_X1    g658(.A1(new_n853), .A2(new_n599), .ZN(new_n860));
  INV_X1    g659(.A(new_n216), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n859), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  OR4_X1    g661(.A1(new_n859), .A2(new_n853), .A3(new_n861), .A4(new_n599), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT60), .ZN(new_n865));
  OAI21_X1  g664(.A(KEYINPUT123), .B1(new_n865), .B2(KEYINPUT122), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n865), .A2(KEYINPUT123), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n867), .B1(new_n860), .B2(G183gat), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n864), .A2(new_n866), .A3(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(new_n869), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n866), .B1(new_n864), .B2(new_n868), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n870), .A2(new_n871), .ZN(G1350gat));
  NOR2_X1   g671(.A1(new_n853), .A2(new_n671), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n873), .A2(new_n209), .ZN(new_n874));
  XOR2_X1   g673(.A(new_n874), .B(KEYINPUT61), .Z(new_n875));
  NAND2_X1  g674(.A1(new_n873), .A2(new_n209), .ZN(new_n876));
  XNOR2_X1  g675(.A(new_n876), .B(KEYINPUT124), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n875), .A2(new_n877), .ZN(G1351gat));
  NAND2_X1  g677(.A1(new_n852), .A2(new_n690), .ZN(new_n879));
  INV_X1    g678(.A(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n837), .A2(new_n880), .ZN(new_n881));
  OAI21_X1  g680(.A(G197gat), .B1(new_n881), .B2(new_n542), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n797), .A2(new_n880), .ZN(new_n883));
  INV_X1    g682(.A(new_n883), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n884), .A2(new_n525), .A3(new_n782), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n882), .A2(new_n885), .ZN(G1352gat));
  NOR3_X1   g685(.A1(new_n883), .A2(G204gat), .A3(new_n640), .ZN(new_n887));
  XNOR2_X1  g686(.A(new_n887), .B(KEYINPUT62), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n837), .A2(new_n618), .A3(new_n880), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(G204gat), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n888), .A2(new_n890), .ZN(G1353gat));
  NAND4_X1  g690(.A1(new_n835), .A2(new_n713), .A3(new_n836), .A4(new_n880), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT126), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT63), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n892), .A2(G211gat), .A3(new_n895), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n893), .A2(new_n894), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n713), .A2(new_n260), .ZN(new_n899));
  OR3_X1    g698(.A1(new_n883), .A2(KEYINPUT125), .A3(new_n899), .ZN(new_n900));
  OAI21_X1  g699(.A(KEYINPUT125), .B1(new_n883), .B2(new_n899), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  INV_X1    g701(.A(new_n897), .ZN(new_n903));
  NAND4_X1  g702(.A1(new_n892), .A2(G211gat), .A3(new_n903), .A4(new_n895), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n898), .A2(new_n902), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(KEYINPUT127), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT127), .ZN(new_n907));
  NAND4_X1  g706(.A1(new_n898), .A2(new_n902), .A3(new_n907), .A4(new_n904), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n906), .A2(new_n908), .ZN(G1354gat));
  NOR3_X1   g708(.A1(new_n881), .A2(new_n261), .A3(new_n671), .ZN(new_n910));
  AOI21_X1  g709(.A(G218gat), .B1(new_n884), .B2(new_n578), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n910), .A2(new_n911), .ZN(G1355gat));
endmodule


