//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 1 0 1 0 0 0 0 0 0 1 0 1 1 0 0 0 1 1 0 1 0 0 0 0 0 1 0 1 1 1 1 1 1 0 0 0 1 0 0 1 1 1 0 1 1 1 0 1 1 0 1 1 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:57 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n731, new_n732, new_n733, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n743, new_n744,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n772, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n834,
    new_n836, new_n837, new_n838, new_n840, new_n841, new_n842, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n896, new_n897, new_n898, new_n899, new_n901, new_n902, new_n903,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n955, new_n956, new_n957, new_n958,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n974,
    new_n975, new_n976;
  INV_X1    g000(.A(KEYINPUT18), .ZN(new_n202));
  INV_X1    g001(.A(G1gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(KEYINPUT16), .ZN(new_n204));
  INV_X1    g003(.A(G15gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G22gat), .ZN(new_n206));
  INV_X1    g005(.A(G22gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(G15gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n204), .A2(new_n206), .A3(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  AOI21_X1  g009(.A(G1gat), .B1(new_n206), .B2(new_n208), .ZN(new_n211));
  NOR3_X1   g010(.A1(new_n210), .A2(new_n211), .A3(G8gat), .ZN(new_n212));
  INV_X1    g011(.A(G8gat), .ZN(new_n213));
  INV_X1    g012(.A(new_n211), .ZN(new_n214));
  AOI21_X1  g013(.A(new_n213), .B1(new_n214), .B2(new_n209), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n212), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(new_n216), .ZN(new_n217));
  XOR2_X1   g016(.A(G43gat), .B(G50gat), .Z(new_n218));
  INV_X1    g017(.A(KEYINPUT15), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(G29gat), .ZN(new_n221));
  INV_X1    g020(.A(G36gat), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT14), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n224), .A2(new_n221), .A3(new_n222), .ZN(new_n225));
  OAI21_X1  g024(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n223), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  XNOR2_X1  g026(.A(G43gat), .B(G50gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(KEYINPUT15), .ZN(new_n229));
  AND3_X1   g028(.A1(new_n220), .A2(new_n227), .A3(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT90), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n225), .A2(KEYINPUT89), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT89), .ZN(new_n234));
  NAND4_X1  g033(.A1(new_n234), .A2(new_n224), .A3(new_n221), .A4(new_n222), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n233), .A2(new_n226), .A3(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(new_n223), .ZN(new_n237));
  AOI211_X1 g036(.A(new_n232), .B(new_n229), .C1(new_n236), .C2(new_n237), .ZN(new_n238));
  NOR3_X1   g037(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n226), .B1(new_n239), .B2(new_n234), .ZN(new_n240));
  INV_X1    g039(.A(new_n235), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n237), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(new_n229), .ZN(new_n243));
  AOI21_X1  g042(.A(KEYINPUT90), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n231), .B1(new_n238), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(KEYINPUT17), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n221), .A2(new_n222), .ZN(new_n247));
  AOI22_X1  g046(.A1(new_n225), .A2(KEYINPUT89), .B1(new_n247), .B2(KEYINPUT14), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n223), .B1(new_n248), .B2(new_n235), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n232), .B1(new_n249), .B2(new_n229), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n242), .A2(KEYINPUT90), .A3(new_n243), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT17), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n252), .A2(new_n253), .A3(new_n231), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n217), .B1(new_n246), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n245), .A2(new_n217), .ZN(new_n256));
  NAND2_X1  g055(.A1(G229gat), .A2(G233gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n202), .B1(new_n255), .B2(new_n258), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n253), .B1(new_n252), .B2(new_n231), .ZN(new_n260));
  AOI211_X1 g059(.A(KEYINPUT17), .B(new_n230), .C1(new_n250), .C2(new_n251), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n216), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  AOI22_X1  g061(.A1(new_n245), .A2(new_n217), .B1(G229gat), .B2(G233gat), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n262), .A2(KEYINPUT18), .A3(new_n263), .ZN(new_n264));
  OAI21_X1  g063(.A(KEYINPUT92), .B1(new_n245), .B2(new_n217), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n230), .B1(new_n250), .B2(new_n251), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT92), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n266), .A2(new_n267), .A3(new_n216), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n265), .A2(new_n268), .A3(new_n256), .ZN(new_n269));
  XNOR2_X1  g068(.A(KEYINPUT91), .B(KEYINPUT13), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n270), .B(new_n257), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n259), .A2(new_n264), .A3(new_n272), .ZN(new_n273));
  XNOR2_X1  g072(.A(G113gat), .B(G141gat), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n274), .B(G197gat), .ZN(new_n275));
  XOR2_X1   g074(.A(KEYINPUT11), .B(G169gat), .Z(new_n276));
  XNOR2_X1  g075(.A(new_n275), .B(new_n276), .ZN(new_n277));
  XOR2_X1   g076(.A(new_n277), .B(KEYINPUT12), .Z(new_n278));
  NAND2_X1  g077(.A1(new_n273), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(new_n278), .ZN(new_n280));
  NAND4_X1  g079(.A1(new_n259), .A2(new_n264), .A3(new_n272), .A4(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(G228gat), .A2(G233gat), .ZN(new_n284));
  XNOR2_X1  g083(.A(G197gat), .B(G204gat), .ZN(new_n285));
  XNOR2_X1  g084(.A(KEYINPUT73), .B(G218gat), .ZN(new_n286));
  INV_X1    g085(.A(G211gat), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n285), .B1(new_n288), .B2(KEYINPUT22), .ZN(new_n289));
  XNOR2_X1  g088(.A(G211gat), .B(G218gat), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  OAI211_X1 g091(.A(new_n285), .B(new_n290), .C1(new_n288), .C2(KEYINPUT22), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT3), .ZN(new_n295));
  XNOR2_X1  g094(.A(G155gat), .B(G162gat), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(G141gat), .B(G148gat), .ZN(new_n298));
  XNOR2_X1  g097(.A(KEYINPUT78), .B(KEYINPUT2), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n297), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  XOR2_X1   g099(.A(G141gat), .B(G148gat), .Z(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(KEYINPUT79), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT79), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n298), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n302), .A2(new_n296), .A3(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT2), .ZN(new_n306));
  XNOR2_X1  g105(.A(KEYINPUT80), .B(G155gat), .ZN(new_n307));
  XNOR2_X1  g106(.A(KEYINPUT81), .B(G162gat), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n306), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  OAI211_X1 g108(.A(new_n295), .B(new_n300), .C1(new_n305), .C2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT29), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT85), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n294), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n310), .A2(KEYINPUT85), .A3(new_n311), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n284), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n300), .B1(new_n305), .B2(new_n309), .ZN(new_n317));
  AOI21_X1  g116(.A(KEYINPUT29), .B1(new_n292), .B2(new_n293), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT84), .ZN(new_n319));
  AND2_X1   g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n295), .B1(new_n318), .B2(new_n319), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n317), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n317), .B1(new_n318), .B2(KEYINPUT3), .ZN(new_n323));
  INV_X1    g122(.A(new_n294), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n312), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  XOR2_X1   g125(.A(new_n284), .B(KEYINPUT83), .Z(new_n327));
  AOI22_X1  g126(.A1(new_n316), .A2(new_n322), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT86), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n316), .A2(new_n322), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n326), .A2(new_n327), .ZN(new_n333));
  AOI21_X1  g132(.A(KEYINPUT86), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  XNOR2_X1  g133(.A(G78gat), .B(G106gat), .ZN(new_n335));
  XNOR2_X1  g134(.A(KEYINPUT31), .B(G50gat), .ZN(new_n336));
  XOR2_X1   g135(.A(new_n335), .B(new_n336), .Z(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  OAI21_X1  g137(.A(G22gat), .B1(new_n334), .B2(new_n338), .ZN(new_n339));
  OAI211_X1 g138(.A(new_n207), .B(new_n337), .C1(new_n328), .C2(KEYINPUT86), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n331), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n339), .A2(new_n331), .A3(new_n340), .ZN(new_n343));
  XNOR2_X1  g142(.A(G15gat), .B(G43gat), .ZN(new_n344));
  XNOR2_X1  g143(.A(G71gat), .B(G99gat), .ZN(new_n345));
  XNOR2_X1  g144(.A(new_n344), .B(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(G169gat), .A2(G176gat), .ZN(new_n347));
  INV_X1    g146(.A(G169gat), .ZN(new_n348));
  INV_X1    g147(.A(G176gat), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(KEYINPUT26), .ZN(new_n351));
  NOR3_X1   g150(.A1(new_n350), .A2(KEYINPUT67), .A3(KEYINPUT26), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT67), .ZN(new_n353));
  NOR2_X1   g152(.A1(G169gat), .A2(G176gat), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT26), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n353), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  OAI211_X1 g155(.A(new_n347), .B(new_n351), .C1(new_n352), .C2(new_n356), .ZN(new_n357));
  AND2_X1   g156(.A1(G183gat), .A2(G190gat), .ZN(new_n358));
  XNOR2_X1  g157(.A(KEYINPUT27), .B(G183gat), .ZN(new_n359));
  INV_X1    g158(.A(G190gat), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n358), .B1(new_n361), .B2(KEYINPUT28), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT28), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n359), .A2(new_n363), .A3(new_n360), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n357), .A2(new_n362), .A3(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n354), .B1(KEYINPUT23), .B2(new_n347), .ZN(new_n366));
  AND2_X1   g165(.A1(new_n354), .A2(KEYINPUT23), .ZN(new_n367));
  OR2_X1    g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g167(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n369), .B1(G183gat), .B2(G190gat), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT24), .ZN(new_n371));
  OR2_X1    g170(.A1(new_n371), .A2(KEYINPUT66), .ZN(new_n372));
  AOI22_X1  g171(.A1(new_n371), .A2(KEYINPUT66), .B1(G183gat), .B2(G190gat), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n370), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  OAI21_X1  g173(.A(KEYINPUT25), .B1(new_n368), .B2(new_n374), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n366), .A2(KEYINPUT25), .ZN(new_n376));
  XNOR2_X1  g175(.A(KEYINPUT65), .B(G176gat), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n377), .A2(KEYINPUT23), .A3(new_n348), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT64), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n369), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n369), .A2(new_n379), .ZN(new_n381));
  OAI21_X1  g180(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n381), .B1(new_n383), .B2(new_n358), .ZN(new_n384));
  OAI211_X1 g183(.A(new_n376), .B(new_n378), .C1(new_n380), .C2(new_n384), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n365), .A2(new_n375), .A3(new_n385), .ZN(new_n386));
  XNOR2_X1  g185(.A(G127gat), .B(G134gat), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n387), .B1(KEYINPUT68), .B2(KEYINPUT1), .ZN(new_n388));
  XNOR2_X1  g187(.A(G113gat), .B(G120gat), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n389), .A2(KEYINPUT1), .ZN(new_n390));
  XNOR2_X1  g189(.A(new_n388), .B(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n386), .A2(new_n391), .ZN(new_n392));
  XOR2_X1   g191(.A(new_n388), .B(new_n390), .Z(new_n393));
  NAND4_X1  g192(.A1(new_n393), .A2(new_n365), .A3(new_n375), .A4(new_n385), .ZN(new_n394));
  AND2_X1   g193(.A1(G227gat), .A2(G233gat), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n392), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(KEYINPUT69), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT69), .ZN(new_n398));
  NAND4_X1  g197(.A1(new_n392), .A2(new_n394), .A3(new_n398), .A4(new_n395), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n346), .B1(new_n400), .B2(KEYINPUT32), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT33), .ZN(new_n402));
  AOI21_X1  g201(.A(KEYINPUT70), .B1(new_n400), .B2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT70), .ZN(new_n404));
  AOI211_X1 g203(.A(new_n404), .B(KEYINPUT33), .C1(new_n397), .C2(new_n399), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n401), .B1(new_n403), .B2(new_n405), .ZN(new_n406));
  OAI211_X1 g205(.A(new_n400), .B(KEYINPUT32), .C1(new_n402), .C2(new_n346), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT72), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n395), .B1(new_n392), .B2(new_n394), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT71), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n408), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  OR2_X1    g210(.A1(new_n411), .A2(KEYINPUT34), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n411), .A2(KEYINPUT34), .ZN(new_n413));
  OR2_X1    g212(.A1(new_n409), .A2(new_n408), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n412), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n406), .A2(new_n407), .A3(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n415), .B1(new_n406), .B2(new_n407), .ZN(new_n418));
  OAI211_X1 g217(.A(new_n342), .B(new_n343), .C1(new_n417), .C2(new_n418), .ZN(new_n419));
  XNOR2_X1  g218(.A(G8gat), .B(G36gat), .ZN(new_n420));
  XNOR2_X1  g219(.A(G64gat), .B(G92gat), .ZN(new_n421));
  XNOR2_X1  g220(.A(new_n420), .B(new_n421), .ZN(new_n422));
  XNOR2_X1  g221(.A(KEYINPUT76), .B(KEYINPUT77), .ZN(new_n423));
  XOR2_X1   g222(.A(new_n422), .B(new_n423), .Z(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(G226gat), .ZN(new_n426));
  INV_X1    g225(.A(G233gat), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  AND3_X1   g228(.A1(new_n365), .A2(new_n375), .A3(new_n385), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT74), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n386), .A2(KEYINPUT74), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n428), .A2(KEYINPUT29), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  OAI221_X1 g235(.A(new_n324), .B1(new_n386), .B2(new_n429), .C1(new_n434), .C2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT75), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n429), .B1(new_n432), .B2(new_n433), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n430), .A2(new_n436), .ZN(new_n440));
  OAI211_X1 g239(.A(new_n438), .B(new_n294), .C1(new_n439), .C2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n437), .A2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n440), .ZN(new_n443));
  XNOR2_X1  g242(.A(new_n386), .B(new_n431), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n443), .B1(new_n444), .B2(new_n429), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n438), .B1(new_n445), .B2(new_n294), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n425), .B1(new_n442), .B2(new_n446), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n439), .A2(new_n440), .ZN(new_n448));
  OAI21_X1  g247(.A(KEYINPUT75), .B1(new_n448), .B2(new_n324), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n449), .A2(new_n437), .A3(new_n441), .A4(new_n424), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n447), .A2(new_n450), .A3(KEYINPUT30), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n442), .A2(new_n446), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT30), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n452), .A2(new_n453), .A3(new_n424), .ZN(new_n454));
  NAND2_X1  g253(.A1(G225gat), .A2(G233gat), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  OR2_X1    g255(.A1(new_n305), .A2(new_n309), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n391), .B1(new_n457), .B2(new_n300), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n393), .A2(new_n317), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n456), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(KEYINPUT5), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n317), .A2(KEYINPUT3), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n462), .A2(new_n310), .A3(new_n393), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT4), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n464), .B1(new_n393), .B2(new_n317), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n457), .A2(KEYINPUT4), .A3(new_n300), .A4(new_n391), .ZN(new_n466));
  NAND4_X1  g265(.A1(new_n463), .A2(new_n455), .A3(new_n465), .A4(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n461), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n465), .A2(new_n466), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n470), .A2(KEYINPUT5), .A3(new_n455), .A4(new_n463), .ZN(new_n471));
  XNOR2_X1  g270(.A(G1gat), .B(G29gat), .ZN(new_n472));
  XNOR2_X1  g271(.A(new_n472), .B(KEYINPUT0), .ZN(new_n473));
  XNOR2_X1  g272(.A(G57gat), .B(G85gat), .ZN(new_n474));
  XOR2_X1   g273(.A(new_n473), .B(new_n474), .Z(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n468), .A2(new_n471), .A3(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT6), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n468), .A2(new_n471), .ZN(new_n481));
  AOI21_X1  g280(.A(KEYINPUT6), .B1(new_n481), .B2(new_n475), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n477), .A2(KEYINPUT82), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT82), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n468), .A2(new_n471), .A3(new_n484), .A4(new_n476), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n482), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  AOI22_X1  g285(.A1(new_n451), .A2(new_n454), .B1(new_n480), .B2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  OAI21_X1  g287(.A(KEYINPUT35), .B1(new_n419), .B2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(new_n343), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n490), .A2(new_n341), .ZN(new_n491));
  INV_X1    g290(.A(new_n418), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(new_n416), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n451), .A2(new_n454), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n479), .B1(new_n477), .B2(new_n482), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n495), .A2(KEYINPUT35), .ZN(new_n496));
  NAND4_X1  g295(.A1(new_n491), .A2(new_n493), .A3(new_n494), .A4(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n489), .A2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT36), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n499), .B1(new_n417), .B2(new_n418), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n492), .A2(KEYINPUT36), .A3(new_n416), .ZN(new_n501));
  AND2_X1   g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(new_n477), .ZN(new_n503));
  INV_X1    g302(.A(new_n463), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n456), .B1(new_n504), .B2(new_n469), .ZN(new_n505));
  OR2_X1    g304(.A1(new_n458), .A2(new_n459), .ZN(new_n506));
  OAI211_X1 g305(.A(new_n505), .B(KEYINPUT39), .C1(new_n456), .C2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT39), .ZN(new_n508));
  OAI211_X1 g307(.A(new_n508), .B(new_n456), .C1(new_n504), .C2(new_n469), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT87), .ZN(new_n510));
  AND3_X1   g309(.A1(new_n509), .A2(new_n510), .A3(new_n475), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n510), .B1(new_n509), .B2(new_n475), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n507), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT40), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n503), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  OAI211_X1 g314(.A(KEYINPUT40), .B(new_n507), .C1(new_n511), .C2(new_n512), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n515), .A2(new_n451), .A3(new_n454), .A4(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT88), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n518), .B1(new_n445), .B2(new_n294), .ZN(new_n519));
  OAI22_X1  g318(.A1(new_n434), .A2(new_n436), .B1(new_n386), .B2(new_n429), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(new_n294), .ZN(new_n521));
  INV_X1    g320(.A(new_n439), .ZN(new_n522));
  NAND4_X1  g321(.A1(new_n522), .A2(KEYINPUT88), .A3(new_n324), .A4(new_n443), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n519), .A2(new_n521), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(KEYINPUT37), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT38), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n449), .A2(new_n437), .A3(new_n441), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n425), .B1(new_n528), .B2(KEYINPUT37), .ZN(new_n529));
  OAI211_X1 g328(.A(new_n450), .B(new_n495), .C1(new_n527), .C2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT37), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n424), .B1(new_n452), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n528), .A2(KEYINPUT37), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n526), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  OAI211_X1 g333(.A(new_n491), .B(new_n517), .C1(new_n530), .C2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n342), .A2(new_n343), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n488), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n502), .A2(new_n535), .A3(new_n537), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n283), .B1(new_n498), .B2(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(G190gat), .B(G218gat), .ZN(new_n540));
  XNOR2_X1  g339(.A(G99gat), .B(G106gat), .ZN(new_n541));
  NAND2_X1  g340(.A1(G85gat), .A2(G92gat), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT7), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n545));
  AND2_X1   g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(G99gat), .A2(G106gat), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(KEYINPUT8), .ZN(new_n548));
  INV_X1    g347(.A(G85gat), .ZN(new_n549));
  INV_X1    g348(.A(G92gat), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  AND2_X1   g350(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n541), .B1(new_n546), .B2(new_n552), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n548), .A2(new_n544), .A3(new_n551), .A4(new_n545), .ZN(new_n554));
  INV_X1    g353(.A(new_n541), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n553), .A2(new_n556), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n557), .B1(new_n246), .B2(new_n254), .ZN(new_n558));
  AND2_X1   g357(.A1(G232gat), .A2(G233gat), .ZN(new_n559));
  AOI22_X1  g358(.A1(new_n245), .A2(new_n557), .B1(KEYINPUT41), .B2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n540), .B1(new_n558), .B2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT96), .ZN(new_n563));
  OR2_X1    g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n562), .A2(new_n563), .ZN(new_n565));
  INV_X1    g364(.A(new_n557), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n566), .B1(new_n260), .B2(new_n261), .ZN(new_n567));
  INV_X1    g366(.A(new_n540), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n567), .A2(new_n568), .A3(new_n560), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n559), .A2(KEYINPUT41), .ZN(new_n570));
  XNOR2_X1  g369(.A(G134gat), .B(G162gat), .ZN(new_n571));
  XOR2_X1   g370(.A(new_n570), .B(new_n571), .Z(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  AND2_X1   g372(.A1(new_n569), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n564), .A2(new_n565), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n562), .A2(new_n569), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(new_n572), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n577), .A2(KEYINPUT95), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n573), .B1(new_n562), .B2(new_n569), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT95), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n575), .A2(new_n578), .A3(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(G71gat), .A2(G78gat), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT9), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  OR2_X1    g385(.A1(G57gat), .A2(G64gat), .ZN(new_n587));
  NAND2_X1  g386(.A1(G57gat), .A2(G64gat), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT93), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(G71gat), .B(G78gat), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n589), .A2(new_n590), .A3(new_n592), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n596), .A2(KEYINPUT21), .ZN(new_n597));
  NAND2_X1  g396(.A1(G231gat), .A2(G233gat), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n597), .B(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(G127gat), .B(G155gat), .ZN(new_n600));
  XOR2_X1   g399(.A(new_n600), .B(KEYINPUT20), .Z(new_n601));
  XNOR2_X1  g400(.A(new_n599), .B(new_n601), .ZN(new_n602));
  XOR2_X1   g401(.A(G183gat), .B(G211gat), .Z(new_n603));
  OR2_X1    g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n602), .A2(new_n603), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n217), .B1(KEYINPUT21), .B2(new_n596), .ZN(new_n607));
  XNOR2_X1  g406(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n606), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n604), .A2(new_n609), .A3(new_n605), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n583), .A2(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(G120gat), .B(G148gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(G176gat), .B(G204gat), .ZN(new_n616));
  XOR2_X1   g415(.A(new_n615), .B(new_n616), .Z(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  OAI211_X1 g417(.A(new_n594), .B(new_n595), .C1(new_n553), .C2(new_n556), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n552), .A2(new_n546), .A3(new_n541), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n554), .A2(new_n555), .ZN(new_n621));
  AND3_X1   g420(.A1(new_n589), .A2(new_n590), .A3(new_n592), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n592), .B1(new_n589), .B2(new_n590), .ZN(new_n623));
  OAI211_X1 g422(.A(new_n620), .B(new_n621), .C1(new_n622), .C2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT10), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n619), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n557), .A2(new_n596), .A3(KEYINPUT10), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(G230gat), .A2(G233gat), .ZN(new_n629));
  XOR2_X1   g428(.A(new_n629), .B(KEYINPUT98), .Z(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n628), .A2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT99), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n628), .A2(KEYINPUT99), .A3(new_n631), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n619), .A2(new_n624), .ZN(new_n637));
  INV_X1    g436(.A(new_n629), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n618), .B1(new_n636), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n641), .A2(KEYINPUT100), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT100), .ZN(new_n643));
  OAI211_X1 g442(.A(new_n643), .B(new_n618), .C1(new_n636), .C2(new_n640), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT97), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n628), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n626), .A2(KEYINPUT97), .A3(new_n627), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n647), .A2(new_n648), .A3(new_n629), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n649), .A2(new_n639), .A3(new_n617), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n645), .A2(new_n650), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n614), .A2(new_n651), .ZN(new_n652));
  AND2_X1   g451(.A1(new_n539), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n486), .A2(new_n480), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(G1gat), .ZN(G1324gat));
  INV_X1    g456(.A(new_n494), .ZN(new_n658));
  AND2_X1   g457(.A1(new_n653), .A2(new_n658), .ZN(new_n659));
  XOR2_X1   g458(.A(KEYINPUT16), .B(G8gat), .Z(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n661), .B1(new_n213), .B2(new_n659), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n662), .A2(KEYINPUT42), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT42), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n663), .A2(new_n665), .ZN(G1325gat));
  AOI21_X1  g465(.A(G15gat), .B1(new_n653), .B2(new_n493), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n502), .A2(new_n205), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(KEYINPUT101), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n667), .B1(new_n653), .B2(new_n669), .ZN(G1326gat));
  AND2_X1   g469(.A1(new_n539), .A2(new_n536), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n671), .A2(new_n652), .ZN(new_n672));
  XNOR2_X1  g471(.A(KEYINPUT43), .B(G22gat), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n672), .B(new_n673), .ZN(G1327gat));
  NOR3_X1   g473(.A1(new_n583), .A2(new_n613), .A3(new_n651), .ZN(new_n675));
  AND2_X1   g474(.A1(new_n539), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n676), .A2(new_n221), .A3(new_n655), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(KEYINPUT45), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n498), .A2(new_n538), .ZN(new_n679));
  AND2_X1   g478(.A1(new_n582), .A2(KEYINPUT44), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n613), .B(KEYINPUT103), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  AND3_X1   g482(.A1(new_n279), .A2(KEYINPUT102), .A3(new_n281), .ZN(new_n684));
  AOI21_X1  g483(.A(KEYINPUT102), .B1(new_n279), .B2(new_n281), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NOR3_X1   g485(.A1(new_n683), .A2(new_n651), .A3(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT104), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n488), .A2(new_n536), .A3(new_n688), .ZN(new_n689));
  OAI21_X1  g488(.A(KEYINPUT104), .B1(new_n491), .B2(new_n487), .ZN(new_n690));
  NAND4_X1  g489(.A1(new_n502), .A2(new_n535), .A3(new_n689), .A4(new_n690), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n583), .B1(new_n691), .B2(new_n498), .ZN(new_n692));
  OAI211_X1 g491(.A(new_n681), .B(new_n687), .C1(new_n692), .C2(KEYINPUT44), .ZN(new_n693));
  OAI21_X1  g492(.A(G29gat), .B1(new_n693), .B2(new_n654), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n678), .A2(new_n694), .ZN(G1328gat));
  INV_X1    g494(.A(KEYINPUT106), .ZN(new_n696));
  NAND4_X1  g495(.A1(new_n539), .A2(new_n222), .A3(new_n658), .A4(new_n675), .ZN(new_n697));
  OR2_X1    g496(.A1(new_n697), .A2(KEYINPUT105), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(KEYINPUT105), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n696), .B1(new_n700), .B2(KEYINPUT46), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT46), .ZN(new_n702));
  NAND4_X1  g501(.A1(new_n698), .A2(KEYINPUT106), .A3(new_n702), .A4(new_n699), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  OR2_X1    g503(.A1(new_n693), .A2(new_n494), .ZN(new_n705));
  AOI22_X1  g504(.A1(new_n700), .A2(KEYINPUT46), .B1(new_n705), .B2(G36gat), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n704), .A2(new_n706), .ZN(G1329gat));
  OAI21_X1  g506(.A(G43gat), .B1(new_n693), .B2(new_n502), .ZN(new_n708));
  INV_X1    g507(.A(G43gat), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n676), .A2(new_n709), .A3(new_n493), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g510(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n711), .B(new_n712), .ZN(G1330gat));
  OAI21_X1  g512(.A(G50gat), .B1(new_n693), .B2(new_n491), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT108), .ZN(new_n715));
  AOI21_X1  g514(.A(KEYINPUT48), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(G50gat), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n671), .A2(new_n717), .A3(new_n675), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n714), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n716), .B(new_n719), .ZN(G1331gat));
  INV_X1    g519(.A(KEYINPUT102), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n282), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n279), .A2(KEYINPUT102), .A3(new_n281), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n724), .B1(new_n691), .B2(new_n498), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(new_n651), .ZN(new_n727));
  NOR3_X1   g526(.A1(new_n726), .A2(new_n614), .A3(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(new_n655), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g529(.A1(new_n728), .A2(new_n658), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n731), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n732));
  XOR2_X1   g531(.A(KEYINPUT49), .B(G64gat), .Z(new_n733));
  OAI21_X1  g532(.A(new_n732), .B1(new_n731), .B2(new_n733), .ZN(G1333gat));
  INV_X1    g533(.A(G71gat), .ZN(new_n735));
  AND3_X1   g534(.A1(new_n728), .A2(new_n735), .A3(new_n493), .ZN(new_n736));
  INV_X1    g535(.A(new_n502), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n735), .B1(new_n728), .B2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT50), .ZN(new_n739));
  OR3_X1    g538(.A1(new_n736), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n739), .B1(new_n736), .B2(new_n738), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(new_n741), .ZN(G1334gat));
  NAND2_X1  g541(.A1(new_n728), .A2(new_n536), .ZN(new_n743));
  XNOR2_X1  g542(.A(KEYINPUT109), .B(G78gat), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n743), .B(new_n744), .ZN(G1335gat));
  NOR3_X1   g544(.A1(new_n724), .A2(new_n727), .A3(new_n613), .ZN(new_n746));
  OAI211_X1 g545(.A(new_n681), .B(new_n746), .C1(new_n692), .C2(KEYINPUT44), .ZN(new_n747));
  OAI21_X1  g546(.A(G85gat), .B1(new_n747), .B2(new_n654), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT51), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n583), .A2(new_n613), .ZN(new_n750));
  AND3_X1   g549(.A1(new_n725), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n749), .B1(new_n725), .B2(new_n750), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(new_n753), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n655), .A2(new_n549), .A3(new_n651), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n748), .B1(new_n754), .B2(new_n755), .ZN(G1336gat));
  NOR3_X1   g555(.A1(new_n494), .A2(new_n727), .A3(G92gat), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n753), .A2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT52), .ZN(new_n759));
  OAI21_X1  g558(.A(G92gat), .B1(new_n747), .B2(new_n494), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n758), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n691), .A2(new_n498), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n749), .A2(KEYINPUT110), .ZN(new_n763));
  AND4_X1   g562(.A1(new_n762), .A2(new_n686), .A3(new_n750), .A4(new_n763), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n763), .B1(new_n725), .B2(new_n750), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n757), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n760), .A2(new_n766), .ZN(new_n767));
  AOI21_X1  g566(.A(KEYINPUT111), .B1(new_n767), .B2(KEYINPUT52), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT111), .ZN(new_n769));
  AOI211_X1 g568(.A(new_n769), .B(new_n759), .C1(new_n760), .C2(new_n766), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n761), .B1(new_n768), .B2(new_n770), .ZN(G1337gat));
  OAI21_X1  g570(.A(G99gat), .B1(new_n747), .B2(new_n502), .ZN(new_n772));
  INV_X1    g571(.A(G99gat), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n493), .A2(new_n773), .A3(new_n651), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n772), .B1(new_n754), .B2(new_n774), .ZN(G1338gat));
  OAI21_X1  g574(.A(G106gat), .B1(new_n747), .B2(new_n491), .ZN(new_n776));
  NOR3_X1   g575(.A1(new_n491), .A2(G106gat), .A3(new_n727), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n777), .B1(new_n764), .B2(new_n765), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(KEYINPUT53), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT112), .ZN(new_n781));
  AOI21_X1  g580(.A(KEYINPUT53), .B1(new_n753), .B2(new_n777), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n781), .B1(new_n782), .B2(new_n776), .ZN(new_n783));
  INV_X1    g582(.A(new_n752), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n725), .A2(new_n749), .A3(new_n750), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n784), .A2(new_n785), .A3(new_n777), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT53), .ZN(new_n787));
  AND4_X1   g586(.A1(new_n781), .A2(new_n786), .A3(new_n776), .A4(new_n787), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n780), .B1(new_n783), .B2(new_n788), .ZN(G1339gat));
  NOR3_X1   g588(.A1(new_n614), .A2(new_n651), .A3(new_n724), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT114), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n257), .B1(new_n262), .B2(new_n256), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n269), .A2(new_n271), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n277), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(new_n281), .ZN(new_n795));
  INV_X1    g594(.A(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n582), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n626), .A2(new_n627), .A3(new_n630), .ZN(new_n798));
  AND2_X1   g597(.A1(new_n798), .A2(KEYINPUT54), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n649), .A2(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT54), .ZN(new_n801));
  AOI21_X1  g600(.A(KEYINPUT99), .B1(new_n628), .B2(new_n631), .ZN(new_n802));
  AOI211_X1 g601(.A(new_n633), .B(new_n630), .C1(new_n626), .C2(new_n627), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n801), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n800), .A2(new_n804), .A3(KEYINPUT55), .A4(new_n618), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(new_n650), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(KEYINPUT113), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT113), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n805), .A2(new_n808), .A3(new_n650), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n800), .A2(new_n804), .A3(new_n618), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT55), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n807), .A2(new_n809), .A3(new_n812), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n791), .B1(new_n797), .B2(new_n813), .ZN(new_n814));
  AND3_X1   g613(.A1(new_n805), .A2(new_n808), .A3(new_n650), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n808), .B1(new_n805), .B2(new_n650), .ZN(new_n816));
  AND2_X1   g615(.A1(new_n810), .A2(new_n811), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n815), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n818), .A2(new_n582), .A3(KEYINPUT114), .A4(new_n796), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n814), .A2(new_n819), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n795), .B1(new_n645), .B2(new_n650), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n821), .B1(new_n724), .B2(new_n818), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT115), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n583), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n651), .A2(new_n796), .ZN(new_n825));
  OAI211_X1 g624(.A(new_n825), .B(new_n823), .C1(new_n686), .C2(new_n813), .ZN(new_n826));
  INV_X1    g625(.A(new_n826), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n820), .B1(new_n824), .B2(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n790), .B1(new_n828), .B2(new_n682), .ZN(new_n829));
  NOR4_X1   g628(.A1(new_n829), .A2(new_n654), .A3(new_n658), .A4(new_n419), .ZN(new_n830));
  AOI21_X1  g629(.A(G113gat), .B1(new_n830), .B2(new_n724), .ZN(new_n831));
  AND2_X1   g630(.A1(new_n282), .A2(G113gat), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n831), .B1(new_n830), .B2(new_n832), .ZN(G1340gat));
  NAND2_X1  g632(.A1(new_n830), .A2(new_n651), .ZN(new_n834));
  XNOR2_X1  g633(.A(new_n834), .B(G120gat), .ZN(G1341gat));
  INV_X1    g634(.A(G127gat), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n830), .A2(new_n836), .A3(new_n613), .ZN(new_n837));
  AND2_X1   g636(.A1(new_n830), .A2(new_n683), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n837), .B1(new_n838), .B2(new_n836), .ZN(G1342gat));
  AOI21_X1  g638(.A(new_n583), .B1(KEYINPUT56), .B2(G134gat), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n830), .A2(new_n840), .ZN(new_n841));
  NOR2_X1   g640(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n842));
  XOR2_X1   g641(.A(new_n841), .B(new_n842), .Z(G1343gat));
  INV_X1    g642(.A(KEYINPUT57), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n825), .B1(new_n686), .B2(new_n813), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(KEYINPUT115), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n846), .A2(new_n583), .A3(new_n826), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n683), .B1(new_n847), .B2(new_n820), .ZN(new_n848));
  OAI211_X1 g647(.A(new_n844), .B(new_n536), .C1(new_n848), .C2(new_n790), .ZN(new_n849));
  NOR3_X1   g648(.A1(new_n737), .A2(new_n654), .A3(new_n658), .ZN(new_n850));
  XOR2_X1   g649(.A(KEYINPUT116), .B(KEYINPUT55), .Z(new_n851));
  NAND2_X1  g650(.A1(new_n810), .A2(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT117), .ZN(new_n853));
  NAND4_X1  g652(.A1(new_n852), .A2(new_n853), .A3(new_n650), .A4(new_n805), .ZN(new_n854));
  AND2_X1   g653(.A1(new_n854), .A2(new_n282), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n852), .A2(new_n650), .A3(new_n805), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(KEYINPUT117), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n821), .B1(new_n855), .B2(new_n857), .ZN(new_n858));
  OAI211_X1 g657(.A(new_n814), .B(new_n819), .C1(new_n858), .C2(new_n582), .ZN(new_n859));
  INV_X1    g658(.A(new_n613), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n790), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(KEYINPUT57), .B1(new_n861), .B2(new_n491), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n849), .A2(new_n850), .A3(new_n862), .ZN(new_n863));
  OAI21_X1  g662(.A(G141gat), .B1(new_n863), .B2(new_n283), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT58), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n502), .A2(new_n494), .A3(new_n536), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n283), .A2(G141gat), .ZN(new_n867));
  INV_X1    g666(.A(new_n867), .ZN(new_n868));
  NOR4_X1   g667(.A1(new_n829), .A2(new_n654), .A3(new_n866), .A4(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(new_n869), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n864), .A2(new_n865), .A3(new_n870), .ZN(new_n871));
  NAND4_X1  g670(.A1(new_n849), .A2(new_n724), .A3(new_n850), .A4(new_n862), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(G141gat), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(new_n870), .ZN(new_n874));
  AOI21_X1  g673(.A(KEYINPUT118), .B1(new_n874), .B2(KEYINPUT58), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n869), .B1(new_n872), .B2(G141gat), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT118), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n876), .A2(new_n877), .A3(new_n865), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n871), .B1(new_n875), .B2(new_n878), .ZN(G1344gat));
  NOR3_X1   g678(.A1(new_n829), .A2(new_n654), .A3(new_n866), .ZN(new_n880));
  INV_X1    g679(.A(G148gat), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n880), .A2(new_n881), .A3(new_n651), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT59), .ZN(new_n883));
  OAI21_X1  g682(.A(KEYINPUT57), .B1(new_n829), .B2(new_n491), .ZN(new_n884));
  OR2_X1    g683(.A1(new_n858), .A2(new_n582), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n818), .A2(new_n582), .A3(new_n796), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n613), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n614), .A2(new_n282), .A3(new_n651), .ZN(new_n888));
  OAI211_X1 g687(.A(new_n844), .B(new_n536), .C1(new_n887), .C2(new_n888), .ZN(new_n889));
  AND2_X1   g688(.A1(new_n884), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n890), .A2(new_n651), .A3(new_n850), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n883), .B1(new_n891), .B2(G148gat), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n863), .A2(new_n727), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n893), .A2(KEYINPUT59), .A3(new_n881), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n882), .B1(new_n892), .B2(new_n894), .ZN(G1345gat));
  NAND2_X1  g694(.A1(new_n683), .A2(new_n307), .ZN(new_n896));
  XNOR2_X1  g695(.A(new_n896), .B(KEYINPUT119), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n863), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n307), .B1(new_n880), .B2(new_n613), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n898), .A2(new_n899), .ZN(G1346gat));
  INV_X1    g699(.A(new_n308), .ZN(new_n901));
  NOR3_X1   g700(.A1(new_n863), .A2(new_n901), .A3(new_n583), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n308), .B1(new_n880), .B2(new_n582), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n902), .A2(new_n903), .ZN(G1347gat));
  INV_X1    g703(.A(new_n829), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n658), .A2(new_n654), .ZN(new_n906));
  XNOR2_X1  g705(.A(new_n906), .B(KEYINPUT121), .ZN(new_n907));
  AND3_X1   g706(.A1(new_n907), .A2(new_n491), .A3(new_n493), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n905), .A2(new_n908), .ZN(new_n909));
  OAI21_X1  g708(.A(G169gat), .B1(new_n909), .B2(new_n283), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT120), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n829), .A2(new_n655), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n419), .A2(new_n494), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  INV_X1    g713(.A(new_n914), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n686), .A2(G169gat), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n911), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NOR4_X1   g716(.A1(new_n914), .A2(KEYINPUT120), .A3(G169gat), .A4(new_n686), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n910), .B1(new_n917), .B2(new_n918), .ZN(G1348gat));
  NOR3_X1   g718(.A1(new_n909), .A2(new_n377), .A3(new_n727), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n915), .A2(new_n651), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n920), .B1(new_n921), .B2(new_n349), .ZN(G1349gat));
  OAI211_X1 g721(.A(new_n908), .B(new_n683), .C1(new_n848), .C2(new_n790), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT122), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND4_X1  g724(.A1(new_n905), .A2(KEYINPUT122), .A3(new_n683), .A4(new_n908), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n925), .A2(new_n926), .A3(G183gat), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n613), .A2(new_n359), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n927), .B1(new_n914), .B2(new_n928), .ZN(new_n929));
  XNOR2_X1  g728(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n930));
  INV_X1    g729(.A(new_n930), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  OAI211_X1 g731(.A(new_n927), .B(new_n930), .C1(new_n914), .C2(new_n928), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(G1350gat));
  INV_X1    g733(.A(KEYINPUT124), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n583), .A2(G190gat), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n935), .B1(new_n915), .B2(new_n936), .ZN(new_n937));
  NOR4_X1   g736(.A1(new_n914), .A2(KEYINPUT124), .A3(G190gat), .A4(new_n583), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT61), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n905), .A2(new_n582), .A3(new_n908), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n939), .B1(new_n940), .B2(G190gat), .ZN(new_n941));
  AND3_X1   g740(.A1(new_n940), .A2(new_n939), .A3(G190gat), .ZN(new_n942));
  OAI22_X1  g741(.A1(new_n937), .A2(new_n938), .B1(new_n941), .B2(new_n942), .ZN(G1351gat));
  AND2_X1   g742(.A1(new_n907), .A2(new_n502), .ZN(new_n944));
  AND2_X1   g743(.A1(new_n890), .A2(new_n944), .ZN(new_n945));
  INV_X1    g744(.A(G197gat), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n283), .A2(new_n946), .ZN(new_n947));
  NOR3_X1   g746(.A1(new_n737), .A2(new_n494), .A3(new_n491), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n912), .A2(KEYINPUT125), .A3(new_n948), .ZN(new_n949));
  OAI211_X1 g748(.A(new_n948), .B(new_n654), .C1(new_n848), .C2(new_n790), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT125), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n949), .A2(new_n724), .A3(new_n952), .ZN(new_n953));
  AOI22_X1  g752(.A1(new_n945), .A2(new_n947), .B1(new_n946), .B2(new_n953), .ZN(G1352gat));
  NAND3_X1  g753(.A1(new_n890), .A2(new_n651), .A3(new_n944), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n955), .A2(G204gat), .ZN(new_n956));
  NOR3_X1   g755(.A1(new_n950), .A2(G204gat), .A3(new_n727), .ZN(new_n957));
  XNOR2_X1  g756(.A(new_n957), .B(KEYINPUT62), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n956), .A2(new_n958), .ZN(G1353gat));
  INV_X1    g758(.A(KEYINPUT127), .ZN(new_n960));
  OR2_X1    g759(.A1(new_n960), .A2(KEYINPUT63), .ZN(new_n961));
  NAND4_X1  g760(.A1(new_n884), .A2(new_n889), .A3(new_n613), .A4(new_n944), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n960), .A2(KEYINPUT63), .ZN(new_n963));
  AND3_X1   g762(.A1(new_n962), .A2(G211gat), .A3(new_n963), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n963), .B1(new_n962), .B2(G211gat), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n961), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n860), .A2(G211gat), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n949), .A2(new_n952), .A3(new_n967), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT126), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND4_X1  g769(.A1(new_n949), .A2(KEYINPUT126), .A3(new_n952), .A4(new_n967), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n966), .A2(new_n972), .ZN(G1354gat));
  NOR2_X1   g772(.A1(new_n583), .A2(new_n286), .ZN(new_n974));
  INV_X1    g773(.A(G218gat), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n949), .A2(new_n582), .A3(new_n952), .ZN(new_n976));
  AOI22_X1  g775(.A1(new_n945), .A2(new_n974), .B1(new_n975), .B2(new_n976), .ZN(G1355gat));
endmodule


