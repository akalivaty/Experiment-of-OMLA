//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 0 0 0 0 0 0 1 1 0 1 1 0 1 0 1 0 0 1 0 1 1 0 0 0 0 1 1 0 1 0 0 0 0 0 1 0 0 0 1 0 1 0 0 1 1 0 0 1 1 0 0 0 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:24 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n677, new_n678, new_n679, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n695, new_n696, new_n697, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n729, new_n730, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n890, new_n891,
    new_n892, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  XNOR2_X1  g002(.A(KEYINPUT26), .B(G101), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n189), .B(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT68), .B(G237), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n193), .A2(G953), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G210), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(KEYINPUT70), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT70), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n194), .A2(new_n197), .A3(G210), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n192), .A2(new_n196), .A3(new_n198), .ZN(new_n199));
  AND3_X1   g013(.A1(new_n194), .A2(new_n197), .A3(G210), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n197), .B1(new_n194), .B2(G210), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n191), .B1(new_n200), .B2(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n199), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT71), .ZN(new_n204));
  XNOR2_X1  g018(.A(new_n203), .B(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT28), .ZN(new_n206));
  INV_X1    g020(.A(G146), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G143), .ZN(new_n208));
  INV_X1    g022(.A(G143), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G146), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n208), .A2(KEYINPUT1), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n211), .A2(new_n212), .A3(G128), .ZN(new_n213));
  INV_X1    g027(.A(G128), .ZN(new_n214));
  OAI211_X1 g028(.A(new_n208), .B(new_n210), .C1(KEYINPUT1), .C2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(G137), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n218), .A2(KEYINPUT11), .A3(G134), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT11), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G137), .ZN(new_n221));
  AND2_X1   g035(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  NOR2_X1   g036(.A1(KEYINPUT65), .A2(G134), .ZN(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n218), .A2(KEYINPUT11), .ZN(new_n225));
  NAND2_X1  g039(.A1(KEYINPUT65), .A2(G134), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G131), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n222), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n228), .B1(G134), .B2(G137), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n224), .A2(new_n226), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n230), .B1(new_n231), .B2(G137), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n217), .A2(new_n229), .A3(new_n232), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n220), .A2(G137), .ZN(new_n234));
  AND2_X1   g048(.A1(KEYINPUT65), .A2(G134), .ZN(new_n235));
  NOR3_X1   g049(.A1(new_n234), .A2(new_n235), .A3(new_n223), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n219), .A2(new_n221), .ZN(new_n237));
  OAI21_X1  g051(.A(G131), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(new_n229), .ZN(new_n239));
  AND2_X1   g053(.A1(KEYINPUT0), .A2(G128), .ZN(new_n240));
  XNOR2_X1  g054(.A(G143), .B(G146), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n240), .B1(new_n241), .B2(KEYINPUT64), .ZN(new_n242));
  NOR2_X1   g056(.A1(KEYINPUT0), .A2(G128), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n240), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT64), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n211), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  AND2_X1   g060(.A1(new_n242), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n239), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n233), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(G116), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n250), .A2(G119), .ZN(new_n251));
  INV_X1    g065(.A(G119), .ZN(new_n252));
  OAI21_X1  g066(.A(KEYINPUT66), .B1(new_n252), .B2(G116), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT66), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n254), .A2(new_n250), .A3(G119), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n251), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  XOR2_X1   g070(.A(KEYINPUT2), .B(G113), .Z(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n256), .A2(new_n257), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n206), .B1(new_n249), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n249), .A2(new_n262), .ZN(new_n264));
  AND2_X1   g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  AND3_X1   g079(.A1(new_n217), .A2(new_n229), .A3(new_n232), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT67), .ZN(new_n267));
  NOR3_X1   g081(.A1(new_n236), .A2(G131), .A3(new_n237), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n228), .B1(new_n222), .B2(new_n227), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n242), .A2(new_n246), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n267), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n239), .A2(KEYINPUT67), .A3(new_n247), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n266), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n274), .A2(KEYINPUT28), .A3(new_n261), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n205), .B1(new_n265), .B2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT30), .ZN(new_n278));
  AND3_X1   g092(.A1(new_n233), .A2(new_n248), .A3(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n280), .B1(new_n274), .B2(new_n278), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(new_n262), .ZN(new_n282));
  AND2_X1   g096(.A1(new_n199), .A2(new_n202), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n283), .B1(new_n274), .B2(new_n261), .ZN(new_n284));
  AOI21_X1  g098(.A(KEYINPUT31), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  AND3_X1   g099(.A1(new_n239), .A2(KEYINPUT67), .A3(new_n247), .ZN(new_n286));
  AOI21_X1  g100(.A(KEYINPUT67), .B1(new_n239), .B2(new_n247), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n233), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n279), .B1(new_n288), .B2(KEYINPUT30), .ZN(new_n289));
  OAI211_X1 g103(.A(new_n284), .B(KEYINPUT31), .C1(new_n289), .C2(new_n261), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n277), .B1(new_n285), .B2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT72), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n284), .B1(new_n289), .B2(new_n261), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT31), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(new_n290), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n298), .A2(KEYINPUT72), .A3(new_n277), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n188), .B1(new_n294), .B2(new_n299), .ZN(new_n300));
  OAI21_X1  g114(.A(KEYINPUT73), .B1(new_n300), .B2(KEYINPUT32), .ZN(new_n301));
  INV_X1    g115(.A(G472), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n274), .A2(new_n261), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n282), .A2(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(KEYINPUT29), .B1(new_n304), .B2(new_n283), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n265), .A2(new_n205), .A3(new_n275), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT74), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND4_X1  g122(.A1(new_n265), .A2(new_n205), .A3(KEYINPUT74), .A4(new_n275), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n305), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n288), .A2(new_n262), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n303), .A2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT75), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n313), .A2(new_n314), .A3(KEYINPUT28), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n206), .B1(new_n303), .B2(new_n312), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n263), .A2(KEYINPUT75), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n315), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  AND2_X1   g132(.A1(new_n203), .A2(KEYINPUT29), .ZN(new_n319));
  AOI21_X1  g133(.A(G902), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n302), .B1(new_n311), .B2(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n321), .B1(new_n300), .B2(KEYINPUT32), .ZN(new_n322));
  AOI21_X1  g136(.A(KEYINPUT72), .B1(new_n298), .B2(new_n277), .ZN(new_n323));
  AOI211_X1 g137(.A(new_n293), .B(new_n276), .C1(new_n297), .C2(new_n290), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n187), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT73), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT32), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n325), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n301), .A2(new_n322), .A3(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(G217), .ZN(new_n330));
  INV_X1    g144(.A(G902), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n330), .B1(G234), .B2(new_n331), .ZN(new_n332));
  XNOR2_X1  g146(.A(G125), .B(G140), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(KEYINPUT16), .ZN(new_n334));
  INV_X1    g148(.A(G125), .ZN(new_n335));
  OR3_X1    g149(.A1(new_n335), .A2(KEYINPUT16), .A3(G140), .ZN(new_n336));
  AND3_X1   g150(.A1(new_n334), .A2(G146), .A3(new_n336), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n337), .B1(new_n207), .B2(new_n333), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n214), .A2(G119), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n252), .A2(G128), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  XNOR2_X1  g155(.A(KEYINPUT24), .B(G110), .ZN(new_n342));
  AND2_X1   g156(.A1(new_n342), .A2(KEYINPUT76), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n342), .A2(KEYINPUT76), .ZN(new_n344));
  OAI211_X1 g158(.A(KEYINPUT78), .B(new_n341), .C1(new_n343), .C2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT23), .ZN(new_n346));
  AND2_X1   g160(.A1(new_n346), .A2(KEYINPUT77), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n346), .A2(KEYINPUT77), .ZN(new_n348));
  OAI211_X1 g162(.A(G119), .B(new_n214), .C1(new_n347), .C2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(G110), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n339), .B1(KEYINPUT77), .B2(new_n346), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n349), .A2(new_n350), .A3(new_n340), .A4(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n345), .A2(new_n352), .ZN(new_n353));
  XNOR2_X1  g167(.A(new_n342), .B(KEYINPUT76), .ZN(new_n354));
  AOI21_X1  g168(.A(KEYINPUT78), .B1(new_n354), .B2(new_n341), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n338), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n334), .A2(new_n336), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(new_n207), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n334), .A2(G146), .A3(new_n336), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n349), .A2(new_n340), .A3(new_n351), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(G110), .ZN(new_n362));
  OAI211_X1 g176(.A(new_n360), .B(new_n362), .C1(new_n341), .C2(new_n354), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n356), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT80), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n356), .A2(KEYINPUT80), .A3(new_n363), .ZN(new_n367));
  INV_X1    g181(.A(G953), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n368), .A2(G221), .A3(G234), .ZN(new_n369));
  XNOR2_X1  g183(.A(new_n369), .B(KEYINPUT79), .ZN(new_n370));
  XNOR2_X1  g184(.A(KEYINPUT22), .B(G137), .ZN(new_n371));
  XNOR2_X1  g185(.A(new_n370), .B(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n366), .A2(new_n367), .A3(new_n373), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n364), .A2(new_n365), .A3(new_n372), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  AOI21_X1  g190(.A(KEYINPUT25), .B1(new_n376), .B2(new_n331), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT25), .ZN(new_n378));
  AOI211_X1 g192(.A(new_n378), .B(G902), .C1(new_n374), .C2(new_n375), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n332), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n332), .A2(G902), .ZN(new_n381));
  XNOR2_X1  g195(.A(new_n381), .B(KEYINPUT81), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n376), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n380), .A2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(G210), .B1(G237), .B2(G902), .ZN(new_n386));
  XOR2_X1   g200(.A(new_n386), .B(KEYINPUT89), .Z(new_n387));
  NAND2_X1  g201(.A1(new_n252), .A2(G116), .ZN(new_n388));
  OAI21_X1  g202(.A(G113), .B1(new_n388), .B2(KEYINPUT5), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n389), .B1(new_n256), .B2(KEYINPUT5), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(G104), .ZN(new_n392));
  OAI21_X1  g206(.A(KEYINPUT3), .B1(new_n392), .B2(G107), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT3), .ZN(new_n394));
  INV_X1    g208(.A(G107), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n394), .A2(new_n395), .A3(G104), .ZN(new_n396));
  INV_X1    g210(.A(G101), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n392), .A2(G107), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n393), .A2(new_n396), .A3(new_n397), .A4(new_n398), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n392), .A2(G107), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n395), .A2(G104), .ZN(new_n401));
  OAI21_X1  g215(.A(G101), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n399), .A2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n391), .A2(new_n258), .A3(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n393), .A2(new_n396), .A3(new_n398), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(G101), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT83), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  AND2_X1   g223(.A1(new_n399), .A2(KEYINPUT4), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n406), .A2(KEYINPUT83), .A3(G101), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n409), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT4), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n406), .A2(new_n414), .A3(G101), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n415), .B1(new_n259), .B2(new_n260), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n405), .B1(new_n413), .B2(new_n416), .ZN(new_n417));
  XNOR2_X1  g231(.A(G110), .B(G122), .ZN(new_n418));
  XNOR2_X1  g232(.A(new_n418), .B(KEYINPUT86), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n417), .A2(new_n420), .ZN(new_n421));
  OAI211_X1 g235(.A(new_n405), .B(new_n419), .C1(new_n413), .C2(new_n416), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n421), .A2(KEYINPUT6), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n216), .A2(new_n335), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(KEYINPUT87), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n271), .A2(G125), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT87), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n216), .A2(new_n427), .A3(new_n335), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n425), .A2(new_n426), .A3(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(G224), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n430), .A2(G953), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n429), .B(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT6), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n417), .A2(new_n433), .A3(new_n420), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n423), .A2(new_n432), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(new_n331), .ZN(new_n436));
  AND2_X1   g250(.A1(new_n428), .A2(new_n426), .ZN(new_n437));
  INV_X1    g251(.A(new_n431), .ZN(new_n438));
  NAND4_X1  g252(.A1(new_n437), .A2(KEYINPUT7), .A3(new_n438), .A4(new_n425), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(KEYINPUT7), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n429), .A2(new_n440), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n403), .B1(new_n259), .B2(new_n390), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n405), .A2(new_n442), .ZN(new_n443));
  XNOR2_X1  g257(.A(new_n419), .B(KEYINPUT8), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT88), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n439), .A2(new_n441), .A3(new_n445), .A4(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(new_n422), .ZN(new_n448));
  AOI22_X1  g262(.A1(new_n429), .A2(new_n440), .B1(new_n443), .B2(new_n444), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n446), .B1(new_n449), .B2(new_n439), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n387), .B1(new_n436), .B2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT90), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n439), .A2(new_n441), .A3(new_n445), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(KEYINPUT88), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n455), .A2(new_n422), .A3(new_n447), .ZN(new_n456));
  INV_X1    g270(.A(new_n387), .ZN(new_n457));
  NAND4_X1  g271(.A1(new_n456), .A2(new_n331), .A3(new_n457), .A4(new_n435), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n452), .A2(new_n453), .A3(new_n458), .ZN(new_n459));
  OAI211_X1 g273(.A(KEYINPUT90), .B(new_n387), .C1(new_n436), .C2(new_n451), .ZN(new_n460));
  OAI21_X1  g274(.A(G214), .B1(G237), .B2(G902), .ZN(new_n461));
  XNOR2_X1  g275(.A(new_n461), .B(KEYINPUT85), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n459), .A2(new_n460), .A3(new_n463), .ZN(new_n464));
  XNOR2_X1  g278(.A(KEYINPUT9), .B(G234), .ZN(new_n465));
  OAI21_X1  g279(.A(G221), .B1(new_n465), .B2(G902), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n466), .B(KEYINPUT82), .ZN(new_n467));
  INV_X1    g281(.A(G469), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n468), .A2(new_n331), .ZN(new_n469));
  NAND4_X1  g283(.A1(new_n213), .A2(new_n215), .A3(new_n399), .A4(new_n402), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n470), .B(KEYINPUT10), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n412), .A2(new_n247), .A3(new_n415), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n471), .A2(new_n472), .A3(new_n270), .ZN(new_n473));
  XNOR2_X1  g287(.A(G110), .B(G140), .ZN(new_n474));
  INV_X1    g288(.A(G227), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n475), .A2(G953), .ZN(new_n476));
  XNOR2_X1  g290(.A(new_n474), .B(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n473), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n270), .B1(new_n471), .B2(new_n472), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  OR2_X1    g295(.A1(KEYINPUT84), .A2(KEYINPUT12), .ZN(new_n482));
  INV_X1    g296(.A(new_n470), .ZN(new_n483));
  AOI22_X1  g297(.A1(new_n213), .A2(new_n215), .B1(new_n399), .B2(new_n402), .ZN(new_n484));
  OAI211_X1 g298(.A(new_n239), .B(new_n482), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n216), .A2(new_n403), .ZN(new_n486));
  AOI22_X1  g300(.A1(new_n486), .A2(new_n470), .B1(new_n229), .B2(new_n238), .ZN(new_n487));
  XOR2_X1   g301(.A(KEYINPUT84), .B(KEYINPUT12), .Z(new_n488));
  OAI21_X1  g302(.A(new_n485), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n478), .B1(new_n473), .B2(new_n489), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n481), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n469), .B1(new_n491), .B2(G469), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n471), .A2(new_n472), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(new_n239), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n478), .B1(new_n494), .B2(new_n473), .ZN(new_n495));
  AND3_X1   g309(.A1(new_n473), .A2(new_n489), .A3(new_n478), .ZN(new_n496));
  OAI211_X1 g310(.A(new_n468), .B(new_n331), .C1(new_n495), .C2(new_n496), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n467), .B1(new_n492), .B2(new_n497), .ZN(new_n498));
  OR2_X1    g312(.A1(new_n333), .A2(KEYINPUT19), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n333), .A2(KEYINPUT19), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(new_n207), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(KEYINPUT92), .ZN(new_n503));
  AOI21_X1  g317(.A(G146), .B1(new_n499), .B2(new_n500), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT92), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n337), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  XOR2_X1   g320(.A(KEYINPUT68), .B(G237), .Z(new_n507));
  NAND3_X1  g321(.A1(new_n507), .A2(G214), .A3(new_n368), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(new_n209), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n194), .A2(G143), .A3(G214), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n509), .A2(new_n228), .A3(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n228), .B1(new_n509), .B2(new_n510), .ZN(new_n513));
  OAI211_X1 g327(.A(new_n503), .B(new_n506), .C1(new_n512), .C2(new_n513), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n508), .A2(new_n209), .ZN(new_n515));
  AOI21_X1  g329(.A(G143), .B1(new_n194), .B2(G214), .ZN(new_n516));
  OAI211_X1 g330(.A(KEYINPUT18), .B(G131), .C1(new_n515), .C2(new_n516), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n333), .B(new_n207), .ZN(new_n518));
  NAND2_X1  g332(.A1(KEYINPUT18), .A2(G131), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n509), .A2(new_n510), .A3(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n517), .A2(new_n518), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n514), .A2(new_n521), .ZN(new_n522));
  XNOR2_X1  g336(.A(G113), .B(G122), .ZN(new_n523));
  XNOR2_X1  g337(.A(new_n523), .B(new_n392), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n522), .A2(new_n525), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n360), .B1(new_n513), .B2(KEYINPUT17), .ZN(new_n527));
  OAI21_X1  g341(.A(G131), .B1(new_n515), .B2(new_n516), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(new_n511), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n527), .B1(new_n529), .B2(KEYINPUT17), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n530), .A2(new_n524), .A3(new_n521), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n526), .A2(new_n531), .ZN(new_n532));
  NOR2_X1   g346(.A1(G475), .A2(G902), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  XNOR2_X1  g348(.A(KEYINPUT91), .B(KEYINPUT20), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT20), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n532), .A2(new_n538), .A3(new_n533), .ZN(new_n539));
  INV_X1    g353(.A(new_n531), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n524), .B1(new_n530), .B2(new_n521), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n331), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  XOR2_X1   g356(.A(KEYINPUT93), .B(G475), .Z(new_n543));
  AOI22_X1  g357(.A1(new_n537), .A2(new_n539), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  XNOR2_X1  g358(.A(G116), .B(G122), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n545), .B(new_n395), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n209), .A2(G128), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT13), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n214), .A2(G143), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n547), .A2(new_n548), .ZN(new_n552));
  OAI21_X1  g366(.A(G134), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n547), .A2(new_n550), .ZN(new_n554));
  OAI211_X1 g368(.A(new_n546), .B(new_n553), .C1(new_n231), .C2(new_n554), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n231), .B(new_n554), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n545), .A2(new_n395), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n250), .A2(KEYINPUT14), .A3(G122), .ZN(new_n558));
  INV_X1    g372(.A(new_n545), .ZN(new_n559));
  OAI211_X1 g373(.A(G107), .B(new_n558), .C1(new_n559), .C2(KEYINPUT14), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n556), .A2(new_n557), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n555), .A2(new_n561), .ZN(new_n562));
  NOR3_X1   g376(.A1(new_n465), .A2(new_n330), .A3(G953), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n563), .B1(new_n555), .B2(new_n561), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n567), .A2(G902), .ZN(new_n568));
  INV_X1    g382(.A(G478), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n569), .A2(KEYINPUT15), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n568), .B(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(G234), .A2(G237), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n573), .A2(G952), .A3(new_n368), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n573), .A2(G902), .A3(G953), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  XNOR2_X1  g391(.A(KEYINPUT21), .B(G898), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n575), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n572), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n498), .A2(new_n544), .A3(new_n580), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n464), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n329), .A2(new_n385), .A3(new_n582), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n583), .B(G101), .ZN(G3));
  OAI21_X1  g398(.A(new_n331), .B1(new_n323), .B2(new_n324), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(G472), .ZN(new_n586));
  INV_X1    g400(.A(new_n498), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n384), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n586), .A2(new_n325), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(KEYINPUT94), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n300), .B1(new_n585), .B2(G472), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT94), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n591), .A2(new_n592), .A3(new_n588), .ZN(new_n593));
  INV_X1    g407(.A(new_n461), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n594), .B1(new_n452), .B2(new_n458), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n533), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n597), .B1(new_n526), .B2(new_n531), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n539), .B1(new_n535), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n542), .A2(new_n543), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  AOI21_X1  g415(.A(KEYINPUT95), .B1(new_n555), .B2(new_n561), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT33), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n567), .A2(new_n604), .ZN(new_n605));
  OAI22_X1  g419(.A1(new_n565), .A2(new_n566), .B1(new_n603), .B2(new_n602), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n605), .A2(new_n606), .A3(G478), .A4(new_n331), .ZN(new_n607));
  XOR2_X1   g421(.A(KEYINPUT96), .B(G478), .Z(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n609), .B1(new_n567), .B2(G902), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n601), .A2(new_n611), .ZN(new_n612));
  NOR3_X1   g426(.A1(new_n596), .A2(new_n612), .A3(new_n579), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n590), .A2(new_n593), .A3(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n614), .B(G104), .ZN(new_n615));
  XOR2_X1   g429(.A(KEYINPUT97), .B(KEYINPUT34), .Z(new_n616));
  XNOR2_X1  g430(.A(new_n615), .B(new_n616), .ZN(G6));
  AOI21_X1  g431(.A(KEYINPUT98), .B1(new_n534), .B2(new_n536), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n618), .B1(new_n536), .B2(new_n534), .ZN(new_n619));
  AND2_X1   g433(.A1(new_n572), .A2(new_n600), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n598), .A2(KEYINPUT98), .A3(new_n535), .ZN(new_n621));
  AND3_X1   g435(.A1(new_n619), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT100), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n579), .B(KEYINPUT99), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n622), .A2(new_n623), .A3(new_n595), .A4(new_n624), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n619), .A2(new_n620), .A3(new_n624), .A4(new_n621), .ZN(new_n626));
  OAI21_X1  g440(.A(KEYINPUT100), .B1(new_n626), .B2(new_n596), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n590), .A2(new_n593), .A3(new_n628), .ZN(new_n629));
  XOR2_X1   g443(.A(KEYINPUT35), .B(G107), .Z(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(G9));
  INV_X1    g445(.A(KEYINPUT101), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n364), .B(new_n632), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n373), .A2(KEYINPUT36), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(new_n382), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n380), .A2(new_n636), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n582), .A2(new_n586), .A3(new_n325), .A4(new_n637), .ZN(new_n638));
  XOR2_X1   g452(.A(KEYINPUT37), .B(G110), .Z(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G12));
  NOR2_X1   g454(.A1(new_n534), .A2(new_n536), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n618), .B(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(new_n620), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n637), .A2(new_n595), .ZN(new_n644));
  XNOR2_X1  g458(.A(KEYINPUT102), .B(G900), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n577), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(new_n574), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  NOR4_X1   g462(.A1(new_n643), .A2(new_n644), .A3(new_n587), .A4(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(new_n329), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(G128), .ZN(G30));
  XNOR2_X1  g465(.A(new_n568), .B(new_n570), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n652), .B1(new_n599), .B2(new_n600), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n653), .A2(new_n461), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT40), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n647), .B(KEYINPUT39), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n498), .A2(KEYINPUT104), .A3(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  AOI21_X1  g472(.A(KEYINPUT104), .B1(new_n498), .B2(new_n656), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n655), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(new_n659), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n661), .A2(KEYINPUT40), .A3(new_n657), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n654), .B1(new_n660), .B2(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(new_n637), .ZN(new_n664));
  INV_X1    g478(.A(new_n205), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(new_n313), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(new_n295), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n302), .B1(new_n667), .B2(new_n331), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n668), .B1(new_n300), .B2(KEYINPUT32), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n301), .A2(new_n669), .A3(new_n328), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n459), .A2(new_n460), .ZN(new_n671));
  XNOR2_X1  g485(.A(KEYINPUT103), .B(KEYINPUT38), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n663), .A2(new_n664), .A3(new_n670), .A4(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G143), .ZN(G45));
  AND2_X1   g490(.A1(new_n607), .A2(new_n610), .ZN(new_n677));
  NOR3_X1   g491(.A1(new_n544), .A2(new_n677), .A3(new_n648), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n679), .A2(new_n644), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n329), .A2(new_n498), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G146), .ZN(G48));
  OAI21_X1  g496(.A(new_n331), .B1(new_n495), .B2(new_n496), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(G469), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(new_n497), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n685), .A2(new_n467), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n329), .A2(new_n385), .A3(new_n613), .A4(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT105), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(KEYINPUT41), .B(G113), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n689), .B(new_n690), .ZN(G15));
  NAND4_X1  g505(.A1(new_n329), .A2(new_n628), .A3(new_n385), .A4(new_n686), .ZN(new_n692));
  XOR2_X1   g506(.A(KEYINPUT106), .B(G116), .Z(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(G18));
  NAND3_X1  g508(.A1(new_n686), .A2(new_n544), .A3(new_n580), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n644), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n329), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G119), .ZN(G21));
  AND4_X1   g512(.A1(new_n595), .A2(new_n686), .A3(new_n653), .A4(new_n624), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n318), .A2(KEYINPUT107), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT107), .ZN(new_n701));
  OAI211_X1 g515(.A(new_n315), .B(new_n701), .C1(new_n316), .C2(new_n317), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n700), .A2(new_n665), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(new_n298), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(new_n187), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n699), .A2(new_n586), .A3(new_n705), .A4(new_n385), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G122), .ZN(G24));
  NAND2_X1  g521(.A1(new_n586), .A2(new_n705), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n708), .A2(new_n664), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n595), .A2(new_n686), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n679), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G125), .ZN(G27));
  XNOR2_X1  g527(.A(new_n498), .B(KEYINPUT108), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n671), .A2(new_n461), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n329), .A2(new_n385), .A3(new_n678), .A4(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT42), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n325), .A2(new_n327), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n384), .B1(new_n322), .B2(new_n720), .ZN(new_n721));
  NOR3_X1   g535(.A1(new_n714), .A2(new_n679), .A3(new_n715), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n721), .A2(new_n722), .A3(KEYINPUT42), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n719), .A2(KEYINPUT109), .A3(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(new_n724), .ZN(new_n725));
  AOI21_X1  g539(.A(KEYINPUT109), .B1(new_n719), .B2(new_n723), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G131), .ZN(G33));
  NOR2_X1   g542(.A1(new_n643), .A2(new_n648), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n329), .A2(new_n385), .A3(new_n729), .A4(new_n716), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G134), .ZN(G36));
  INV_X1    g545(.A(KEYINPUT44), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT43), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n544), .A2(new_n733), .A3(new_n611), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n599), .A2(new_n600), .A3(new_n611), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(KEYINPUT43), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n734), .A2(new_n736), .A3(new_n637), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n732), .B1(new_n591), .B2(new_n737), .ZN(new_n738));
  AND3_X1   g552(.A1(new_n734), .A2(new_n736), .A3(new_n637), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n294), .A2(new_n299), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n302), .B1(new_n740), .B2(new_n331), .ZN(new_n741));
  OAI211_X1 g555(.A(new_n739), .B(KEYINPUT44), .C1(new_n300), .C2(new_n741), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n594), .B1(new_n459), .B2(new_n460), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n738), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT111), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(new_n656), .ZN(new_n747));
  INV_X1    g561(.A(new_n497), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT45), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n749), .B1(new_n481), .B2(new_n490), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n473), .A2(new_n489), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(new_n477), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n494), .A2(new_n478), .A3(new_n473), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n752), .A2(new_n753), .A3(KEYINPUT45), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n750), .A2(G469), .A3(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT110), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n752), .A2(new_n753), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n468), .B1(new_n758), .B2(new_n749), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n759), .A2(KEYINPUT110), .A3(new_n754), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n469), .B1(new_n757), .B2(new_n760), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n748), .B1(new_n761), .B2(KEYINPUT46), .ZN(new_n762));
  AOI21_X1  g576(.A(KEYINPUT110), .B1(new_n759), .B2(new_n754), .ZN(new_n763));
  AND4_X1   g577(.A1(KEYINPUT110), .A2(new_n750), .A3(G469), .A4(new_n754), .ZN(new_n764));
  OAI22_X1  g578(.A1(new_n763), .A2(new_n764), .B1(new_n468), .B2(new_n331), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT46), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  AOI211_X1 g581(.A(new_n467), .B(new_n747), .C1(new_n762), .C2(new_n767), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n738), .A2(new_n742), .A3(KEYINPUT111), .A4(new_n743), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n746), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G137), .ZN(G39));
  AND3_X1   g585(.A1(new_n743), .A2(new_n384), .A3(new_n678), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n772), .A2(new_n301), .A3(new_n322), .A4(new_n328), .ZN(new_n773));
  INV_X1    g587(.A(new_n467), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n497), .B1(new_n765), .B2(new_n766), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n761), .A2(KEYINPUT46), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n774), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT47), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  OAI211_X1 g593(.A(KEYINPUT47), .B(new_n774), .C1(new_n775), .C2(new_n776), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n773), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  XOR2_X1   g595(.A(new_n781), .B(G140), .Z(G42));
  NAND3_X1  g596(.A1(new_n385), .A2(new_n463), .A3(new_n774), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(KEYINPUT112), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n685), .B(KEYINPUT49), .ZN(new_n785));
  OR2_X1    g599(.A1(new_n785), .A2(new_n735), .ZN(new_n786));
  OR4_X1    g600(.A1(new_n670), .A2(new_n784), .A3(new_n674), .A4(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT54), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n459), .A2(new_n460), .A3(new_n463), .A4(new_n624), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n789), .A2(new_n612), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n590), .A2(new_n593), .A3(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT113), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n791), .A2(new_n583), .A3(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n544), .A2(new_n572), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n789), .A2(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n590), .A2(new_n593), .A3(new_n795), .ZN(new_n796));
  AND2_X1   g610(.A1(new_n638), .A2(new_n706), .ZN(new_n797));
  AND4_X1   g611(.A1(new_n692), .A2(new_n796), .A3(new_n697), .A4(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n791), .A2(new_n583), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(KEYINPUT113), .ZN(new_n800));
  AND4_X1   g614(.A1(new_n689), .A2(new_n793), .A3(new_n798), .A4(new_n800), .ZN(new_n801));
  AOI22_X1  g615(.A1(new_n709), .A2(new_n711), .B1(new_n649), .B2(new_n329), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n595), .A2(new_n653), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n587), .A2(new_n648), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n670), .A2(new_n664), .A3(new_n803), .A4(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n802), .A2(new_n681), .A3(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT52), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n802), .A2(KEYINPUT52), .A3(new_n681), .A4(new_n805), .ZN(new_n809));
  AND3_X1   g623(.A1(new_n652), .A2(new_n600), .A3(new_n647), .ZN(new_n810));
  AND4_X1   g624(.A1(new_n642), .A2(new_n743), .A3(new_n637), .A4(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n329), .A2(new_n498), .A3(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n709), .A2(new_n722), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT114), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n730), .A2(new_n812), .A3(new_n813), .A4(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n730), .A2(new_n813), .A3(new_n812), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(KEYINPUT114), .ZN(new_n817));
  AOI22_X1  g631(.A1(new_n808), .A2(new_n809), .B1(new_n815), .B2(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n801), .A2(new_n818), .A3(new_n727), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT53), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n820), .B1(new_n802), .B2(new_n807), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n801), .A2(new_n818), .A3(new_n822), .A4(new_n727), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n788), .B1(new_n821), .B2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT115), .ZN(new_n825));
  OAI21_X1  g639(.A(KEYINPUT53), .B1(new_n802), .B2(new_n807), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n826), .B1(new_n719), .B2(new_n723), .ZN(new_n827));
  AND2_X1   g641(.A1(new_n818), .A2(new_n827), .ZN(new_n828));
  AOI22_X1  g642(.A1(new_n801), .A2(new_n828), .B1(new_n819), .B2(new_n820), .ZN(new_n829));
  AOI22_X1  g643(.A1(new_n824), .A2(new_n825), .B1(new_n829), .B2(new_n788), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n821), .A2(new_n823), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n831), .A2(KEYINPUT54), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n832), .A2(KEYINPUT115), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n734), .A2(new_n736), .ZN(new_n834));
  INV_X1    g648(.A(new_n834), .ZN(new_n835));
  AND3_X1   g649(.A1(new_n743), .A2(new_n575), .A3(new_n686), .ZN(new_n836));
  AND3_X1   g650(.A1(new_n709), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  NOR4_X1   g651(.A1(new_n708), .A2(new_n384), .A3(new_n574), .A4(new_n834), .ZN(new_n838));
  INV_X1    g652(.A(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n673), .A2(new_n594), .A3(new_n686), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  OR2_X1    g655(.A1(new_n841), .A2(KEYINPUT50), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(KEYINPUT50), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n837), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n779), .A2(new_n780), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n685), .A2(new_n774), .ZN(new_n846));
  OAI211_X1 g660(.A(new_n838), .B(new_n743), .C1(new_n845), .C2(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n836), .A2(new_n385), .ZN(new_n848));
  OR2_X1    g662(.A1(new_n848), .A2(new_n670), .ZN(new_n849));
  XNOR2_X1  g663(.A(new_n849), .B(KEYINPUT116), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n544), .A2(new_n677), .ZN(new_n851));
  OAI211_X1 g665(.A(new_n844), .B(new_n847), .C1(new_n850), .C2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT51), .ZN(new_n853));
  AND2_X1   g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n852), .A2(new_n853), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n850), .A2(new_n612), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n721), .A2(new_n835), .A3(new_n836), .ZN(new_n857));
  XOR2_X1   g671(.A(KEYINPUT117), .B(KEYINPUT48), .Z(new_n858));
  NOR2_X1   g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n857), .A2(new_n858), .ZN(new_n860));
  OAI211_X1 g674(.A(G952), .B(new_n368), .C1(new_n839), .C2(new_n710), .ZN(new_n861));
  OR4_X1    g675(.A1(new_n856), .A2(new_n859), .A3(new_n860), .A4(new_n861), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n854), .A2(new_n855), .A3(new_n862), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n830), .A2(new_n833), .A3(new_n863), .ZN(new_n864));
  NOR2_X1   g678(.A1(G952), .A2(G953), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n787), .B1(new_n864), .B2(new_n865), .ZN(G75));
  NOR2_X1   g680(.A1(new_n368), .A2(G952), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT56), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n801), .A2(new_n818), .A3(new_n827), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n821), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n870), .A2(G902), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n868), .B1(new_n871), .B2(new_n457), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n423), .A2(new_n434), .ZN(new_n873));
  XNOR2_X1  g687(.A(new_n873), .B(new_n432), .ZN(new_n874));
  XNOR2_X1  g688(.A(KEYINPUT118), .B(KEYINPUT55), .ZN(new_n875));
  XOR2_X1   g689(.A(new_n874), .B(new_n875), .Z(new_n876));
  INV_X1    g690(.A(new_n876), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n867), .B1(new_n872), .B2(new_n877), .ZN(new_n878));
  OAI211_X1 g692(.A(new_n868), .B(new_n876), .C1(new_n871), .C2(new_n457), .ZN(new_n879));
  AND2_X1   g693(.A1(new_n878), .A2(new_n879), .ZN(G51));
  XNOR2_X1  g694(.A(new_n469), .B(KEYINPUT119), .ZN(new_n881));
  XOR2_X1   g695(.A(new_n881), .B(KEYINPUT57), .Z(new_n882));
  NOR2_X1   g696(.A1(new_n870), .A2(KEYINPUT54), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n788), .B1(new_n821), .B2(new_n869), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n882), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n885), .B1(new_n495), .B2(new_n496), .ZN(new_n886));
  INV_X1    g700(.A(new_n871), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n887), .A2(new_n757), .A3(new_n760), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n867), .B1(new_n886), .B2(new_n888), .ZN(G54));
  AND2_X1   g703(.A1(KEYINPUT58), .A2(G475), .ZN(new_n890));
  AND3_X1   g704(.A1(new_n887), .A2(new_n532), .A3(new_n890), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n532), .B1(new_n887), .B2(new_n890), .ZN(new_n892));
  NOR3_X1   g706(.A1(new_n891), .A2(new_n892), .A3(new_n867), .ZN(G60));
  NAND2_X1  g707(.A1(new_n605), .A2(new_n606), .ZN(new_n894));
  XOR2_X1   g708(.A(new_n894), .B(KEYINPUT120), .Z(new_n895));
  NAND2_X1  g709(.A1(G478), .A2(G902), .ZN(new_n896));
  XOR2_X1   g710(.A(new_n896), .B(KEYINPUT59), .Z(new_n897));
  NOR2_X1   g711(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n898), .B1(new_n883), .B2(new_n884), .ZN(new_n899));
  INV_X1    g713(.A(new_n867), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n830), .A2(new_n833), .ZN(new_n902));
  INV_X1    g716(.A(new_n897), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n901), .B1(new_n904), .B2(new_n895), .ZN(G63));
  NAND2_X1  g719(.A1(G217), .A2(G902), .ZN(new_n906));
  XOR2_X1   g720(.A(new_n906), .B(KEYINPUT60), .Z(new_n907));
  NAND2_X1  g721(.A1(new_n870), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n908), .A2(new_n375), .A3(new_n374), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n870), .A2(new_n635), .A3(new_n907), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n909), .A2(new_n900), .A3(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT61), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n909), .A2(KEYINPUT61), .A3(new_n900), .A4(new_n910), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n913), .A2(new_n914), .ZN(G66));
  OAI21_X1  g729(.A(G953), .B1(new_n578), .B2(new_n430), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n916), .B1(new_n801), .B2(G953), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n873), .B1(G898), .B2(new_n368), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n917), .B(new_n918), .ZN(G69));
  XNOR2_X1  g733(.A(new_n289), .B(new_n501), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n920), .B1(G900), .B2(G953), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n681), .A2(new_n712), .A3(new_n650), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n768), .A2(new_n721), .A3(new_n803), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(new_n730), .ZN(new_n924));
  NOR3_X1   g738(.A1(new_n922), .A2(new_n924), .A3(new_n781), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n719), .A2(new_n723), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT109), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n925), .A2(new_n928), .A3(new_n724), .A4(new_n770), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n921), .B1(new_n929), .B2(G953), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n802), .A2(new_n675), .A3(new_n681), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(KEYINPUT62), .ZN(new_n932));
  AND2_X1   g746(.A1(new_n794), .A2(new_n612), .ZN(new_n933));
  NOR3_X1   g747(.A1(new_n933), .A2(new_n659), .A3(new_n658), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n329), .A2(new_n385), .A3(new_n743), .A4(new_n934), .ZN(new_n935));
  OR2_X1    g749(.A1(new_n935), .A2(KEYINPUT121), .ZN(new_n936));
  INV_X1    g750(.A(new_n781), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n935), .A2(KEYINPUT121), .ZN(new_n938));
  AND3_X1   g752(.A1(new_n936), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n939), .A2(new_n770), .ZN(new_n940));
  OAI21_X1  g754(.A(KEYINPUT122), .B1(new_n932), .B2(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT62), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n931), .B(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT122), .ZN(new_n944));
  NAND4_X1  g758(.A1(new_n943), .A2(new_n944), .A3(new_n770), .A4(new_n939), .ZN(new_n945));
  AOI21_X1  g759(.A(G953), .B1(new_n941), .B2(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(new_n920), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n930), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  AND2_X1   g762(.A1(new_n947), .A2(KEYINPUT123), .ZN(new_n949));
  AOI211_X1 g763(.A(new_n368), .B(new_n949), .C1(G227), .C2(G900), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n948), .B(new_n950), .ZN(G72));
  NAND3_X1  g765(.A1(new_n941), .A2(new_n945), .A3(new_n801), .ZN(new_n952));
  NAND2_X1  g766(.A1(G472), .A2(G902), .ZN(new_n953));
  XOR2_X1   g767(.A(new_n953), .B(KEYINPUT63), .Z(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(KEYINPUT124), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n952), .A2(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n283), .B1(new_n282), .B2(new_n303), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n304), .A2(new_n203), .ZN(new_n958));
  INV_X1    g772(.A(new_n954), .ZN(new_n959));
  NOR3_X1   g773(.A1(new_n958), .A2(new_n959), .A3(new_n957), .ZN(new_n960));
  AOI22_X1  g774(.A1(new_n956), .A2(new_n957), .B1(new_n831), .B2(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT125), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n689), .A2(new_n798), .A3(new_n793), .A4(new_n800), .ZN(new_n963));
  OAI211_X1 g777(.A(new_n962), .B(new_n955), .C1(new_n929), .C2(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(new_n958), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n922), .A2(new_n781), .ZN(new_n966));
  INV_X1    g780(.A(new_n924), .ZN(new_n967));
  AND3_X1   g781(.A1(new_n966), .A2(new_n770), .A3(new_n967), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n801), .A2(new_n727), .A3(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n962), .B1(new_n969), .B2(new_n955), .ZN(new_n970));
  OAI211_X1 g784(.A(KEYINPUT126), .B(new_n900), .C1(new_n965), .C2(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(new_n971), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n955), .B1(new_n929), .B2(new_n963), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n973), .A2(KEYINPUT125), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n974), .A2(new_n958), .A3(new_n964), .ZN(new_n975));
  AOI21_X1  g789(.A(KEYINPUT126), .B1(new_n975), .B2(new_n900), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n961), .B1(new_n972), .B2(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT127), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  OAI211_X1 g793(.A(KEYINPUT127), .B(new_n961), .C1(new_n972), .C2(new_n976), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n979), .A2(new_n980), .ZN(G57));
endmodule


