//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 0 1 0 0 0 0 0 0 1 0 0 1 0 1 0 1 0 1 1 1 1 1 0 1 1 0 0 0 0 0 1 0 0 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:08 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n722, new_n723, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n741, new_n742, new_n743,
    new_n744, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n758, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n904, new_n905,
    new_n906, new_n907, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n926, new_n927, new_n928, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987;
  INV_X1    g000(.A(G475), .ZN(new_n187));
  XNOR2_X1  g001(.A(G113), .B(G122), .ZN(new_n188));
  INV_X1    g002(.A(G104), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n188), .B(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G237), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT70), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n193), .A2(G953), .ZN(new_n194));
  INV_X1    g008(.A(G953), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n195), .A2(KEYINPUT70), .ZN(new_n196));
  OAI211_X1 g010(.A(G214), .B(new_n192), .C1(new_n194), .C2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G143), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n195), .A2(KEYINPUT70), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n193), .A2(G953), .ZN(new_n201));
  AOI21_X1  g015(.A(G237), .B1(new_n200), .B2(new_n201), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n202), .A2(G143), .A3(G214), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n199), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G131), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT17), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT89), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n209), .B1(new_n204), .B2(G131), .ZN(new_n210));
  AOI211_X1 g024(.A(KEYINPUT89), .B(new_n206), .C1(new_n199), .C2(new_n203), .ZN(new_n211));
  OAI211_X1 g025(.A(new_n207), .B(new_n208), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n210), .A2(new_n211), .ZN(new_n213));
  AOI22_X1  g027(.A1(new_n212), .A2(KEYINPUT92), .B1(new_n213), .B2(KEYINPUT17), .ZN(new_n214));
  INV_X1    g028(.A(G140), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G125), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n216), .A2(KEYINPUT16), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n215), .A2(KEYINPUT76), .A3(G125), .ZN(new_n219));
  INV_X1    g033(.A(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT76), .ZN(new_n221));
  XNOR2_X1  g035(.A(G125), .B(G140), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n220), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT16), .ZN(new_n224));
  OAI211_X1 g038(.A(G146), .B(new_n218), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(G146), .ZN(new_n226));
  INV_X1    g040(.A(G125), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(G140), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n216), .A2(new_n228), .A3(new_n221), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n224), .B1(new_n229), .B2(new_n219), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n226), .B1(new_n230), .B2(new_n217), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n225), .A2(new_n231), .A3(KEYINPUT77), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT77), .ZN(new_n233));
  OAI211_X1 g047(.A(new_n233), .B(new_n226), .C1(new_n230), .C2(new_n217), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(KEYINPUT91), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT91), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n232), .A2(new_n237), .A3(new_n234), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT92), .ZN(new_n240));
  NOR4_X1   g054(.A1(new_n210), .A2(new_n211), .A3(new_n240), .A4(new_n208), .ZN(new_n241));
  NOR3_X1   g055(.A1(new_n214), .A2(new_n239), .A3(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT18), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n205), .B1(new_n243), .B2(new_n206), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n222), .A2(new_n226), .ZN(new_n245));
  INV_X1    g059(.A(new_n223), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n245), .B1(new_n246), .B2(new_n226), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n200), .A2(new_n201), .ZN(new_n248));
  AND4_X1   g062(.A1(G143), .A2(new_n248), .A3(G214), .A4(new_n192), .ZN(new_n249));
  AOI21_X1  g063(.A(G143), .B1(new_n202), .B2(G214), .ZN(new_n250));
  OAI21_X1  g064(.A(G131), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  OAI211_X1 g065(.A(new_n244), .B(new_n247), .C1(new_n243), .C2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(new_n252), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n191), .B1(new_n242), .B2(new_n253), .ZN(new_n254));
  NOR3_X1   g068(.A1(new_n210), .A2(new_n211), .A3(new_n208), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(KEYINPUT92), .ZN(new_n256));
  AND3_X1   g070(.A1(new_n232), .A2(new_n237), .A3(new_n234), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n237), .B1(new_n232), .B2(new_n234), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n204), .A2(G131), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n251), .A2(KEYINPUT89), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n204), .A2(new_n209), .A3(G131), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n260), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n240), .B1(new_n263), .B2(new_n208), .ZN(new_n264));
  OAI211_X1 g078(.A(new_n256), .B(new_n259), .C1(new_n264), .C2(new_n255), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n265), .A2(new_n190), .A3(new_n252), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n254), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(G902), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n187), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n223), .A2(KEYINPUT19), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT19), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n222), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  MUX2_X1   g087(.A(new_n270), .B(new_n273), .S(KEYINPUT90), .Z(new_n274));
  OAI21_X1  g088(.A(new_n225), .B1(new_n274), .B2(G146), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n252), .B1(new_n275), .B2(new_n263), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(new_n191), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n266), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n278), .A2(new_n187), .A3(new_n268), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(KEYINPUT20), .ZN(new_n280));
  AOI21_X1  g094(.A(G475), .B1(new_n266), .B2(new_n277), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT20), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n281), .A2(new_n282), .A3(new_n268), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n269), .B1(new_n280), .B2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(G478), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n285), .A2(KEYINPUT15), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  XNOR2_X1  g101(.A(KEYINPUT9), .B(G234), .ZN(new_n288));
  XOR2_X1   g102(.A(new_n288), .B(KEYINPUT79), .Z(new_n289));
  INV_X1    g103(.A(G217), .ZN(new_n290));
  NOR3_X1   g104(.A1(new_n289), .A2(new_n290), .A3(G953), .ZN(new_n291));
  XOR2_X1   g105(.A(KEYINPUT68), .B(G116), .Z(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(G122), .ZN(new_n293));
  INV_X1    g107(.A(G122), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(G116), .ZN(new_n295));
  AND3_X1   g109(.A1(new_n293), .A2(KEYINPUT93), .A3(new_n295), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n293), .A2(KEYINPUT93), .ZN(new_n297));
  OAI21_X1  g111(.A(G107), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  OR2_X1    g112(.A1(new_n293), .A2(KEYINPUT93), .ZN(new_n299));
  INV_X1    g113(.A(G107), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n293), .A2(KEYINPUT93), .A3(new_n295), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n299), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  XNOR2_X1  g116(.A(KEYINPUT65), .B(G128), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n303), .A2(new_n198), .ZN(new_n304));
  OAI21_X1  g118(.A(G134), .B1(new_n304), .B2(KEYINPUT13), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n198), .A2(G128), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n306), .B1(new_n303), .B2(new_n198), .ZN(new_n307));
  AND2_X1   g121(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n305), .A2(new_n307), .ZN(new_n309));
  OAI211_X1 g123(.A(new_n298), .B(new_n302), .C1(new_n308), .C2(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n300), .B1(new_n295), .B2(KEYINPUT14), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n312), .B1(new_n296), .B2(new_n297), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n299), .A2(new_n301), .A3(new_n311), .ZN(new_n314));
  INV_X1    g128(.A(G134), .ZN(new_n315));
  OR2_X1    g129(.A1(new_n307), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n307), .A2(new_n315), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n313), .A2(new_n314), .A3(new_n316), .A4(new_n317), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n291), .B1(new_n310), .B2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n310), .A2(new_n318), .A3(new_n291), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n287), .B1(new_n322), .B2(new_n268), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n322), .A2(new_n268), .A3(new_n287), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  XNOR2_X1  g141(.A(KEYINPUT70), .B(G953), .ZN(new_n328));
  NAND2_X1  g142(.A1(G234), .A2(G237), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n328), .A2(G902), .A3(new_n329), .ZN(new_n330));
  XNOR2_X1  g144(.A(new_n330), .B(KEYINPUT95), .ZN(new_n331));
  XNOR2_X1  g145(.A(KEYINPUT21), .B(G898), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  XNOR2_X1  g147(.A(KEYINPUT94), .B(G952), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n334), .A2(G953), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(new_n329), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n333), .A2(new_n336), .ZN(new_n337));
  XOR2_X1   g151(.A(new_n337), .B(KEYINPUT96), .Z(new_n338));
  NAND3_X1  g152(.A1(new_n284), .A2(new_n327), .A3(new_n338), .ZN(new_n339));
  OAI21_X1  g153(.A(KEYINPUT3), .B1(new_n189), .B2(G107), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT3), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n341), .A2(new_n300), .A3(G104), .ZN(new_n342));
  INV_X1    g156(.A(G101), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n189), .A2(G107), .ZN(new_n344));
  NAND4_X1  g158(.A1(new_n340), .A2(new_n342), .A3(new_n343), .A4(new_n344), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n300), .A2(G104), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n189), .A2(G107), .ZN(new_n347));
  OAI21_X1  g161(.A(G101), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  XNOR2_X1  g163(.A(new_n349), .B(KEYINPUT83), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n226), .A2(G143), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n198), .A2(G146), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(G128), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(KEYINPUT65), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT65), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(G128), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT1), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n359), .B1(G143), .B2(new_n226), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n353), .B1(new_n358), .B2(new_n360), .ZN(new_n361));
  XNOR2_X1  g175(.A(G143), .B(G146), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n362), .A2(new_n359), .A3(G128), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n350), .A2(KEYINPUT10), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n315), .A2(G137), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT11), .ZN(new_n367));
  INV_X1    g181(.A(G137), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n367), .B1(G134), .B2(new_n368), .ZN(new_n369));
  NOR3_X1   g183(.A1(new_n315), .A2(KEYINPUT11), .A3(G137), .ZN(new_n370));
  OAI211_X1 g184(.A(new_n206), .B(new_n366), .C1(new_n369), .C2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  OAI21_X1  g186(.A(KEYINPUT11), .B1(new_n315), .B2(G137), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n367), .A2(new_n368), .A3(G134), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n206), .B1(new_n375), .B2(new_n366), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n372), .A2(new_n376), .ZN(new_n377));
  AND2_X1   g191(.A1(new_n345), .A2(new_n348), .ZN(new_n378));
  AND4_X1   g192(.A1(new_n359), .A2(new_n351), .A3(new_n352), .A4(G128), .ZN(new_n379));
  OAI21_X1  g193(.A(KEYINPUT1), .B1(new_n198), .B2(G146), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n362), .B1(G128), .B2(new_n380), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n378), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT10), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n340), .A2(new_n342), .A3(new_n344), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(G101), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n386), .A2(KEYINPUT82), .A3(KEYINPUT4), .A4(new_n345), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT0), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n388), .A2(new_n354), .ZN(new_n389));
  NOR2_X1   g203(.A1(KEYINPUT0), .A2(G128), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n353), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n362), .B1(new_n388), .B2(new_n354), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(KEYINPUT82), .A2(KEYINPUT4), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n385), .A2(G101), .A3(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n387), .A2(new_n393), .A3(new_n395), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n365), .A2(new_n377), .A3(new_n384), .A4(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n248), .A2(G227), .ZN(new_n398));
  XNOR2_X1  g212(.A(new_n398), .B(new_n215), .ZN(new_n399));
  XNOR2_X1  g213(.A(KEYINPUT81), .B(G110), .ZN(new_n400));
  XNOR2_X1  g214(.A(new_n399), .B(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n397), .A2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT85), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n349), .A2(new_n361), .A3(new_n363), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n382), .A2(KEYINPUT84), .A3(new_n405), .ZN(new_n406));
  OR2_X1    g220(.A1(new_n405), .A2(KEYINPUT84), .ZN(new_n407));
  INV_X1    g221(.A(new_n377), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT12), .ZN(new_n410));
  OR2_X1    g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n409), .A2(new_n410), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n397), .A2(KEYINPUT85), .A3(new_n401), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n404), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(new_n401), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n365), .A2(new_n384), .A3(new_n396), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(new_n408), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(new_n397), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n416), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n415), .A2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(G469), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n422), .A2(new_n423), .A3(new_n268), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n413), .A2(new_n397), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(new_n416), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n419), .A2(new_n402), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n426), .A2(G469), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(G469), .A2(G902), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n424), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(new_n289), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(new_n268), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(G221), .ZN(new_n434));
  XNOR2_X1  g248(.A(new_n434), .B(KEYINPUT80), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n431), .A2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT69), .ZN(new_n437));
  INV_X1    g251(.A(G119), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(G116), .ZN(new_n439));
  XNOR2_X1  g253(.A(KEYINPUT68), .B(G116), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n439), .B1(new_n440), .B2(new_n438), .ZN(new_n441));
  XNOR2_X1  g255(.A(KEYINPUT2), .B(G113), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n437), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n292), .A2(G119), .ZN(new_n444));
  INV_X1    g258(.A(new_n442), .ZN(new_n445));
  NAND4_X1  g259(.A1(new_n444), .A2(KEYINPUT69), .A3(new_n439), .A4(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n443), .A2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT5), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n448), .A2(new_n438), .A3(G116), .ZN(new_n449));
  OAI211_X1 g263(.A(G113), .B(new_n449), .C1(new_n441), .C2(new_n448), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n447), .A2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT83), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n349), .B(new_n452), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n442), .B(KEYINPUT67), .ZN(new_n454));
  AOI22_X1  g268(.A1(new_n443), .A2(new_n446), .B1(new_n454), .B2(new_n441), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n387), .A2(new_n395), .ZN(new_n456));
  OAI22_X1  g270(.A1(new_n451), .A2(new_n453), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  XOR2_X1   g271(.A(G110), .B(G122), .Z(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(new_n458), .ZN(new_n460));
  OAI221_X1 g274(.A(new_n460), .B1(new_n455), .B2(new_n456), .C1(new_n451), .C2(new_n453), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n459), .A2(new_n461), .A3(KEYINPUT6), .ZN(new_n462));
  INV_X1    g276(.A(G224), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n463), .A2(G953), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n391), .A2(new_n392), .A3(G125), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n466), .B1(new_n364), .B2(G125), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(KEYINPUT86), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT86), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n465), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n468), .A2(new_n465), .A3(new_n470), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n472), .A2(KEYINPUT87), .A3(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT87), .ZN(new_n475));
  INV_X1    g289(.A(new_n473), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n475), .B1(new_n476), .B2(new_n471), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT6), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n457), .A2(new_n478), .A3(new_n458), .ZN(new_n479));
  NAND4_X1  g293(.A1(new_n462), .A2(new_n474), .A3(new_n477), .A4(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n476), .A2(KEYINPUT7), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT7), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n467), .B1(new_n482), .B2(new_n464), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n451), .A2(new_n378), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n458), .A2(KEYINPUT8), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n447), .A2(new_n349), .A3(new_n450), .ZN(new_n486));
  OR2_X1    g300(.A1(new_n458), .A2(KEYINPUT8), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n484), .A2(new_n485), .A3(new_n486), .A4(new_n487), .ZN(new_n488));
  NAND4_X1  g302(.A1(new_n481), .A2(new_n461), .A3(new_n483), .A4(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n480), .A2(new_n268), .A3(new_n489), .ZN(new_n490));
  OAI21_X1  g304(.A(G210), .B1(G237), .B2(G902), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n480), .A2(new_n268), .A3(new_n491), .A4(new_n489), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n493), .A2(KEYINPUT88), .A3(new_n494), .ZN(new_n495));
  OAI21_X1  g309(.A(G214), .B1(G237), .B2(G902), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT88), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n490), .A2(new_n497), .A3(new_n492), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n495), .A2(new_n496), .A3(new_n498), .ZN(new_n499));
  NOR3_X1   g313(.A1(new_n339), .A2(new_n436), .A3(new_n499), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n303), .A2(new_n438), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n501), .B1(new_n438), .B2(G128), .ZN(new_n502));
  XOR2_X1   g316(.A(KEYINPUT24), .B(G110), .Z(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n501), .A2(KEYINPUT23), .ZN(new_n505));
  OAI21_X1  g319(.A(KEYINPUT23), .B1(new_n354), .B2(G119), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(KEYINPUT75), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT75), .ZN(new_n508));
  OAI211_X1 g322(.A(new_n508), .B(KEYINPUT23), .C1(new_n354), .C2(G119), .ZN(new_n509));
  OAI211_X1 g323(.A(new_n507), .B(new_n509), .C1(new_n438), .C2(G128), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n505), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(G110), .ZN(new_n512));
  NAND4_X1  g326(.A1(new_n232), .A2(new_n234), .A3(new_n504), .A4(new_n512), .ZN(new_n513));
  OAI22_X1  g327(.A1(new_n511), .A2(G110), .B1(new_n502), .B2(new_n503), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n514), .A2(new_n225), .A3(new_n245), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n248), .A2(G221), .A3(G234), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n517), .B(G137), .ZN(new_n518));
  XNOR2_X1  g332(.A(KEYINPUT78), .B(KEYINPUT22), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n518), .B(new_n519), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n516), .B(new_n520), .ZN(new_n521));
  OR3_X1    g335(.A1(new_n521), .A2(KEYINPUT25), .A3(G902), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n290), .B1(G234), .B2(new_n268), .ZN(new_n523));
  OAI21_X1  g337(.A(KEYINPUT25), .B1(new_n521), .B2(G902), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  OR3_X1    g339(.A1(new_n521), .A2(G902), .A3(new_n523), .ZN(new_n526));
  AND2_X1   g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  NOR2_X1   g342(.A1(G472), .A2(G902), .ZN(new_n529));
  XNOR2_X1  g343(.A(new_n529), .B(KEYINPUT74), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n454), .A2(new_n441), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n447), .A2(new_n532), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n393), .B1(new_n372), .B2(new_n376), .ZN(new_n534));
  OAI21_X1  g348(.A(KEYINPUT64), .B1(new_n368), .B2(G134), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT64), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n536), .A2(new_n315), .A3(G137), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n368), .A2(G134), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n535), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(G131), .ZN(new_n540));
  AOI22_X1  g354(.A1(new_n303), .A2(new_n380), .B1(new_n351), .B2(new_n352), .ZN(new_n541));
  OAI211_X1 g355(.A(new_n540), .B(new_n371), .C1(new_n541), .C2(new_n379), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n534), .A2(KEYINPUT30), .A3(new_n542), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n366), .B1(new_n369), .B2(new_n370), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(G131), .ZN(new_n545));
  AOI22_X1  g359(.A1(new_n545), .A2(new_n371), .B1(new_n391), .B2(new_n392), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n542), .A2(KEYINPUT66), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT66), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n364), .A2(new_n548), .A3(new_n371), .A4(new_n540), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n546), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  OAI211_X1 g364(.A(new_n533), .B(new_n543), .C1(new_n550), .C2(KEYINPUT30), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n455), .A2(new_n534), .A3(new_n542), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n202), .A2(G210), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n553), .B(G101), .ZN(new_n554));
  XNOR2_X1  g368(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n554), .B(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n551), .A2(new_n552), .A3(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT71), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n551), .A2(KEYINPUT71), .A3(new_n552), .A4(new_n556), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(KEYINPUT31), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n557), .A2(KEYINPUT31), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(KEYINPUT72), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT31), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n566), .B1(new_n559), .B2(new_n560), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT72), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT28), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n534), .A2(new_n542), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n569), .B1(new_n533), .B2(new_n570), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n455), .A2(KEYINPUT28), .A3(new_n534), .A4(new_n542), .ZN(new_n572));
  OAI211_X1 g386(.A(new_n571), .B(new_n572), .C1(new_n455), .C2(new_n550), .ZN(new_n573));
  INV_X1    g387(.A(new_n556), .ZN(new_n574));
  AOI21_X1  g388(.A(KEYINPUT73), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  AND3_X1   g389(.A1(new_n573), .A2(KEYINPUT73), .A3(new_n574), .ZN(new_n576));
  OAI22_X1  g390(.A1(new_n567), .A2(new_n568), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n531), .B1(new_n565), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(KEYINPUT32), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n576), .A2(new_n575), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n580), .B1(new_n562), .B2(KEYINPUT72), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n568), .B1(new_n567), .B2(new_n563), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT32), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n583), .A2(new_n584), .A3(new_n531), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n579), .A2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(G472), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n551), .A2(new_n552), .ZN(new_n588));
  AOI21_X1  g402(.A(KEYINPUT29), .B1(new_n588), .B2(new_n574), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n589), .B1(new_n574), .B2(new_n573), .ZN(new_n590));
  AND2_X1   g404(.A1(new_n571), .A2(new_n572), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n533), .A2(new_n570), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n556), .A2(KEYINPUT29), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n268), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n587), .B1(new_n590), .B2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n528), .B1(new_n586), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n500), .A2(new_n599), .ZN(new_n600));
  XOR2_X1   g414(.A(KEYINPUT97), .B(G101), .Z(new_n601));
  XNOR2_X1  g415(.A(new_n600), .B(new_n601), .ZN(G3));
  INV_X1    g416(.A(KEYINPUT98), .ZN(new_n603));
  OAI211_X1 g417(.A(new_n603), .B(new_n268), .C1(new_n565), .C2(new_n577), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(G472), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n603), .B1(new_n583), .B2(new_n268), .ZN(new_n606));
  OAI211_X1 g420(.A(new_n578), .B(new_n527), .C1(new_n605), .C2(new_n606), .ZN(new_n607));
  OAI21_X1  g421(.A(KEYINPUT99), .B1(new_n607), .B2(new_n436), .ZN(new_n608));
  INV_X1    g422(.A(new_n578), .ZN(new_n609));
  AOI21_X1  g423(.A(G902), .B1(new_n581), .B2(new_n582), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n587), .B1(new_n610), .B2(new_n603), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n268), .B1(new_n565), .B2(new_n577), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(KEYINPUT98), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n609), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT99), .ZN(new_n615));
  INV_X1    g429(.A(new_n436), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n614), .A2(new_n615), .A3(new_n527), .A4(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n321), .ZN(new_n618));
  OAI21_X1  g432(.A(KEYINPUT33), .B1(new_n618), .B2(new_n319), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT33), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n320), .A2(new_n620), .A3(new_n321), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n619), .A2(new_n621), .A3(G478), .ZN(new_n622));
  NAND2_X1  g436(.A1(G478), .A2(G902), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n322), .A2(new_n285), .A3(new_n268), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n622), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT100), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n284), .A2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT101), .ZN(new_n629));
  INV_X1    g443(.A(new_n496), .ZN(new_n630));
  INV_X1    g444(.A(new_n338), .ZN(new_n631));
  AOI211_X1 g445(.A(new_n630), .B(new_n631), .C1(new_n493), .C2(new_n494), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n628), .A2(new_n629), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n267), .A2(new_n268), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(G475), .ZN(new_n635));
  INV_X1    g449(.A(new_n283), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n282), .B1(new_n281), .B2(new_n268), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n635), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n625), .B(KEYINPUT100), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n638), .A2(new_n639), .A3(new_n632), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(KEYINPUT101), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n633), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n608), .A2(new_n617), .A3(new_n642), .ZN(new_n643));
  XOR2_X1   g457(.A(KEYINPUT34), .B(G104), .Z(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G6));
  NAND2_X1  g459(.A1(new_n608), .A2(new_n617), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT103), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT102), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n648), .B1(new_n636), .B2(new_n637), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n280), .A2(KEYINPUT102), .A3(new_n283), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n269), .A2(new_n327), .ZN(new_n652));
  AND4_X1   g466(.A1(new_n647), .A2(new_n651), .A3(new_n632), .A4(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n635), .A2(new_n326), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n654), .B1(new_n649), .B2(new_n650), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n647), .B1(new_n655), .B2(new_n632), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n646), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(KEYINPUT35), .B(G107), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G9));
  OR2_X1    g474(.A1(new_n520), .A2(KEYINPUT36), .ZN(new_n661));
  XOR2_X1   g475(.A(new_n661), .B(new_n516), .Z(new_n662));
  OAI211_X1 g476(.A(new_n662), .B(new_n268), .C1(new_n290), .C2(G234), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n525), .A2(new_n663), .ZN(new_n664));
  OAI211_X1 g478(.A(new_n578), .B(new_n664), .C1(new_n605), .C2(new_n606), .ZN(new_n665));
  INV_X1    g479(.A(KEYINPUT104), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n613), .A2(G472), .A3(new_n604), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n668), .A2(KEYINPUT104), .A3(new_n578), .A4(new_n664), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n667), .A2(new_n500), .A3(new_n669), .ZN(new_n670));
  XOR2_X1   g484(.A(KEYINPUT37), .B(G110), .Z(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G12));
  AOI21_X1  g486(.A(new_n584), .B1(new_n583), .B2(new_n531), .ZN(new_n673));
  AOI211_X1 g487(.A(KEYINPUT32), .B(new_n530), .C1(new_n581), .C2(new_n582), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n598), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n630), .B1(new_n493), .B2(new_n494), .ZN(new_n676));
  INV_X1    g490(.A(new_n664), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n436), .A2(new_n677), .ZN(new_n678));
  AND3_X1   g492(.A1(new_n675), .A2(new_n676), .A3(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(new_n336), .ZN(new_n680));
  INV_X1    g494(.A(G900), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n680), .B1(new_n331), .B2(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n655), .A2(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n679), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G128), .ZN(G30));
  XNOR2_X1  g501(.A(new_n682), .B(KEYINPUT39), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n436), .A2(new_n688), .ZN(new_n689));
  OR2_X1    g503(.A1(new_n689), .A2(KEYINPUT40), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n689), .A2(KEYINPUT40), .ZN(new_n691));
  AOI211_X1 g505(.A(new_n630), .B(new_n664), .C1(new_n690), .C2(new_n691), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n556), .B1(new_n552), .B2(new_n592), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n693), .B1(new_n559), .B2(new_n560), .ZN(new_n694));
  OAI21_X1  g508(.A(G472), .B1(new_n694), .B2(G902), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n586), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n495), .A2(new_n498), .ZN(new_n697));
  XOR2_X1   g511(.A(new_n697), .B(KEYINPUT38), .Z(new_n698));
  NOR2_X1   g512(.A1(new_n284), .A2(new_n327), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n692), .A2(new_n696), .A3(new_n698), .A4(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G143), .ZN(G45));
  NOR3_X1   g515(.A1(new_n284), .A2(new_n627), .A3(new_n682), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n675), .A2(new_n702), .A3(new_n676), .A4(new_n678), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT105), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g519(.A(new_n676), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n706), .B1(new_n586), .B2(new_n598), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n707), .A2(KEYINPUT105), .A3(new_n678), .A4(new_n702), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n705), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G146), .ZN(G48));
  AOI21_X1  g524(.A(new_n597), .B1(new_n579), .B2(new_n585), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n422), .A2(new_n268), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(G469), .ZN(new_n713));
  AND3_X1   g527(.A1(new_n713), .A2(new_n424), .A3(new_n434), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  NOR3_X1   g529(.A1(new_n711), .A2(new_n528), .A3(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n642), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(KEYINPUT41), .B(G113), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n717), .B(new_n718), .ZN(G15));
  OAI21_X1  g533(.A(new_n716), .B1(new_n653), .B2(new_n656), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G116), .ZN(G18));
  NOR2_X1   g535(.A1(new_n339), .A2(new_n715), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n707), .A2(new_n664), .A3(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G119), .ZN(G21));
  NOR2_X1   g538(.A1(new_n567), .A2(new_n563), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n593), .A2(new_n574), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n530), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  INV_X1    g541(.A(new_n727), .ZN(new_n728));
  OAI211_X1 g542(.A(new_n527), .B(new_n728), .C1(new_n610), .C2(new_n587), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n729), .A2(new_n715), .ZN(new_n730));
  NOR4_X1   g544(.A1(new_n284), .A2(new_n706), .A3(new_n327), .A4(new_n631), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT106), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n730), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n727), .B1(new_n612), .B2(G472), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n734), .A2(new_n527), .A3(new_n714), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n638), .A2(new_n676), .A3(new_n326), .A4(new_n338), .ZN(new_n736));
  OAI21_X1  g550(.A(KEYINPUT106), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n733), .A2(new_n737), .ZN(new_n738));
  XOR2_X1   g552(.A(KEYINPUT107), .B(G122), .Z(new_n739));
  XNOR2_X1  g553(.A(new_n738), .B(new_n739), .ZN(G24));
  NAND3_X1  g554(.A1(new_n638), .A2(new_n639), .A3(new_n683), .ZN(new_n741));
  OAI211_X1 g555(.A(new_n664), .B(new_n728), .C1(new_n610), .C2(new_n587), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n714), .A2(new_n676), .ZN(new_n743));
  NOR3_X1   g557(.A1(new_n741), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(new_n227), .ZN(G27));
  AOI21_X1  g559(.A(new_n630), .B1(new_n495), .B2(new_n498), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT108), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n429), .A2(new_n747), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n426), .A2(KEYINPUT108), .A3(new_n428), .A4(G469), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n748), .A2(new_n424), .A3(new_n430), .A4(new_n749), .ZN(new_n750));
  AND3_X1   g564(.A1(new_n746), .A2(new_n434), .A3(new_n750), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n675), .A2(new_n751), .A3(new_n702), .A4(new_n527), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT42), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n599), .A2(KEYINPUT42), .A3(new_n702), .A4(new_n751), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G131), .ZN(G33));
  NAND3_X1  g571(.A1(new_n685), .A2(new_n599), .A3(new_n751), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G134), .ZN(G36));
  NAND2_X1  g573(.A1(new_n284), .A2(new_n639), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT43), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n760), .B(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(new_n614), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n762), .A2(KEYINPUT44), .A3(new_n763), .A4(new_n664), .ZN(new_n764));
  AND2_X1   g578(.A1(new_n764), .A2(new_n746), .ZN(new_n765));
  INV_X1    g579(.A(new_n424), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n426), .A2(KEYINPUT45), .A3(new_n428), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT45), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n401), .B1(new_n413), .B2(new_n397), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n768), .B1(new_n769), .B2(new_n427), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n767), .A2(G469), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(new_n430), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT46), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n766), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n771), .A2(KEYINPUT46), .A3(new_n430), .ZN(new_n775));
  AOI22_X1  g589(.A1(new_n774), .A2(new_n775), .B1(G221), .B2(new_n433), .ZN(new_n776));
  INV_X1    g590(.A(new_n776), .ZN(new_n777));
  OR2_X1    g591(.A1(new_n777), .A2(new_n688), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n762), .A2(new_n763), .A3(new_n664), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT44), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n778), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n765), .A2(new_n781), .ZN(new_n782));
  XOR2_X1   g596(.A(KEYINPUT109), .B(G137), .Z(new_n783));
  XNOR2_X1  g597(.A(new_n782), .B(new_n783), .ZN(G39));
  XOR2_X1   g598(.A(KEYINPUT110), .B(KEYINPUT47), .Z(new_n785));
  INV_X1    g599(.A(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n776), .A2(new_n786), .ZN(new_n787));
  NOR2_X1   g601(.A1(KEYINPUT110), .A2(KEYINPUT47), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n787), .B1(new_n776), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n711), .A2(new_n528), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n702), .A2(new_n746), .ZN(new_n791));
  NOR3_X1   g605(.A1(new_n789), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(new_n215), .ZN(G42));
  INV_X1    g607(.A(KEYINPUT54), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n744), .B1(new_n679), .B2(new_n685), .ZN(new_n795));
  NOR4_X1   g609(.A1(new_n284), .A2(new_n706), .A3(new_n327), .A4(new_n682), .ZN(new_n796));
  AND2_X1   g610(.A1(new_n677), .A2(new_n750), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n696), .A2(new_n796), .A3(new_n434), .A4(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n709), .A2(new_n795), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(KEYINPUT52), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT52), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n709), .A2(new_n795), .A3(new_n801), .A4(new_n798), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(new_n742), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n804), .A2(new_n751), .A3(new_n702), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n805), .A2(KEYINPUT112), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT112), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n804), .A2(new_n751), .A3(new_n702), .A4(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  AND3_X1   g623(.A1(new_n678), .A2(new_n683), .A3(new_n746), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT111), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n326), .B(new_n811), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n812), .B1(new_n649), .B2(new_n650), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n810), .A2(new_n813), .A3(new_n675), .A4(new_n635), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n756), .A2(new_n809), .A3(new_n758), .A4(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n720), .A2(new_n717), .A3(new_n738), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n670), .A2(new_n600), .A3(new_n723), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n638), .A2(new_n639), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n284), .A2(new_n812), .ZN(new_n819));
  AOI211_X1 g633(.A(new_n499), .B(new_n631), .C1(new_n818), .C2(new_n819), .ZN(new_n820));
  AND3_X1   g634(.A1(new_n608), .A2(new_n617), .A3(new_n820), .ZN(new_n821));
  NOR4_X1   g635(.A1(new_n815), .A2(new_n816), .A3(new_n817), .A4(new_n821), .ZN(new_n822));
  AOI21_X1  g636(.A(KEYINPUT53), .B1(new_n803), .B2(new_n822), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n816), .A2(new_n817), .A3(new_n821), .ZN(new_n824));
  AND4_X1   g638(.A1(new_n756), .A2(new_n809), .A3(new_n758), .A4(new_n814), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n824), .A2(new_n800), .A3(new_n825), .A4(new_n802), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT53), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n794), .B1(new_n823), .B2(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n803), .A2(new_n822), .A3(KEYINPUT53), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n826), .A2(new_n827), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n830), .A2(new_n831), .A3(KEYINPUT54), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n829), .A2(new_n832), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n762), .A2(new_n680), .ZN(new_n834));
  INV_X1    g648(.A(new_n746), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n835), .A2(new_n715), .ZN(new_n836));
  AND3_X1   g650(.A1(new_n834), .A2(new_n599), .A3(new_n836), .ZN(new_n837));
  OR3_X1    g651(.A1(new_n837), .A2(KEYINPUT114), .A3(KEYINPUT48), .ZN(new_n838));
  INV_X1    g652(.A(new_n729), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n834), .A2(new_n839), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n715), .A2(new_n706), .ZN(new_n841));
  AOI211_X1 g655(.A(G953), .B(new_n334), .C1(new_n840), .C2(new_n841), .ZN(new_n842));
  AND2_X1   g656(.A1(new_n838), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n837), .A2(KEYINPUT114), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(KEYINPUT48), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n837), .A2(KEYINPUT114), .ZN(new_n846));
  OR2_X1    g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT115), .ZN(new_n848));
  INV_X1    g662(.A(new_n696), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n849), .A2(new_n527), .A3(new_n680), .A4(new_n836), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n850), .A2(new_n818), .ZN(new_n851));
  INV_X1    g665(.A(new_n851), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n843), .A2(new_n847), .A3(new_n848), .A4(new_n852), .ZN(new_n853));
  OAI211_X1 g667(.A(new_n838), .B(new_n842), .C1(new_n845), .C2(new_n846), .ZN(new_n854));
  OAI21_X1  g668(.A(KEYINPUT115), .B1(new_n854), .B2(new_n851), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT50), .ZN(new_n856));
  AOI211_X1 g670(.A(new_n496), .B(new_n698), .C1(KEYINPUT113), .C2(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n840), .A2(new_n714), .A3(new_n857), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n856), .A2(KEYINPUT113), .ZN(new_n859));
  OR2_X1    g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n834), .A2(new_n804), .A3(new_n836), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n858), .A2(new_n859), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n850), .A2(new_n638), .A3(new_n639), .ZN(new_n863));
  AND2_X1   g677(.A1(new_n713), .A2(new_n424), .ZN(new_n864));
  INV_X1    g678(.A(new_n435), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n835), .B1(new_n789), .B2(new_n866), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n863), .B1(new_n840), .B2(new_n867), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n860), .A2(new_n861), .A3(new_n862), .A4(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT51), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n833), .A2(new_n853), .A3(new_n855), .A4(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n869), .A2(new_n870), .ZN(new_n873));
  OAI22_X1  g687(.A1(new_n872), .A2(new_n873), .B1(G952), .B2(G953), .ZN(new_n874));
  INV_X1    g688(.A(new_n864), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n528), .B1(new_n875), .B2(KEYINPUT49), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n876), .B1(KEYINPUT49), .B2(new_n875), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n877), .A2(new_n630), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n698), .A2(new_n696), .A3(new_n760), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n878), .A2(new_n879), .A3(new_n435), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n874), .A2(new_n880), .ZN(G75));
  AOI21_X1  g695(.A(new_n268), .B1(new_n830), .B2(new_n831), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(G210), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n462), .A2(new_n479), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n477), .A2(new_n474), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n886), .A2(new_n480), .ZN(new_n887));
  XOR2_X1   g701(.A(new_n887), .B(KEYINPUT55), .Z(new_n888));
  XNOR2_X1  g702(.A(KEYINPUT116), .B(KEYINPUT56), .ZN(new_n889));
  AND3_X1   g703(.A1(new_n883), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT56), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n888), .B1(new_n883), .B2(new_n891), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n248), .A2(G952), .ZN(new_n893));
  NOR3_X1   g707(.A1(new_n890), .A2(new_n892), .A3(new_n893), .ZN(G51));
  XOR2_X1   g708(.A(new_n430), .B(KEYINPUT57), .Z(new_n895));
  NAND3_X1  g709(.A1(new_n829), .A2(new_n832), .A3(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT117), .ZN(new_n897));
  AND3_X1   g711(.A1(new_n896), .A2(new_n897), .A3(new_n422), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n897), .B1(new_n896), .B2(new_n422), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(new_n771), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n882), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n893), .B1(new_n900), .B2(new_n902), .ZN(G54));
  NAND3_X1  g717(.A1(new_n882), .A2(KEYINPUT58), .A3(G475), .ZN(new_n904));
  INV_X1    g718(.A(new_n278), .ZN(new_n905));
  AND2_X1   g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n904), .A2(new_n905), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n906), .A2(new_n907), .A3(new_n893), .ZN(G60));
  INV_X1    g722(.A(new_n833), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n619), .A2(new_n621), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n623), .B(KEYINPUT118), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n911), .B(KEYINPUT59), .ZN(new_n912));
  AND3_X1   g726(.A1(new_n909), .A2(new_n910), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n910), .B1(new_n909), .B2(new_n912), .ZN(new_n914));
  NOR3_X1   g728(.A1(new_n913), .A2(new_n914), .A3(new_n893), .ZN(G63));
  NAND2_X1  g729(.A1(new_n830), .A2(new_n831), .ZN(new_n916));
  XNOR2_X1  g730(.A(KEYINPUT119), .B(KEYINPUT60), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n290), .A2(new_n268), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n917), .B(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n916), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n893), .B1(new_n920), .B2(new_n521), .ZN(new_n921));
  INV_X1    g735(.A(new_n662), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n921), .B1(new_n922), .B2(new_n920), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT61), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n923), .B(new_n924), .ZN(G66));
  OAI21_X1  g739(.A(G953), .B1(new_n332), .B2(new_n463), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n926), .B1(new_n824), .B2(new_n328), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n884), .B1(G898), .B2(new_n248), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n927), .B(new_n928), .ZN(G69));
  AND2_X1   g743(.A1(new_n709), .A2(new_n795), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(new_n700), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT123), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT62), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  OR2_X1    g748(.A1(new_n931), .A2(new_n934), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n932), .A2(new_n933), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n936), .B1(new_n931), .B2(new_n934), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n818), .A2(new_n819), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n599), .A2(new_n689), .A3(new_n746), .A4(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n792), .B1(new_n765), .B2(new_n781), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n935), .A2(new_n937), .A3(new_n939), .A4(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(new_n248), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n543), .B1(new_n550), .B2(KEYINPUT30), .ZN(new_n943));
  XOR2_X1   g757(.A(KEYINPUT120), .B(KEYINPUT121), .Z(new_n944));
  XNOR2_X1  g758(.A(new_n943), .B(new_n944), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n945), .B(new_n274), .Z(new_n946));
  INV_X1    g760(.A(KEYINPUT122), .ZN(new_n947));
  OR2_X1    g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n946), .A2(new_n947), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n942), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(KEYINPUT125), .ZN(new_n951));
  NAND2_X1  g765(.A1(G227), .A2(G900), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n951), .A2(new_n328), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n709), .A2(new_n795), .ZN(new_n954));
  AOI211_X1 g768(.A(new_n792), .B(new_n954), .C1(new_n765), .C2(new_n781), .ZN(new_n955));
  AND2_X1   g769(.A1(new_n756), .A2(new_n758), .ZN(new_n956));
  INV_X1    g770(.A(new_n778), .ZN(new_n957));
  NAND4_X1  g771(.A1(new_n957), .A2(new_n599), .A3(new_n676), .A4(new_n699), .ZN(new_n958));
  NAND4_X1  g772(.A1(new_n955), .A2(KEYINPUT124), .A3(new_n956), .A4(new_n958), .ZN(new_n959));
  NAND4_X1  g773(.A1(new_n940), .A2(new_n956), .A3(new_n930), .A4(new_n958), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT124), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n959), .A2(new_n962), .A3(new_n248), .ZN(new_n963));
  OAI211_X1 g777(.A(new_n963), .B(new_n946), .C1(new_n681), .C2(new_n248), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n953), .A2(new_n950), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n964), .A2(new_n950), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n966), .A2(new_n328), .A3(new_n951), .A4(new_n952), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n965), .A2(new_n967), .ZN(G72));
  NAND3_X1  g782(.A1(new_n959), .A2(new_n962), .A3(new_n824), .ZN(new_n969));
  XNOR2_X1  g783(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n970));
  NAND2_X1  g784(.A1(G472), .A2(G902), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n970), .B(new_n971), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n556), .B1(new_n969), .B2(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(new_n588), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(new_n893), .ZN(new_n976));
  INV_X1    g790(.A(new_n824), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n972), .B1(new_n941), .B2(new_n977), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n978), .A2(new_n588), .A3(new_n556), .ZN(new_n979));
  AND2_X1   g793(.A1(new_n916), .A2(new_n972), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n561), .B1(new_n974), .B2(new_n556), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND4_X1  g796(.A1(new_n975), .A2(new_n976), .A3(new_n979), .A4(new_n982), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n983), .A2(KEYINPUT127), .ZN(new_n984));
  AOI22_X1  g798(.A1(new_n973), .A2(new_n974), .B1(new_n980), .B2(new_n981), .ZN(new_n985));
  INV_X1    g799(.A(KEYINPUT127), .ZN(new_n986));
  NAND4_X1  g800(.A1(new_n985), .A2(new_n986), .A3(new_n976), .A4(new_n979), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n984), .A2(new_n987), .ZN(G57));
endmodule


