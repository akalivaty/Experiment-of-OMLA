

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U550 ( .A(KEYINPUT31), .ZN(n696) );
  XNOR2_X1 U551 ( .A(n696), .B(KEYINPUT106), .ZN(n697) );
  XNOR2_X1 U552 ( .A(n698), .B(n697), .ZN(n743) );
  NOR2_X2 U553 ( .A1(n772), .A2(n685), .ZN(n714) );
  INV_X1 U554 ( .A(n714), .ZN(n730) );
  NAND2_X1 U555 ( .A1(G8), .A2(n730), .ZN(n765) );
  NOR2_X1 U556 ( .A1(G1384), .A2(G164), .ZN(n684) );
  NOR2_X2 U557 ( .A1(G2104), .A2(G2105), .ZN(n514) );
  NOR2_X1 U558 ( .A1(G651), .A2(n621), .ZN(n639) );
  NOR2_X1 U559 ( .A1(n522), .A2(n521), .ZN(G164) );
  XOR2_X2 U560 ( .A(KEYINPUT17), .B(n514), .Z(n874) );
  NAND2_X1 U561 ( .A1(G138), .A2(n874), .ZN(n516) );
  INV_X1 U562 ( .A(G2105), .ZN(n518) );
  AND2_X1 U563 ( .A1(n518), .A2(G2104), .ZN(n875) );
  NAND2_X1 U564 ( .A1(G102), .A2(n875), .ZN(n515) );
  NAND2_X1 U565 ( .A1(n516), .A2(n515), .ZN(n517) );
  XNOR2_X1 U566 ( .A(n517), .B(KEYINPUT88), .ZN(n522) );
  AND2_X1 U567 ( .A1(G2104), .A2(G2105), .ZN(n878) );
  NAND2_X1 U568 ( .A1(G114), .A2(n878), .ZN(n520) );
  NOR2_X1 U569 ( .A1(G2104), .A2(n518), .ZN(n879) );
  NAND2_X1 U570 ( .A1(G126), .A2(n879), .ZN(n519) );
  NAND2_X1 U571 ( .A1(n520), .A2(n519), .ZN(n521) );
  XNOR2_X1 U572 ( .A(KEYINPUT67), .B(G651), .ZN(n527) );
  NOR2_X1 U573 ( .A1(G543), .A2(n527), .ZN(n523) );
  XOR2_X1 U574 ( .A(KEYINPUT1), .B(n523), .Z(n640) );
  NAND2_X1 U575 ( .A1(n640), .A2(G64), .ZN(n526) );
  XOR2_X1 U576 ( .A(G543), .B(KEYINPUT0), .Z(n524) );
  XNOR2_X1 U577 ( .A(KEYINPUT66), .B(n524), .ZN(n621) );
  NAND2_X1 U578 ( .A1(n639), .A2(G52), .ZN(n525) );
  AND2_X1 U579 ( .A1(n526), .A2(n525), .ZN(n533) );
  XNOR2_X1 U580 ( .A(KEYINPUT9), .B(KEYINPUT70), .ZN(n531) );
  NOR2_X1 U581 ( .A1(G543), .A2(G651), .ZN(n635) );
  NAND2_X1 U582 ( .A1(G90), .A2(n635), .ZN(n529) );
  NOR2_X1 U583 ( .A1(n621), .A2(n527), .ZN(n636) );
  NAND2_X1 U584 ( .A1(G77), .A2(n636), .ZN(n528) );
  NAND2_X1 U585 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U586 ( .A(n531), .B(n530), .ZN(n532) );
  NAND2_X1 U587 ( .A1(n533), .A2(n532), .ZN(G301) );
  INV_X1 U588 ( .A(G301), .ZN(G171) );
  XNOR2_X1 U589 ( .A(G2451), .B(G2443), .ZN(n543) );
  XOR2_X1 U590 ( .A(G2446), .B(G2454), .Z(n535) );
  XNOR2_X1 U591 ( .A(KEYINPUT110), .B(G2435), .ZN(n534) );
  XNOR2_X1 U592 ( .A(n535), .B(n534), .ZN(n539) );
  XOR2_X1 U593 ( .A(KEYINPUT111), .B(G2438), .Z(n537) );
  XNOR2_X1 U594 ( .A(G1341), .B(G1348), .ZN(n536) );
  XNOR2_X1 U595 ( .A(n537), .B(n536), .ZN(n538) );
  XOR2_X1 U596 ( .A(n539), .B(n538), .Z(n541) );
  XNOR2_X1 U597 ( .A(G2430), .B(G2427), .ZN(n540) );
  XNOR2_X1 U598 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U599 ( .A(n543), .B(n542), .ZN(n544) );
  AND2_X1 U600 ( .A1(n544), .A2(G14), .ZN(G401) );
  AND2_X1 U601 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U602 ( .A1(G99), .A2(n875), .ZN(n546) );
  NAND2_X1 U603 ( .A1(G111), .A2(n878), .ZN(n545) );
  NAND2_X1 U604 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U605 ( .A(KEYINPUT80), .B(n547), .ZN(n550) );
  NAND2_X1 U606 ( .A1(n879), .A2(G123), .ZN(n548) );
  XOR2_X1 U607 ( .A(KEYINPUT18), .B(n548), .Z(n549) );
  NOR2_X1 U608 ( .A1(n550), .A2(n549), .ZN(n552) );
  NAND2_X1 U609 ( .A1(n874), .A2(G135), .ZN(n551) );
  NAND2_X1 U610 ( .A1(n552), .A2(n551), .ZN(n964) );
  XNOR2_X1 U611 ( .A(G2096), .B(n964), .ZN(n553) );
  OR2_X1 U612 ( .A1(G2100), .A2(n553), .ZN(G156) );
  INV_X1 U613 ( .A(G132), .ZN(G219) );
  INV_X1 U614 ( .A(G57), .ZN(G237) );
  NAND2_X1 U615 ( .A1(G88), .A2(n635), .ZN(n555) );
  NAND2_X1 U616 ( .A1(G75), .A2(n636), .ZN(n554) );
  NAND2_X1 U617 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U618 ( .A(KEYINPUT82), .B(n556), .ZN(n560) );
  NAND2_X1 U619 ( .A1(n639), .A2(G50), .ZN(n558) );
  NAND2_X1 U620 ( .A1(G62), .A2(n640), .ZN(n557) );
  NAND2_X1 U621 ( .A1(n558), .A2(n557), .ZN(n559) );
  NOR2_X1 U622 ( .A1(n560), .A2(n559), .ZN(G166) );
  NAND2_X1 U623 ( .A1(n639), .A2(G51), .ZN(n562) );
  NAND2_X1 U624 ( .A1(G63), .A2(n640), .ZN(n561) );
  NAND2_X1 U625 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U626 ( .A(KEYINPUT6), .B(n563), .ZN(n570) );
  NAND2_X1 U627 ( .A1(n635), .A2(G89), .ZN(n564) );
  XNOR2_X1 U628 ( .A(n564), .B(KEYINPUT4), .ZN(n566) );
  NAND2_X1 U629 ( .A1(G76), .A2(n636), .ZN(n565) );
  NAND2_X1 U630 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U631 ( .A(KEYINPUT5), .B(n567), .Z(n568) );
  XNOR2_X1 U632 ( .A(KEYINPUT76), .B(n568), .ZN(n569) );
  NOR2_X1 U633 ( .A1(n570), .A2(n569), .ZN(n571) );
  XOR2_X1 U634 ( .A(KEYINPUT7), .B(n571), .Z(G168) );
  XOR2_X1 U635 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U636 ( .A1(G7), .A2(G661), .ZN(n572) );
  XNOR2_X1 U637 ( .A(n572), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U638 ( .A(G223), .ZN(n828) );
  NAND2_X1 U639 ( .A1(n828), .A2(G567), .ZN(n573) );
  XOR2_X1 U640 ( .A(KEYINPUT11), .B(n573), .Z(G234) );
  NAND2_X1 U641 ( .A1(G56), .A2(n640), .ZN(n574) );
  XNOR2_X1 U642 ( .A(n574), .B(KEYINPUT14), .ZN(n576) );
  NAND2_X1 U643 ( .A1(G43), .A2(n639), .ZN(n575) );
  NAND2_X1 U644 ( .A1(n576), .A2(n575), .ZN(n584) );
  XOR2_X1 U645 ( .A(KEYINPUT12), .B(KEYINPUT74), .Z(n578) );
  NAND2_X1 U646 ( .A1(G81), .A2(n635), .ZN(n577) );
  XNOR2_X1 U647 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U648 ( .A(KEYINPUT73), .B(n579), .ZN(n581) );
  NAND2_X1 U649 ( .A1(G68), .A2(n636), .ZN(n580) );
  NAND2_X1 U650 ( .A1(n581), .A2(n580), .ZN(n582) );
  XOR2_X1 U651 ( .A(KEYINPUT13), .B(n582), .Z(n583) );
  NOR2_X1 U652 ( .A1(n584), .A2(n583), .ZN(n999) );
  NAND2_X1 U653 ( .A1(G860), .A2(n999), .ZN(n585) );
  XOR2_X1 U654 ( .A(KEYINPUT75), .B(n585), .Z(G153) );
  NAND2_X1 U655 ( .A1(G868), .A2(G301), .ZN(n594) );
  NAND2_X1 U656 ( .A1(n639), .A2(G54), .ZN(n587) );
  NAND2_X1 U657 ( .A1(G66), .A2(n640), .ZN(n586) );
  NAND2_X1 U658 ( .A1(n587), .A2(n586), .ZN(n591) );
  NAND2_X1 U659 ( .A1(G92), .A2(n635), .ZN(n589) );
  NAND2_X1 U660 ( .A1(G79), .A2(n636), .ZN(n588) );
  NAND2_X1 U661 ( .A1(n589), .A2(n588), .ZN(n590) );
  NOR2_X1 U662 ( .A1(n591), .A2(n590), .ZN(n592) );
  XOR2_X1 U663 ( .A(KEYINPUT15), .B(n592), .Z(n834) );
  INV_X1 U664 ( .A(n834), .ZN(n987) );
  INV_X1 U665 ( .A(G868), .ZN(n658) );
  NAND2_X1 U666 ( .A1(n987), .A2(n658), .ZN(n593) );
  NAND2_X1 U667 ( .A1(n594), .A2(n593), .ZN(G284) );
  NAND2_X1 U668 ( .A1(G91), .A2(n635), .ZN(n596) );
  NAND2_X1 U669 ( .A1(G78), .A2(n636), .ZN(n595) );
  NAND2_X1 U670 ( .A1(n596), .A2(n595), .ZN(n597) );
  XNOR2_X1 U671 ( .A(KEYINPUT71), .B(n597), .ZN(n601) );
  NAND2_X1 U672 ( .A1(n640), .A2(G65), .ZN(n599) );
  NAND2_X1 U673 ( .A1(n639), .A2(G53), .ZN(n598) );
  AND2_X1 U674 ( .A1(n599), .A2(n598), .ZN(n600) );
  NAND2_X1 U675 ( .A1(n601), .A2(n600), .ZN(G299) );
  NOR2_X1 U676 ( .A1(G286), .A2(n658), .ZN(n602) );
  XOR2_X1 U677 ( .A(KEYINPUT77), .B(n602), .Z(n605) );
  NOR2_X1 U678 ( .A1(G868), .A2(G299), .ZN(n603) );
  XNOR2_X1 U679 ( .A(KEYINPUT78), .B(n603), .ZN(n604) );
  NOR2_X1 U680 ( .A1(n605), .A2(n604), .ZN(G297) );
  INV_X1 U681 ( .A(G559), .ZN(n606) );
  NOR2_X1 U682 ( .A1(G860), .A2(n606), .ZN(n607) );
  XNOR2_X1 U683 ( .A(KEYINPUT79), .B(n607), .ZN(n608) );
  NAND2_X1 U684 ( .A1(n608), .A2(n834), .ZN(n609) );
  XNOR2_X1 U685 ( .A(n609), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U686 ( .A1(n834), .A2(G868), .ZN(n610) );
  NOR2_X1 U687 ( .A1(G559), .A2(n610), .ZN(n612) );
  AND2_X1 U688 ( .A1(n658), .A2(n999), .ZN(n611) );
  NOR2_X1 U689 ( .A1(n612), .A2(n611), .ZN(G282) );
  NAND2_X1 U690 ( .A1(n639), .A2(G55), .ZN(n614) );
  NAND2_X1 U691 ( .A1(G67), .A2(n640), .ZN(n613) );
  NAND2_X1 U692 ( .A1(n614), .A2(n613), .ZN(n618) );
  NAND2_X1 U693 ( .A1(G93), .A2(n635), .ZN(n616) );
  NAND2_X1 U694 ( .A1(G80), .A2(n636), .ZN(n615) );
  NAND2_X1 U695 ( .A1(n616), .A2(n615), .ZN(n617) );
  OR2_X1 U696 ( .A1(n618), .A2(n617), .ZN(n657) );
  NAND2_X1 U697 ( .A1(n834), .A2(G559), .ZN(n655) );
  XOR2_X1 U698 ( .A(n999), .B(n655), .Z(n619) );
  NOR2_X1 U699 ( .A1(G860), .A2(n619), .ZN(n620) );
  XOR2_X1 U700 ( .A(n657), .B(n620), .Z(G145) );
  NAND2_X1 U701 ( .A1(G49), .A2(n639), .ZN(n623) );
  NAND2_X1 U702 ( .A1(G87), .A2(n621), .ZN(n622) );
  NAND2_X1 U703 ( .A1(n623), .A2(n622), .ZN(n624) );
  NOR2_X1 U704 ( .A1(n640), .A2(n624), .ZN(n626) );
  NAND2_X1 U705 ( .A1(G651), .A2(G74), .ZN(n625) );
  NAND2_X1 U706 ( .A1(n626), .A2(n625), .ZN(G288) );
  NAND2_X1 U707 ( .A1(n636), .A2(G73), .ZN(n627) );
  XNOR2_X1 U708 ( .A(n627), .B(KEYINPUT2), .ZN(n634) );
  NAND2_X1 U709 ( .A1(n635), .A2(G86), .ZN(n629) );
  NAND2_X1 U710 ( .A1(G61), .A2(n640), .ZN(n628) );
  NAND2_X1 U711 ( .A1(n629), .A2(n628), .ZN(n632) );
  NAND2_X1 U712 ( .A1(G48), .A2(n639), .ZN(n630) );
  XNOR2_X1 U713 ( .A(KEYINPUT81), .B(n630), .ZN(n631) );
  NOR2_X1 U714 ( .A1(n632), .A2(n631), .ZN(n633) );
  NAND2_X1 U715 ( .A1(n634), .A2(n633), .ZN(G305) );
  NAND2_X1 U716 ( .A1(G85), .A2(n635), .ZN(n638) );
  NAND2_X1 U717 ( .A1(G72), .A2(n636), .ZN(n637) );
  NAND2_X1 U718 ( .A1(n638), .A2(n637), .ZN(n645) );
  NAND2_X1 U719 ( .A1(n639), .A2(G47), .ZN(n642) );
  NAND2_X1 U720 ( .A1(G60), .A2(n640), .ZN(n641) );
  NAND2_X1 U721 ( .A1(n642), .A2(n641), .ZN(n643) );
  XNOR2_X1 U722 ( .A(KEYINPUT68), .B(n643), .ZN(n644) );
  NOR2_X1 U723 ( .A1(n645), .A2(n644), .ZN(n646) );
  XNOR2_X1 U724 ( .A(n646), .B(KEYINPUT69), .ZN(G290) );
  INV_X1 U725 ( .A(G299), .ZN(n706) );
  XOR2_X1 U726 ( .A(KEYINPUT83), .B(KEYINPUT19), .Z(n647) );
  XNOR2_X1 U727 ( .A(G288), .B(n647), .ZN(n648) );
  XOR2_X1 U728 ( .A(n657), .B(n648), .Z(n650) );
  XNOR2_X1 U729 ( .A(G305), .B(n999), .ZN(n649) );
  XNOR2_X1 U730 ( .A(n650), .B(n649), .ZN(n651) );
  XNOR2_X1 U731 ( .A(n706), .B(n651), .ZN(n653) );
  XNOR2_X1 U732 ( .A(G290), .B(G166), .ZN(n652) );
  XNOR2_X1 U733 ( .A(n653), .B(n652), .ZN(n835) );
  XOR2_X1 U734 ( .A(n835), .B(KEYINPUT84), .Z(n654) );
  XNOR2_X1 U735 ( .A(n655), .B(n654), .ZN(n656) );
  NAND2_X1 U736 ( .A1(n656), .A2(G868), .ZN(n660) );
  NAND2_X1 U737 ( .A1(n658), .A2(n657), .ZN(n659) );
  NAND2_X1 U738 ( .A1(n660), .A2(n659), .ZN(G295) );
  NAND2_X1 U739 ( .A1(G2084), .A2(G2078), .ZN(n661) );
  XOR2_X1 U740 ( .A(KEYINPUT20), .B(n661), .Z(n662) );
  NAND2_X1 U741 ( .A1(G2090), .A2(n662), .ZN(n664) );
  XOR2_X1 U742 ( .A(KEYINPUT21), .B(KEYINPUT85), .Z(n663) );
  XNOR2_X1 U743 ( .A(n664), .B(n663), .ZN(n665) );
  NAND2_X1 U744 ( .A1(G2072), .A2(n665), .ZN(G158) );
  XNOR2_X1 U745 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U746 ( .A(KEYINPUT72), .B(G82), .Z(G220) );
  NAND2_X1 U747 ( .A1(G108), .A2(G120), .ZN(n666) );
  NOR2_X1 U748 ( .A1(G237), .A2(n666), .ZN(n667) );
  NAND2_X1 U749 ( .A1(G69), .A2(n667), .ZN(n832) );
  NAND2_X1 U750 ( .A1(n832), .A2(G567), .ZN(n673) );
  NOR2_X1 U751 ( .A1(G220), .A2(G219), .ZN(n668) );
  XNOR2_X1 U752 ( .A(KEYINPUT22), .B(n668), .ZN(n669) );
  NAND2_X1 U753 ( .A1(n669), .A2(G96), .ZN(n670) );
  NOR2_X1 U754 ( .A1(G218), .A2(n670), .ZN(n671) );
  XOR2_X1 U755 ( .A(KEYINPUT86), .B(n671), .Z(n833) );
  NAND2_X1 U756 ( .A1(G2106), .A2(n833), .ZN(n672) );
  NAND2_X1 U757 ( .A1(n673), .A2(n672), .ZN(n905) );
  NAND2_X1 U758 ( .A1(G483), .A2(G661), .ZN(n674) );
  NOR2_X1 U759 ( .A1(n905), .A2(n674), .ZN(n675) );
  XOR2_X1 U760 ( .A(KEYINPUT87), .B(n675), .Z(n831) );
  NAND2_X1 U761 ( .A1(n831), .A2(G36), .ZN(G176) );
  NAND2_X1 U762 ( .A1(G101), .A2(n875), .ZN(n676) );
  XOR2_X1 U763 ( .A(KEYINPUT23), .B(n676), .Z(n679) );
  NAND2_X1 U764 ( .A1(n874), .A2(G137), .ZN(n677) );
  XOR2_X1 U765 ( .A(KEYINPUT65), .B(n677), .Z(n678) );
  NAND2_X1 U766 ( .A1(n679), .A2(n678), .ZN(n683) );
  NAND2_X1 U767 ( .A1(G113), .A2(n878), .ZN(n681) );
  NAND2_X1 U768 ( .A1(G125), .A2(n879), .ZN(n680) );
  NAND2_X1 U769 ( .A1(n681), .A2(n680), .ZN(n682) );
  NOR2_X1 U770 ( .A1(n683), .A2(n682), .ZN(G160) );
  INV_X1 U771 ( .A(G166), .ZN(G303) );
  NAND2_X1 U772 ( .A1(G160), .A2(G40), .ZN(n772) );
  XNOR2_X1 U773 ( .A(n684), .B(KEYINPUT64), .ZN(n771) );
  INV_X1 U774 ( .A(n771), .ZN(n685) );
  NOR2_X1 U775 ( .A1(G1976), .A2(G288), .ZN(n751) );
  NAND2_X1 U776 ( .A1(n751), .A2(KEYINPUT33), .ZN(n686) );
  NOR2_X1 U777 ( .A1(n765), .A2(n686), .ZN(n756) );
  NAND2_X1 U778 ( .A1(G1976), .A2(G288), .ZN(n990) );
  INV_X1 U779 ( .A(n990), .ZN(n687) );
  NOR2_X1 U780 ( .A1(n687), .A2(n765), .ZN(n753) );
  XNOR2_X1 U781 ( .A(G2078), .B(KEYINPUT25), .ZN(n913) );
  NOR2_X1 U782 ( .A1(n730), .A2(n913), .ZN(n689) );
  XOR2_X1 U783 ( .A(KEYINPUT100), .B(G1961), .Z(n929) );
  NOR2_X1 U784 ( .A1(n714), .A2(n929), .ZN(n688) );
  NOR2_X1 U785 ( .A1(n689), .A2(n688), .ZN(n699) );
  OR2_X1 U786 ( .A1(G171), .A2(n699), .ZN(n690) );
  XNOR2_X1 U787 ( .A(n690), .B(KEYINPUT105), .ZN(n695) );
  NOR2_X1 U788 ( .A1(G1966), .A2(n765), .ZN(n745) );
  NOR2_X1 U789 ( .A1(G2084), .A2(n730), .ZN(n741) );
  NOR2_X1 U790 ( .A1(n745), .A2(n741), .ZN(n691) );
  NAND2_X1 U791 ( .A1(G8), .A2(n691), .ZN(n692) );
  XNOR2_X1 U792 ( .A(n692), .B(KEYINPUT30), .ZN(n693) );
  NOR2_X1 U793 ( .A1(n693), .A2(G168), .ZN(n694) );
  NOR2_X1 U794 ( .A1(n695), .A2(n694), .ZN(n698) );
  NAND2_X1 U795 ( .A1(n699), .A2(G171), .ZN(n728) );
  NAND2_X1 U796 ( .A1(n714), .A2(G2072), .ZN(n700) );
  XNOR2_X1 U797 ( .A(n700), .B(KEYINPUT27), .ZN(n702) );
  INV_X1 U798 ( .A(G1956), .ZN(n930) );
  NOR2_X1 U799 ( .A1(n930), .A2(n714), .ZN(n701) );
  NOR2_X1 U800 ( .A1(n702), .A2(n701), .ZN(n705) );
  NOR2_X1 U801 ( .A1(n706), .A2(n705), .ZN(n704) );
  XNOR2_X1 U802 ( .A(KEYINPUT28), .B(KEYINPUT101), .ZN(n703) );
  XNOR2_X1 U803 ( .A(n704), .B(n703), .ZN(n724) );
  NAND2_X1 U804 ( .A1(n706), .A2(n705), .ZN(n722) );
  NAND2_X1 U805 ( .A1(n730), .A2(G1341), .ZN(n707) );
  XNOR2_X1 U806 ( .A(n707), .B(KEYINPUT102), .ZN(n708) );
  NAND2_X1 U807 ( .A1(n708), .A2(n999), .ZN(n711) );
  NAND2_X1 U808 ( .A1(G1996), .A2(n714), .ZN(n709) );
  XOR2_X1 U809 ( .A(KEYINPUT26), .B(n709), .Z(n710) );
  NOR2_X1 U810 ( .A1(n711), .A2(n710), .ZN(n712) );
  OR2_X1 U811 ( .A1(n834), .A2(n712), .ZN(n720) );
  NAND2_X1 U812 ( .A1(n834), .A2(n712), .ZN(n718) );
  AND2_X1 U813 ( .A1(n730), .A2(G1348), .ZN(n713) );
  XNOR2_X1 U814 ( .A(n713), .B(KEYINPUT103), .ZN(n716) );
  NAND2_X1 U815 ( .A1(n714), .A2(G2067), .ZN(n715) );
  NAND2_X1 U816 ( .A1(n716), .A2(n715), .ZN(n717) );
  NAND2_X1 U817 ( .A1(n718), .A2(n717), .ZN(n719) );
  NAND2_X1 U818 ( .A1(n720), .A2(n719), .ZN(n721) );
  NAND2_X1 U819 ( .A1(n722), .A2(n721), .ZN(n723) );
  NAND2_X1 U820 ( .A1(n724), .A2(n723), .ZN(n726) );
  XOR2_X1 U821 ( .A(KEYINPUT29), .B(KEYINPUT104), .Z(n725) );
  XNOR2_X1 U822 ( .A(n726), .B(n725), .ZN(n727) );
  NAND2_X1 U823 ( .A1(n728), .A2(n727), .ZN(n742) );
  NOR2_X1 U824 ( .A1(G1971), .A2(n765), .ZN(n729) );
  XNOR2_X1 U825 ( .A(KEYINPUT107), .B(n729), .ZN(n733) );
  NOR2_X1 U826 ( .A1(G2090), .A2(n730), .ZN(n731) );
  NOR2_X1 U827 ( .A1(G166), .A2(n731), .ZN(n732) );
  NAND2_X1 U828 ( .A1(n733), .A2(n732), .ZN(n735) );
  AND2_X1 U829 ( .A1(n742), .A2(n735), .ZN(n734) );
  NAND2_X1 U830 ( .A1(n743), .A2(n734), .ZN(n738) );
  INV_X1 U831 ( .A(n735), .ZN(n736) );
  OR2_X1 U832 ( .A1(n736), .A2(G286), .ZN(n737) );
  AND2_X1 U833 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U834 ( .A1(n739), .A2(G8), .ZN(n740) );
  XNOR2_X1 U835 ( .A(n740), .B(KEYINPUT32), .ZN(n749) );
  NAND2_X1 U836 ( .A1(G8), .A2(n741), .ZN(n747) );
  AND2_X1 U837 ( .A1(n743), .A2(n742), .ZN(n744) );
  NOR2_X1 U838 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U839 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U840 ( .A1(n749), .A2(n748), .ZN(n764) );
  NOR2_X1 U841 ( .A1(G1971), .A2(G303), .ZN(n750) );
  NOR2_X1 U842 ( .A1(n751), .A2(n750), .ZN(n995) );
  NAND2_X1 U843 ( .A1(n764), .A2(n995), .ZN(n752) );
  AND2_X1 U844 ( .A1(n753), .A2(n752), .ZN(n754) );
  NOR2_X1 U845 ( .A1(KEYINPUT33), .A2(n754), .ZN(n755) );
  NOR2_X1 U846 ( .A1(n756), .A2(n755), .ZN(n758) );
  XOR2_X1 U847 ( .A(KEYINPUT108), .B(G1981), .Z(n757) );
  XNOR2_X1 U848 ( .A(G305), .B(n757), .ZN(n1002) );
  NAND2_X1 U849 ( .A1(n758), .A2(n1002), .ZN(n770) );
  NOR2_X1 U850 ( .A1(G1981), .A2(G305), .ZN(n759) );
  XOR2_X1 U851 ( .A(n759), .B(KEYINPUT24), .Z(n760) );
  NOR2_X1 U852 ( .A1(n765), .A2(n760), .ZN(n761) );
  XNOR2_X1 U853 ( .A(KEYINPUT99), .B(n761), .ZN(n768) );
  NOR2_X1 U854 ( .A1(G2090), .A2(G303), .ZN(n762) );
  NAND2_X1 U855 ( .A1(G8), .A2(n762), .ZN(n763) );
  NAND2_X1 U856 ( .A1(n764), .A2(n763), .ZN(n766) );
  NAND2_X1 U857 ( .A1(n766), .A2(n765), .ZN(n767) );
  AND2_X1 U858 ( .A1(n768), .A2(n767), .ZN(n769) );
  NAND2_X1 U859 ( .A1(n770), .A2(n769), .ZN(n811) );
  NOR2_X1 U860 ( .A1(n772), .A2(n771), .ZN(n823) );
  XNOR2_X1 U861 ( .A(G2067), .B(KEYINPUT37), .ZN(n820) );
  NAND2_X1 U862 ( .A1(n879), .A2(G128), .ZN(n773) );
  XOR2_X1 U863 ( .A(KEYINPUT91), .B(n773), .Z(n775) );
  NAND2_X1 U864 ( .A1(n878), .A2(G116), .ZN(n774) );
  NAND2_X1 U865 ( .A1(n775), .A2(n774), .ZN(n776) );
  XNOR2_X1 U866 ( .A(n776), .B(KEYINPUT35), .ZN(n782) );
  NAND2_X1 U867 ( .A1(n874), .A2(G140), .ZN(n777) );
  XNOR2_X1 U868 ( .A(n777), .B(KEYINPUT90), .ZN(n779) );
  NAND2_X1 U869 ( .A1(G104), .A2(n875), .ZN(n778) );
  NAND2_X1 U870 ( .A1(n779), .A2(n778), .ZN(n780) );
  XOR2_X1 U871 ( .A(KEYINPUT34), .B(n780), .Z(n781) );
  NAND2_X1 U872 ( .A1(n782), .A2(n781), .ZN(n783) );
  XOR2_X1 U873 ( .A(n783), .B(KEYINPUT36), .Z(n891) );
  OR2_X1 U874 ( .A1(n820), .A2(n891), .ZN(n784) );
  XOR2_X1 U875 ( .A(KEYINPUT92), .B(n784), .Z(n974) );
  NAND2_X1 U876 ( .A1(n823), .A2(n974), .ZN(n818) );
  NAND2_X1 U877 ( .A1(G131), .A2(n874), .ZN(n786) );
  NAND2_X1 U878 ( .A1(G95), .A2(n875), .ZN(n785) );
  NAND2_X1 U879 ( .A1(n786), .A2(n785), .ZN(n791) );
  NAND2_X1 U880 ( .A1(G107), .A2(n878), .ZN(n788) );
  NAND2_X1 U881 ( .A1(G119), .A2(n879), .ZN(n787) );
  NAND2_X1 U882 ( .A1(n788), .A2(n787), .ZN(n789) );
  XOR2_X1 U883 ( .A(KEYINPUT93), .B(n789), .Z(n790) );
  NOR2_X1 U884 ( .A1(n791), .A2(n790), .ZN(n792) );
  XOR2_X1 U885 ( .A(KEYINPUT94), .B(n792), .Z(n894) );
  NAND2_X1 U886 ( .A1(G1991), .A2(n894), .ZN(n804) );
  NAND2_X1 U887 ( .A1(n879), .A2(G129), .ZN(n793) );
  XOR2_X1 U888 ( .A(KEYINPUT95), .B(n793), .Z(n795) );
  NAND2_X1 U889 ( .A1(n878), .A2(G117), .ZN(n794) );
  NAND2_X1 U890 ( .A1(n795), .A2(n794), .ZN(n796) );
  XNOR2_X1 U891 ( .A(KEYINPUT96), .B(n796), .ZN(n799) );
  NAND2_X1 U892 ( .A1(n875), .A2(G105), .ZN(n797) );
  XOR2_X1 U893 ( .A(KEYINPUT38), .B(n797), .Z(n798) );
  NOR2_X1 U894 ( .A1(n799), .A2(n798), .ZN(n801) );
  NAND2_X1 U895 ( .A1(n874), .A2(G141), .ZN(n800) );
  NAND2_X1 U896 ( .A1(n801), .A2(n800), .ZN(n887) );
  NAND2_X1 U897 ( .A1(G1996), .A2(n887), .ZN(n802) );
  XOR2_X1 U898 ( .A(KEYINPUT97), .B(n802), .Z(n803) );
  NAND2_X1 U899 ( .A1(n804), .A2(n803), .ZN(n805) );
  XOR2_X1 U900 ( .A(KEYINPUT98), .B(n805), .Z(n971) );
  INV_X1 U901 ( .A(n971), .ZN(n806) );
  NAND2_X1 U902 ( .A1(n823), .A2(n806), .ZN(n812) );
  NAND2_X1 U903 ( .A1(n818), .A2(n812), .ZN(n809) );
  XOR2_X1 U904 ( .A(G1986), .B(KEYINPUT89), .Z(n807) );
  XNOR2_X1 U905 ( .A(G290), .B(n807), .ZN(n997) );
  AND2_X1 U906 ( .A1(n997), .A2(n823), .ZN(n808) );
  NOR2_X1 U907 ( .A1(n809), .A2(n808), .ZN(n810) );
  NAND2_X1 U908 ( .A1(n811), .A2(n810), .ZN(n826) );
  NOR2_X1 U909 ( .A1(G1996), .A2(n887), .ZN(n967) );
  INV_X1 U910 ( .A(n812), .ZN(n815) );
  NOR2_X1 U911 ( .A1(G1991), .A2(n894), .ZN(n963) );
  NOR2_X1 U912 ( .A1(G1986), .A2(G290), .ZN(n813) );
  NOR2_X1 U913 ( .A1(n963), .A2(n813), .ZN(n814) );
  NOR2_X1 U914 ( .A1(n815), .A2(n814), .ZN(n816) );
  NOR2_X1 U915 ( .A1(n967), .A2(n816), .ZN(n817) );
  XNOR2_X1 U916 ( .A(n817), .B(KEYINPUT39), .ZN(n819) );
  NAND2_X1 U917 ( .A1(n819), .A2(n818), .ZN(n821) );
  NAND2_X1 U918 ( .A1(n820), .A2(n891), .ZN(n960) );
  NAND2_X1 U919 ( .A1(n821), .A2(n960), .ZN(n822) );
  XOR2_X1 U920 ( .A(KEYINPUT109), .B(n822), .Z(n824) );
  NAND2_X1 U921 ( .A1(n824), .A2(n823), .ZN(n825) );
  NAND2_X1 U922 ( .A1(n826), .A2(n825), .ZN(n827) );
  XNOR2_X1 U923 ( .A(KEYINPUT40), .B(n827), .ZN(G329) );
  NAND2_X1 U924 ( .A1(G2106), .A2(n828), .ZN(G217) );
  AND2_X1 U925 ( .A1(G15), .A2(G2), .ZN(n829) );
  NAND2_X1 U926 ( .A1(G661), .A2(n829), .ZN(G259) );
  NAND2_X1 U927 ( .A1(G3), .A2(G1), .ZN(n830) );
  NAND2_X1 U928 ( .A1(n831), .A2(n830), .ZN(G188) );
  XOR2_X1 U929 ( .A(G120), .B(KEYINPUT112), .Z(G236) );
  XNOR2_X1 U930 ( .A(G96), .B(KEYINPUT113), .ZN(G221) );
  INV_X1 U932 ( .A(G108), .ZN(G238) );
  NOR2_X1 U933 ( .A1(n833), .A2(n832), .ZN(G325) );
  INV_X1 U934 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U935 ( .A(n834), .B(G286), .ZN(n836) );
  XNOR2_X1 U936 ( .A(n836), .B(n835), .ZN(n837) );
  XNOR2_X1 U937 ( .A(n837), .B(G171), .ZN(n838) );
  NOR2_X1 U938 ( .A1(G37), .A2(n838), .ZN(G397) );
  XOR2_X1 U939 ( .A(G2096), .B(KEYINPUT114), .Z(n840) );
  XNOR2_X1 U940 ( .A(G2072), .B(KEYINPUT43), .ZN(n839) );
  XNOR2_X1 U941 ( .A(n840), .B(n839), .ZN(n841) );
  XOR2_X1 U942 ( .A(n841), .B(KEYINPUT42), .Z(n843) );
  XNOR2_X1 U943 ( .A(G2067), .B(G2090), .ZN(n842) );
  XNOR2_X1 U944 ( .A(n843), .B(n842), .ZN(n847) );
  XOR2_X1 U945 ( .A(G2678), .B(G2100), .Z(n845) );
  XNOR2_X1 U946 ( .A(G2084), .B(G2078), .ZN(n844) );
  XNOR2_X1 U947 ( .A(n845), .B(n844), .ZN(n846) );
  XNOR2_X1 U948 ( .A(n847), .B(n846), .ZN(G227) );
  XOR2_X1 U949 ( .A(G1956), .B(G1966), .Z(n849) );
  XNOR2_X1 U950 ( .A(G1981), .B(G1971), .ZN(n848) );
  XNOR2_X1 U951 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U952 ( .A(n850), .B(G2474), .Z(n852) );
  XNOR2_X1 U953 ( .A(G1996), .B(G1991), .ZN(n851) );
  XNOR2_X1 U954 ( .A(n852), .B(n851), .ZN(n856) );
  XOR2_X1 U955 ( .A(KEYINPUT41), .B(G1961), .Z(n854) );
  XNOR2_X1 U956 ( .A(G1986), .B(G1976), .ZN(n853) );
  XNOR2_X1 U957 ( .A(n854), .B(n853), .ZN(n855) );
  XNOR2_X1 U958 ( .A(n856), .B(n855), .ZN(G229) );
  NAND2_X1 U959 ( .A1(G124), .A2(n879), .ZN(n857) );
  XNOR2_X1 U960 ( .A(n857), .B(KEYINPUT44), .ZN(n860) );
  NAND2_X1 U961 ( .A1(G136), .A2(n874), .ZN(n858) );
  XOR2_X1 U962 ( .A(KEYINPUT115), .B(n858), .Z(n859) );
  NAND2_X1 U963 ( .A1(n860), .A2(n859), .ZN(n864) );
  NAND2_X1 U964 ( .A1(G100), .A2(n875), .ZN(n862) );
  NAND2_X1 U965 ( .A1(G112), .A2(n878), .ZN(n861) );
  NAND2_X1 U966 ( .A1(n862), .A2(n861), .ZN(n863) );
  NOR2_X1 U967 ( .A1(n864), .A2(n863), .ZN(G162) );
  NAND2_X1 U968 ( .A1(G118), .A2(n878), .ZN(n866) );
  NAND2_X1 U969 ( .A1(G130), .A2(n879), .ZN(n865) );
  NAND2_X1 U970 ( .A1(n866), .A2(n865), .ZN(n872) );
  NAND2_X1 U971 ( .A1(G142), .A2(n874), .ZN(n868) );
  NAND2_X1 U972 ( .A1(G106), .A2(n875), .ZN(n867) );
  NAND2_X1 U973 ( .A1(n868), .A2(n867), .ZN(n869) );
  XOR2_X1 U974 ( .A(KEYINPUT116), .B(n869), .Z(n870) );
  XNOR2_X1 U975 ( .A(KEYINPUT45), .B(n870), .ZN(n871) );
  NOR2_X1 U976 ( .A1(n872), .A2(n871), .ZN(n873) );
  XOR2_X1 U977 ( .A(n873), .B(G162), .Z(n886) );
  NAND2_X1 U978 ( .A1(G139), .A2(n874), .ZN(n877) );
  NAND2_X1 U979 ( .A1(G103), .A2(n875), .ZN(n876) );
  NAND2_X1 U980 ( .A1(n877), .A2(n876), .ZN(n884) );
  NAND2_X1 U981 ( .A1(G115), .A2(n878), .ZN(n881) );
  NAND2_X1 U982 ( .A1(G127), .A2(n879), .ZN(n880) );
  NAND2_X1 U983 ( .A1(n881), .A2(n880), .ZN(n882) );
  XOR2_X1 U984 ( .A(KEYINPUT47), .B(n882), .Z(n883) );
  NOR2_X1 U985 ( .A1(n884), .A2(n883), .ZN(n955) );
  XNOR2_X1 U986 ( .A(G160), .B(n955), .ZN(n885) );
  XNOR2_X1 U987 ( .A(n886), .B(n885), .ZN(n890) );
  XNOR2_X1 U988 ( .A(KEYINPUT48), .B(n887), .ZN(n888) );
  XNOR2_X1 U989 ( .A(n888), .B(n964), .ZN(n889) );
  XOR2_X1 U990 ( .A(n890), .B(n889), .Z(n893) );
  XOR2_X1 U991 ( .A(n891), .B(KEYINPUT46), .Z(n892) );
  XNOR2_X1 U992 ( .A(n893), .B(n892), .ZN(n896) );
  XNOR2_X1 U993 ( .A(n894), .B(G164), .ZN(n895) );
  XNOR2_X1 U994 ( .A(n896), .B(n895), .ZN(n897) );
  NOR2_X1 U995 ( .A1(G37), .A2(n897), .ZN(G395) );
  NOR2_X1 U996 ( .A1(G401), .A2(n905), .ZN(n902) );
  NOR2_X1 U997 ( .A1(G227), .A2(G229), .ZN(n898) );
  XOR2_X1 U998 ( .A(KEYINPUT49), .B(n898), .Z(n899) );
  XNOR2_X1 U999 ( .A(n899), .B(KEYINPUT117), .ZN(n900) );
  NOR2_X1 U1000 ( .A1(G397), .A2(n900), .ZN(n901) );
  NAND2_X1 U1001 ( .A1(n902), .A2(n901), .ZN(n903) );
  NOR2_X1 U1002 ( .A1(n903), .A2(G395), .ZN(n904) );
  XNOR2_X1 U1003 ( .A(n904), .B(KEYINPUT118), .ZN(G308) );
  INV_X1 U1004 ( .A(G308), .ZN(G225) );
  INV_X1 U1005 ( .A(n905), .ZN(G319) );
  INV_X1 U1006 ( .A(G69), .ZN(G235) );
  INV_X1 U1007 ( .A(KEYINPUT55), .ZN(n979) );
  XNOR2_X1 U1008 ( .A(G2090), .B(G35), .ZN(n921) );
  XNOR2_X1 U1009 ( .A(KEYINPUT121), .B(G2067), .ZN(n906) );
  XNOR2_X1 U1010 ( .A(n906), .B(G26), .ZN(n912) );
  XOR2_X1 U1011 ( .A(G1991), .B(G25), .Z(n907) );
  NAND2_X1 U1012 ( .A1(n907), .A2(G28), .ZN(n910) );
  XNOR2_X1 U1013 ( .A(KEYINPUT122), .B(G2072), .ZN(n908) );
  XNOR2_X1 U1014 ( .A(G33), .B(n908), .ZN(n909) );
  NOR2_X1 U1015 ( .A1(n910), .A2(n909), .ZN(n911) );
  NAND2_X1 U1016 ( .A1(n912), .A2(n911), .ZN(n918) );
  XOR2_X1 U1017 ( .A(G1996), .B(G32), .Z(n915) );
  XNOR2_X1 U1018 ( .A(n913), .B(G27), .ZN(n914) );
  NAND2_X1 U1019 ( .A1(n915), .A2(n914), .ZN(n916) );
  XOR2_X1 U1020 ( .A(KEYINPUT123), .B(n916), .Z(n917) );
  NOR2_X1 U1021 ( .A1(n918), .A2(n917), .ZN(n919) );
  XNOR2_X1 U1022 ( .A(KEYINPUT53), .B(n919), .ZN(n920) );
  NOR2_X1 U1023 ( .A1(n921), .A2(n920), .ZN(n924) );
  XOR2_X1 U1024 ( .A(G2084), .B(G34), .Z(n922) );
  XNOR2_X1 U1025 ( .A(KEYINPUT54), .B(n922), .ZN(n923) );
  NAND2_X1 U1026 ( .A1(n924), .A2(n923), .ZN(n925) );
  XNOR2_X1 U1027 ( .A(n979), .B(n925), .ZN(n927) );
  INV_X1 U1028 ( .A(G29), .ZN(n926) );
  NAND2_X1 U1029 ( .A1(n927), .A2(n926), .ZN(n928) );
  NAND2_X1 U1030 ( .A1(G11), .A2(n928), .ZN(n954) );
  XNOR2_X1 U1031 ( .A(n929), .B(G5), .ZN(n950) );
  XNOR2_X1 U1032 ( .A(G20), .B(n930), .ZN(n934) );
  XNOR2_X1 U1033 ( .A(G1981), .B(G6), .ZN(n932) );
  XNOR2_X1 U1034 ( .A(G1341), .B(G19), .ZN(n931) );
  NOR2_X1 U1035 ( .A1(n932), .A2(n931), .ZN(n933) );
  NAND2_X1 U1036 ( .A1(n934), .A2(n933), .ZN(n937) );
  XOR2_X1 U1037 ( .A(KEYINPUT59), .B(G1348), .Z(n935) );
  XNOR2_X1 U1038 ( .A(G4), .B(n935), .ZN(n936) );
  NOR2_X1 U1039 ( .A1(n937), .A2(n936), .ZN(n938) );
  XOR2_X1 U1040 ( .A(KEYINPUT60), .B(n938), .Z(n940) );
  XNOR2_X1 U1041 ( .A(G1966), .B(G21), .ZN(n939) );
  NOR2_X1 U1042 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1043 ( .A(KEYINPUT127), .B(n941), .ZN(n948) );
  XNOR2_X1 U1044 ( .A(G1976), .B(G23), .ZN(n943) );
  XNOR2_X1 U1045 ( .A(G1971), .B(G22), .ZN(n942) );
  NOR2_X1 U1046 ( .A1(n943), .A2(n942), .ZN(n945) );
  XOR2_X1 U1047 ( .A(G1986), .B(G24), .Z(n944) );
  NAND2_X1 U1048 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1049 ( .A(KEYINPUT58), .B(n946), .ZN(n947) );
  NOR2_X1 U1050 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1051 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1052 ( .A(KEYINPUT61), .B(n951), .ZN(n952) );
  NOR2_X1 U1053 ( .A1(G16), .A2(n952), .ZN(n953) );
  NOR2_X1 U1054 ( .A1(n954), .A2(n953), .ZN(n983) );
  XOR2_X1 U1055 ( .A(G2072), .B(n955), .Z(n956) );
  XNOR2_X1 U1056 ( .A(KEYINPUT120), .B(n956), .ZN(n958) );
  XOR2_X1 U1057 ( .A(G164), .B(G2078), .Z(n957) );
  NOR2_X1 U1058 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1059 ( .A(n959), .B(KEYINPUT50), .ZN(n961) );
  NAND2_X1 U1060 ( .A1(n961), .A2(n960), .ZN(n977) );
  XOR2_X1 U1061 ( .A(G160), .B(G2084), .Z(n962) );
  NOR2_X1 U1062 ( .A1(n963), .A2(n962), .ZN(n965) );
  NAND2_X1 U1063 ( .A1(n965), .A2(n964), .ZN(n970) );
  XOR2_X1 U1064 ( .A(G2090), .B(G162), .Z(n966) );
  NOR2_X1 U1065 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1066 ( .A(n968), .B(KEYINPUT51), .ZN(n969) );
  NOR2_X1 U1067 ( .A1(n970), .A2(n969), .ZN(n972) );
  NAND2_X1 U1068 ( .A1(n972), .A2(n971), .ZN(n973) );
  NOR2_X1 U1069 ( .A1(n974), .A2(n973), .ZN(n975) );
  XNOR2_X1 U1070 ( .A(n975), .B(KEYINPUT119), .ZN(n976) );
  NOR2_X1 U1071 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1072 ( .A(KEYINPUT52), .B(n978), .ZN(n980) );
  NAND2_X1 U1073 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1074 ( .A1(n981), .A2(G29), .ZN(n982) );
  NAND2_X1 U1075 ( .A1(n983), .A2(n982), .ZN(n1011) );
  XOR2_X1 U1076 ( .A(G16), .B(KEYINPUT124), .Z(n984) );
  XNOR2_X1 U1077 ( .A(KEYINPUT56), .B(n984), .ZN(n1009) );
  XNOR2_X1 U1078 ( .A(G1961), .B(G171), .ZN(n986) );
  NAND2_X1 U1079 ( .A1(G1971), .A2(G303), .ZN(n985) );
  NAND2_X1 U1080 ( .A1(n986), .A2(n985), .ZN(n993) );
  XNOR2_X1 U1081 ( .A(G299), .B(G1956), .ZN(n989) );
  XNOR2_X1 U1082 ( .A(n987), .B(G1348), .ZN(n988) );
  NOR2_X1 U1083 ( .A1(n989), .A2(n988), .ZN(n991) );
  NAND2_X1 U1084 ( .A1(n991), .A2(n990), .ZN(n992) );
  NOR2_X1 U1085 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1086 ( .A1(n995), .A2(n994), .ZN(n996) );
  NOR2_X1 U1087 ( .A1(n997), .A2(n996), .ZN(n998) );
  XOR2_X1 U1088 ( .A(KEYINPUT125), .B(n998), .Z(n1001) );
  XNOR2_X1 U1089 ( .A(n999), .B(G1341), .ZN(n1000) );
  NAND2_X1 U1090 ( .A1(n1001), .A2(n1000), .ZN(n1006) );
  XNOR2_X1 U1091 ( .A(G168), .B(G1966), .ZN(n1003) );
  NAND2_X1 U1092 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XOR2_X1 U1093 ( .A(KEYINPUT57), .B(n1004), .Z(n1005) );
  NOR2_X1 U1094 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1095 ( .A(n1007), .B(KEYINPUT126), .ZN(n1008) );
  NOR2_X1 U1096 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NOR2_X1 U1097 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1098 ( .A(n1012), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1099 ( .A(G311), .ZN(G150) );
endmodule

