//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 0 0 0 1 0 0 0 1 0 0 0 1 0 0 0 1 0 1 0 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 1 1 0 0 1 1 0 0 1 0 0 0 0 1 1 0 1 1 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:02 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n741, new_n742, new_n743, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n776, new_n777,
    new_n778, new_n779, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n792, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n816, new_n817,
    new_n818, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n869,
    new_n871, new_n873, new_n874, new_n875, new_n876, new_n877, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n931, new_n932, new_n933, new_n935, new_n936, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n955, new_n956,
    new_n957, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n967, new_n968, new_n969, new_n970, new_n971, new_n973,
    new_n974, new_n975, new_n976, new_n978, new_n979;
  XOR2_X1   g000(.A(G1gat), .B(G29gat), .Z(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT90), .B(KEYINPUT0), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(G57gat), .B(G85gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(G225gat), .A2(G233gat), .ZN(new_n208));
  OR2_X1    g007(.A1(KEYINPUT72), .A2(KEYINPUT1), .ZN(new_n209));
  XNOR2_X1  g008(.A(G127gat), .B(G134gat), .ZN(new_n210));
  XNOR2_X1  g009(.A(G113gat), .B(G120gat), .ZN(new_n211));
  OAI211_X1 g010(.A(new_n209), .B(new_n210), .C1(new_n211), .C2(KEYINPUT1), .ZN(new_n212));
  INV_X1    g011(.A(G120gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(G113gat), .ZN(new_n214));
  INV_X1    g013(.A(G113gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(G120gat), .ZN(new_n216));
  AOI21_X1  g015(.A(KEYINPUT1), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  AND2_X1   g016(.A1(G127gat), .A2(G134gat), .ZN(new_n218));
  NOR2_X1   g017(.A1(G127gat), .A2(G134gat), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n209), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n217), .A2(new_n220), .ZN(new_n221));
  AND2_X1   g020(.A1(new_n212), .A2(new_n221), .ZN(new_n222));
  XOR2_X1   g021(.A(G141gat), .B(G148gat), .Z(new_n223));
  NAND2_X1  g022(.A1(G155gat), .A2(G162gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(KEYINPUT2), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(G155gat), .ZN(new_n227));
  INV_X1    g026(.A(G162gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n229), .A2(KEYINPUT81), .A3(new_n224), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT81), .ZN(new_n231));
  AND2_X1   g030(.A1(G155gat), .A2(G162gat), .ZN(new_n232));
  NOR2_X1   g031(.A1(G155gat), .A2(G162gat), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n231), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n226), .A2(new_n230), .A3(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT85), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT82), .ZN(new_n238));
  NOR3_X1   g037(.A1(new_n232), .A2(new_n233), .A3(new_n238), .ZN(new_n239));
  AOI21_X1  g038(.A(KEYINPUT82), .B1(new_n229), .B2(new_n224), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n223), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT2), .ZN(new_n242));
  XOR2_X1   g041(.A(KEYINPUT83), .B(G155gat), .Z(new_n243));
  XNOR2_X1  g042(.A(KEYINPUT84), .B(G162gat), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n242), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n237), .B1(new_n241), .B2(new_n245), .ZN(new_n246));
  XOR2_X1   g045(.A(KEYINPUT84), .B(G162gat), .Z(new_n247));
  XNOR2_X1  g046(.A(KEYINPUT83), .B(G155gat), .ZN(new_n248));
  OAI21_X1  g047(.A(KEYINPUT2), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(G141gat), .B(G148gat), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n238), .B1(new_n232), .B2(new_n233), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n229), .A2(KEYINPUT82), .A3(new_n224), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n250), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n249), .A2(new_n253), .A3(KEYINPUT85), .ZN(new_n254));
  AOI211_X1 g053(.A(new_n222), .B(new_n236), .C1(new_n246), .C2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(KEYINPUT4), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n236), .B1(new_n246), .B2(new_n254), .ZN(new_n257));
  INV_X1    g056(.A(new_n222), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT4), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n256), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT88), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT86), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT3), .ZN(new_n266));
  NOR3_X1   g065(.A1(new_n257), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(KEYINPUT87), .B(KEYINPUT3), .ZN(new_n268));
  AND3_X1   g067(.A1(new_n249), .A2(new_n253), .A3(KEYINPUT85), .ZN(new_n269));
  AOI21_X1  g068(.A(KEYINPUT85), .B1(new_n249), .B2(new_n253), .ZN(new_n270));
  OAI211_X1 g069(.A(new_n235), .B(new_n268), .C1(new_n269), .C2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(new_n222), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n267), .A2(new_n272), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n265), .B1(new_n257), .B2(new_n266), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n264), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n258), .B1(new_n257), .B2(new_n268), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n235), .B1(new_n269), .B2(new_n270), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n277), .A2(KEYINPUT86), .A3(KEYINPUT3), .ZN(new_n278));
  NAND4_X1  g077(.A1(new_n274), .A2(new_n276), .A3(new_n278), .A4(new_n264), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  OAI211_X1 g079(.A(new_n208), .B(new_n263), .C1(new_n275), .C2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(new_n208), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n257), .A2(new_n258), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n282), .B1(new_n283), .B2(new_n255), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT89), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  OAI211_X1 g085(.A(KEYINPUT89), .B(new_n282), .C1(new_n283), .C2(new_n255), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n286), .A2(new_n287), .A3(KEYINPUT5), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n281), .A2(new_n289), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n274), .A2(new_n276), .A3(new_n278), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(KEYINPUT88), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(new_n279), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT5), .ZN(new_n294));
  NAND4_X1  g093(.A1(new_n293), .A2(new_n294), .A3(new_n208), .A4(new_n263), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n207), .B1(new_n290), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(KEYINPUT6), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n290), .A2(new_n207), .A3(new_n295), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT6), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n297), .B1(new_n300), .B2(new_n296), .ZN(new_n301));
  NAND2_X1  g100(.A1(G183gat), .A2(G190gat), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT66), .ZN(new_n303));
  AOI21_X1  g102(.A(KEYINPUT24), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n304), .B1(new_n303), .B2(new_n302), .ZN(new_n305));
  XNOR2_X1  g104(.A(KEYINPUT68), .B(G183gat), .ZN(new_n306));
  INV_X1    g105(.A(G190gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g107(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n309));
  OR2_X1    g108(.A1(new_n309), .A2(KEYINPUT67), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(KEYINPUT67), .ZN(new_n311));
  NAND4_X1  g110(.A1(new_n305), .A2(new_n308), .A3(new_n310), .A4(new_n311), .ZN(new_n312));
  NOR2_X1   g111(.A1(G169gat), .A2(G176gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(KEYINPUT23), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(KEYINPUT25), .ZN(new_n315));
  NAND2_X1  g114(.A1(G169gat), .A2(G176gat), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n313), .B1(KEYINPUT23), .B2(new_n316), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n312), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(KEYINPUT69), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT69), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n312), .A2(new_n321), .A3(new_n318), .ZN(new_n322));
  INV_X1    g121(.A(new_n317), .ZN(new_n323));
  OR2_X1    g122(.A1(G183gat), .A2(G190gat), .ZN(new_n324));
  INV_X1    g123(.A(new_n302), .ZN(new_n325));
  OAI211_X1 g124(.A(new_n309), .B(new_n324), .C1(new_n325), .C2(KEYINPUT24), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n314), .A2(KEYINPUT65), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT65), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n328), .B1(new_n313), .B2(KEYINPUT23), .ZN(new_n329));
  OAI211_X1 g128(.A(new_n323), .B(new_n326), .C1(new_n327), .C2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT25), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n320), .A2(new_n322), .A3(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n316), .ZN(new_n334));
  NOR3_X1   g133(.A1(new_n334), .A2(new_n313), .A3(KEYINPUT26), .ZN(new_n335));
  AND2_X1   g134(.A1(new_n313), .A2(KEYINPUT26), .ZN(new_n336));
  NOR3_X1   g135(.A1(new_n335), .A2(new_n336), .A3(new_n325), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(KEYINPUT71), .B(KEYINPUT28), .ZN(new_n339));
  INV_X1    g138(.A(new_n306), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT27), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(G183gat), .ZN(new_n343));
  AOI21_X1  g142(.A(G190gat), .B1(new_n343), .B2(KEYINPUT70), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n344), .B1(KEYINPUT70), .B2(new_n343), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n339), .B1(new_n342), .B2(new_n345), .ZN(new_n346));
  XNOR2_X1  g145(.A(KEYINPUT27), .B(G183gat), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n347), .A2(KEYINPUT28), .A3(new_n307), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n338), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  AOI21_X1  g149(.A(KEYINPUT29), .B1(new_n333), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(G226gat), .A2(G233gat), .ZN(new_n352));
  XNOR2_X1  g151(.A(new_n352), .B(KEYINPUT75), .ZN(new_n353));
  OAI21_X1  g152(.A(KEYINPUT77), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  XNOR2_X1  g153(.A(G197gat), .B(G204gat), .ZN(new_n355));
  INV_X1    g154(.A(G211gat), .ZN(new_n356));
  INV_X1    g155(.A(G218gat), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n355), .B1(KEYINPUT22), .B2(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(G211gat), .B(G218gat), .ZN(new_n360));
  XNOR2_X1  g159(.A(new_n359), .B(new_n360), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n361), .B(KEYINPUT74), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n333), .A2(new_n350), .ZN(new_n363));
  XNOR2_X1  g162(.A(new_n353), .B(KEYINPUT76), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT77), .ZN(new_n366));
  INV_X1    g165(.A(new_n353), .ZN(new_n367));
  AOI22_X1  g166(.A1(new_n319), .A2(KEYINPUT69), .B1(new_n331), .B2(new_n330), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n349), .B1(new_n368), .B2(new_n322), .ZN(new_n369));
  OAI211_X1 g168(.A(new_n366), .B(new_n367), .C1(new_n369), .C2(KEYINPUT29), .ZN(new_n370));
  NAND4_X1  g169(.A1(new_n354), .A2(new_n362), .A3(new_n365), .A4(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n362), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT29), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n364), .B1(new_n363), .B2(new_n373), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n369), .A2(new_n367), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n372), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  XOR2_X1   g175(.A(G8gat), .B(G36gat), .Z(new_n377));
  XNOR2_X1  g176(.A(new_n377), .B(KEYINPUT78), .ZN(new_n378));
  XNOR2_X1  g177(.A(G64gat), .B(G92gat), .ZN(new_n379));
  XNOR2_X1  g178(.A(new_n378), .B(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  AND2_X1   g180(.A1(new_n381), .A2(KEYINPUT30), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n371), .A2(new_n376), .A3(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT79), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND4_X1  g184(.A1(new_n371), .A2(new_n376), .A3(KEYINPUT79), .A4(new_n382), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n371), .A2(new_n376), .A3(new_n381), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n381), .B1(new_n371), .B2(new_n376), .ZN(new_n389));
  XNOR2_X1  g188(.A(KEYINPUT80), .B(KEYINPUT30), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n388), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n387), .A2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n301), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n363), .A2(new_n258), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n369), .A2(new_n222), .ZN(new_n398));
  NAND2_X1  g197(.A1(G227gat), .A2(G233gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n399), .B(KEYINPUT64), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n397), .A2(new_n398), .A3(new_n400), .ZN(new_n401));
  XOR2_X1   g200(.A(G71gat), .B(G99gat), .Z(new_n402));
  XNOR2_X1  g201(.A(G15gat), .B(G43gat), .ZN(new_n403));
  XNOR2_X1  g202(.A(new_n402), .B(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(KEYINPUT33), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n401), .A2(KEYINPUT32), .A3(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT73), .ZN(new_n407));
  XNOR2_X1  g206(.A(new_n406), .B(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n397), .A2(new_n398), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(new_n399), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(KEYINPUT34), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n400), .A2(KEYINPUT34), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n409), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n401), .A2(KEYINPUT32), .ZN(new_n416));
  INV_X1    g215(.A(new_n401), .ZN(new_n417));
  OAI211_X1 g216(.A(new_n416), .B(new_n404), .C1(new_n417), .C2(KEYINPUT33), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n408), .A2(new_n415), .A3(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n415), .B1(new_n408), .B2(new_n418), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(G22gat), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n362), .B1(new_n373), .B2(new_n271), .ZN(new_n424));
  INV_X1    g223(.A(new_n361), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n277), .A2(new_n373), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n277), .A2(KEYINPUT3), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n426), .A2(new_n427), .A3(G228gat), .A4(G233gat), .ZN(new_n428));
  OR2_X1    g227(.A1(new_n424), .A2(new_n428), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n426), .B1(new_n257), .B2(new_n268), .ZN(new_n430));
  INV_X1    g229(.A(G228gat), .ZN(new_n431));
  INV_X1    g230(.A(G233gat), .ZN(new_n432));
  OAI22_X1  g231(.A1(new_n424), .A2(new_n430), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n423), .B1(new_n429), .B2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n429), .A2(new_n433), .A3(new_n423), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  XNOR2_X1  g236(.A(G78gat), .B(G106gat), .ZN(new_n438));
  XNOR2_X1  g237(.A(KEYINPUT31), .B(G50gat), .ZN(new_n439));
  XNOR2_X1  g238(.A(new_n438), .B(new_n439), .ZN(new_n440));
  XOR2_X1   g239(.A(new_n440), .B(KEYINPUT91), .Z(new_n441));
  NAND2_X1  g240(.A1(new_n437), .A2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT92), .ZN(new_n443));
  OAI211_X1 g242(.A(new_n440), .B(new_n436), .C1(new_n434), .C2(new_n443), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n435), .A2(KEYINPUT92), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n442), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  AND2_X1   g245(.A1(new_n422), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n396), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(KEYINPUT35), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT97), .ZN(new_n450));
  AOI211_X1 g249(.A(new_n299), .B(new_n207), .C1(new_n290), .C2(new_n295), .ZN(new_n451));
  AOI211_X1 g250(.A(new_n282), .B(new_n262), .C1(new_n292), .C2(new_n279), .ZN(new_n452));
  OAI211_X1 g251(.A(new_n295), .B(KEYINPUT94), .C1(new_n452), .C2(new_n288), .ZN(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(KEYINPUT94), .B1(new_n290), .B2(new_n295), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n206), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(new_n300), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n451), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n387), .A2(KEYINPUT93), .A3(new_n392), .ZN(new_n459));
  INV_X1    g258(.A(new_n459), .ZN(new_n460));
  AOI21_X1  g259(.A(KEYINPUT93), .B1(new_n387), .B2(new_n392), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n450), .B1(new_n458), .B2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT35), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT94), .ZN(new_n465));
  INV_X1    g264(.A(new_n295), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n262), .B1(new_n292), .B2(new_n279), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n288), .B1(new_n467), .B2(new_n208), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n465), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n207), .B1(new_n469), .B2(new_n453), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n297), .B1(new_n470), .B2(new_n300), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT93), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n393), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(new_n459), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n471), .A2(KEYINPUT97), .A3(new_n474), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n463), .A2(new_n464), .A3(new_n447), .A4(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(new_n446), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n374), .A2(new_n375), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n478), .A2(KEYINPUT96), .A3(new_n362), .ZN(new_n479));
  OAI221_X1 g278(.A(new_n362), .B1(new_n369), .B2(new_n367), .C1(new_n351), .C2(new_n364), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT96), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n479), .A2(new_n482), .ZN(new_n483));
  AND2_X1   g282(.A1(new_n370), .A2(new_n365), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n362), .B1(new_n484), .B2(new_n354), .ZN(new_n485));
  OAI21_X1  g284(.A(KEYINPUT37), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT38), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT37), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n381), .A2(new_n488), .ZN(new_n489));
  OAI211_X1 g288(.A(new_n486), .B(new_n487), .C1(new_n389), .C2(new_n489), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n389), .A2(new_n489), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n488), .B1(new_n371), .B2(new_n376), .ZN(new_n492));
  OAI21_X1  g291(.A(KEYINPUT38), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  AND3_X1   g292(.A1(new_n490), .A2(new_n388), .A3(new_n493), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n477), .B1(new_n458), .B2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(new_n467), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT39), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n496), .A2(new_n497), .A3(new_n282), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n283), .A2(new_n255), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n497), .B1(new_n499), .B2(new_n208), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n500), .B1(new_n467), .B2(new_n208), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n498), .A2(new_n207), .A3(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT40), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n498), .A2(new_n501), .A3(KEYINPUT40), .A4(new_n207), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n506), .A2(new_n470), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n507), .A2(KEYINPUT95), .A3(new_n462), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT95), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n456), .A2(new_n505), .A3(new_n504), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n509), .B1(new_n510), .B2(new_n474), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n495), .A2(new_n508), .A3(new_n511), .ZN(new_n512));
  OAI21_X1  g311(.A(KEYINPUT36), .B1(new_n420), .B2(new_n421), .ZN(new_n513));
  INV_X1    g312(.A(new_n421), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT36), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n514), .A2(new_n515), .A3(new_n419), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n513), .A2(new_n516), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n517), .B1(new_n395), .B2(new_n477), .ZN(new_n518));
  AOI22_X1  g317(.A1(new_n449), .A2(new_n476), .B1(new_n512), .B2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT106), .ZN(new_n520));
  XNOR2_X1  g319(.A(G15gat), .B(G22gat), .ZN(new_n521));
  INV_X1    g320(.A(G1gat), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n521), .A2(KEYINPUT16), .A3(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT101), .ZN(new_n524));
  OR2_X1    g323(.A1(new_n524), .A2(G8gat), .ZN(new_n525));
  OAI211_X1 g324(.A(new_n523), .B(new_n525), .C1(new_n522), .C2(new_n521), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n524), .A2(G8gat), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n526), .B(new_n527), .ZN(new_n528));
  XNOR2_X1  g327(.A(G43gat), .B(G50gat), .ZN(new_n529));
  AND2_X1   g328(.A1(new_n529), .A2(KEYINPUT15), .ZN(new_n530));
  NAND2_X1  g329(.A1(G29gat), .A2(G36gat), .ZN(new_n531));
  NOR3_X1   g330(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n532));
  OAI21_X1  g331(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(KEYINPUT98), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT98), .ZN(new_n535));
  OAI211_X1 g334(.A(new_n535), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n532), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n531), .B1(new_n537), .B2(KEYINPUT99), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT99), .ZN(new_n539));
  AOI211_X1 g338(.A(new_n539), .B(new_n532), .C1(new_n534), .C2(new_n536), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n530), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  AOI22_X1  g340(.A1(new_n529), .A2(KEYINPUT15), .B1(G29gat), .B2(G36gat), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT100), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n532), .B(new_n543), .ZN(new_n544));
  AND2_X1   g343(.A1(new_n534), .A2(new_n536), .ZN(new_n545));
  OAI221_X1 g344(.A(new_n542), .B1(KEYINPUT15), .B2(new_n529), .C1(new_n544), .C2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n541), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n528), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(G229gat), .A2(G233gat), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n541), .A2(new_n546), .A3(KEYINPUT17), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(KEYINPUT102), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT102), .ZN(new_n554));
  NAND4_X1  g353(.A1(new_n541), .A2(new_n546), .A3(new_n554), .A4(KEYINPUT17), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT103), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT17), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n528), .B1(new_n558), .B2(new_n547), .ZN(new_n559));
  AND3_X1   g358(.A1(new_n556), .A2(new_n557), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n557), .B1(new_n556), .B2(new_n559), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n551), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT105), .ZN(new_n563));
  XNOR2_X1  g362(.A(KEYINPUT104), .B(KEYINPUT18), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n562), .A2(new_n563), .A3(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n528), .B(new_n547), .ZN(new_n568));
  XOR2_X1   g367(.A(new_n549), .B(KEYINPUT13), .Z(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(G113gat), .B(G141gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n571), .B(G197gat), .ZN(new_n572));
  XOR2_X1   g371(.A(KEYINPUT11), .B(G169gat), .Z(new_n573));
  XNOR2_X1  g372(.A(new_n572), .B(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n574), .B(KEYINPUT12), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT18), .ZN(new_n576));
  OAI211_X1 g375(.A(new_n570), .B(new_n575), .C1(new_n562), .C2(new_n576), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n563), .B1(new_n562), .B2(new_n565), .ZN(new_n578));
  NOR3_X1   g377(.A1(new_n567), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n556), .A2(new_n559), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n580), .A2(KEYINPUT103), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n556), .A2(new_n559), .A3(new_n557), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n550), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  AOI22_X1  g382(.A1(new_n583), .A2(KEYINPUT18), .B1(new_n568), .B2(new_n569), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n562), .A2(new_n565), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n575), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n520), .B1(new_n579), .B2(new_n586), .ZN(new_n587));
  OAI21_X1  g386(.A(KEYINPUT105), .B1(new_n583), .B2(new_n564), .ZN(new_n588));
  NAND4_X1  g387(.A1(new_n584), .A2(new_n588), .A3(new_n575), .A4(new_n566), .ZN(new_n589));
  INV_X1    g388(.A(new_n575), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n570), .B1(new_n562), .B2(new_n576), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n583), .A2(new_n564), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n590), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n589), .A2(new_n593), .A3(KEYINPUT106), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n587), .A2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n519), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(G85gat), .A2(G92gat), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n598), .B(KEYINPUT7), .ZN(new_n599));
  NOR2_X1   g398(.A1(G85gat), .A2(G92gat), .ZN(new_n600));
  NAND2_X1  g399(.A1(G99gat), .A2(G106gat), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n600), .B1(KEYINPUT8), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n599), .A2(new_n602), .ZN(new_n603));
  XOR2_X1   g402(.A(G99gat), .B(G106gat), .Z(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n603), .A2(new_n604), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(KEYINPUT109), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT109), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n610), .B1(new_n606), .B2(new_n607), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n547), .ZN(new_n613));
  OAI211_X1 g412(.A(new_n556), .B(new_n612), .C1(KEYINPUT17), .C2(new_n613), .ZN(new_n614));
  XOR2_X1   g413(.A(G190gat), .B(G218gat), .Z(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  AND2_X1   g415(.A1(G232gat), .A2(G233gat), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n617), .A2(KEYINPUT41), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n618), .B1(new_n612), .B2(new_n613), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  AND3_X1   g419(.A1(new_n614), .A2(new_n616), .A3(new_n620), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n616), .B1(new_n614), .B2(new_n620), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n617), .A2(KEYINPUT41), .ZN(new_n623));
  XNOR2_X1  g422(.A(G134gat), .B(G162gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n623), .B(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  OR3_X1    g425(.A1(new_n621), .A2(new_n622), .A3(new_n626), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n626), .B1(new_n621), .B2(new_n622), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  XOR2_X1   g428(.A(G71gat), .B(G78gat), .Z(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT9), .ZN(new_n632));
  INV_X1    g431(.A(G71gat), .ZN(new_n633));
  INV_X1    g432(.A(G78gat), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n632), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  XOR2_X1   g434(.A(G57gat), .B(G64gat), .Z(new_n636));
  NAND3_X1  g435(.A1(new_n631), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n635), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n638), .A2(new_n630), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT21), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g441(.A(KEYINPUT108), .B(KEYINPUT19), .Z(new_n643));
  XOR2_X1   g442(.A(new_n642), .B(new_n643), .Z(new_n644));
  INV_X1    g443(.A(new_n528), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n645), .B1(new_n641), .B2(new_n640), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n644), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(G127gat), .B(G155gat), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n648), .B(KEYINPUT20), .ZN(new_n649));
  NAND2_X1  g448(.A1(G231gat), .A2(G233gat), .ZN(new_n650));
  XOR2_X1   g449(.A(new_n650), .B(KEYINPUT107), .Z(new_n651));
  XNOR2_X1  g450(.A(new_n649), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(G183gat), .B(G211gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n647), .B(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n629), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(G230gat), .A2(G233gat), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n640), .B1(new_n606), .B2(new_n607), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(KEYINPUT110), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n640), .A2(new_n607), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n606), .A2(KEYINPUT111), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT111), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n605), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n661), .A2(new_n662), .A3(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT10), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT110), .ZN(new_n667));
  OAI211_X1 g466(.A(new_n667), .B(new_n640), .C1(new_n606), .C2(new_n607), .ZN(new_n668));
  NAND4_X1  g467(.A1(new_n660), .A2(new_n665), .A3(new_n666), .A4(new_n668), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n640), .A2(new_n666), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n609), .A2(new_n611), .A3(new_n670), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n658), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n660), .A2(new_n665), .A3(new_n668), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n672), .B1(new_n658), .B2(new_n673), .ZN(new_n674));
  XNOR2_X1  g473(.A(G120gat), .B(G148gat), .ZN(new_n675));
  XNOR2_X1  g474(.A(G176gat), .B(G204gat), .ZN(new_n676));
  XOR2_X1   g475(.A(new_n675), .B(new_n676), .Z(new_n677));
  OR2_X1    g476(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n669), .A2(new_n671), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n679), .A2(new_n657), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n673), .A2(new_n658), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n680), .A2(new_n681), .A3(new_n677), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n678), .A2(new_n682), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n656), .A2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT112), .ZN(new_n685));
  OR2_X1    g484(.A1(new_n301), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n301), .A2(new_n685), .ZN(new_n687));
  AND2_X1   g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n597), .A2(new_n684), .A3(new_n688), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(G1gat), .ZN(G1324gat));
  NAND3_X1  g489(.A1(new_n597), .A2(new_n684), .A3(new_n462), .ZN(new_n691));
  AND2_X1   g490(.A1(new_n691), .A2(G8gat), .ZN(new_n692));
  XNOR2_X1  g491(.A(KEYINPUT16), .B(G8gat), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  OAI21_X1  g493(.A(KEYINPUT42), .B1(new_n692), .B2(new_n694), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n695), .B1(KEYINPUT42), .B2(new_n694), .ZN(G1325gat));
  INV_X1    g495(.A(G15gat), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n476), .A2(new_n449), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n512), .A2(new_n518), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(new_n595), .ZN(new_n701));
  INV_X1    g500(.A(new_n684), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n697), .B1(new_n703), .B2(new_n517), .ZN(new_n704));
  INV_X1    g503(.A(new_n422), .ZN(new_n705));
  NOR4_X1   g504(.A1(new_n701), .A2(G15gat), .A3(new_n702), .A4(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT113), .ZN(new_n707));
  OR3_X1    g506(.A1(new_n704), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n707), .B1(new_n704), .B2(new_n706), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(G1326gat));
  NAND2_X1  g509(.A1(new_n703), .A2(new_n477), .ZN(new_n711));
  XNOR2_X1  g510(.A(KEYINPUT43), .B(G22gat), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n711), .B(new_n712), .ZN(G1327gat));
  INV_X1    g512(.A(KEYINPUT44), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n714), .B1(new_n519), .B2(new_n629), .ZN(new_n715));
  INV_X1    g514(.A(new_n629), .ZN(new_n716));
  AND2_X1   g515(.A1(new_n513), .A2(new_n516), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n717), .B1(new_n396), .B2(new_n446), .ZN(new_n718));
  AOI21_X1  g517(.A(KEYINPUT95), .B1(new_n507), .B2(new_n462), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n490), .A2(new_n388), .A3(new_n493), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n446), .B1(new_n471), .B2(new_n720), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n718), .B1(new_n722), .B2(new_n508), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n422), .A2(new_n464), .A3(new_n446), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n471), .A2(new_n474), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n724), .B1(new_n725), .B2(new_n450), .ZN(new_n726));
  AOI22_X1  g525(.A1(new_n726), .A2(new_n475), .B1(new_n448), .B2(KEYINPUT35), .ZN(new_n727));
  OAI211_X1 g526(.A(KEYINPUT44), .B(new_n716), .C1(new_n723), .C2(new_n727), .ZN(new_n728));
  AND2_X1   g527(.A1(new_n715), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n579), .A2(new_n586), .ZN(new_n730));
  NOR3_X1   g529(.A1(new_n730), .A2(new_n655), .A3(new_n683), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(new_n688), .ZN(new_n733));
  OAI21_X1  g532(.A(G29gat), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n683), .A2(new_n655), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n716), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n736), .A2(G29gat), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n597), .A2(new_n688), .A3(new_n737), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(KEYINPUT45), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n734), .A2(new_n739), .ZN(G1328gat));
  NOR4_X1   g539(.A1(new_n701), .A2(G36gat), .A3(new_n474), .A4(new_n736), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(KEYINPUT46), .ZN(new_n742));
  OAI21_X1  g541(.A(G36gat), .B1(new_n732), .B2(new_n474), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(G1329gat));
  NOR2_X1   g543(.A1(new_n736), .A2(G43gat), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n700), .A2(new_n422), .A3(new_n595), .A4(new_n745), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(KEYINPUT114), .ZN(new_n747));
  INV_X1    g546(.A(new_n747), .ZN(new_n748));
  NAND4_X1  g547(.A1(new_n715), .A2(new_n517), .A3(new_n728), .A4(new_n731), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(G43gat), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n748), .A2(KEYINPUT47), .A3(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT47), .ZN(new_n752));
  INV_X1    g551(.A(new_n750), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n752), .B1(new_n753), .B2(new_n747), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n751), .A2(new_n754), .ZN(G1330gat));
  OR2_X1    g554(.A1(new_n446), .A2(G50gat), .ZN(new_n756));
  INV_X1    g555(.A(new_n756), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n736), .B1(new_n757), .B2(KEYINPUT115), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n758), .B1(KEYINPUT115), .B2(new_n757), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n701), .A2(new_n759), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n715), .A2(new_n477), .A3(new_n728), .A4(new_n731), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n760), .B1(new_n761), .B2(G50gat), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT48), .ZN(new_n763));
  AND3_X1   g562(.A1(new_n762), .A2(KEYINPUT116), .A3(new_n763), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n763), .A2(KEYINPUT116), .ZN(new_n765));
  AND2_X1   g564(.A1(new_n763), .A2(KEYINPUT116), .ZN(new_n766));
  NOR3_X1   g565(.A1(new_n762), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n764), .A2(new_n767), .ZN(G1331gat));
  INV_X1    g567(.A(new_n730), .ZN(new_n769));
  INV_X1    g568(.A(new_n683), .ZN(new_n770));
  NOR3_X1   g569(.A1(new_n769), .A2(new_n656), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n700), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n772), .A2(new_n733), .ZN(new_n773));
  XOR2_X1   g572(.A(KEYINPUT117), .B(G57gat), .Z(new_n774));
  XNOR2_X1  g573(.A(new_n773), .B(new_n774), .ZN(G1332gat));
  NOR2_X1   g574(.A1(new_n772), .A2(new_n474), .ZN(new_n776));
  NOR2_X1   g575(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n777));
  AND2_X1   g576(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n776), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n779), .B1(new_n776), .B2(new_n777), .ZN(G1333gat));
  INV_X1    g579(.A(new_n772), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT118), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n781), .A2(new_n782), .A3(new_n422), .ZN(new_n783));
  OAI21_X1  g582(.A(KEYINPUT118), .B1(new_n772), .B2(new_n705), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n783), .A2(new_n633), .A3(new_n784), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n781), .A2(G71gat), .A3(new_n517), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(KEYINPUT50), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT50), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n785), .A2(new_n789), .A3(new_n786), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n788), .A2(new_n790), .ZN(G1334gat));
  NOR2_X1   g590(.A1(new_n772), .A2(new_n446), .ZN(new_n792));
  XNOR2_X1  g591(.A(new_n792), .B(new_n634), .ZN(G1335gat));
  AOI21_X1  g592(.A(new_n629), .B1(new_n698), .B2(new_n699), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n769), .A2(new_n655), .ZN(new_n795));
  AOI21_X1  g594(.A(KEYINPUT51), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT51), .ZN(new_n797));
  INV_X1    g596(.A(new_n795), .ZN(new_n798));
  NOR4_X1   g597(.A1(new_n519), .A2(new_n797), .A3(new_n629), .A4(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT119), .ZN(new_n800));
  OR3_X1    g599(.A1(new_n796), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n800), .B1(new_n796), .B2(new_n799), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n733), .A2(G85gat), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n801), .A2(new_n683), .A3(new_n802), .A4(new_n803), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n798), .A2(new_n770), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n729), .A2(new_n805), .ZN(new_n806));
  OAI21_X1  g605(.A(G85gat), .B1(new_n806), .B2(new_n733), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n804), .A2(new_n807), .ZN(G1336gat));
  NAND4_X1  g607(.A1(new_n715), .A2(new_n462), .A3(new_n728), .A4(new_n805), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(G92gat), .ZN(new_n810));
  NOR3_X1   g609(.A1(new_n474), .A2(G92gat), .A3(new_n770), .ZN(new_n811));
  XNOR2_X1  g610(.A(new_n811), .B(KEYINPUT120), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n812), .B1(new_n796), .B2(new_n799), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n810), .A2(new_n813), .ZN(new_n814));
  XNOR2_X1  g613(.A(new_n814), .B(KEYINPUT52), .ZN(G1337gat));
  NOR2_X1   g614(.A1(new_n705), .A2(G99gat), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n801), .A2(new_n683), .A3(new_n802), .A4(new_n816), .ZN(new_n817));
  OAI21_X1  g616(.A(G99gat), .B1(new_n806), .B2(new_n717), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(G1338gat));
  NOR2_X1   g618(.A1(new_n770), .A2(G106gat), .ZN(new_n820));
  OAI211_X1 g619(.A(new_n477), .B(new_n820), .C1(new_n796), .C2(new_n799), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n715), .A2(new_n477), .A3(new_n728), .A4(new_n805), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(G106gat), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT121), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n821), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n824), .A2(new_n826), .A3(KEYINPUT53), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT53), .ZN(new_n828));
  OAI211_X1 g627(.A(new_n821), .B(new_n823), .C1(new_n825), .C2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n827), .A2(new_n829), .ZN(G1339gat));
  INV_X1    g629(.A(KEYINPUT122), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n669), .A2(new_n671), .A3(new_n658), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n680), .A2(KEYINPUT54), .A3(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT54), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n677), .B1(new_n672), .B2(new_n834), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n833), .A2(KEYINPUT55), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(new_n682), .ZN(new_n837));
  AOI21_X1  g636(.A(KEYINPUT55), .B1(new_n833), .B2(new_n835), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n831), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(new_n838), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n840), .A2(KEYINPUT122), .A3(new_n682), .A4(new_n836), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n730), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n581), .A2(new_n582), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n549), .B1(new_n844), .B2(new_n548), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n568), .A2(new_n569), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n574), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  AND3_X1   g646(.A1(new_n589), .A2(new_n683), .A3(new_n847), .ZN(new_n848));
  OAI21_X1  g647(.A(KEYINPUT123), .B1(new_n843), .B2(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(new_n848), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT123), .ZN(new_n851));
  OAI211_X1 g650(.A(new_n850), .B(new_n851), .C1(new_n730), .C2(new_n842), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n849), .A2(new_n852), .A3(new_n629), .ZN(new_n853));
  INV_X1    g652(.A(new_n842), .ZN(new_n854));
  AND2_X1   g653(.A1(new_n589), .A2(new_n847), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n854), .A2(new_n716), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n655), .B1(new_n853), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n684), .A2(new_n730), .ZN(new_n858));
  INV_X1    g657(.A(new_n858), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(new_n447), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n733), .A2(new_n462), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NOR3_X1   g663(.A1(new_n864), .A2(new_n215), .A3(new_n596), .ZN(new_n865));
  INV_X1    g664(.A(new_n864), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(new_n769), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n865), .B1(new_n215), .B2(new_n867), .ZN(G1340gat));
  NOR2_X1   g667(.A1(new_n864), .A2(new_n770), .ZN(new_n869));
  XNOR2_X1  g668(.A(new_n869), .B(new_n213), .ZN(G1341gat));
  NAND2_X1  g669(.A1(new_n866), .A2(new_n655), .ZN(new_n871));
  XNOR2_X1  g670(.A(new_n871), .B(G127gat), .ZN(G1342gat));
  NOR2_X1   g671(.A1(new_n462), .A2(new_n629), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n733), .A2(G134gat), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n862), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  XOR2_X1   g674(.A(new_n875), .B(KEYINPUT56), .Z(new_n876));
  OAI21_X1  g675(.A(G134gat), .B1(new_n864), .B2(new_n629), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(G1343gat));
  OAI21_X1  g677(.A(new_n477), .B1(new_n857), .B2(new_n859), .ZN(new_n879));
  INV_X1    g678(.A(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n863), .A2(new_n717), .ZN(new_n881));
  INV_X1    g680(.A(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(G141gat), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n595), .A2(new_n884), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  XNOR2_X1  g685(.A(KEYINPUT124), .B(KEYINPUT57), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n879), .A2(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT57), .ZN(new_n889));
  INV_X1    g688(.A(new_n655), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n837), .A2(new_n838), .ZN(new_n891));
  AND3_X1   g690(.A1(new_n589), .A2(KEYINPUT106), .A3(new_n593), .ZN(new_n892));
  AOI21_X1  g691(.A(KEYINPUT106), .B1(new_n589), .B2(new_n593), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n891), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n716), .B1(new_n894), .B2(new_n850), .ZN(new_n895));
  INV_X1    g694(.A(new_n856), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n890), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  AOI211_X1 g696(.A(new_n889), .B(new_n446), .C1(new_n897), .C2(new_n858), .ZN(new_n898));
  INV_X1    g697(.A(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n888), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n900), .A2(new_n769), .A3(new_n882), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n886), .B1(new_n901), .B2(G141gat), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT58), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n881), .B1(new_n888), .B2(new_n899), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n884), .B1(new_n904), .B2(new_n595), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n903), .B1(new_n883), .B2(new_n885), .ZN(new_n906));
  OAI22_X1  g705(.A1(new_n902), .A2(new_n903), .B1(new_n905), .B2(new_n906), .ZN(G1344gat));
  OR3_X1    g706(.A1(new_n883), .A2(G148gat), .A3(new_n770), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT59), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT125), .ZN(new_n910));
  NOR3_X1   g709(.A1(new_n629), .A2(new_n838), .A3(new_n837), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n911), .A2(new_n855), .ZN(new_n912));
  INV_X1    g711(.A(new_n912), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n890), .B1(new_n895), .B2(new_n913), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n702), .A2(new_n595), .ZN(new_n915));
  INV_X1    g714(.A(new_n915), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n446), .B1(new_n914), .B2(new_n916), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n910), .B1(new_n917), .B2(KEYINPUT57), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n848), .B1(new_n595), .B2(new_n891), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n912), .B1(new_n919), .B2(new_n716), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n915), .B1(new_n920), .B2(new_n890), .ZN(new_n921));
  OAI211_X1 g720(.A(KEYINPUT125), .B(new_n889), .C1(new_n921), .C2(new_n446), .ZN(new_n922));
  INV_X1    g721(.A(new_n887), .ZN(new_n923));
  OAI211_X1 g722(.A(new_n477), .B(new_n923), .C1(new_n857), .C2(new_n859), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n918), .A2(new_n922), .A3(new_n924), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n925), .A2(new_n683), .A3(new_n882), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n909), .B1(new_n926), .B2(G148gat), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n909), .A2(G148gat), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n928), .B1(new_n904), .B2(new_n683), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n908), .B1(new_n927), .B2(new_n929), .ZN(G1345gat));
  INV_X1    g729(.A(new_n904), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n243), .B1(new_n931), .B2(new_n890), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n655), .A2(new_n248), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n932), .B1(new_n883), .B2(new_n933), .ZN(G1346gat));
  OAI21_X1  g733(.A(new_n244), .B1(new_n931), .B2(new_n629), .ZN(new_n935));
  NAND4_X1  g734(.A1(new_n688), .A2(new_n247), .A3(new_n717), .A4(new_n873), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n935), .B1(new_n879), .B2(new_n936), .ZN(G1347gat));
  NAND2_X1  g736(.A1(new_n733), .A2(new_n462), .ZN(new_n938));
  NOR3_X1   g737(.A1(new_n860), .A2(new_n861), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g738(.A(G169gat), .B1(new_n939), .B2(new_n769), .ZN(new_n940));
  AND2_X1   g739(.A1(new_n595), .A2(G169gat), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n940), .B1(new_n939), .B2(new_n941), .ZN(G1348gat));
  NAND2_X1  g741(.A1(new_n939), .A2(new_n683), .ZN(new_n943));
  XNOR2_X1  g742(.A(new_n943), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g743(.A1(new_n939), .A2(new_n655), .ZN(new_n945));
  OR2_X1    g744(.A1(new_n306), .A2(KEYINPUT126), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n347), .B1(new_n340), .B2(KEYINPUT126), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n939), .A2(new_n655), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT60), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n947), .A2(KEYINPUT60), .A3(new_n949), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n952), .A2(new_n953), .ZN(G1350gat));
  NOR2_X1   g753(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n955), .B1(new_n939), .B2(new_n716), .ZN(new_n956));
  NAND2_X1  g755(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n957));
  XOR2_X1   g756(.A(new_n956), .B(new_n957), .Z(G1351gat));
  NOR2_X1   g757(.A1(new_n938), .A2(new_n517), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n880), .A2(new_n959), .ZN(new_n960));
  INV_X1    g759(.A(new_n960), .ZN(new_n961));
  XOR2_X1   g760(.A(KEYINPUT127), .B(G197gat), .Z(new_n962));
  NAND3_X1  g761(.A1(new_n961), .A2(new_n769), .A3(new_n962), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n925), .A2(new_n959), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n964), .A2(new_n596), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n963), .B1(new_n965), .B2(new_n962), .ZN(G1352gat));
  OAI21_X1  g765(.A(G204gat), .B1(new_n964), .B2(new_n770), .ZN(new_n967));
  NOR2_X1   g766(.A1(new_n770), .A2(G204gat), .ZN(new_n968));
  INV_X1    g767(.A(new_n968), .ZN(new_n969));
  OAI21_X1  g768(.A(KEYINPUT62), .B1(new_n960), .B2(new_n969), .ZN(new_n970));
  OR3_X1    g769(.A1(new_n960), .A2(KEYINPUT62), .A3(new_n969), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n967), .A2(new_n970), .A3(new_n971), .ZN(G1353gat));
  NAND3_X1  g771(.A1(new_n961), .A2(new_n356), .A3(new_n655), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n925), .A2(new_n655), .A3(new_n959), .ZN(new_n974));
  AND3_X1   g773(.A1(new_n974), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n975));
  AOI21_X1  g774(.A(KEYINPUT63), .B1(new_n974), .B2(G211gat), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n973), .B1(new_n975), .B2(new_n976), .ZN(G1354gat));
  OAI21_X1  g776(.A(G218gat), .B1(new_n964), .B2(new_n629), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n961), .A2(new_n357), .A3(new_n716), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n978), .A2(new_n979), .ZN(G1355gat));
endmodule


