

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X1 U554 ( .A1(n733), .A2(n732), .ZN(n736) );
  NOR2_X1 U555 ( .A1(n542), .A2(n541), .ZN(G160) );
  XNOR2_X1 U556 ( .A(n716), .B(KEYINPUT31), .ZN(n717) );
  XNOR2_X1 U557 ( .A(n718), .B(n717), .ZN(n747) );
  INV_X1 U558 ( .A(KEYINPUT97), .ZN(n764) );
  NAND2_X1 U559 ( .A1(G8), .A2(n751), .ZN(n789) );
  NOR2_X1 U560 ( .A1(G651), .A2(G543), .ZN(n639) );
  NOR2_X1 U561 ( .A1(n531), .A2(n530), .ZN(G164) );
  INV_X1 U562 ( .A(G2104), .ZN(n526) );
  NOR2_X4 U563 ( .A1(G2105), .A2(n526), .ZN(n898) );
  NAND2_X1 U564 ( .A1(G102), .A2(n898), .ZN(n522) );
  AND2_X1 U565 ( .A1(G2104), .A2(G2105), .ZN(n893) );
  NAND2_X1 U566 ( .A1(G114), .A2(n893), .ZN(n521) );
  NAND2_X1 U567 ( .A1(n522), .A2(n521), .ZN(n531) );
  XNOR2_X1 U568 ( .A(KEYINPUT67), .B(KEYINPUT17), .ZN(n524) );
  NOR2_X1 U569 ( .A1(G2104), .A2(G2105), .ZN(n523) );
  XNOR2_X2 U570 ( .A(n524), .B(n523), .ZN(n896) );
  NAND2_X1 U571 ( .A1(G138), .A2(n896), .ZN(n525) );
  XNOR2_X1 U572 ( .A(n525), .B(KEYINPUT84), .ZN(n529) );
  AND2_X1 U573 ( .A1(n526), .A2(G2105), .ZN(n892) );
  NAND2_X1 U574 ( .A1(G126), .A2(n892), .ZN(n527) );
  XOR2_X1 U575 ( .A(KEYINPUT83), .B(n527), .Z(n528) );
  NAND2_X1 U576 ( .A1(n529), .A2(n528), .ZN(n530) );
  NAND2_X1 U577 ( .A1(n893), .A2(G113), .ZN(n532) );
  XNOR2_X1 U578 ( .A(n532), .B(KEYINPUT66), .ZN(n534) );
  NAND2_X1 U579 ( .A1(G137), .A2(n896), .ZN(n533) );
  NAND2_X1 U580 ( .A1(n534), .A2(n533), .ZN(n542) );
  INV_X1 U581 ( .A(KEYINPUT65), .ZN(n540) );
  INV_X1 U582 ( .A(KEYINPUT23), .ZN(n536) );
  NAND2_X1 U583 ( .A1(n898), .A2(G101), .ZN(n535) );
  XNOR2_X1 U584 ( .A(n536), .B(n535), .ZN(n538) );
  NAND2_X1 U585 ( .A1(n892), .A2(G125), .ZN(n537) );
  NAND2_X1 U586 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U587 ( .A(n540), .B(n539), .ZN(n541) );
  NAND2_X1 U588 ( .A1(G85), .A2(n639), .ZN(n546) );
  INV_X1 U589 ( .A(G651), .ZN(n547) );
  NOR2_X1 U590 ( .A1(G543), .A2(n547), .ZN(n543) );
  XOR2_X1 U591 ( .A(KEYINPUT1), .B(n543), .Z(n544) );
  XNOR2_X1 U592 ( .A(KEYINPUT68), .B(n544), .ZN(n652) );
  NAND2_X1 U593 ( .A1(G60), .A2(n652), .ZN(n545) );
  NAND2_X1 U594 ( .A1(n546), .A2(n545), .ZN(n552) );
  XOR2_X1 U595 ( .A(KEYINPUT0), .B(G543), .Z(n646) );
  NOR2_X1 U596 ( .A1(n646), .A2(n547), .ZN(n636) );
  NAND2_X1 U597 ( .A1(G72), .A2(n636), .ZN(n550) );
  NOR2_X1 U598 ( .A1(G651), .A2(n646), .ZN(n548) );
  XNOR2_X1 U599 ( .A(KEYINPUT64), .B(n548), .ZN(n648) );
  NAND2_X1 U600 ( .A1(G47), .A2(n648), .ZN(n549) );
  NAND2_X1 U601 ( .A1(n550), .A2(n549), .ZN(n551) );
  OR2_X1 U602 ( .A1(n552), .A2(n551), .ZN(G290) );
  AND2_X1 U603 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U604 ( .A(G57), .ZN(G237) );
  INV_X1 U605 ( .A(G132), .ZN(G219) );
  INV_X1 U606 ( .A(G82), .ZN(G220) );
  NAND2_X1 U607 ( .A1(G88), .A2(n639), .ZN(n554) );
  NAND2_X1 U608 ( .A1(G75), .A2(n636), .ZN(n553) );
  NAND2_X1 U609 ( .A1(n554), .A2(n553), .ZN(n558) );
  NAND2_X1 U610 ( .A1(G62), .A2(n652), .ZN(n556) );
  NAND2_X1 U611 ( .A1(G50), .A2(n648), .ZN(n555) );
  NAND2_X1 U612 ( .A1(n556), .A2(n555), .ZN(n557) );
  NOR2_X1 U613 ( .A1(n558), .A2(n557), .ZN(G166) );
  NAND2_X1 U614 ( .A1(G63), .A2(n652), .ZN(n560) );
  NAND2_X1 U615 ( .A1(G51), .A2(n648), .ZN(n559) );
  NAND2_X1 U616 ( .A1(n560), .A2(n559), .ZN(n562) );
  XOR2_X1 U617 ( .A(KEYINPUT73), .B(KEYINPUT6), .Z(n561) );
  XNOR2_X1 U618 ( .A(n562), .B(n561), .ZN(n569) );
  NAND2_X1 U619 ( .A1(n639), .A2(G89), .ZN(n563) );
  XOR2_X1 U620 ( .A(KEYINPUT4), .B(n563), .Z(n566) );
  NAND2_X1 U621 ( .A1(n636), .A2(G76), .ZN(n564) );
  XOR2_X1 U622 ( .A(KEYINPUT72), .B(n564), .Z(n565) );
  NOR2_X1 U623 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U624 ( .A(n567), .B(KEYINPUT5), .ZN(n568) );
  NOR2_X1 U625 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U626 ( .A(KEYINPUT7), .B(n570), .Z(G168) );
  XOR2_X1 U627 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U628 ( .A1(G7), .A2(G661), .ZN(n571) );
  XNOR2_X1 U629 ( .A(n571), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U630 ( .A(KEYINPUT11), .B(KEYINPUT70), .Z(n573) );
  INV_X1 U631 ( .A(G223), .ZN(n824) );
  NAND2_X1 U632 ( .A1(G567), .A2(n824), .ZN(n572) );
  XNOR2_X1 U633 ( .A(n573), .B(n572), .ZN(G234) );
  NAND2_X1 U634 ( .A1(n652), .A2(G56), .ZN(n574) );
  XOR2_X1 U635 ( .A(KEYINPUT14), .B(n574), .Z(n580) );
  NAND2_X1 U636 ( .A1(n639), .A2(G81), .ZN(n575) );
  XNOR2_X1 U637 ( .A(n575), .B(KEYINPUT12), .ZN(n577) );
  NAND2_X1 U638 ( .A1(G68), .A2(n636), .ZN(n576) );
  NAND2_X1 U639 ( .A1(n577), .A2(n576), .ZN(n578) );
  XOR2_X1 U640 ( .A(KEYINPUT13), .B(n578), .Z(n579) );
  NOR2_X1 U641 ( .A1(n580), .A2(n579), .ZN(n582) );
  NAND2_X1 U642 ( .A1(G43), .A2(n648), .ZN(n581) );
  NAND2_X1 U643 ( .A1(n582), .A2(n581), .ZN(n923) );
  INV_X1 U644 ( .A(G860), .ZN(n627) );
  OR2_X1 U645 ( .A1(n923), .A2(n627), .ZN(G153) );
  NAND2_X1 U646 ( .A1(n636), .A2(G77), .ZN(n583) );
  XOR2_X1 U647 ( .A(KEYINPUT69), .B(n583), .Z(n585) );
  NAND2_X1 U648 ( .A1(n639), .A2(G90), .ZN(n584) );
  NAND2_X1 U649 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U650 ( .A(KEYINPUT9), .B(n586), .ZN(n590) );
  NAND2_X1 U651 ( .A1(n652), .A2(G64), .ZN(n588) );
  NAND2_X1 U652 ( .A1(n648), .A2(G52), .ZN(n587) );
  AND2_X1 U653 ( .A1(n588), .A2(n587), .ZN(n589) );
  NAND2_X1 U654 ( .A1(n590), .A2(n589), .ZN(G301) );
  NAND2_X1 U655 ( .A1(G868), .A2(G301), .ZN(n600) );
  NAND2_X1 U656 ( .A1(G54), .A2(n648), .ZN(n597) );
  NAND2_X1 U657 ( .A1(G79), .A2(n636), .ZN(n592) );
  NAND2_X1 U658 ( .A1(G66), .A2(n652), .ZN(n591) );
  NAND2_X1 U659 ( .A1(n592), .A2(n591), .ZN(n595) );
  NAND2_X1 U660 ( .A1(G92), .A2(n639), .ZN(n593) );
  XNOR2_X1 U661 ( .A(KEYINPUT71), .B(n593), .ZN(n594) );
  NOR2_X1 U662 ( .A1(n595), .A2(n594), .ZN(n596) );
  NAND2_X1 U663 ( .A1(n597), .A2(n596), .ZN(n598) );
  XOR2_X1 U664 ( .A(KEYINPUT15), .B(n598), .Z(n933) );
  INV_X1 U665 ( .A(G868), .ZN(n666) );
  NAND2_X1 U666 ( .A1(n933), .A2(n666), .ZN(n599) );
  NAND2_X1 U667 ( .A1(n600), .A2(n599), .ZN(G284) );
  NAND2_X1 U668 ( .A1(G65), .A2(n652), .ZN(n602) );
  NAND2_X1 U669 ( .A1(G53), .A2(n648), .ZN(n601) );
  NAND2_X1 U670 ( .A1(n602), .A2(n601), .ZN(n606) );
  NAND2_X1 U671 ( .A1(G91), .A2(n639), .ZN(n604) );
  NAND2_X1 U672 ( .A1(G78), .A2(n636), .ZN(n603) );
  NAND2_X1 U673 ( .A1(n604), .A2(n603), .ZN(n605) );
  NOR2_X1 U674 ( .A1(n606), .A2(n605), .ZN(n922) );
  INV_X1 U675 ( .A(n922), .ZN(G299) );
  NOR2_X1 U676 ( .A1(G286), .A2(n666), .ZN(n608) );
  NOR2_X1 U677 ( .A1(G868), .A2(G299), .ZN(n607) );
  NOR2_X1 U678 ( .A1(n608), .A2(n607), .ZN(G297) );
  NAND2_X1 U679 ( .A1(n627), .A2(G559), .ZN(n609) );
  INV_X1 U680 ( .A(n933), .ZN(n625) );
  NAND2_X1 U681 ( .A1(n609), .A2(n625), .ZN(n610) );
  XNOR2_X1 U682 ( .A(n610), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U683 ( .A1(n625), .A2(G868), .ZN(n611) );
  NOR2_X1 U684 ( .A1(G559), .A2(n611), .ZN(n612) );
  XOR2_X1 U685 ( .A(KEYINPUT75), .B(n612), .Z(n615) );
  NOR2_X1 U686 ( .A1(G868), .A2(n923), .ZN(n613) );
  XNOR2_X1 U687 ( .A(KEYINPUT74), .B(n613), .ZN(n614) );
  NOR2_X1 U688 ( .A1(n615), .A2(n614), .ZN(G282) );
  NAND2_X1 U689 ( .A1(n892), .A2(G123), .ZN(n616) );
  XNOR2_X1 U690 ( .A(n616), .B(KEYINPUT18), .ZN(n618) );
  NAND2_X1 U691 ( .A1(G111), .A2(n893), .ZN(n617) );
  NAND2_X1 U692 ( .A1(n618), .A2(n617), .ZN(n622) );
  NAND2_X1 U693 ( .A1(G99), .A2(n898), .ZN(n620) );
  NAND2_X1 U694 ( .A1(G135), .A2(n896), .ZN(n619) );
  NAND2_X1 U695 ( .A1(n620), .A2(n619), .ZN(n621) );
  NOR2_X1 U696 ( .A1(n622), .A2(n621), .ZN(n975) );
  XOR2_X1 U697 ( .A(G2096), .B(n975), .Z(n623) );
  NOR2_X1 U698 ( .A1(G2100), .A2(n623), .ZN(n624) );
  XOR2_X1 U699 ( .A(KEYINPUT76), .B(n624), .Z(G156) );
  NAND2_X1 U700 ( .A1(G559), .A2(n625), .ZN(n626) );
  XOR2_X1 U701 ( .A(n923), .B(n626), .Z(n663) );
  NAND2_X1 U702 ( .A1(n627), .A2(n663), .ZN(n635) );
  NAND2_X1 U703 ( .A1(G93), .A2(n639), .ZN(n629) );
  NAND2_X1 U704 ( .A1(G80), .A2(n636), .ZN(n628) );
  NAND2_X1 U705 ( .A1(n629), .A2(n628), .ZN(n634) );
  NAND2_X1 U706 ( .A1(G67), .A2(n652), .ZN(n631) );
  NAND2_X1 U707 ( .A1(G55), .A2(n648), .ZN(n630) );
  NAND2_X1 U708 ( .A1(n631), .A2(n630), .ZN(n632) );
  XOR2_X1 U709 ( .A(KEYINPUT77), .B(n632), .Z(n633) );
  NOR2_X1 U710 ( .A1(n634), .A2(n633), .ZN(n665) );
  XOR2_X1 U711 ( .A(n635), .B(n665), .Z(G145) );
  XOR2_X1 U712 ( .A(KEYINPUT2), .B(KEYINPUT80), .Z(n638) );
  NAND2_X1 U713 ( .A1(G73), .A2(n636), .ZN(n637) );
  XNOR2_X1 U714 ( .A(n638), .B(n637), .ZN(n643) );
  NAND2_X1 U715 ( .A1(G86), .A2(n639), .ZN(n641) );
  NAND2_X1 U716 ( .A1(G61), .A2(n652), .ZN(n640) );
  NAND2_X1 U717 ( .A1(n641), .A2(n640), .ZN(n642) );
  NOR2_X1 U718 ( .A1(n643), .A2(n642), .ZN(n645) );
  NAND2_X1 U719 ( .A1(G48), .A2(n648), .ZN(n644) );
  NAND2_X1 U720 ( .A1(n645), .A2(n644), .ZN(G305) );
  NAND2_X1 U721 ( .A1(G87), .A2(n646), .ZN(n647) );
  XNOR2_X1 U722 ( .A(n647), .B(KEYINPUT78), .ZN(n654) );
  NAND2_X1 U723 ( .A1(G651), .A2(G74), .ZN(n650) );
  NAND2_X1 U724 ( .A1(G49), .A2(n648), .ZN(n649) );
  NAND2_X1 U725 ( .A1(n650), .A2(n649), .ZN(n651) );
  NOR2_X1 U726 ( .A1(n652), .A2(n651), .ZN(n653) );
  NAND2_X1 U727 ( .A1(n654), .A2(n653), .ZN(n655) );
  XOR2_X1 U728 ( .A(KEYINPUT79), .B(n655), .Z(G288) );
  XNOR2_X1 U729 ( .A(n665), .B(G305), .ZN(n656) );
  XNOR2_X1 U730 ( .A(n656), .B(G288), .ZN(n660) );
  XNOR2_X1 U731 ( .A(KEYINPUT81), .B(KEYINPUT19), .ZN(n658) );
  XNOR2_X1 U732 ( .A(G290), .B(KEYINPUT82), .ZN(n657) );
  XNOR2_X1 U733 ( .A(n658), .B(n657), .ZN(n659) );
  XOR2_X1 U734 ( .A(n660), .B(n659), .Z(n662) );
  XNOR2_X1 U735 ( .A(n922), .B(G166), .ZN(n661) );
  XNOR2_X1 U736 ( .A(n662), .B(n661), .ZN(n909) );
  XOR2_X1 U737 ( .A(n909), .B(n663), .Z(n664) );
  NOR2_X1 U738 ( .A1(n666), .A2(n664), .ZN(n668) );
  AND2_X1 U739 ( .A1(n666), .A2(n665), .ZN(n667) );
  NOR2_X1 U740 ( .A1(n668), .A2(n667), .ZN(G295) );
  NAND2_X1 U741 ( .A1(G2084), .A2(G2078), .ZN(n669) );
  XOR2_X1 U742 ( .A(KEYINPUT20), .B(n669), .Z(n670) );
  NAND2_X1 U743 ( .A1(G2090), .A2(n670), .ZN(n671) );
  XNOR2_X1 U744 ( .A(KEYINPUT21), .B(n671), .ZN(n672) );
  NAND2_X1 U745 ( .A1(n672), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U746 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U747 ( .A1(G220), .A2(G219), .ZN(n673) );
  XOR2_X1 U748 ( .A(KEYINPUT22), .B(n673), .Z(n674) );
  NOR2_X1 U749 ( .A1(G218), .A2(n674), .ZN(n675) );
  NAND2_X1 U750 ( .A1(G96), .A2(n675), .ZN(n829) );
  NAND2_X1 U751 ( .A1(n829), .A2(G2106), .ZN(n679) );
  NAND2_X1 U752 ( .A1(G69), .A2(G120), .ZN(n676) );
  NOR2_X1 U753 ( .A1(G237), .A2(n676), .ZN(n677) );
  NAND2_X1 U754 ( .A1(G108), .A2(n677), .ZN(n830) );
  NAND2_X1 U755 ( .A1(n830), .A2(G567), .ZN(n678) );
  NAND2_X1 U756 ( .A1(n679), .A2(n678), .ZN(n920) );
  NAND2_X1 U757 ( .A1(G483), .A2(G661), .ZN(n680) );
  NOR2_X1 U758 ( .A1(n920), .A2(n680), .ZN(n828) );
  NAND2_X1 U759 ( .A1(n828), .A2(G36), .ZN(G176) );
  INV_X1 U760 ( .A(G166), .ZN(G303) );
  NAND2_X1 U761 ( .A1(n892), .A2(G119), .ZN(n687) );
  NAND2_X1 U762 ( .A1(G107), .A2(n893), .ZN(n682) );
  NAND2_X1 U763 ( .A1(G131), .A2(n896), .ZN(n681) );
  NAND2_X1 U764 ( .A1(n682), .A2(n681), .ZN(n685) );
  NAND2_X1 U765 ( .A1(n898), .A2(G95), .ZN(n683) );
  XOR2_X1 U766 ( .A(KEYINPUT88), .B(n683), .Z(n684) );
  NOR2_X1 U767 ( .A1(n685), .A2(n684), .ZN(n686) );
  NAND2_X1 U768 ( .A1(n687), .A2(n686), .ZN(n688) );
  XOR2_X1 U769 ( .A(KEYINPUT89), .B(n688), .Z(n874) );
  NAND2_X1 U770 ( .A1(G1991), .A2(n874), .ZN(n689) );
  XOR2_X1 U771 ( .A(KEYINPUT90), .B(n689), .Z(n700) );
  NAND2_X1 U772 ( .A1(n892), .A2(G129), .ZN(n696) );
  NAND2_X1 U773 ( .A1(G117), .A2(n893), .ZN(n691) );
  NAND2_X1 U774 ( .A1(G141), .A2(n896), .ZN(n690) );
  NAND2_X1 U775 ( .A1(n691), .A2(n690), .ZN(n694) );
  NAND2_X1 U776 ( .A1(n898), .A2(G105), .ZN(n692) );
  XOR2_X1 U777 ( .A(KEYINPUT38), .B(n692), .Z(n693) );
  NOR2_X1 U778 ( .A1(n694), .A2(n693), .ZN(n695) );
  NAND2_X1 U779 ( .A1(n696), .A2(n695), .ZN(n697) );
  XOR2_X1 U780 ( .A(KEYINPUT91), .B(n697), .Z(n873) );
  INV_X1 U781 ( .A(n873), .ZN(n698) );
  INV_X1 U782 ( .A(G1996), .ZN(n724) );
  NOR2_X1 U783 ( .A1(n698), .A2(n724), .ZN(n699) );
  NOR2_X1 U784 ( .A1(n700), .A2(n699), .ZN(n986) );
  NOR2_X1 U785 ( .A1(G164), .A2(G1384), .ZN(n706) );
  NAND2_X1 U786 ( .A1(G160), .A2(G40), .ZN(n705) );
  NOR2_X1 U787 ( .A1(n706), .A2(n705), .ZN(n819) );
  INV_X1 U788 ( .A(n819), .ZN(n701) );
  NOR2_X1 U789 ( .A1(n986), .A2(n701), .ZN(n810) );
  INV_X1 U790 ( .A(n810), .ZN(n704) );
  XNOR2_X1 U791 ( .A(G1986), .B(G290), .ZN(n925) );
  NAND2_X1 U792 ( .A1(n925), .A2(n819), .ZN(n702) );
  XOR2_X1 U793 ( .A(KEYINPUT85), .B(n702), .Z(n703) );
  NAND2_X1 U794 ( .A1(n704), .A2(n703), .ZN(n795) );
  XOR2_X1 U795 ( .A(G1981), .B(G305), .Z(n938) );
  INV_X1 U796 ( .A(n705), .ZN(n707) );
  NAND2_X1 U797 ( .A1(n707), .A2(n706), .ZN(n751) );
  NAND2_X1 U798 ( .A1(G1961), .A2(n751), .ZN(n709) );
  INV_X1 U799 ( .A(n751), .ZN(n729) );
  XOR2_X1 U800 ( .A(KEYINPUT25), .B(G2078), .Z(n950) );
  NAND2_X1 U801 ( .A1(n729), .A2(n950), .ZN(n708) );
  NAND2_X1 U802 ( .A1(n709), .A2(n708), .ZN(n743) );
  NAND2_X1 U803 ( .A1(G301), .A2(n743), .ZN(n710) );
  XNOR2_X1 U804 ( .A(n710), .B(KEYINPUT93), .ZN(n715) );
  NOR2_X1 U805 ( .A1(G2084), .A2(n751), .ZN(n766) );
  NOR2_X1 U806 ( .A1(G1966), .A2(n789), .ZN(n762) );
  NOR2_X1 U807 ( .A1(n766), .A2(n762), .ZN(n711) );
  NAND2_X1 U808 ( .A1(n711), .A2(G8), .ZN(n712) );
  XNOR2_X1 U809 ( .A(KEYINPUT30), .B(n712), .ZN(n713) );
  NOR2_X1 U810 ( .A1(n713), .A2(G168), .ZN(n714) );
  NOR2_X1 U811 ( .A1(n715), .A2(n714), .ZN(n718) );
  XOR2_X1 U812 ( .A(KEYINPUT94), .B(KEYINPUT95), .Z(n716) );
  NAND2_X1 U813 ( .A1(n729), .A2(G2072), .ZN(n719) );
  XNOR2_X1 U814 ( .A(n719), .B(KEYINPUT27), .ZN(n721) );
  XOR2_X1 U815 ( .A(KEYINPUT92), .B(G1956), .Z(n1002) );
  NOR2_X1 U816 ( .A1(n729), .A2(n1002), .ZN(n720) );
  NOR2_X1 U817 ( .A1(n721), .A2(n720), .ZN(n737) );
  NOR2_X1 U818 ( .A1(n922), .A2(n737), .ZN(n723) );
  INV_X1 U819 ( .A(KEYINPUT28), .ZN(n722) );
  XNOR2_X1 U820 ( .A(n723), .B(n722), .ZN(n741) );
  NOR2_X1 U821 ( .A1(n751), .A2(n724), .ZN(n725) );
  XOR2_X1 U822 ( .A(n725), .B(KEYINPUT26), .Z(n727) );
  NAND2_X1 U823 ( .A1(n751), .A2(G1341), .ZN(n726) );
  NAND2_X1 U824 ( .A1(n727), .A2(n726), .ZN(n728) );
  NOR2_X1 U825 ( .A1(n923), .A2(n728), .ZN(n733) );
  NAND2_X1 U826 ( .A1(G1348), .A2(n751), .ZN(n731) );
  NAND2_X1 U827 ( .A1(n729), .A2(G2067), .ZN(n730) );
  NAND2_X1 U828 ( .A1(n731), .A2(n730), .ZN(n734) );
  NOR2_X1 U829 ( .A1(n933), .A2(n734), .ZN(n732) );
  NAND2_X1 U830 ( .A1(n933), .A2(n734), .ZN(n735) );
  NAND2_X1 U831 ( .A1(n736), .A2(n735), .ZN(n739) );
  NAND2_X1 U832 ( .A1(n922), .A2(n737), .ZN(n738) );
  NAND2_X1 U833 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U834 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U835 ( .A(n742), .B(KEYINPUT29), .ZN(n745) );
  NOR2_X1 U836 ( .A1(G301), .A2(n743), .ZN(n744) );
  NOR2_X1 U837 ( .A1(n745), .A2(n744), .ZN(n746) );
  NOR2_X1 U838 ( .A1(n747), .A2(n746), .ZN(n748) );
  XNOR2_X1 U839 ( .A(n748), .B(KEYINPUT96), .ZN(n763) );
  INV_X1 U840 ( .A(n763), .ZN(n750) );
  AND2_X1 U841 ( .A1(G286), .A2(G8), .ZN(n749) );
  NAND2_X1 U842 ( .A1(n750), .A2(n749), .ZN(n760) );
  INV_X1 U843 ( .A(G8), .ZN(n758) );
  NOR2_X1 U844 ( .A1(G1971), .A2(n789), .ZN(n753) );
  NOR2_X1 U845 ( .A1(G2090), .A2(n751), .ZN(n752) );
  NOR2_X1 U846 ( .A1(n753), .A2(n752), .ZN(n754) );
  XOR2_X1 U847 ( .A(KEYINPUT98), .B(n754), .Z(n755) );
  NOR2_X1 U848 ( .A1(G166), .A2(n755), .ZN(n756) );
  XNOR2_X1 U849 ( .A(n756), .B(KEYINPUT99), .ZN(n757) );
  OR2_X1 U850 ( .A1(n758), .A2(n757), .ZN(n759) );
  AND2_X1 U851 ( .A1(n760), .A2(n759), .ZN(n761) );
  XNOR2_X1 U852 ( .A(KEYINPUT32), .B(n761), .ZN(n770) );
  NOR2_X1 U853 ( .A1(n763), .A2(n762), .ZN(n765) );
  XNOR2_X1 U854 ( .A(n765), .B(n764), .ZN(n768) );
  NAND2_X1 U855 ( .A1(G8), .A2(n766), .ZN(n767) );
  NAND2_X1 U856 ( .A1(n768), .A2(n767), .ZN(n769) );
  NAND2_X1 U857 ( .A1(n770), .A2(n769), .ZN(n784) );
  NOR2_X1 U858 ( .A1(G1976), .A2(G288), .ZN(n937) );
  NOR2_X1 U859 ( .A1(G1971), .A2(G303), .ZN(n771) );
  NOR2_X1 U860 ( .A1(n937), .A2(n771), .ZN(n772) );
  XNOR2_X1 U861 ( .A(n772), .B(KEYINPUT100), .ZN(n773) );
  NAND2_X1 U862 ( .A1(n784), .A2(n773), .ZN(n776) );
  NAND2_X1 U863 ( .A1(G1976), .A2(G288), .ZN(n935) );
  INV_X1 U864 ( .A(n935), .ZN(n774) );
  NOR2_X1 U865 ( .A1(n789), .A2(n774), .ZN(n775) );
  AND2_X1 U866 ( .A1(n776), .A2(n775), .ZN(n777) );
  NOR2_X1 U867 ( .A1(KEYINPUT33), .A2(n777), .ZN(n780) );
  NAND2_X1 U868 ( .A1(n937), .A2(KEYINPUT33), .ZN(n778) );
  NOR2_X1 U869 ( .A1(n789), .A2(n778), .ZN(n779) );
  NOR2_X1 U870 ( .A1(n780), .A2(n779), .ZN(n781) );
  NAND2_X1 U871 ( .A1(n938), .A2(n781), .ZN(n793) );
  NOR2_X1 U872 ( .A1(G2090), .A2(G303), .ZN(n782) );
  XOR2_X1 U873 ( .A(KEYINPUT101), .B(n782), .Z(n783) );
  NAND2_X1 U874 ( .A1(G8), .A2(n783), .ZN(n785) );
  NAND2_X1 U875 ( .A1(n785), .A2(n784), .ZN(n786) );
  AND2_X1 U876 ( .A1(n786), .A2(n789), .ZN(n791) );
  NOR2_X1 U877 ( .A1(G1981), .A2(G305), .ZN(n787) );
  XOR2_X1 U878 ( .A(n787), .B(KEYINPUT24), .Z(n788) );
  NOR2_X1 U879 ( .A1(n789), .A2(n788), .ZN(n790) );
  NOR2_X1 U880 ( .A1(n791), .A2(n790), .ZN(n792) );
  AND2_X1 U881 ( .A1(n793), .A2(n792), .ZN(n794) );
  NOR2_X1 U882 ( .A1(n795), .A2(n794), .ZN(n807) );
  XNOR2_X1 U883 ( .A(KEYINPUT86), .B(KEYINPUT87), .ZN(n800) );
  NAND2_X1 U884 ( .A1(G128), .A2(n892), .ZN(n797) );
  NAND2_X1 U885 ( .A1(G116), .A2(n893), .ZN(n796) );
  NAND2_X1 U886 ( .A1(n797), .A2(n796), .ZN(n798) );
  XNOR2_X1 U887 ( .A(n798), .B(KEYINPUT35), .ZN(n799) );
  XNOR2_X1 U888 ( .A(n800), .B(n799), .ZN(n805) );
  NAND2_X1 U889 ( .A1(G104), .A2(n898), .ZN(n802) );
  NAND2_X1 U890 ( .A1(G140), .A2(n896), .ZN(n801) );
  NAND2_X1 U891 ( .A1(n802), .A2(n801), .ZN(n803) );
  XNOR2_X1 U892 ( .A(KEYINPUT34), .B(n803), .ZN(n804) );
  NOR2_X1 U893 ( .A1(n805), .A2(n804), .ZN(n806) );
  XNOR2_X1 U894 ( .A(KEYINPUT36), .B(n806), .ZN(n906) );
  XNOR2_X1 U895 ( .A(G2067), .B(KEYINPUT37), .ZN(n816) );
  NOR2_X1 U896 ( .A1(n906), .A2(n816), .ZN(n992) );
  NAND2_X1 U897 ( .A1(n992), .A2(n819), .ZN(n814) );
  NAND2_X1 U898 ( .A1(n807), .A2(n814), .ZN(n821) );
  NOR2_X1 U899 ( .A1(G1996), .A2(n873), .ZN(n971) );
  NOR2_X1 U900 ( .A1(G1986), .A2(G290), .ZN(n808) );
  NOR2_X1 U901 ( .A1(G1991), .A2(n874), .ZN(n977) );
  NOR2_X1 U902 ( .A1(n808), .A2(n977), .ZN(n809) );
  NOR2_X1 U903 ( .A1(n810), .A2(n809), .ZN(n811) );
  XNOR2_X1 U904 ( .A(n811), .B(KEYINPUT102), .ZN(n812) );
  NOR2_X1 U905 ( .A1(n971), .A2(n812), .ZN(n813) );
  XNOR2_X1 U906 ( .A(KEYINPUT39), .B(n813), .ZN(n815) );
  NAND2_X1 U907 ( .A1(n815), .A2(n814), .ZN(n817) );
  NAND2_X1 U908 ( .A1(n906), .A2(n816), .ZN(n990) );
  NAND2_X1 U909 ( .A1(n817), .A2(n990), .ZN(n818) );
  NAND2_X1 U910 ( .A1(n819), .A2(n818), .ZN(n820) );
  NAND2_X1 U911 ( .A1(n821), .A2(n820), .ZN(n823) );
  XOR2_X1 U912 ( .A(KEYINPUT40), .B(KEYINPUT103), .Z(n822) );
  XNOR2_X1 U913 ( .A(n823), .B(n822), .ZN(G329) );
  NAND2_X1 U914 ( .A1(G2106), .A2(n824), .ZN(G217) );
  AND2_X1 U915 ( .A1(G15), .A2(G2), .ZN(n825) );
  NAND2_X1 U916 ( .A1(G661), .A2(n825), .ZN(G259) );
  NAND2_X1 U917 ( .A1(G3), .A2(G1), .ZN(n826) );
  XOR2_X1 U918 ( .A(KEYINPUT109), .B(n826), .Z(n827) );
  NAND2_X1 U919 ( .A1(n828), .A2(n827), .ZN(G188) );
  INV_X1 U921 ( .A(G120), .ZN(G236) );
  INV_X1 U922 ( .A(G96), .ZN(G221) );
  INV_X1 U923 ( .A(G69), .ZN(G235) );
  NOR2_X1 U924 ( .A1(n830), .A2(n829), .ZN(G325) );
  INV_X1 U925 ( .A(G325), .ZN(G261) );
  XOR2_X1 U926 ( .A(G2438), .B(G2430), .Z(n832) );
  XNOR2_X1 U927 ( .A(G1341), .B(G1348), .ZN(n831) );
  XNOR2_X1 U928 ( .A(n832), .B(n831), .ZN(n842) );
  XOR2_X1 U929 ( .A(KEYINPUT107), .B(KEYINPUT104), .Z(n834) );
  XNOR2_X1 U930 ( .A(G2446), .B(G2443), .ZN(n833) );
  XNOR2_X1 U931 ( .A(n834), .B(n833), .ZN(n838) );
  XOR2_X1 U932 ( .A(KEYINPUT106), .B(G2451), .Z(n836) );
  XNOR2_X1 U933 ( .A(G2454), .B(G2435), .ZN(n835) );
  XNOR2_X1 U934 ( .A(n836), .B(n835), .ZN(n837) );
  XOR2_X1 U935 ( .A(n838), .B(n837), .Z(n840) );
  XNOR2_X1 U936 ( .A(KEYINPUT105), .B(G2427), .ZN(n839) );
  XNOR2_X1 U937 ( .A(n840), .B(n839), .ZN(n841) );
  XNOR2_X1 U938 ( .A(n842), .B(n841), .ZN(n843) );
  NAND2_X1 U939 ( .A1(n843), .A2(G14), .ZN(n844) );
  XOR2_X1 U940 ( .A(KEYINPUT108), .B(n844), .Z(G401) );
  XOR2_X1 U941 ( .A(G2100), .B(G2096), .Z(n846) );
  XNOR2_X1 U942 ( .A(KEYINPUT42), .B(G2678), .ZN(n845) );
  XNOR2_X1 U943 ( .A(n846), .B(n845), .ZN(n850) );
  XOR2_X1 U944 ( .A(KEYINPUT43), .B(G2090), .Z(n848) );
  XNOR2_X1 U945 ( .A(G2067), .B(G2072), .ZN(n847) );
  XNOR2_X1 U946 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U947 ( .A(n850), .B(n849), .Z(n852) );
  XNOR2_X1 U948 ( .A(G2084), .B(G2078), .ZN(n851) );
  XNOR2_X1 U949 ( .A(n852), .B(n851), .ZN(G227) );
  XOR2_X1 U950 ( .A(KEYINPUT41), .B(G1991), .Z(n854) );
  XNOR2_X1 U951 ( .A(G1996), .B(G1956), .ZN(n853) );
  XNOR2_X1 U952 ( .A(n854), .B(n853), .ZN(n855) );
  XOR2_X1 U953 ( .A(n855), .B(KEYINPUT111), .Z(n857) );
  XNOR2_X1 U954 ( .A(G1971), .B(G1986), .ZN(n856) );
  XNOR2_X1 U955 ( .A(n857), .B(n856), .ZN(n861) );
  XOR2_X1 U956 ( .A(G1976), .B(G1981), .Z(n859) );
  XNOR2_X1 U957 ( .A(G1966), .B(G1961), .ZN(n858) );
  XNOR2_X1 U958 ( .A(n859), .B(n858), .ZN(n860) );
  XOR2_X1 U959 ( .A(n861), .B(n860), .Z(n863) );
  XNOR2_X1 U960 ( .A(G2474), .B(KEYINPUT110), .ZN(n862) );
  XNOR2_X1 U961 ( .A(n863), .B(n862), .ZN(G229) );
  NAND2_X1 U962 ( .A1(G112), .A2(n893), .ZN(n864) );
  XNOR2_X1 U963 ( .A(n864), .B(KEYINPUT112), .ZN(n867) );
  NAND2_X1 U964 ( .A1(G100), .A2(n898), .ZN(n865) );
  XOR2_X1 U965 ( .A(KEYINPUT113), .B(n865), .Z(n866) );
  NAND2_X1 U966 ( .A1(n867), .A2(n866), .ZN(n872) );
  NAND2_X1 U967 ( .A1(n892), .A2(G124), .ZN(n868) );
  XNOR2_X1 U968 ( .A(n868), .B(KEYINPUT44), .ZN(n870) );
  NAND2_X1 U969 ( .A1(G136), .A2(n896), .ZN(n869) );
  NAND2_X1 U970 ( .A1(n870), .A2(n869), .ZN(n871) );
  NOR2_X1 U971 ( .A1(n872), .A2(n871), .ZN(G162) );
  XNOR2_X1 U972 ( .A(G160), .B(n873), .ZN(n875) );
  XNOR2_X1 U973 ( .A(n875), .B(n874), .ZN(n879) );
  XOR2_X1 U974 ( .A(KEYINPUT48), .B(KEYINPUT117), .Z(n877) );
  XNOR2_X1 U975 ( .A(KEYINPUT46), .B(KEYINPUT115), .ZN(n876) );
  XNOR2_X1 U976 ( .A(n877), .B(n876), .ZN(n878) );
  XOR2_X1 U977 ( .A(n879), .B(n878), .Z(n891) );
  NAND2_X1 U978 ( .A1(G103), .A2(n898), .ZN(n881) );
  NAND2_X1 U979 ( .A1(G139), .A2(n896), .ZN(n880) );
  NAND2_X1 U980 ( .A1(n881), .A2(n880), .ZN(n886) );
  NAND2_X1 U981 ( .A1(G127), .A2(n892), .ZN(n883) );
  NAND2_X1 U982 ( .A1(G115), .A2(n893), .ZN(n882) );
  NAND2_X1 U983 ( .A1(n883), .A2(n882), .ZN(n884) );
  XOR2_X1 U984 ( .A(KEYINPUT47), .B(n884), .Z(n885) );
  NOR2_X1 U985 ( .A1(n886), .A2(n885), .ZN(n887) );
  XNOR2_X1 U986 ( .A(KEYINPUT116), .B(n887), .ZN(n980) );
  XOR2_X1 U987 ( .A(G164), .B(G162), .Z(n888) );
  XNOR2_X1 U988 ( .A(n980), .B(n888), .ZN(n889) );
  XNOR2_X1 U989 ( .A(n975), .B(n889), .ZN(n890) );
  XNOR2_X1 U990 ( .A(n891), .B(n890), .ZN(n905) );
  NAND2_X1 U991 ( .A1(G130), .A2(n892), .ZN(n895) );
  NAND2_X1 U992 ( .A1(G118), .A2(n893), .ZN(n894) );
  NAND2_X1 U993 ( .A1(n895), .A2(n894), .ZN(n903) );
  NAND2_X1 U994 ( .A1(n896), .A2(G142), .ZN(n897) );
  XNOR2_X1 U995 ( .A(n897), .B(KEYINPUT114), .ZN(n900) );
  NAND2_X1 U996 ( .A1(G106), .A2(n898), .ZN(n899) );
  NAND2_X1 U997 ( .A1(n900), .A2(n899), .ZN(n901) );
  XOR2_X1 U998 ( .A(n901), .B(KEYINPUT45), .Z(n902) );
  NOR2_X1 U999 ( .A1(n903), .A2(n902), .ZN(n904) );
  XOR2_X1 U1000 ( .A(n905), .B(n904), .Z(n907) );
  XNOR2_X1 U1001 ( .A(n907), .B(n906), .ZN(n908) );
  NOR2_X1 U1002 ( .A1(G37), .A2(n908), .ZN(G395) );
  INV_X1 U1003 ( .A(G301), .ZN(G171) );
  XNOR2_X1 U1004 ( .A(n909), .B(KEYINPUT118), .ZN(n911) );
  XNOR2_X1 U1005 ( .A(n923), .B(G286), .ZN(n910) );
  XNOR2_X1 U1006 ( .A(n911), .B(n910), .ZN(n913) );
  XNOR2_X1 U1007 ( .A(n933), .B(G171), .ZN(n912) );
  XNOR2_X1 U1008 ( .A(n913), .B(n912), .ZN(n914) );
  NOR2_X1 U1009 ( .A1(G37), .A2(n914), .ZN(G397) );
  OR2_X1 U1010 ( .A1(n920), .A2(G401), .ZN(n917) );
  NOR2_X1 U1011 ( .A1(G227), .A2(G229), .ZN(n915) );
  XNOR2_X1 U1012 ( .A(KEYINPUT49), .B(n915), .ZN(n916) );
  NOR2_X1 U1013 ( .A1(n917), .A2(n916), .ZN(n919) );
  NOR2_X1 U1014 ( .A1(G395), .A2(G397), .ZN(n918) );
  NAND2_X1 U1015 ( .A1(n919), .A2(n918), .ZN(G225) );
  INV_X1 U1016 ( .A(G225), .ZN(G308) );
  INV_X1 U1017 ( .A(n920), .ZN(G319) );
  INV_X1 U1018 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1019 ( .A(G16), .B(KEYINPUT56), .Z(n921) );
  XNOR2_X1 U1020 ( .A(KEYINPUT124), .B(n921), .ZN(n946) );
  XNOR2_X1 U1021 ( .A(G171), .B(G1961), .ZN(n932) );
  XNOR2_X1 U1022 ( .A(n922), .B(G1956), .ZN(n927) );
  XNOR2_X1 U1023 ( .A(G1341), .B(n923), .ZN(n924) );
  NOR2_X1 U1024 ( .A1(n925), .A2(n924), .ZN(n926) );
  NAND2_X1 U1025 ( .A1(n927), .A2(n926), .ZN(n930) );
  XOR2_X1 U1026 ( .A(G1971), .B(G303), .Z(n928) );
  XNOR2_X1 U1027 ( .A(KEYINPUT125), .B(n928), .ZN(n929) );
  NOR2_X1 U1028 ( .A1(n930), .A2(n929), .ZN(n931) );
  NAND2_X1 U1029 ( .A1(n932), .A2(n931), .ZN(n944) );
  XOR2_X1 U1030 ( .A(G1348), .B(n933), .Z(n934) );
  NAND2_X1 U1031 ( .A1(n935), .A2(n934), .ZN(n936) );
  NOR2_X1 U1032 ( .A1(n937), .A2(n936), .ZN(n942) );
  XNOR2_X1 U1033 ( .A(G1966), .B(G168), .ZN(n939) );
  NAND2_X1 U1034 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1035 ( .A(n940), .B(KEYINPUT57), .ZN(n941) );
  NAND2_X1 U1036 ( .A1(n942), .A2(n941), .ZN(n943) );
  NOR2_X1 U1037 ( .A1(n944), .A2(n943), .ZN(n945) );
  NOR2_X1 U1038 ( .A1(n946), .A2(n945), .ZN(n968) );
  INV_X1 U1039 ( .A(KEYINPUT55), .ZN(n997) );
  XNOR2_X1 U1040 ( .A(G2090), .B(G35), .ZN(n959) );
  XOR2_X1 U1041 ( .A(G1991), .B(G25), .Z(n947) );
  NAND2_X1 U1042 ( .A1(n947), .A2(G28), .ZN(n956) );
  XNOR2_X1 U1043 ( .A(G2067), .B(G26), .ZN(n949) );
  XNOR2_X1 U1044 ( .A(G33), .B(G2072), .ZN(n948) );
  NOR2_X1 U1045 ( .A1(n949), .A2(n948), .ZN(n954) );
  XNOR2_X1 U1046 ( .A(n950), .B(G27), .ZN(n952) );
  XNOR2_X1 U1047 ( .A(G1996), .B(G32), .ZN(n951) );
  NOR2_X1 U1048 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1049 ( .A1(n954), .A2(n953), .ZN(n955) );
  NOR2_X1 U1050 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1051 ( .A(KEYINPUT53), .B(n957), .ZN(n958) );
  NOR2_X1 U1052 ( .A1(n959), .A2(n958), .ZN(n962) );
  XOR2_X1 U1053 ( .A(G2084), .B(G34), .Z(n960) );
  XNOR2_X1 U1054 ( .A(KEYINPUT54), .B(n960), .ZN(n961) );
  NAND2_X1 U1055 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1056 ( .A(n997), .B(n963), .ZN(n965) );
  INV_X1 U1057 ( .A(G29), .ZN(n964) );
  NAND2_X1 U1058 ( .A1(n965), .A2(n964), .ZN(n966) );
  NAND2_X1 U1059 ( .A1(G11), .A2(n966), .ZN(n967) );
  NOR2_X1 U1060 ( .A1(n968), .A2(n967), .ZN(n1001) );
  XOR2_X1 U1061 ( .A(KEYINPUT51), .B(KEYINPUT120), .Z(n973) );
  XNOR2_X1 U1062 ( .A(G2090), .B(G162), .ZN(n969) );
  XNOR2_X1 U1063 ( .A(n969), .B(KEYINPUT119), .ZN(n970) );
  NOR2_X1 U1064 ( .A1(n971), .A2(n970), .ZN(n972) );
  XOR2_X1 U1065 ( .A(n973), .B(n972), .Z(n974) );
  NOR2_X1 U1066 ( .A1(n975), .A2(n974), .ZN(n979) );
  XOR2_X1 U1067 ( .A(G2084), .B(G160), .Z(n976) );
  NOR2_X1 U1068 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1069 ( .A1(n979), .A2(n978), .ZN(n989) );
  XNOR2_X1 U1070 ( .A(G2072), .B(KEYINPUT121), .ZN(n981) );
  XNOR2_X1 U1071 ( .A(n981), .B(n980), .ZN(n983) );
  XOR2_X1 U1072 ( .A(G164), .B(G2078), .Z(n982) );
  NOR2_X1 U1073 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1074 ( .A(n984), .B(KEYINPUT50), .ZN(n985) );
  XNOR2_X1 U1075 ( .A(n985), .B(KEYINPUT122), .ZN(n987) );
  NAND2_X1 U1076 ( .A1(n987), .A2(n986), .ZN(n988) );
  NOR2_X1 U1077 ( .A1(n989), .A2(n988), .ZN(n994) );
  INV_X1 U1078 ( .A(n990), .ZN(n991) );
  NOR2_X1 U1079 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1080 ( .A1(n994), .A2(n993), .ZN(n995) );
  XNOR2_X1 U1081 ( .A(KEYINPUT52), .B(n995), .ZN(n996) );
  XNOR2_X1 U1082 ( .A(KEYINPUT123), .B(n996), .ZN(n998) );
  NAND2_X1 U1083 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1084 ( .A1(n999), .A2(G29), .ZN(n1000) );
  NAND2_X1 U1085 ( .A1(n1001), .A2(n1000), .ZN(n1027) );
  XNOR2_X1 U1086 ( .A(n1002), .B(G20), .ZN(n1006) );
  XNOR2_X1 U1087 ( .A(G1341), .B(G19), .ZN(n1004) );
  XNOR2_X1 U1088 ( .A(G1981), .B(G6), .ZN(n1003) );
  NOR2_X1 U1089 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1090 ( .A1(n1006), .A2(n1005), .ZN(n1009) );
  XOR2_X1 U1091 ( .A(KEYINPUT59), .B(G1348), .Z(n1007) );
  XNOR2_X1 U1092 ( .A(G4), .B(n1007), .ZN(n1008) );
  NOR2_X1 U1093 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1094 ( .A(KEYINPUT60), .B(n1010), .ZN(n1014) );
  XNOR2_X1 U1095 ( .A(G1966), .B(G21), .ZN(n1012) );
  XNOR2_X1 U1096 ( .A(G5), .B(G1961), .ZN(n1011) );
  NOR2_X1 U1097 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1098 ( .A1(n1014), .A2(n1013), .ZN(n1022) );
  XNOR2_X1 U1099 ( .A(G1976), .B(G23), .ZN(n1016) );
  XNOR2_X1 U1100 ( .A(G1986), .B(G24), .ZN(n1015) );
  NOR2_X1 U1101 ( .A1(n1016), .A2(n1015), .ZN(n1019) );
  XNOR2_X1 U1102 ( .A(G1971), .B(KEYINPUT127), .ZN(n1017) );
  XNOR2_X1 U1103 ( .A(n1017), .B(G22), .ZN(n1018) );
  NAND2_X1 U1104 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1105 ( .A(KEYINPUT58), .B(n1020), .ZN(n1021) );
  NOR2_X1 U1106 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XOR2_X1 U1107 ( .A(KEYINPUT61), .B(n1023), .Z(n1025) );
  XNOR2_X1 U1108 ( .A(KEYINPUT126), .B(G16), .ZN(n1024) );
  NOR2_X1 U1109 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NOR2_X1 U1110 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XNOR2_X1 U1111 ( .A(n1028), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1112 ( .A(G311), .ZN(G150) );
endmodule

