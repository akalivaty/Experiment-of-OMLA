//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 1 0 1 0 1 1 1 1 0 0 0 1 1 0 1 0 1 1 1 1 0 0 0 1 0 1 1 1 1 0 1 1 1 0 1 0 0 1 0 0 1 0 0 0 1 1 1 0 0 1 1 1 0 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:22 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n720, new_n721,
    new_n722, new_n724, new_n725, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n778, new_n779, new_n780, new_n781, new_n783, new_n784, new_n785,
    new_n786, new_n788, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n813, new_n814, new_n815, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n873, new_n874, new_n875, new_n877, new_n878,
    new_n879, new_n880, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n940, new_n941, new_n943, new_n944, new_n945,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n973, new_n974, new_n975, new_n976, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n986, new_n987,
    new_n988, new_n989, new_n991, new_n992, new_n993;
  NAND2_X1  g000(.A1(G232gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT41), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  XOR2_X1   g003(.A(new_n204), .B(KEYINPUT97), .Z(new_n205));
  XNOR2_X1  g004(.A(G134gat), .B(G162gat), .ZN(new_n206));
  XOR2_X1   g005(.A(new_n205), .B(new_n206), .Z(new_n207));
  NOR2_X1   g006(.A1(new_n207), .A2(KEYINPUT102), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT101), .ZN(new_n209));
  XNOR2_X1  g008(.A(G43gat), .B(G50gat), .ZN(new_n210));
  AND2_X1   g009(.A1(new_n210), .A2(KEYINPUT15), .ZN(new_n211));
  NOR2_X1   g010(.A1(G29gat), .A2(G36gat), .ZN(new_n212));
  XNOR2_X1  g011(.A(new_n212), .B(KEYINPUT14), .ZN(new_n213));
  NAND2_X1  g012(.A1(G29gat), .A2(G36gat), .ZN(new_n214));
  XNOR2_X1  g013(.A(new_n214), .B(KEYINPUT89), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n211), .B1(new_n213), .B2(new_n215), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n211), .A2(new_n215), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n217), .B1(KEYINPUT15), .B2(new_n210), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT90), .ZN(new_n219));
  XNOR2_X1  g018(.A(new_n213), .B(new_n219), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n216), .B1(new_n218), .B2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT91), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI211_X1 g022(.A(KEYINPUT91), .B(new_n216), .C1(new_n218), .C2(new_n220), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT92), .ZN(new_n226));
  OR3_X1    g025(.A1(new_n225), .A2(new_n226), .A3(KEYINPUT17), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n226), .B1(new_n225), .B2(KEYINPUT17), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(G85gat), .A2(G92gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(KEYINPUT98), .A2(KEYINPUT7), .ZN(new_n231));
  XOR2_X1   g030(.A(new_n230), .B(new_n231), .Z(new_n232));
  NAND2_X1  g031(.A1(G99gat), .A2(G106gat), .ZN(new_n233));
  INV_X1    g032(.A(G85gat), .ZN(new_n234));
  INV_X1    g033(.A(G92gat), .ZN(new_n235));
  AOI22_X1  g034(.A1(KEYINPUT8), .A2(new_n233), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n232), .A2(new_n236), .ZN(new_n237));
  XNOR2_X1  g036(.A(G99gat), .B(G106gat), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n237), .B(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(new_n221), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n239), .B1(new_n240), .B2(KEYINPUT17), .ZN(new_n241));
  INV_X1    g040(.A(new_n239), .ZN(new_n242));
  OAI22_X1  g041(.A1(new_n225), .A2(new_n242), .B1(new_n203), .B2(new_n202), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT99), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  OAI221_X1 g044(.A(KEYINPUT99), .B1(new_n203), .B2(new_n202), .C1(new_n225), .C2(new_n242), .ZN(new_n246));
  AOI22_X1  g045(.A1(new_n229), .A2(new_n241), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(G190gat), .B(G218gat), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n209), .B1(new_n247), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n229), .A2(new_n241), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n245), .A2(new_n246), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n253), .A2(KEYINPUT101), .A3(new_n248), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n208), .B1(new_n250), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n207), .A2(KEYINPUT102), .ZN(new_n256));
  OAI21_X1  g055(.A(KEYINPUT100), .B1(new_n253), .B2(new_n248), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT100), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n247), .A2(new_n258), .A3(new_n249), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n255), .A2(new_n256), .A3(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n256), .B1(new_n255), .B2(new_n260), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(G57gat), .B(G64gat), .ZN(new_n265));
  AOI21_X1  g064(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(G71gat), .B(G78gat), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n267), .B(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT21), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  XNOR2_X1  g070(.A(G127gat), .B(G155gat), .ZN(new_n272));
  XOR2_X1   g071(.A(new_n271), .B(new_n272), .Z(new_n273));
  XNOR2_X1  g072(.A(G15gat), .B(G22gat), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT16), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n274), .B1(new_n275), .B2(G1gat), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n276), .B1(G1gat), .B2(new_n274), .ZN(new_n277));
  INV_X1    g076(.A(G8gat), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n277), .B(new_n278), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n279), .B1(new_n269), .B2(new_n270), .ZN(new_n280));
  XOR2_X1   g079(.A(new_n273), .B(new_n280), .Z(new_n281));
  NAND2_X1  g080(.A1(G231gat), .A2(G233gat), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n282), .B(KEYINPUT96), .ZN(new_n283));
  XOR2_X1   g082(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n284));
  XNOR2_X1  g083(.A(new_n283), .B(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(G183gat), .B(G211gat), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n285), .B(new_n286), .ZN(new_n287));
  XOR2_X1   g086(.A(new_n281), .B(new_n287), .Z(new_n288));
  XNOR2_X1  g087(.A(new_n239), .B(new_n269), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT10), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  OR3_X1    g090(.A1(new_n242), .A2(new_n290), .A3(new_n269), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(G230gat), .A2(G233gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(KEYINPUT103), .ZN(new_n296));
  INV_X1    g095(.A(new_n289), .ZN(new_n297));
  INV_X1    g096(.A(new_n294), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(G120gat), .B(G148gat), .ZN(new_n300));
  XNOR2_X1  g099(.A(G176gat), .B(G204gat), .ZN(new_n301));
  XOR2_X1   g100(.A(new_n300), .B(new_n301), .Z(new_n302));
  AOI21_X1  g101(.A(new_n298), .B1(new_n291), .B2(new_n292), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT103), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND4_X1  g104(.A1(new_n296), .A2(new_n299), .A3(new_n302), .A4(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(new_n302), .ZN(new_n307));
  INV_X1    g106(.A(new_n299), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n307), .B1(new_n308), .B2(new_n303), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n306), .A2(new_n309), .ZN(new_n310));
  NOR3_X1   g109(.A1(new_n264), .A2(new_n288), .A3(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT17), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n279), .B1(new_n221), .B2(new_n312), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n313), .B1(new_n227), .B2(new_n228), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT18), .ZN(new_n315));
  NAND2_X1  g114(.A1(G229gat), .A2(G233gat), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n225), .A2(new_n279), .ZN(new_n318));
  NOR4_X1   g117(.A1(new_n314), .A2(new_n315), .A3(new_n317), .A4(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n318), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n225), .A2(new_n279), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n320), .A2(KEYINPUT94), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(KEYINPUT94), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(new_n318), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  XOR2_X1   g124(.A(new_n316), .B(KEYINPUT13), .Z(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n319), .A2(new_n328), .ZN(new_n329));
  OR2_X1    g128(.A1(new_n314), .A2(new_n318), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n315), .B1(new_n330), .B2(new_n317), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  NOR3_X1   g131(.A1(new_n314), .A2(new_n317), .A3(new_n318), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(KEYINPUT18), .ZN(new_n334));
  INV_X1    g133(.A(new_n328), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT93), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  XNOR2_X1  g136(.A(G113gat), .B(G141gat), .ZN(new_n338));
  INV_X1    g137(.A(G197gat), .ZN(new_n339));
  XNOR2_X1  g138(.A(new_n338), .B(new_n339), .ZN(new_n340));
  XNOR2_X1  g139(.A(KEYINPUT11), .B(G169gat), .ZN(new_n341));
  XNOR2_X1  g140(.A(new_n340), .B(new_n341), .ZN(new_n342));
  XNOR2_X1  g141(.A(KEYINPUT88), .B(KEYINPUT12), .ZN(new_n343));
  XOR2_X1   g142(.A(new_n342), .B(new_n343), .Z(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n332), .A2(new_n337), .A3(new_n345), .ZN(new_n346));
  OAI211_X1 g145(.A(new_n329), .B(new_n331), .C1(new_n336), .C2(new_n344), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT35), .ZN(new_n349));
  INV_X1    g148(.A(G227gat), .ZN(new_n350));
  INV_X1    g149(.A(G233gat), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT71), .ZN(new_n354));
  XNOR2_X1  g153(.A(KEYINPUT70), .B(KEYINPUT1), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  XNOR2_X1  g155(.A(G127gat), .B(G134gat), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(G113gat), .ZN(new_n359));
  OAI21_X1  g158(.A(KEYINPUT67), .B1(new_n359), .B2(G120gat), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT67), .ZN(new_n361));
  INV_X1    g160(.A(G120gat), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n361), .A2(new_n362), .A3(G113gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n360), .A2(new_n363), .ZN(new_n364));
  AND2_X1   g163(.A1(KEYINPUT68), .A2(G113gat), .ZN(new_n365));
  NOR2_X1   g164(.A1(KEYINPUT68), .A2(G113gat), .ZN(new_n366));
  NOR3_X1   g165(.A1(new_n365), .A2(new_n366), .A3(new_n362), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT69), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n364), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  OR2_X1    g168(.A1(KEYINPUT68), .A2(G113gat), .ZN(new_n370));
  NAND2_X1  g169(.A1(KEYINPUT68), .A2(G113gat), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n370), .A2(G120gat), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(KEYINPUT69), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n358), .B1(new_n369), .B2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT1), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n362), .A2(G113gat), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n359), .A2(G120gat), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n357), .B1(new_n375), .B2(new_n378), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n354), .B1(new_n374), .B2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n357), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n381), .A2(new_n355), .ZN(new_n382));
  NAND4_X1  g181(.A1(new_n370), .A2(new_n368), .A3(G120gat), .A4(new_n371), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n383), .A2(new_n360), .A3(new_n363), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n365), .A2(new_n366), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n368), .B1(new_n385), .B2(G120gat), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n382), .B1(new_n384), .B2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n379), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n387), .A2(KEYINPUT71), .A3(new_n388), .ZN(new_n389));
  NOR2_X1   g188(.A1(G169gat), .A2(G176gat), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT26), .ZN(new_n392));
  NAND2_X1  g191(.A1(G169gat), .A2(G176gat), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n391), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  AOI22_X1  g193(.A1(new_n390), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT66), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(G183gat), .ZN(new_n397));
  AOI21_X1  g196(.A(G190gat), .B1(new_n397), .B2(KEYINPUT27), .ZN(new_n398));
  INV_X1    g197(.A(G183gat), .ZN(new_n399));
  OR3_X1    g198(.A1(new_n399), .A2(KEYINPUT66), .A3(KEYINPUT27), .ZN(new_n400));
  AOI21_X1  g199(.A(KEYINPUT28), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  XNOR2_X1  g200(.A(KEYINPUT27), .B(G183gat), .ZN(new_n402));
  INV_X1    g201(.A(G190gat), .ZN(new_n403));
  AND3_X1   g202(.A1(new_n402), .A2(KEYINPUT28), .A3(new_n403), .ZN(new_n404));
  OAI211_X1 g203(.A(new_n394), .B(new_n395), .C1(new_n401), .C2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(G183gat), .A2(G190gat), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(KEYINPUT24), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT24), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n408), .A2(G183gat), .A3(G190gat), .ZN(new_n409));
  AOI22_X1  g208(.A1(new_n407), .A2(new_n409), .B1(new_n399), .B2(new_n403), .ZN(new_n410));
  INV_X1    g209(.A(G169gat), .ZN(new_n411));
  INV_X1    g210(.A(G176gat), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n411), .A2(new_n412), .A3(KEYINPUT23), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(new_n393), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT25), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n415), .B1(new_n390), .B2(KEYINPUT23), .ZN(new_n416));
  NOR3_X1   g215(.A1(new_n410), .A2(new_n414), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n407), .A2(new_n409), .ZN(new_n418));
  OAI21_X1  g217(.A(KEYINPUT65), .B1(G183gat), .B2(G190gat), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT65), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n420), .A2(new_n399), .A3(new_n403), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n418), .A2(new_n419), .A3(new_n421), .ZN(new_n422));
  OR2_X1    g221(.A1(new_n390), .A2(KEYINPUT23), .ZN(new_n423));
  AOI21_X1  g222(.A(KEYINPUT64), .B1(new_n413), .B2(new_n393), .ZN(new_n424));
  AND3_X1   g223(.A1(new_n413), .A2(KEYINPUT64), .A3(new_n393), .ZN(new_n425));
  OAI211_X1 g224(.A(new_n422), .B(new_n423), .C1(new_n424), .C2(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n417), .B1(new_n426), .B2(KEYINPUT25), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n380), .A2(new_n389), .A3(new_n405), .A4(new_n427), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n425), .A2(new_n424), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n399), .A2(KEYINPUT24), .ZN(new_n430));
  AOI22_X1  g229(.A1(new_n430), .A2(G190gat), .B1(KEYINPUT24), .B2(new_n406), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n421), .A2(new_n419), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n423), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  OAI21_X1  g232(.A(KEYINPUT25), .B1(new_n429), .B2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n417), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n434), .A2(new_n405), .A3(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(new_n364), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n373), .A2(new_n437), .A3(new_n383), .ZN(new_n438));
  AOI211_X1 g237(.A(new_n354), .B(new_n379), .C1(new_n438), .C2(new_n382), .ZN(new_n439));
  AOI21_X1  g238(.A(KEYINPUT71), .B1(new_n387), .B2(new_n388), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n436), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n353), .B1(new_n428), .B2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT32), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  XNOR2_X1  g243(.A(G15gat), .B(G43gat), .ZN(new_n445));
  XNOR2_X1  g244(.A(G71gat), .B(G99gat), .ZN(new_n446));
  XNOR2_X1  g245(.A(new_n445), .B(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(KEYINPUT33), .ZN(new_n449));
  AND2_X1   g248(.A1(new_n444), .A2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT72), .ZN(new_n452));
  NOR3_X1   g251(.A1(new_n436), .A2(new_n439), .A3(new_n440), .ZN(new_n453));
  AOI22_X1  g252(.A1(new_n380), .A2(new_n389), .B1(new_n427), .B2(new_n405), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n352), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n447), .B1(new_n455), .B2(KEYINPUT32), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT33), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n452), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n448), .B1(new_n442), .B2(new_n443), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n428), .A2(new_n441), .ZN(new_n461));
  AOI21_X1  g260(.A(KEYINPUT33), .B1(new_n461), .B2(new_n352), .ZN(new_n462));
  NOR3_X1   g261(.A1(new_n460), .A2(KEYINPUT72), .A3(new_n462), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n451), .B1(new_n459), .B2(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n428), .A2(new_n441), .A3(new_n353), .ZN(new_n465));
  XNOR2_X1  g264(.A(KEYINPUT73), .B(KEYINPUT34), .ZN(new_n466));
  XNOR2_X1  g265(.A(new_n465), .B(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n464), .A2(KEYINPUT74), .A3(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT74), .ZN(new_n469));
  OAI21_X1  g268(.A(KEYINPUT72), .B1(new_n460), .B2(new_n462), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n455), .A2(KEYINPUT32), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n471), .A2(new_n458), .A3(new_n452), .A4(new_n448), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n450), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n467), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n469), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n473), .A2(new_n474), .ZN(new_n476));
  XOR2_X1   g275(.A(G141gat), .B(G148gat), .Z(new_n477));
  INV_X1    g276(.A(G155gat), .ZN(new_n478));
  INV_X1    g277(.A(G162gat), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(G155gat), .A2(G162gat), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(KEYINPUT2), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n477), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  XNOR2_X1  g283(.A(G141gat), .B(G148gat), .ZN(new_n485));
  OAI211_X1 g284(.A(new_n481), .B(new_n480), .C1(new_n485), .C2(KEYINPUT2), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT22), .ZN(new_n488));
  INV_X1    g287(.A(G211gat), .ZN(new_n489));
  INV_X1    g288(.A(G218gat), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n488), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(KEYINPUT76), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT76), .ZN(new_n493));
  OAI211_X1 g292(.A(new_n493), .B(new_n488), .C1(new_n489), .C2(new_n490), .ZN(new_n494));
  XNOR2_X1  g293(.A(G197gat), .B(G204gat), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n492), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  XOR2_X1   g295(.A(G211gat), .B(G218gat), .Z(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(new_n497), .ZN(new_n499));
  NAND4_X1  g298(.A1(new_n499), .A2(new_n492), .A3(new_n494), .A4(new_n495), .ZN(new_n500));
  AOI21_X1  g299(.A(KEYINPUT29), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n487), .B1(new_n501), .B2(KEYINPUT3), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n498), .A2(new_n500), .ZN(new_n503));
  INV_X1    g302(.A(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT29), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n505), .B1(new_n487), .B2(KEYINPUT3), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n502), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(G228gat), .A2(G233gat), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n509), .B1(new_n507), .B2(KEYINPUT83), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT83), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n504), .A2(new_n512), .A3(new_n506), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(new_n487), .ZN(new_n515));
  INV_X1    g314(.A(new_n501), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT82), .ZN(new_n517));
  AOI21_X1  g316(.A(KEYINPUT3), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n501), .A2(KEYINPUT82), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n515), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n510), .B1(new_n514), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(G22gat), .ZN(new_n522));
  INV_X1    g321(.A(G22gat), .ZN(new_n523));
  OAI211_X1 g322(.A(new_n523), .B(new_n510), .C1(new_n514), .C2(new_n520), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g324(.A(KEYINPUT84), .B1(new_n521), .B2(G22gat), .ZN(new_n526));
  XNOR2_X1  g325(.A(G78gat), .B(G106gat), .ZN(new_n527));
  XNOR2_X1  g326(.A(KEYINPUT31), .B(G50gat), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n527), .B(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(new_n529), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n525), .B1(new_n526), .B2(new_n530), .ZN(new_n531));
  NAND4_X1  g330(.A1(new_n522), .A2(KEYINPUT84), .A3(new_n524), .A4(new_n529), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n468), .A2(new_n475), .A3(new_n476), .A4(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(G226gat), .A2(G233gat), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n537), .B1(new_n436), .B2(new_n505), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n536), .B1(new_n427), .B2(new_n405), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n504), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT77), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n436), .A2(new_n537), .ZN(new_n542));
  AOI21_X1  g341(.A(KEYINPUT29), .B1(new_n427), .B2(new_n405), .ZN(new_n543));
  OAI211_X1 g342(.A(new_n542), .B(new_n503), .C1(new_n543), .C2(new_n537), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n540), .A2(new_n541), .A3(new_n544), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n538), .A2(new_n539), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n546), .A2(KEYINPUT77), .A3(new_n503), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(G8gat), .B(G36gat), .ZN(new_n549));
  XNOR2_X1  g348(.A(G64gat), .B(G92gat), .ZN(new_n550));
  XOR2_X1   g349(.A(new_n549), .B(new_n550), .Z(new_n551));
  NAND2_X1  g350(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n551), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n545), .A2(new_n547), .A3(new_n553), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n552), .A2(KEYINPUT30), .A3(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT30), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n548), .A2(new_n556), .A3(new_n551), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT6), .ZN(new_n560));
  XOR2_X1   g359(.A(G1gat), .B(G29gat), .Z(new_n561));
  XNOR2_X1  g360(.A(KEYINPUT78), .B(KEYINPUT0), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n561), .B(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(G57gat), .B(G85gat), .ZN(new_n564));
  XOR2_X1   g363(.A(new_n563), .B(new_n564), .Z(new_n565));
  NAND4_X1  g364(.A1(new_n380), .A2(KEYINPUT4), .A3(new_n389), .A4(new_n515), .ZN(new_n566));
  NAND2_X1  g365(.A1(G225gat), .A2(G233gat), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT3), .ZN(new_n569));
  AND3_X1   g368(.A1(new_n484), .A2(new_n486), .A3(new_n569), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n569), .B1(new_n484), .B2(new_n486), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n387), .A2(new_n388), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n568), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n379), .B1(new_n438), .B2(new_n382), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(new_n515), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT4), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n566), .A2(new_n574), .A3(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT5), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n573), .A2(new_n487), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(new_n576), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n580), .B1(new_n582), .B2(new_n568), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n579), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n380), .A2(new_n389), .A3(new_n515), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n585), .A2(new_n577), .ZN(new_n586));
  NOR3_X1   g385(.A1(new_n573), .A2(new_n577), .A3(new_n487), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  AOI211_X1 g387(.A(KEYINPUT5), .B(new_n568), .C1(new_n572), .C2(new_n573), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n586), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  AOI211_X1 g389(.A(new_n560), .B(new_n565), .C1(new_n584), .C2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n584), .A2(new_n590), .ZN(new_n592));
  INV_X1    g391(.A(new_n565), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT80), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n565), .B1(new_n584), .B2(new_n590), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n597), .A2(KEYINPUT80), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n584), .A2(new_n590), .A3(new_n565), .ZN(new_n599));
  AND3_X1   g398(.A1(new_n599), .A2(KEYINPUT79), .A3(new_n560), .ZN(new_n600));
  AOI21_X1  g399(.A(KEYINPUT79), .B1(new_n599), .B2(new_n560), .ZN(new_n601));
  OAI211_X1 g400(.A(new_n596), .B(new_n598), .C1(new_n600), .C2(new_n601), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n591), .B1(new_n602), .B2(KEYINPUT81), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n599), .A2(new_n560), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT79), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n599), .A2(KEYINPUT79), .A3(new_n560), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n597), .B(new_n595), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT81), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n559), .B1(new_n603), .B2(new_n611), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n349), .B1(new_n535), .B2(new_n612), .ZN(new_n613));
  AND2_X1   g412(.A1(new_n599), .A2(new_n560), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n591), .B1(new_n614), .B2(new_n594), .ZN(new_n615));
  NOR3_X1   g414(.A1(new_n559), .A2(KEYINPUT35), .A3(new_n615), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n464), .A2(new_n467), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n473), .A2(new_n474), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n616), .A2(new_n619), .A3(new_n533), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n613), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT36), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n623), .B1(new_n473), .B2(new_n474), .ZN(new_n624));
  NAND4_X1  g423(.A1(new_n475), .A2(new_n468), .A3(new_n624), .A4(KEYINPUT75), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n623), .B1(new_n617), .B2(new_n618), .ZN(new_n626));
  AND2_X1   g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n475), .A2(new_n468), .A3(new_n624), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT75), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n602), .A2(KEYINPUT81), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n597), .A2(KEYINPUT6), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n631), .A2(new_n611), .A3(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n533), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n633), .A2(new_n634), .A3(new_n558), .ZN(new_n635));
  XOR2_X1   g434(.A(KEYINPUT87), .B(KEYINPUT37), .Z(new_n636));
  NAND2_X1  g435(.A1(new_n548), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT86), .ZN(new_n638));
  AND2_X1   g437(.A1(new_n540), .A2(new_n544), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT37), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n638), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n640), .B1(new_n540), .B2(new_n544), .ZN(new_n642));
  AOI21_X1  g441(.A(KEYINPUT38), .B1(new_n642), .B2(KEYINPUT86), .ZN(new_n643));
  NAND4_X1  g442(.A1(new_n637), .A2(new_n641), .A3(new_n643), .A4(new_n553), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n615), .A2(new_n644), .A3(new_n552), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT38), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n551), .B1(new_n548), .B2(new_n636), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n545), .A2(new_n547), .A3(KEYINPUT37), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n646), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n582), .A2(new_n568), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT39), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NOR3_X1   g451(.A1(new_n575), .A2(new_n570), .A3(new_n571), .ZN(new_n653));
  AOI211_X1 g452(.A(new_n653), .B(new_n587), .C1(new_n585), .C2(new_n577), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n652), .B1(new_n654), .B2(new_n567), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n586), .A2(new_n588), .ZN(new_n656));
  OAI211_X1 g455(.A(new_n651), .B(new_n568), .C1(new_n656), .C2(new_n653), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n655), .A2(new_n565), .A3(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT85), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n659), .A2(KEYINPUT40), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n660), .ZN(new_n662));
  NAND4_X1  g461(.A1(new_n655), .A2(new_n657), .A3(new_n565), .A4(new_n662), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n661), .A2(new_n594), .A3(new_n663), .ZN(new_n664));
  OAI22_X1  g463(.A1(new_n645), .A2(new_n649), .B1(new_n558), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n665), .A2(new_n533), .ZN(new_n666));
  AOI22_X1  g465(.A1(new_n627), .A2(new_n630), .B1(new_n635), .B2(new_n666), .ZN(new_n667));
  OAI211_X1 g466(.A(KEYINPUT95), .B(new_n348), .C1(new_n622), .C2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  AND3_X1   g468(.A1(new_n630), .A2(new_n626), .A3(new_n625), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n587), .B1(new_n585), .B2(new_n577), .ZN(new_n671));
  AOI22_X1  g470(.A1(new_n579), .A2(new_n583), .B1(new_n671), .B2(new_n589), .ZN(new_n672));
  OAI211_X1 g471(.A(new_n599), .B(new_n560), .C1(new_n672), .C2(new_n565), .ZN(new_n673));
  AND3_X1   g472(.A1(new_n673), .A2(new_n632), .A3(new_n552), .ZN(new_n674));
  AND2_X1   g473(.A1(new_n647), .A2(new_n648), .ZN(new_n675));
  OAI211_X1 g474(.A(new_n674), .B(new_n644), .C1(new_n675), .C2(new_n646), .ZN(new_n676));
  AND2_X1   g475(.A1(new_n663), .A2(new_n594), .ZN(new_n677));
  NAND4_X1  g476(.A1(new_n677), .A2(new_n557), .A3(new_n555), .A4(new_n661), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n634), .B1(new_n676), .B2(new_n678), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n679), .B1(new_n612), .B2(new_n634), .ZN(new_n680));
  OAI22_X1  g479(.A1(new_n670), .A2(new_n680), .B1(new_n613), .B2(new_n621), .ZN(new_n681));
  AOI21_X1  g480(.A(KEYINPUT95), .B1(new_n681), .B2(new_n348), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n311), .B1(new_n669), .B2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(KEYINPUT104), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT95), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n633), .A2(new_n558), .ZN(new_n686));
  OAI21_X1  g485(.A(KEYINPUT35), .B1(new_n686), .B2(new_n534), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n635), .A2(new_n666), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n630), .A2(new_n626), .A3(new_n625), .ZN(new_n689));
  AOI22_X1  g488(.A1(new_n687), .A2(new_n620), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(new_n348), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n685), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(new_n668), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT104), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n693), .A2(new_n694), .A3(new_n311), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n684), .A2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(new_n633), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g498(.A(KEYINPUT16), .B(G8gat), .Z(new_n700));
  AOI21_X1  g499(.A(new_n694), .B1(new_n693), .B2(new_n311), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n264), .A2(new_n288), .ZN(new_n702));
  INV_X1    g501(.A(new_n310), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  AOI211_X1 g503(.A(KEYINPUT104), .B(new_n704), .C1(new_n692), .C2(new_n668), .ZN(new_n705));
  OAI221_X1 g504(.A(new_n559), .B1(KEYINPUT42), .B2(new_n700), .C1(new_n701), .C2(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n278), .A2(KEYINPUT42), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT105), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n558), .B1(new_n684), .B2(new_n695), .ZN(new_n710));
  AND2_X1   g509(.A1(new_n700), .A2(KEYINPUT42), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n709), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  OAI211_X1 g511(.A(new_n559), .B(new_n711), .C1(new_n701), .C2(new_n705), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n713), .A2(KEYINPUT105), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n708), .B1(new_n712), .B2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT106), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  OAI211_X1 g516(.A(new_n708), .B(KEYINPUT106), .C1(new_n712), .C2(new_n714), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(G1325gat));
  INV_X1    g518(.A(G15gat), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n696), .A2(new_n720), .A3(new_n619), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n689), .B1(new_n684), .B2(new_n695), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n721), .B1(new_n722), .B2(new_n720), .ZN(G1326gat));
  NAND2_X1  g522(.A1(new_n696), .A2(new_n634), .ZN(new_n724));
  XNOR2_X1  g523(.A(KEYINPUT43), .B(G22gat), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n724), .B(new_n725), .ZN(G1327gat));
  INV_X1    g525(.A(new_n264), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n703), .A2(new_n288), .ZN(new_n728));
  AOI211_X1 g527(.A(new_n727), .B(new_n728), .C1(new_n692), .C2(new_n668), .ZN(new_n729));
  INV_X1    g528(.A(G29gat), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n729), .A2(new_n730), .A3(new_n697), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(KEYINPUT45), .ZN(new_n732));
  AND2_X1   g531(.A1(KEYINPUT107), .A2(KEYINPUT44), .ZN(new_n733));
  NOR2_X1   g532(.A1(KEYINPUT107), .A2(KEYINPUT44), .ZN(new_n734));
  OAI211_X1 g533(.A(new_n681), .B(new_n264), .C1(new_n733), .C2(new_n734), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n690), .A2(new_n727), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n735), .B1(new_n736), .B2(new_n734), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n691), .A2(new_n728), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  OAI21_X1  g538(.A(G29gat), .B1(new_n739), .B2(new_n633), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n732), .A2(new_n740), .ZN(G1328gat));
  INV_X1    g540(.A(G36gat), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n729), .A2(new_n742), .A3(new_n559), .ZN(new_n743));
  OR2_X1    g542(.A1(new_n743), .A2(KEYINPUT46), .ZN(new_n744));
  OAI21_X1  g543(.A(G36gat), .B1(new_n739), .B2(new_n558), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n743), .A2(KEYINPUT46), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n744), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(KEYINPUT108), .ZN(G1329gat));
  INV_X1    g547(.A(KEYINPUT109), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n739), .A2(new_n689), .ZN(new_n750));
  INV_X1    g549(.A(G43gat), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  AND3_X1   g551(.A1(new_n729), .A2(new_n751), .A3(new_n619), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n749), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g554(.A(KEYINPUT48), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n729), .A2(KEYINPUT110), .ZN(new_n757));
  INV_X1    g556(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n533), .A2(G50gat), .ZN(new_n759));
  INV_X1    g558(.A(new_n759), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n760), .B1(new_n729), .B2(KEYINPUT110), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n758), .A2(KEYINPUT111), .A3(new_n761), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n737), .A2(new_n634), .A3(new_n738), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(G50gat), .ZN(new_n764));
  INV_X1    g563(.A(new_n761), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n764), .B1(new_n765), .B2(new_n757), .ZN(new_n766));
  OAI211_X1 g565(.A(new_n756), .B(new_n762), .C1(new_n766), .C2(KEYINPUT111), .ZN(new_n767));
  NOR3_X1   g566(.A1(new_n766), .A2(KEYINPUT112), .A3(new_n756), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT112), .ZN(new_n769));
  AOI22_X1  g568(.A1(new_n758), .A2(new_n761), .B1(G50gat), .B2(new_n763), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n769), .B1(new_n770), .B2(KEYINPUT48), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n767), .B1(new_n768), .B2(new_n771), .ZN(G1331gat));
  NAND2_X1  g571(.A1(new_n691), .A2(new_n310), .ZN(new_n773));
  INV_X1    g572(.A(new_n773), .ZN(new_n774));
  AND3_X1   g573(.A1(new_n681), .A2(new_n774), .A3(new_n702), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(new_n697), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g576(.A(new_n558), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n775), .A2(new_n778), .ZN(new_n779));
  XOR2_X1   g578(.A(new_n779), .B(KEYINPUT113), .Z(new_n780));
  NOR2_X1   g579(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n780), .B(new_n781), .ZN(G1333gat));
  NAND2_X1  g581(.A1(new_n775), .A2(new_n670), .ZN(new_n783));
  OR2_X1    g582(.A1(new_n617), .A2(new_n618), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n784), .A2(G71gat), .ZN(new_n785));
  AOI22_X1  g584(.A1(new_n783), .A2(G71gat), .B1(new_n775), .B2(new_n785), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n786), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g586(.A1(new_n775), .A2(new_n634), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n788), .B(G78gat), .ZN(G1335gat));
  INV_X1    g588(.A(new_n288), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT114), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT51), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n790), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n736), .A2(new_n691), .A3(new_n793), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n791), .A2(new_n792), .ZN(new_n795));
  OR2_X1    g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n794), .A2(new_n795), .ZN(new_n797));
  AND2_X1   g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n697), .A2(new_n234), .A3(new_n310), .ZN(new_n800));
  AND3_X1   g599(.A1(new_n737), .A2(new_n288), .A3(new_n774), .ZN(new_n801));
  AND2_X1   g600(.A1(new_n801), .A2(new_n697), .ZN(new_n802));
  OAI22_X1  g601(.A1(new_n799), .A2(new_n800), .B1(new_n802), .B2(new_n234), .ZN(G1336gat));
  NAND4_X1  g602(.A1(new_n798), .A2(new_n235), .A3(new_n559), .A4(new_n310), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n801), .A2(new_n559), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(G92gat), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n804), .A2(KEYINPUT115), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n807), .A2(new_n808), .A3(KEYINPUT52), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT52), .ZN(new_n810));
  OAI211_X1 g609(.A(new_n804), .B(new_n806), .C1(KEYINPUT115), .C2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n809), .A2(new_n811), .ZN(G1337gat));
  INV_X1    g611(.A(G99gat), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n619), .A2(new_n813), .A3(new_n310), .ZN(new_n814));
  AND2_X1   g613(.A1(new_n801), .A2(new_n670), .ZN(new_n815));
  OAI22_X1  g614(.A1(new_n799), .A2(new_n814), .B1(new_n815), .B2(new_n813), .ZN(G1338gat));
  NAND2_X1  g615(.A1(new_n801), .A2(new_n634), .ZN(new_n817));
  XNOR2_X1  g616(.A(KEYINPUT116), .B(G106gat), .ZN(new_n818));
  INV_X1    g617(.A(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  NOR3_X1   g619(.A1(new_n703), .A2(G106gat), .A3(new_n533), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n798), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  OR2_X1    g622(.A1(KEYINPUT117), .A2(KEYINPUT53), .ZN(new_n824));
  NAND2_X1  g623(.A1(KEYINPUT117), .A2(KEYINPUT53), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n823), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  NAND4_X1  g625(.A1(new_n820), .A2(new_n822), .A3(KEYINPUT117), .A4(KEYINPUT53), .ZN(new_n827));
  AND2_X1   g626(.A1(new_n826), .A2(new_n827), .ZN(G1339gat));
  INV_X1    g627(.A(new_n263), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n291), .A2(new_n292), .A3(new_n298), .ZN(new_n830));
  AND2_X1   g629(.A1(new_n830), .A2(KEYINPUT54), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n296), .A2(new_n831), .A3(new_n305), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT54), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n302), .B1(new_n303), .B2(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n832), .A2(new_n834), .A3(KEYINPUT55), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT118), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n835), .A2(new_n836), .A3(new_n306), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n832), .A2(new_n834), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT55), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n837), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n836), .B1(new_n835), .B2(new_n306), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n330), .A2(new_n317), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n325), .A2(new_n327), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(new_n342), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n329), .A2(new_n331), .A3(new_n344), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND4_X1  g648(.A1(new_n829), .A2(new_n843), .A3(new_n849), .A4(new_n261), .ZN(new_n850));
  AOI22_X1  g649(.A1(new_n348), .A2(new_n843), .B1(new_n849), .B2(new_n310), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n850), .B1(new_n851), .B2(new_n264), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(new_n288), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n311), .A2(new_n691), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n633), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(new_n535), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n856), .A2(new_n559), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n857), .A2(new_n385), .A3(new_n348), .ZN(new_n858));
  AOI22_X1  g657(.A1(new_n852), .A2(new_n288), .B1(new_n311), .B2(new_n691), .ZN(new_n859));
  NOR3_X1   g658(.A1(new_n859), .A2(new_n784), .A3(new_n634), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n633), .A2(new_n559), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  OAI21_X1  g661(.A(G113gat), .B1(new_n862), .B2(new_n691), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n858), .A2(new_n863), .ZN(G1340gat));
  NAND2_X1  g663(.A1(new_n310), .A2(new_n362), .ZN(new_n865));
  XNOR2_X1  g664(.A(new_n865), .B(KEYINPUT120), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n857), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n860), .A2(new_n310), .A3(new_n861), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT119), .ZN(new_n869));
  AND3_X1   g668(.A1(new_n868), .A2(new_n869), .A3(G120gat), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n869), .B1(new_n868), .B2(G120gat), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n867), .B1(new_n870), .B2(new_n871), .ZN(G1341gat));
  INV_X1    g671(.A(G127gat), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n857), .A2(new_n873), .A3(new_n790), .ZN(new_n874));
  OAI21_X1  g673(.A(G127gat), .B1(new_n862), .B2(new_n288), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(G1342gat));
  OR4_X1    g675(.A1(G134gat), .A2(new_n856), .A3(new_n559), .A4(new_n727), .ZN(new_n877));
  OR2_X1    g676(.A1(new_n877), .A2(KEYINPUT56), .ZN(new_n878));
  OAI21_X1  g677(.A(G134gat), .B1(new_n862), .B2(new_n727), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n877), .A2(KEYINPUT56), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(G1343gat));
  INV_X1    g680(.A(KEYINPUT123), .ZN(new_n882));
  INV_X1    g681(.A(G141gat), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n689), .A2(new_n861), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT57), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n533), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n847), .A2(new_n848), .A3(new_n310), .ZN(new_n887));
  OR2_X1    g686(.A1(new_n887), .A2(KEYINPUT121), .ZN(new_n888));
  AND3_X1   g687(.A1(new_n840), .A2(new_n306), .A3(new_n835), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n348), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n887), .A2(KEYINPUT121), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n888), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(new_n727), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n790), .B1(new_n893), .B2(new_n850), .ZN(new_n894));
  INV_X1    g693(.A(new_n854), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n886), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n885), .B1(new_n859), .B2(new_n533), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n884), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n883), .B1(new_n898), .B2(new_n348), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n689), .A2(new_n634), .ZN(new_n900));
  INV_X1    g699(.A(new_n900), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n691), .A2(G141gat), .ZN(new_n902));
  NAND4_X1  g701(.A1(new_n855), .A2(new_n558), .A3(new_n901), .A4(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT122), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NOR3_X1   g704(.A1(new_n859), .A2(new_n633), .A3(new_n900), .ZN(new_n906));
  NAND4_X1  g705(.A1(new_n906), .A2(KEYINPUT122), .A3(new_n558), .A4(new_n902), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT58), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n905), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n882), .B1(new_n899), .B2(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(new_n884), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n853), .A2(new_n854), .ZN(new_n912));
  AOI21_X1  g711(.A(KEYINPUT57), .B1(new_n912), .B2(new_n634), .ZN(new_n913));
  INV_X1    g712(.A(new_n886), .ZN(new_n914));
  AOI22_X1  g713(.A1(new_n348), .A2(new_n889), .B1(new_n887), .B2(KEYINPUT121), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n264), .B1(new_n915), .B2(new_n888), .ZN(new_n916));
  INV_X1    g715(.A(new_n850), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n288), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n914), .B1(new_n918), .B2(new_n854), .ZN(new_n919));
  OAI211_X1 g718(.A(new_n348), .B(new_n911), .C1(new_n913), .C2(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(G141gat), .ZN(new_n921));
  INV_X1    g720(.A(new_n903), .ZN(new_n922));
  AOI21_X1  g721(.A(KEYINPUT58), .B1(new_n922), .B2(KEYINPUT122), .ZN(new_n923));
  NAND4_X1  g722(.A1(new_n921), .A2(new_n923), .A3(KEYINPUT123), .A4(new_n905), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n910), .A2(new_n924), .ZN(new_n925));
  OAI21_X1  g724(.A(KEYINPUT58), .B1(new_n899), .B2(new_n922), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n925), .A2(new_n926), .ZN(G1344gat));
  INV_X1    g726(.A(G148gat), .ZN(new_n928));
  NAND4_X1  g727(.A1(new_n906), .A2(new_n928), .A3(new_n558), .A4(new_n310), .ZN(new_n929));
  XOR2_X1   g728(.A(new_n929), .B(KEYINPUT124), .Z(new_n930));
  XOR2_X1   g729(.A(KEYINPUT125), .B(KEYINPUT59), .Z(new_n931));
  NAND2_X1  g730(.A1(new_n918), .A2(new_n854), .ZN(new_n932));
  AOI21_X1  g731(.A(KEYINPUT57), .B1(new_n932), .B2(new_n634), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n859), .A2(new_n914), .ZN(new_n934));
  OR2_X1    g733(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n935), .A2(new_n310), .A3(new_n911), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n931), .B1(new_n936), .B2(G148gat), .ZN(new_n937));
  AOI211_X1 g736(.A(KEYINPUT59), .B(new_n928), .C1(new_n898), .C2(new_n310), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n930), .B1(new_n937), .B2(new_n938), .ZN(G1345gat));
  NAND4_X1  g738(.A1(new_n906), .A2(new_n478), .A3(new_n558), .A4(new_n790), .ZN(new_n940));
  AND2_X1   g739(.A1(new_n898), .A2(new_n790), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n940), .B1(new_n941), .B2(new_n478), .ZN(G1346gat));
  NAND4_X1  g741(.A1(new_n906), .A2(new_n479), .A3(new_n558), .A4(new_n264), .ZN(new_n943));
  XOR2_X1   g742(.A(new_n943), .B(KEYINPUT126), .Z(new_n944));
  AND2_X1   g743(.A1(new_n898), .A2(new_n264), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n944), .B1(new_n479), .B2(new_n945), .ZN(G1347gat));
  NOR2_X1   g745(.A1(new_n697), .A2(new_n558), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n860), .A2(new_n947), .ZN(new_n948));
  NOR3_X1   g747(.A1(new_n948), .A2(new_n411), .A3(new_n691), .ZN(new_n949));
  AOI21_X1  g748(.A(KEYINPUT127), .B1(new_n912), .B2(new_n633), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n950), .A2(new_n558), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n912), .A2(KEYINPUT127), .A3(new_n633), .ZN(new_n952));
  AND2_X1   g751(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n953), .A2(new_n535), .A3(new_n348), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n949), .B1(new_n954), .B2(new_n411), .ZN(G1348gat));
  OAI21_X1  g754(.A(G176gat), .B1(new_n948), .B2(new_n703), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n951), .A2(new_n535), .A3(new_n952), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n310), .A2(new_n412), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n956), .B1(new_n957), .B2(new_n958), .ZN(G1349gat));
  OAI21_X1  g758(.A(G183gat), .B1(new_n948), .B2(new_n288), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n790), .A2(new_n402), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n960), .B1(new_n957), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n962), .A2(KEYINPUT60), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT60), .ZN(new_n964));
  OAI211_X1 g763(.A(new_n964), .B(new_n960), .C1(new_n957), .C2(new_n961), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n963), .A2(new_n965), .ZN(G1350gat));
  NAND3_X1  g765(.A1(new_n860), .A2(new_n264), .A3(new_n947), .ZN(new_n967));
  INV_X1    g766(.A(KEYINPUT61), .ZN(new_n968));
  AND3_X1   g767(.A1(new_n967), .A2(new_n968), .A3(G190gat), .ZN(new_n969));
  AOI21_X1  g768(.A(new_n968), .B1(new_n967), .B2(G190gat), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n264), .A2(new_n403), .ZN(new_n971));
  OAI22_X1  g770(.A1(new_n969), .A2(new_n970), .B1(new_n957), .B2(new_n971), .ZN(G1351gat));
  NAND3_X1  g771(.A1(new_n953), .A2(new_n348), .A3(new_n901), .ZN(new_n973));
  AND2_X1   g772(.A1(new_n689), .A2(new_n947), .ZN(new_n974));
  AND2_X1   g773(.A1(new_n935), .A2(new_n974), .ZN(new_n975));
  NOR2_X1   g774(.A1(new_n691), .A2(new_n339), .ZN(new_n976));
  AOI22_X1  g775(.A1(new_n973), .A2(new_n339), .B1(new_n975), .B2(new_n976), .ZN(G1352gat));
  NAND3_X1  g776(.A1(new_n951), .A2(new_n901), .A3(new_n952), .ZN(new_n978));
  NOR2_X1   g777(.A1(new_n703), .A2(G204gat), .ZN(new_n979));
  INV_X1    g778(.A(new_n979), .ZN(new_n980));
  OR3_X1    g779(.A1(new_n978), .A2(KEYINPUT62), .A3(new_n980), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n935), .A2(new_n310), .A3(new_n974), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n982), .A2(G204gat), .ZN(new_n983));
  OAI21_X1  g782(.A(KEYINPUT62), .B1(new_n978), .B2(new_n980), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n981), .A2(new_n983), .A3(new_n984), .ZN(G1353gat));
  OAI211_X1 g784(.A(new_n790), .B(new_n974), .C1(new_n933), .C2(new_n934), .ZN(new_n986));
  AND3_X1   g785(.A1(new_n986), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n987));
  AOI21_X1  g786(.A(KEYINPUT63), .B1(new_n986), .B2(G211gat), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n790), .A2(new_n489), .ZN(new_n989));
  OAI22_X1  g788(.A1(new_n987), .A2(new_n988), .B1(new_n978), .B2(new_n989), .ZN(G1354gat));
  NAND3_X1  g789(.A1(new_n935), .A2(new_n264), .A3(new_n974), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n991), .A2(G218gat), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n264), .A2(new_n490), .ZN(new_n993));
  OAI21_X1  g792(.A(new_n992), .B1(new_n978), .B2(new_n993), .ZN(G1355gat));
endmodule


