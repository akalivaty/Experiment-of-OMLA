//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1 0 1 1 1 0 1 0 0 1 0 1 1 1 0 0 0 1 0 1 1 0 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 0 1 0 0 1 1 0 0 0 0 1 0 0 1 0 0 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:32 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1231,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1289, new_n1290, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1296;
  XOR2_X1   g0000(.A(KEYINPUT64), .B(G50), .Z(new_n201));
  NOR3_X1   g0001(.A1(new_n201), .A2(G58), .A3(G68), .ZN(new_n202));
  INV_X1    g0002(.A(G77), .ZN(new_n203));
  AND2_X1   g0003(.A1(new_n202), .A2(new_n203), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n207));
  INV_X1    g0007(.A(G68), .ZN(new_n208));
  INV_X1    g0008(.A(G238), .ZN(new_n209));
  INV_X1    g0009(.A(G87), .ZN(new_n210));
  INV_X1    g0010(.A(G250), .ZN(new_n211));
  OAI221_X1 g0011(.A(new_n207), .B1(new_n208), .B2(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n213));
  INV_X1    g0013(.A(G244), .ZN(new_n214));
  INV_X1    g0014(.A(G107), .ZN(new_n215));
  INV_X1    g0015(.A(G264), .ZN(new_n216));
  OAI221_X1 g0016(.A(new_n213), .B1(new_n203), .B2(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n206), .B1(new_n212), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n218), .A2(KEYINPUT1), .ZN(new_n219));
  XOR2_X1   g0019(.A(new_n219), .B(KEYINPUT65), .Z(new_n220));
  NOR2_X1   g0020(.A1(new_n206), .A2(G13), .ZN(new_n221));
  OAI211_X1 g0021(.A(new_n221), .B(G250), .C1(G257), .C2(G264), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT0), .ZN(new_n223));
  OAI21_X1  g0023(.A(G50), .B1(G58), .B2(G68), .ZN(new_n224));
  INV_X1    g0024(.A(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  INV_X1    g0026(.A(G20), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n225), .A2(new_n228), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n223), .B(new_n229), .C1(KEYINPUT1), .C2(new_n218), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n220), .A2(new_n230), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XNOR2_X1  g0039(.A(G68), .B(G77), .ZN(new_n240));
  INV_X1    g0040(.A(G58), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(KEYINPUT66), .B(G50), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XOR2_X1   g0045(.A(G107), .B(G116), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  AND2_X1   g0048(.A1(KEYINPUT3), .A2(G33), .ZN(new_n249));
  NOR2_X1   g0049(.A1(KEYINPUT3), .A2(G33), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n251), .A2(G1698), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(G222), .ZN(new_n253));
  XNOR2_X1  g0053(.A(KEYINPUT3), .B(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(G1698), .ZN(new_n255));
  XOR2_X1   g0055(.A(KEYINPUT67), .B(G223), .Z(new_n256));
  OAI221_X1 g0056(.A(new_n253), .B1(new_n203), .B2(new_n254), .C1(new_n255), .C2(new_n256), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n226), .B1(G33), .B2(G41), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(new_n258), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(G274), .ZN(new_n261));
  INV_X1    g0061(.A(G41), .ZN(new_n262));
  INV_X1    g0062(.A(G45), .ZN(new_n263));
  AOI21_X1  g0063(.A(G1), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n261), .A2(new_n265), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n258), .A2(new_n264), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n266), .B1(G226), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n259), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(G190), .ZN(new_n271));
  INV_X1    g0071(.A(G200), .ZN(new_n272));
  NOR2_X1   g0072(.A1(G20), .A2(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(G150), .ZN(new_n274));
  INV_X1    g0074(.A(G33), .ZN(new_n275));
  OR3_X1    g0075(.A1(new_n275), .A2(KEYINPUT70), .A3(G20), .ZN(new_n276));
  OAI21_X1  g0076(.A(KEYINPUT70), .B1(new_n275), .B2(G20), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  XNOR2_X1  g0078(.A(KEYINPUT8), .B(G58), .ZN(new_n279));
  OAI221_X1 g0079(.A(new_n274), .B1(new_n278), .B2(new_n279), .C1(new_n202), .C2(new_n227), .ZN(new_n280));
  NAND3_X1  g0080(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT68), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND4_X1  g0083(.A1(KEYINPUT68), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n283), .A2(new_n226), .A3(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(KEYINPUT69), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT69), .ZN(new_n287));
  NAND4_X1  g0087(.A1(new_n283), .A2(new_n287), .A3(new_n226), .A4(new_n284), .ZN(new_n288));
  AND2_X1   g0088(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G50), .ZN(new_n290));
  INV_X1    g0090(.A(G13), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n291), .A2(G1), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(G20), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  AOI22_X1  g0094(.A1(new_n280), .A2(new_n289), .B1(new_n290), .B2(new_n294), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n289), .A2(new_n294), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n227), .A2(G1), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n296), .A2(G50), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n295), .A2(new_n299), .ZN(new_n300));
  AND2_X1   g0100(.A1(new_n300), .A2(KEYINPUT9), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n300), .A2(KEYINPUT9), .ZN(new_n302));
  OAI221_X1 g0102(.A(new_n271), .B1(new_n272), .B2(new_n270), .C1(new_n301), .C2(new_n302), .ZN(new_n303));
  XNOR2_X1  g0103(.A(new_n303), .B(KEYINPUT10), .ZN(new_n304));
  INV_X1    g0104(.A(G179), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n270), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(G169), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n269), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n306), .A2(new_n300), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n304), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n296), .A2(G68), .A3(new_n298), .ZN(new_n311));
  AOI22_X1  g0111(.A1(new_n273), .A2(G50), .B1(G20), .B2(new_n208), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n312), .B1(new_n278), .B2(new_n203), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n289), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT11), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n294), .A2(new_n208), .ZN(new_n317));
  XNOR2_X1  g0117(.A(new_n317), .B(KEYINPUT12), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n289), .A2(KEYINPUT11), .A3(new_n313), .ZN(new_n319));
  NAND4_X1  g0119(.A1(new_n311), .A2(new_n316), .A3(new_n318), .A4(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(G274), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n258), .A2(new_n321), .ZN(new_n322));
  AOI22_X1  g0122(.A1(G238), .A2(new_n267), .B1(new_n322), .B2(new_n264), .ZN(new_n323));
  INV_X1    g0123(.A(G1698), .ZN(new_n324));
  OAI211_X1 g0124(.A(G226), .B(new_n324), .C1(new_n249), .C2(new_n250), .ZN(new_n325));
  OAI211_X1 g0125(.A(G232), .B(G1698), .C1(new_n249), .C2(new_n250), .ZN(new_n326));
  NAND2_X1  g0126(.A1(G33), .A2(G97), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n325), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT72), .ZN(new_n329));
  AND3_X1   g0129(.A1(new_n328), .A2(new_n329), .A3(new_n258), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n329), .B1(new_n328), .B2(new_n258), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n323), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT13), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n333), .A2(KEYINPUT73), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n332), .A2(new_n335), .ZN(new_n336));
  OAI211_X1 g0136(.A(new_n323), .B(new_n334), .C1(new_n330), .C2(new_n331), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n305), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT14), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n332), .A2(KEYINPUT13), .ZN(new_n340));
  OAI211_X1 g0140(.A(new_n333), .B(new_n323), .C1(new_n330), .C2(new_n331), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n307), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n338), .B1(new_n339), .B2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT74), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n344), .B1(new_n342), .B2(new_n339), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  NOR3_X1   g0146(.A1(new_n342), .A2(new_n344), .A3(new_n339), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n320), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(G190), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n349), .B1(new_n336), .B2(new_n337), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n272), .B1(new_n340), .B2(new_n341), .ZN(new_n351));
  OR3_X1    g0151(.A1(new_n350), .A2(new_n351), .A3(new_n320), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n348), .A2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT75), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n279), .A2(new_n297), .ZN(new_n356));
  AOI22_X1  g0156(.A1(new_n296), .A2(new_n356), .B1(new_n294), .B2(new_n279), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n275), .A2(KEYINPUT76), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT76), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(G33), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n359), .A2(new_n361), .A3(KEYINPUT3), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n275), .A2(KEYINPUT3), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(KEYINPUT77), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT77), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n362), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT7), .ZN(new_n370));
  AOI21_X1  g0170(.A(G20), .B1(new_n370), .B2(KEYINPUT78), .ZN(new_n371));
  OAI211_X1 g0171(.A(new_n369), .B(new_n371), .C1(KEYINPUT78), .C2(new_n370), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT78), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n367), .B1(new_n362), .B2(new_n364), .ZN(new_n374));
  XNOR2_X1  g0174(.A(KEYINPUT76), .B(G33), .ZN(new_n375));
  AOI21_X1  g0175(.A(KEYINPUT77), .B1(new_n375), .B2(KEYINPUT3), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  OAI211_X1 g0177(.A(new_n373), .B(KEYINPUT7), .C1(new_n377), .C2(G20), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n372), .A2(new_n378), .A3(G68), .ZN(new_n379));
  NAND2_X1  g0179(.A1(G58), .A2(G68), .ZN(new_n380));
  XNOR2_X1  g0180(.A(new_n380), .B(KEYINPUT79), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n381), .B1(G58), .B2(G68), .ZN(new_n382));
  AOI22_X1  g0182(.A1(new_n382), .A2(G20), .B1(G159), .B2(new_n273), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n379), .A2(KEYINPUT16), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n286), .A2(new_n288), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n251), .A2(new_n227), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT3), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n375), .A2(new_n387), .ZN(new_n388));
  NOR3_X1   g0188(.A1(new_n249), .A2(new_n370), .A3(G20), .ZN(new_n389));
  AOI22_X1  g0189(.A1(new_n370), .A2(new_n386), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n383), .B1(new_n208), .B2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT16), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n385), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n358), .B1(new_n384), .B2(new_n393), .ZN(new_n394));
  OR2_X1    g0194(.A1(new_n324), .A2(G226), .ZN(new_n395));
  OAI211_X1 g0195(.A(new_n377), .B(new_n395), .C1(G223), .C2(G1698), .ZN(new_n396));
  NAND2_X1  g0196(.A1(G33), .A2(G87), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n260), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n267), .A2(G232), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n399), .B1(new_n261), .B2(new_n265), .ZN(new_n400));
  NOR3_X1   g0200(.A1(new_n398), .A2(new_n349), .A3(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  OAI21_X1  g0202(.A(G200), .B1(new_n398), .B2(new_n400), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n394), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  OR2_X1    g0204(.A1(KEYINPUT80), .A2(KEYINPUT17), .ZN(new_n405));
  NAND2_X1  g0205(.A1(KEYINPUT80), .A2(KEYINPUT17), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n404), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  NOR3_X1   g0207(.A1(new_n398), .A2(new_n305), .A3(new_n400), .ZN(new_n408));
  INV_X1    g0208(.A(new_n408), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n398), .A2(new_n400), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n409), .B1(new_n307), .B2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT18), .ZN(new_n412));
  INV_X1    g0212(.A(new_n394), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(new_n410), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n408), .B1(new_n415), .B2(G169), .ZN(new_n416));
  OAI21_X1  g0216(.A(KEYINPUT18), .B1(new_n416), .B2(new_n394), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n401), .B1(new_n415), .B2(G200), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n418), .A2(new_n394), .A3(KEYINPUT80), .A4(KEYINPUT17), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n407), .A2(new_n414), .A3(new_n417), .A4(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n266), .B1(G244), .B2(new_n267), .ZN(new_n421));
  OAI22_X1  g0221(.A1(new_n255), .A2(new_n209), .B1(new_n215), .B2(new_n254), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n422), .B1(G232), .B2(new_n252), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n421), .B1(new_n423), .B2(new_n260), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(G200), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n425), .B1(new_n349), .B2(new_n424), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n296), .A2(G77), .A3(new_n298), .ZN(new_n427));
  INV_X1    g0227(.A(new_n279), .ZN(new_n428));
  AOI22_X1  g0228(.A1(new_n428), .A2(new_n273), .B1(G20), .B2(G77), .ZN(new_n429));
  XNOR2_X1  g0229(.A(KEYINPUT15), .B(G87), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n429), .B1(new_n430), .B2(new_n278), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(new_n289), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n294), .A2(new_n203), .ZN(new_n433));
  XNOR2_X1  g0233(.A(new_n433), .B(KEYINPUT71), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n427), .A2(new_n432), .A3(new_n434), .ZN(new_n435));
  OR2_X1    g0235(.A1(new_n426), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n424), .A2(new_n307), .ZN(new_n437));
  OAI211_X1 g0237(.A(new_n435), .B(new_n437), .C1(G179), .C2(new_n424), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  NOR4_X1   g0239(.A1(new_n310), .A2(new_n355), .A3(new_n420), .A4(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n353), .A2(new_n354), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  AND2_X1   g0242(.A1(G257), .A2(G1698), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n363), .B1(new_n375), .B2(KEYINPUT3), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n368), .B(new_n443), .C1(new_n444), .C2(new_n367), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(KEYINPUT84), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n366), .A2(G250), .A3(new_n324), .A4(new_n368), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n359), .A2(new_n361), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(G294), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT84), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n366), .A2(new_n450), .A3(new_n368), .A4(new_n443), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n446), .A2(new_n447), .A3(new_n449), .A4(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(new_n258), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n263), .A2(G1), .ZN(new_n454));
  XNOR2_X1  g0254(.A(KEYINPUT5), .B(G41), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n322), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n454), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(new_n260), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n458), .A2(new_n216), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n453), .A2(new_n305), .A3(new_n456), .A4(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT22), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n227), .A2(G87), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n462), .B1(new_n251), .B2(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n448), .A2(new_n227), .A3(G116), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT82), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n466), .B1(new_n227), .B2(G107), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT23), .ZN(new_n468));
  OR2_X1    g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n467), .A2(new_n468), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n464), .A2(new_n465), .A3(new_n469), .A4(new_n470), .ZN(new_n471));
  NOR3_X1   g0271(.A1(new_n374), .A2(new_n376), .A3(G20), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n462), .A2(new_n210), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n471), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n289), .B1(new_n474), .B2(KEYINPUT24), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n366), .A2(new_n227), .A3(new_n368), .A4(new_n473), .ZN(new_n476));
  AND3_X1   g0276(.A1(new_n465), .A2(new_n469), .A3(new_n470), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n476), .A2(new_n464), .A3(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT24), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(G1), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(G33), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n385), .A2(G107), .A3(new_n293), .A4(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT83), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n293), .A2(G107), .ZN(new_n485));
  XNOR2_X1  g0285(.A(new_n485), .B(KEYINPUT25), .ZN(new_n486));
  AND3_X1   g0286(.A1(new_n483), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n484), .B1(new_n483), .B2(new_n486), .ZN(new_n488));
  OAI22_X1  g0288(.A1(new_n475), .A2(new_n480), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n261), .A2(new_n457), .ZN(new_n490));
  AOI211_X1 g0290(.A(new_n490), .B(new_n459), .C1(new_n452), .C2(new_n258), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n461), .B(new_n489), .C1(new_n491), .C2(G169), .ZN(new_n492));
  INV_X1    g0292(.A(new_n458), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n490), .B1(G257), .B2(new_n493), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n254), .A2(KEYINPUT4), .A3(G244), .A4(new_n324), .ZN(new_n495));
  NAND2_X1  g0295(.A1(G33), .A2(G283), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n254), .A2(G250), .A3(G1698), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n495), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n366), .A2(G244), .A3(new_n324), .A4(new_n368), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT4), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n305), .B(new_n494), .C1(new_n501), .C2(new_n260), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n390), .A2(new_n215), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n273), .A2(G77), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT6), .ZN(new_n505));
  INV_X1    g0305(.A(G97), .ZN(new_n506));
  NOR3_X1   g0306(.A1(new_n505), .A2(new_n506), .A3(G107), .ZN(new_n507));
  XNOR2_X1  g0307(.A(G97), .B(G107), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n507), .B1(new_n505), .B2(new_n508), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n504), .B1(new_n509), .B2(new_n227), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n289), .B1(new_n503), .B2(new_n510), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n385), .A2(G97), .A3(new_n293), .A4(new_n482), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n294), .A2(new_n506), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n511), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(new_n494), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n499), .A2(new_n500), .ZN(new_n516));
  INV_X1    g0316(.A(new_n498), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n515), .B1(new_n518), .B2(new_n258), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n502), .B(new_n514), .C1(new_n519), .C2(G169), .ZN(new_n520));
  INV_X1    g0320(.A(new_n514), .ZN(new_n521));
  OAI211_X1 g0321(.A(G190), .B(new_n494), .C1(new_n501), .C2(new_n260), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n521), .B(new_n522), .C1(new_n519), .C2(new_n272), .ZN(new_n523));
  AND3_X1   g0323(.A1(new_n492), .A2(new_n520), .A3(new_n523), .ZN(new_n524));
  NOR2_X1   g0324(.A1(G238), .A2(G1698), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n525), .B1(new_n214), .B2(G1698), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  NOR3_X1   g0327(.A1(new_n374), .A2(new_n376), .A3(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(G116), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n375), .A2(new_n529), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n258), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n454), .A2(new_n211), .ZN(new_n532));
  AOI22_X1  g0332(.A1(new_n322), .A2(new_n454), .B1(new_n260), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n531), .A2(G179), .A3(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(new_n533), .ZN(new_n535));
  INV_X1    g0335(.A(new_n530), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n536), .B1(new_n369), .B2(new_n527), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n535), .B1(new_n537), .B2(new_n258), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n534), .B1(new_n538), .B2(new_n307), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT81), .ZN(new_n540));
  OR2_X1    g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n377), .A2(new_n227), .A3(G68), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n276), .A2(G97), .A3(new_n277), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT19), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n227), .B1(new_n327), .B2(new_n544), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n210), .A2(new_n506), .A3(new_n215), .ZN(new_n546));
  AOI22_X1  g0346(.A1(new_n543), .A2(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n385), .B1(new_n542), .B2(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(new_n430), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n549), .A2(new_n293), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n296), .A2(new_n482), .A3(new_n549), .ZN(new_n552));
  AOI22_X1  g0352(.A1(new_n539), .A2(new_n540), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  AND4_X1   g0353(.A1(G87), .A2(new_n385), .A3(new_n293), .A4(new_n482), .ZN(new_n554));
  NOR3_X1   g0354(.A1(new_n548), .A2(new_n554), .A3(new_n550), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n272), .B1(new_n531), .B2(new_n533), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n556), .B1(G190), .B2(new_n538), .ZN(new_n557));
  AOI22_X1  g0357(.A1(new_n541), .A2(new_n553), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n227), .A2(G116), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n275), .A2(G97), .ZN(new_n560));
  AOI21_X1  g0360(.A(G20), .B1(G33), .B2(G283), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n559), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(new_n285), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT20), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n562), .A2(new_n285), .A3(KEYINPUT20), .ZN(new_n566));
  AOI22_X1  g0366(.A1(new_n565), .A2(new_n566), .B1(new_n292), .B2(new_n559), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n385), .A2(G116), .A3(new_n293), .A4(new_n482), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(new_n569), .ZN(new_n570));
  NOR2_X1   g0370(.A1(G257), .A2(G1698), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n571), .B1(new_n216), .B2(G1698), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n368), .B(new_n572), .C1(new_n444), .C2(new_n367), .ZN(new_n573));
  INV_X1    g0373(.A(G303), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n254), .A2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(new_n575), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n260), .B1(new_n573), .B2(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(G270), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n456), .B1(new_n578), .B2(new_n458), .ZN(new_n579));
  OAI21_X1  g0379(.A(G200), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n573), .A2(new_n576), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(new_n258), .ZN(new_n582));
  INV_X1    g0382(.A(new_n579), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n570), .B(new_n580), .C1(new_n584), .C2(new_n349), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT21), .ZN(new_n586));
  OAI21_X1  g0386(.A(G169), .B1(new_n577), .B2(new_n579), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n586), .B1(new_n570), .B2(new_n587), .ZN(new_n588));
  NOR3_X1   g0388(.A1(new_n577), .A2(new_n305), .A3(new_n579), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(new_n569), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n584), .A2(KEYINPUT21), .A3(new_n569), .A4(G169), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n585), .A2(new_n588), .A3(new_n590), .A4(new_n591), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n489), .B1(G190), .B2(new_n491), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n453), .A2(new_n456), .A3(new_n460), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(G200), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n592), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n524), .A2(new_n558), .A3(new_n596), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n442), .A2(new_n597), .ZN(G372));
  INV_X1    g0398(.A(new_n309), .ZN(new_n599));
  AND2_X1   g0399(.A1(new_n348), .A2(new_n438), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n407), .A2(new_n352), .A3(new_n419), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n417), .B(new_n414), .C1(new_n600), .C2(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n599), .B1(new_n602), .B2(new_n304), .ZN(new_n603));
  INV_X1    g0403(.A(new_n480), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n385), .B1(new_n478), .B2(new_n479), .ZN(new_n605));
  INV_X1    g0405(.A(new_n488), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n483), .A2(new_n484), .A3(new_n486), .ZN(new_n607));
  AOI22_X1  g0407(.A1(new_n604), .A2(new_n605), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n459), .B1(new_n452), .B2(new_n258), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n609), .A2(G190), .A3(new_n456), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n595), .A2(new_n608), .A3(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(new_n550), .ZN(new_n612));
  AND2_X1   g0412(.A1(new_n542), .A2(new_n547), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n552), .B(new_n612), .C1(new_n613), .C2(new_n385), .ZN(new_n614));
  AOI22_X1  g0414(.A1(new_n557), .A2(new_n555), .B1(new_n539), .B2(new_n614), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n611), .A2(new_n520), .A3(new_n615), .A4(new_n523), .ZN(new_n616));
  AND3_X1   g0416(.A1(new_n588), .A2(new_n590), .A3(new_n591), .ZN(new_n617));
  AND2_X1   g0417(.A1(new_n492), .A2(new_n617), .ZN(new_n618));
  OAI21_X1  g0418(.A(KEYINPUT85), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(new_n556), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n531), .A2(new_n533), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n555), .B(new_n620), .C1(new_n349), .C2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n539), .A2(new_n614), .ZN(new_n623));
  AND4_X1   g0423(.A1(new_n520), .A2(new_n523), .A3(new_n622), .A4(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT85), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n492), .A2(new_n617), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n624), .A2(new_n625), .A3(new_n611), .A4(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n619), .A2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT26), .ZN(new_n629));
  INV_X1    g0429(.A(new_n520), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n629), .B1(new_n558), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n615), .A2(new_n630), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n623), .B1(new_n632), .B2(KEYINPUT26), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  AND2_X1   g0434(.A1(new_n628), .A2(new_n634), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n603), .B1(new_n442), .B2(new_n635), .ZN(G369));
  INV_X1    g0436(.A(new_n617), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n292), .A2(new_n227), .ZN(new_n638));
  OR2_X1    g0438(.A1(new_n638), .A2(KEYINPUT27), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(KEYINPUT27), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n639), .A2(G213), .A3(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(G343), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n570), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n637), .A2(new_n645), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n646), .B1(new_n592), .B2(new_n645), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(G330), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n611), .B1(new_n608), .B2(new_n644), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(new_n492), .ZN(new_n650));
  OR2_X1    g0450(.A1(new_n492), .A2(new_n643), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n648), .A2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n637), .A2(new_n644), .ZN(new_n655));
  OR2_X1    g0455(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n654), .A2(new_n651), .A3(new_n656), .ZN(G399));
  NAND3_X1  g0457(.A1(new_n558), .A2(new_n630), .A3(new_n629), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n632), .A2(KEYINPUT26), .ZN(new_n659));
  AND3_X1   g0459(.A1(new_n658), .A2(new_n623), .A3(new_n659), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n624), .A2(new_n611), .A3(new_n626), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n643), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT29), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n643), .B1(new_n628), .B2(new_n634), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n664), .B1(new_n663), .B2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT30), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n453), .A2(new_n460), .A3(new_n589), .A4(new_n538), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n494), .B1(new_n501), .B2(new_n260), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n667), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  OAI211_X1 g0470(.A(KEYINPUT30), .B(new_n494), .C1(new_n501), .C2(new_n260), .ZN(new_n671));
  OAI21_X1  g0471(.A(KEYINPUT86), .B1(new_n668), .B2(new_n671), .ZN(new_n672));
  AND3_X1   g0472(.A1(new_n584), .A2(new_n305), .A3(new_n621), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n673), .A2(new_n594), .A3(new_n669), .ZN(new_n674));
  INV_X1    g0474(.A(new_n671), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n582), .A2(G179), .A3(new_n583), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n676), .A2(new_n621), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT86), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n675), .A2(new_n677), .A3(new_n678), .A4(new_n609), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n670), .A2(new_n672), .A3(new_n674), .A4(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(new_n643), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT31), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n524), .A2(new_n596), .A3(new_n558), .A4(new_n644), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n680), .A2(KEYINPUT31), .A3(new_n643), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n683), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(G330), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT87), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n686), .A2(KEYINPUT87), .A3(G330), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n666), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(new_n481), .ZN(new_n694));
  INV_X1    g0494(.A(new_n221), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n695), .A2(G41), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n546), .A2(G116), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n697), .A2(G1), .A3(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n699), .B1(new_n224), .B2(new_n697), .ZN(new_n700));
  XNOR2_X1  g0500(.A(new_n700), .B(KEYINPUT28), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n694), .A2(new_n701), .ZN(G364));
  NOR2_X1   g0502(.A1(new_n291), .A2(G20), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n481), .B1(new_n703), .B2(G45), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n696), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n226), .B1(G20), .B2(new_n307), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n227), .A2(G190), .ZN(new_n710));
  NOR2_X1   g0510(.A1(G179), .A2(G200), .ZN(new_n711));
  AND2_X1   g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  OR2_X1    g0512(.A1(new_n712), .A2(KEYINPUT89), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(KEYINPUT89), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  OR2_X1    g0516(.A1(new_n716), .A2(KEYINPUT93), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(KEYINPUT93), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(G329), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n227), .A2(new_n305), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(G200), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n723), .A2(new_n349), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  XNOR2_X1  g0525(.A(KEYINPUT91), .B(G326), .ZN(new_n726));
  INV_X1    g0526(.A(G294), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n227), .B1(new_n711), .B2(G190), .ZN(new_n728));
  OAI22_X1  g0528(.A1(new_n725), .A2(new_n726), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT92), .ZN(new_n730));
  OR2_X1    g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n227), .A2(new_n349), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n305), .A2(G200), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(G322), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n251), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n272), .A2(G179), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n732), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n710), .A2(new_n733), .ZN(new_n739));
  INV_X1    g0539(.A(G311), .ZN(new_n740));
  OAI22_X1  g0540(.A1(new_n738), .A2(new_n574), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n710), .A2(new_n737), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  AOI211_X1 g0543(.A(new_n736), .B(new_n741), .C1(G283), .C2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT90), .ZN(new_n745));
  INV_X1    g0545(.A(new_n723), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n745), .B1(new_n746), .B2(new_n349), .ZN(new_n747));
  NOR3_X1   g0547(.A1(new_n723), .A2(KEYINPUT90), .A3(G190), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  XNOR2_X1  g0550(.A(KEYINPUT33), .B(G317), .ZN(new_n751));
  AOI22_X1  g0551(.A1(new_n750), .A2(new_n751), .B1(new_n730), .B2(new_n729), .ZN(new_n752));
  NAND4_X1  g0552(.A1(new_n721), .A2(new_n731), .A3(new_n744), .A4(new_n752), .ZN(new_n753));
  OAI22_X1  g0553(.A1(new_n725), .A2(new_n290), .B1(new_n728), .B2(new_n506), .ZN(new_n754));
  INV_X1    g0554(.A(new_n739), .ZN(new_n755));
  AOI22_X1  g0555(.A1(G77), .A2(new_n755), .B1(new_n743), .B2(G107), .ZN(new_n756));
  OAI211_X1 g0556(.A(new_n756), .B(new_n254), .C1(new_n210), .C2(new_n738), .ZN(new_n757));
  XNOR2_X1  g0557(.A(new_n734), .B(KEYINPUT88), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  AOI211_X1 g0559(.A(new_n754), .B(new_n757), .C1(G58), .C2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(G159), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n715), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g0562(.A(new_n762), .B(KEYINPUT32), .ZN(new_n763));
  OAI211_X1 g0563(.A(new_n760), .B(new_n763), .C1(new_n208), .C2(new_n749), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n709), .B1(new_n753), .B2(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(G13), .A2(G33), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n767), .A2(G20), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(new_n708), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n244), .A2(G45), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n377), .A2(new_n695), .ZN(new_n771));
  OAI211_X1 g0571(.A(new_n770), .B(new_n771), .C1(G45), .C2(new_n224), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n695), .A2(new_n251), .ZN(new_n773));
  AOI22_X1  g0573(.A1(new_n773), .A2(G355), .B1(new_n529), .B2(new_n695), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  AOI211_X1 g0575(.A(new_n707), .B(new_n765), .C1(new_n769), .C2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n768), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n776), .B1(new_n647), .B2(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n706), .B1(new_n647), .B2(G330), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n779), .B1(G330), .B2(new_n647), .ZN(new_n780));
  AND2_X1   g0580(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(G396));
  NAND3_X1  g0582(.A1(new_n435), .A2(KEYINPUT94), .A3(new_n643), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n435), .A2(new_n643), .ZN(new_n784));
  INV_X1    g0584(.A(KEYINPUT94), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n436), .A2(new_n783), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(new_n438), .ZN(new_n788));
  OR2_X1    g0588(.A1(new_n438), .A2(new_n643), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  XNOR2_X1  g0591(.A(new_n665), .B(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n706), .B1(new_n692), .B2(new_n792), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n793), .B1(new_n692), .B2(new_n792), .ZN(new_n794));
  OAI221_X1 g0594(.A(new_n251), .B1(new_n728), .B2(new_n506), .C1(new_n529), .C2(new_n739), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n743), .A2(G87), .ZN(new_n796));
  OAI221_X1 g0596(.A(new_n796), .B1(new_n215), .B2(new_n738), .C1(new_n727), .C2(new_n734), .ZN(new_n797));
  AOI211_X1 g0597(.A(new_n795), .B(new_n797), .C1(G303), .C2(new_n724), .ZN(new_n798));
  INV_X1    g0598(.A(G283), .ZN(new_n799));
  OAI221_X1 g0599(.A(new_n798), .B1(new_n799), .B2(new_n749), .C1(new_n719), .C2(new_n740), .ZN(new_n800));
  AOI22_X1  g0600(.A1(new_n724), .A2(G137), .B1(new_n755), .B2(G159), .ZN(new_n801));
  INV_X1    g0601(.A(G143), .ZN(new_n802));
  INV_X1    g0602(.A(G150), .ZN(new_n803));
  OAI221_X1 g0603(.A(new_n801), .B1(new_n802), .B2(new_n758), .C1(new_n749), .C2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(KEYINPUT34), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n743), .A2(G68), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n807), .B1(new_n290), .B2(new_n738), .ZN(new_n808));
  INV_X1    g0608(.A(new_n728), .ZN(new_n809));
  AOI211_X1 g0609(.A(new_n369), .B(new_n808), .C1(G58), .C2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(G132), .ZN(new_n811));
  OAI211_X1 g0611(.A(new_n806), .B(new_n810), .C1(new_n719), .C2(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n804), .A2(new_n805), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n800), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n814), .A2(new_n708), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n708), .A2(new_n766), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n707), .B1(new_n203), .B2(new_n816), .ZN(new_n817));
  OAI211_X1 g0617(.A(new_n815), .B(new_n817), .C1(new_n791), .C2(new_n767), .ZN(new_n818));
  AND2_X1   g0618(.A1(new_n794), .A2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(G384));
  INV_X1    g0620(.A(new_n509), .ZN(new_n821));
  OR2_X1    g0621(.A1(new_n821), .A2(KEYINPUT35), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n821), .A2(KEYINPUT35), .ZN(new_n823));
  NAND4_X1  g0623(.A1(new_n822), .A2(G116), .A3(new_n228), .A4(new_n823), .ZN(new_n824));
  XOR2_X1   g0624(.A(new_n824), .B(KEYINPUT36), .Z(new_n825));
  INV_X1    g0625(.A(new_n201), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n826), .A2(G68), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n381), .A2(G77), .A3(new_n225), .ZN(new_n828));
  AOI211_X1 g0628(.A(new_n481), .B(G13), .C1(new_n827), .C2(new_n828), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n825), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n320), .A2(new_n643), .ZN(new_n831));
  XOR2_X1   g0631(.A(new_n831), .B(KEYINPUT96), .Z(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n353), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n348), .A2(new_n352), .A3(new_n832), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n790), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT99), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n681), .A2(new_n837), .A3(new_n682), .ZN(new_n838));
  OAI211_X1 g0638(.A(new_n680), .B(new_n643), .C1(KEYINPUT99), .C2(KEYINPUT31), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n838), .A2(new_n684), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n836), .A2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT37), .ZN(new_n842));
  AOI21_X1  g0642(.A(KEYINPUT16), .B1(new_n379), .B2(new_n383), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT97), .ZN(new_n844));
  OR3_X1    g0644(.A1(new_n843), .A2(new_n844), .A3(new_n385), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n844), .B1(new_n843), .B2(new_n385), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n845), .A2(new_n384), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n847), .A2(new_n357), .ZN(new_n848));
  INV_X1    g0648(.A(new_n641), .ZN(new_n849));
  AOI22_X1  g0649(.A1(new_n848), .A2(new_n849), .B1(new_n394), .B2(new_n418), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n848), .A2(new_n411), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n842), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n404), .B1(new_n394), .B2(new_n416), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n394), .A2(new_n641), .ZN(new_n854));
  NOR3_X1   g0654(.A1(new_n853), .A2(KEYINPUT37), .A3(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT98), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n641), .B1(new_n847), .B2(new_n357), .ZN(new_n857));
  AND3_X1   g0657(.A1(new_n420), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n856), .B1(new_n420), .B2(new_n857), .ZN(new_n859));
  OAI22_X1  g0659(.A1(new_n852), .A2(new_n855), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT38), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  OAI221_X1 g0662(.A(KEYINPUT38), .B1(new_n858), .B2(new_n859), .C1(new_n852), .C2(new_n855), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n841), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  OR2_X1    g0664(.A1(new_n864), .A2(KEYINPUT40), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n420), .A2(new_n854), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n853), .A2(new_n854), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n867), .A2(new_n842), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n866), .B1(new_n868), .B2(new_n855), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n869), .A2(new_n861), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n870), .B1(new_n860), .B2(new_n861), .ZN(new_n871));
  NAND4_X1  g0671(.A1(new_n871), .A2(KEYINPUT40), .A3(new_n840), .A4(new_n836), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n865), .A2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(new_n840), .ZN(new_n874));
  OR3_X1    g0674(.A1(new_n873), .A2(new_n442), .A3(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n873), .B1(new_n442), .B2(new_n874), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n875), .A2(G330), .A3(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT39), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n871), .A2(new_n878), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n348), .A2(new_n643), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n862), .A2(new_n863), .A3(KEYINPUT39), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n834), .A2(new_n835), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  AOI211_X1 g0684(.A(new_n643), .B(new_n790), .C1(new_n628), .C2(new_n634), .ZN(new_n885));
  INV_X1    g0685(.A(new_n789), .ZN(new_n886));
  OAI21_X1  g0686(.A(KEYINPUT95), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n665), .A2(new_n791), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT95), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n888), .A2(new_n889), .A3(new_n789), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n884), .B1(new_n887), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n862), .A2(new_n863), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n414), .A2(new_n417), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n641), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n882), .A2(new_n893), .A3(new_n895), .ZN(new_n896));
  OR2_X1    g0696(.A1(new_n666), .A2(new_n442), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(new_n603), .ZN(new_n898));
  XNOR2_X1  g0698(.A(new_n896), .B(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n877), .A2(new_n899), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n900), .B1(new_n481), .B2(new_n703), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n877), .A2(new_n899), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n830), .B1(new_n901), .B2(new_n902), .ZN(G367));
  INV_X1    g0703(.A(KEYINPUT102), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n520), .A2(new_n644), .ZN(new_n905));
  XNOR2_X1  g0705(.A(new_n905), .B(KEYINPUT103), .ZN(new_n906));
  OAI211_X1 g0706(.A(new_n523), .B(new_n520), .C1(new_n521), .C2(new_n644), .ZN(new_n907));
  AND2_X1   g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  OR3_X1    g0708(.A1(new_n656), .A2(KEYINPUT42), .A3(new_n908), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n520), .B1(new_n908), .B2(new_n492), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(new_n644), .ZN(new_n911));
  OAI21_X1  g0711(.A(KEYINPUT42), .B1(new_n656), .B2(new_n908), .ZN(new_n912));
  AND3_X1   g0712(.A1(new_n911), .A2(new_n912), .A3(KEYINPUT104), .ZN(new_n913));
  AOI21_X1  g0713(.A(KEYINPUT104), .B1(new_n911), .B2(new_n912), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n909), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT105), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  OAI211_X1 g0717(.A(KEYINPUT105), .B(new_n909), .C1(new_n913), .C2(new_n914), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n555), .A2(new_n644), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  AND2_X1   g0721(.A1(new_n615), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n921), .A2(new_n623), .ZN(new_n923));
  OR3_X1    g0723(.A1(new_n922), .A2(KEYINPUT100), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n923), .A2(KEYINPUT100), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n924), .A2(KEYINPUT43), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n904), .B1(new_n919), .B2(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(new_n926), .ZN(new_n929));
  AOI211_X1 g0729(.A(KEYINPUT102), .B(new_n929), .C1(new_n917), .C2(new_n918), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n924), .A2(new_n925), .ZN(new_n932));
  XNOR2_X1  g0732(.A(KEYINPUT101), .B(KEYINPUT43), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n928), .A2(new_n931), .A3(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n934), .B1(new_n927), .B2(new_n930), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n654), .A2(new_n908), .ZN(new_n939));
  INV_X1    g0739(.A(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n936), .A2(new_n937), .A3(new_n939), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n656), .A2(new_n651), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(new_n908), .ZN(new_n944));
  XOR2_X1   g0744(.A(new_n944), .B(KEYINPUT44), .Z(new_n945));
  NOR2_X1   g0745(.A1(new_n943), .A2(new_n908), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n946), .B(KEYINPUT45), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n948), .B(new_n654), .ZN(new_n949));
  AOI21_X1  g0749(.A(KEYINPUT106), .B1(new_n652), .B2(new_n655), .ZN(new_n950));
  XOR2_X1   g0750(.A(new_n950), .B(new_n648), .Z(new_n951));
  XNOR2_X1  g0751(.A(new_n951), .B(new_n656), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n693), .B1(new_n949), .B2(new_n953), .ZN(new_n954));
  XOR2_X1   g0754(.A(new_n696), .B(KEYINPUT41), .Z(new_n955));
  OAI21_X1  g0755(.A(new_n704), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n941), .A2(new_n942), .A3(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n932), .A2(new_n768), .ZN(new_n958));
  AOI22_X1  g0758(.A1(new_n750), .A2(G159), .B1(new_n201), .B2(new_n755), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(KEYINPUT109), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n716), .A2(G137), .ZN(new_n961));
  OAI22_X1  g0761(.A1(new_n725), .A2(new_n802), .B1(new_n728), .B2(new_n208), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n254), .B1(new_n738), .B2(new_n241), .ZN(new_n963));
  OAI22_X1  g0763(.A1(new_n734), .A2(new_n803), .B1(new_n742), .B2(new_n203), .ZN(new_n964));
  NOR3_X1   g0764(.A1(new_n962), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n960), .A2(new_n961), .A3(new_n965), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n959), .A2(KEYINPUT109), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n758), .A2(new_n574), .ZN(new_n968));
  INV_X1    g0768(.A(new_n738), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n969), .A2(KEYINPUT46), .A3(G116), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT46), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n971), .B1(new_n738), .B2(new_n529), .ZN(new_n972));
  OAI211_X1 g0772(.A(new_n970), .B(new_n972), .C1(new_n725), .C2(new_n740), .ZN(new_n973));
  OAI22_X1  g0773(.A1(new_n739), .A2(new_n799), .B1(new_n728), .B2(new_n215), .ZN(new_n974));
  NOR3_X1   g0774(.A1(new_n968), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  XOR2_X1   g0775(.A(KEYINPUT107), .B(G317), .Z(new_n976));
  OAI221_X1 g0776(.A(new_n369), .B1(new_n506), .B2(new_n742), .C1(new_n715), .C2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT108), .ZN(new_n978));
  OAI221_X1 g0778(.A(new_n975), .B1(new_n727), .B2(new_n749), .C1(new_n977), .C2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n977), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n980), .A2(KEYINPUT108), .ZN(new_n981));
  OAI22_X1  g0781(.A1(new_n966), .A2(new_n967), .B1(new_n979), .B2(new_n981), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(KEYINPUT47), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(new_n708), .ZN(new_n984));
  INV_X1    g0784(.A(new_n771), .ZN(new_n985));
  OAI221_X1 g0785(.A(new_n769), .B1(new_n221), .B2(new_n430), .C1(new_n985), .C2(new_n238), .ZN(new_n986));
  NAND4_X1  g0786(.A1(new_n958), .A2(new_n706), .A3(new_n984), .A4(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n957), .A2(new_n987), .ZN(G387));
  OAI221_X1 g0788(.A(new_n369), .B1(new_n529), .B2(new_n742), .C1(new_n715), .C2(new_n726), .ZN(new_n989));
  AOI22_X1  g0789(.A1(new_n724), .A2(G322), .B1(new_n755), .B2(G303), .ZN(new_n990));
  OAI221_X1 g0790(.A(new_n990), .B1(new_n758), .B2(new_n976), .C1(new_n749), .C2(new_n740), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT48), .ZN(new_n992));
  OR2_X1    g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n991), .A2(new_n992), .ZN(new_n994));
  AOI22_X1  g0794(.A1(new_n969), .A2(G294), .B1(new_n809), .B2(G283), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n993), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n989), .B1(new_n997), .B2(KEYINPUT49), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n998), .B1(KEYINPUT49), .B2(new_n997), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n728), .A2(new_n430), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n734), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(G50), .A2(new_n1001), .B1(new_n755), .B2(G68), .ZN(new_n1002));
  OAI221_X1 g0802(.A(new_n1002), .B1(new_n203), .B2(new_n738), .C1(new_n506), .C2(new_n742), .ZN(new_n1003));
  AOI211_X1 g0803(.A(new_n1000), .B(new_n1003), .C1(G159), .C2(new_n724), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n369), .B1(new_n750), .B2(new_n428), .ZN(new_n1005));
  OAI211_X1 g0805(.A(new_n1004), .B(new_n1005), .C1(new_n803), .C2(new_n715), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n709), .B1(new_n999), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n698), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(new_n773), .A2(new_n1008), .B1(new_n215), .B2(new_n695), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n235), .A2(new_n263), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n428), .A2(new_n290), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1011), .B(KEYINPUT50), .ZN(new_n1012));
  OAI211_X1 g0812(.A(new_n698), .B(new_n263), .C1(new_n208), .C2(new_n203), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n771), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1009), .B1(new_n1010), .B2(new_n1014), .ZN(new_n1015));
  AOI211_X1 g0815(.A(new_n707), .B(new_n1007), .C1(new_n769), .C2(new_n1015), .ZN(new_n1016));
  XOR2_X1   g0816(.A(new_n1016), .B(KEYINPUT110), .Z(new_n1017));
  AOI21_X1  g0817(.A(new_n1017), .B1(new_n652), .B2(new_n768), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1018), .B1(new_n953), .B2(new_n705), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n952), .A2(new_n693), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1021), .A2(new_n696), .ZN(new_n1022));
  AND2_X1   g0822(.A1(new_n952), .A2(new_n693), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1019), .B1(new_n1022), .B2(new_n1023), .ZN(G393));
  INV_X1    g0824(.A(new_n949), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1025), .A2(new_n1021), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n697), .B1(new_n949), .B2(new_n1020), .ZN(new_n1027));
  AND2_X1   g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n908), .A2(new_n768), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT111), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n716), .A2(G143), .B1(G68), .B2(new_n969), .ZN(new_n1031));
  OR2_X1    g0831(.A1(new_n1031), .A2(KEYINPUT112), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1031), .A2(KEYINPUT112), .ZN(new_n1033));
  NAND4_X1  g0833(.A1(new_n1032), .A2(new_n377), .A3(new_n1033), .A4(new_n796), .ZN(new_n1034));
  XOR2_X1   g0834(.A(new_n1034), .B(KEYINPUT113), .Z(new_n1035));
  AOI22_X1  g0835(.A1(new_n724), .A2(G150), .B1(new_n1001), .B2(G159), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT51), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n755), .A2(new_n428), .B1(new_n809), .B2(G77), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1038), .B1(new_n749), .B2(new_n826), .ZN(new_n1039));
  NOR3_X1   g0839(.A1(new_n1035), .A2(new_n1037), .A3(new_n1039), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n724), .A2(G317), .B1(new_n1001), .B2(G311), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1041), .B(KEYINPUT52), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n251), .B1(new_n742), .B2(new_n215), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n738), .A2(new_n799), .B1(new_n739), .B2(new_n727), .ZN(new_n1044));
  AOI211_X1 g0844(.A(new_n1043), .B(new_n1044), .C1(G116), .C2(new_n809), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1045), .B1(new_n735), .B2(new_n715), .ZN(new_n1046));
  AOI211_X1 g0846(.A(new_n1042), .B(new_n1046), .C1(G303), .C2(new_n750), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n708), .B1(new_n1040), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n771), .A2(new_n247), .ZN(new_n1049));
  OAI211_X1 g0849(.A(new_n1049), .B(new_n769), .C1(new_n506), .C2(new_n221), .ZN(new_n1050));
  NAND4_X1  g0850(.A1(new_n1030), .A2(new_n706), .A3(new_n1048), .A4(new_n1050), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1051), .B1(new_n1025), .B2(new_n704), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n1028), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n1053), .ZN(G390));
  AOI21_X1  g0854(.A(new_n767), .B1(new_n879), .B2(new_n881), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n816), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n720), .A2(G294), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n734), .A2(new_n529), .B1(new_n728), .B2(new_n203), .ZN(new_n1058));
  XOR2_X1   g0858(.A(new_n1058), .B(KEYINPUT120), .Z(new_n1059));
  NOR2_X1   g0859(.A1(new_n749), .A2(new_n215), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n725), .A2(new_n799), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n254), .B1(new_n969), .B2(G87), .ZN(new_n1062));
  OAI211_X1 g0862(.A(new_n1062), .B(new_n807), .C1(new_n506), .C2(new_n739), .ZN(new_n1063));
  NOR4_X1   g0863(.A1(new_n1059), .A2(new_n1060), .A3(new_n1061), .A4(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n720), .A2(G125), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n724), .A2(G128), .ZN(new_n1066));
  OR3_X1    g0866(.A1(new_n738), .A2(KEYINPUT53), .A3(new_n803), .ZN(new_n1067));
  OAI21_X1  g0867(.A(KEYINPUT53), .B1(new_n738), .B2(new_n803), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n809), .A2(G159), .ZN(new_n1069));
  NAND4_X1  g0869(.A1(new_n1066), .A2(new_n1067), .A3(new_n1068), .A4(new_n1069), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(KEYINPUT54), .B(G143), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n251), .B1(new_n755), .B2(new_n1072), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n1073), .B1(new_n811), .B2(new_n734), .C1(new_n826), .C2(new_n742), .ZN(new_n1074));
  AOI211_X1 g0874(.A(new_n1070), .B(new_n1074), .C1(G137), .C2(new_n750), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n1057), .A2(new_n1064), .B1(new_n1065), .B2(new_n1075), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n706), .B1(new_n428), .B2(new_n1056), .C1(new_n1076), .C2(new_n709), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n1055), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n879), .A2(new_n881), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1079), .B1(new_n891), .B2(new_n880), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n790), .B1(new_n689), .B2(new_n690), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1081), .A2(new_n883), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n662), .A2(new_n788), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1083), .A2(new_n789), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n880), .B1(new_n1084), .B2(new_n883), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(new_n871), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1080), .A2(new_n1082), .A3(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n887), .A2(new_n890), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1088), .A2(new_n883), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n880), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n1091), .A2(new_n1079), .B1(new_n871), .B2(new_n1085), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n836), .A2(G330), .A3(new_n840), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1093), .A2(KEYINPUT114), .ZN(new_n1094));
  INV_X1    g0894(.A(KEYINPUT114), .ZN(new_n1095));
  NAND4_X1  g0895(.A1(new_n836), .A2(new_n1095), .A3(G330), .A4(new_n840), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1097), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n1087), .B(new_n705), .C1(new_n1092), .C2(new_n1098), .ZN(new_n1099));
  OR2_X1    g0899(.A1(new_n1099), .A2(KEYINPUT119), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1099), .A2(KEYINPUT119), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1078), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n840), .A2(G330), .A3(new_n791), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(new_n884), .ZN(new_n1104));
  AND4_X1   g0904(.A1(new_n789), .A2(new_n1082), .A3(new_n1083), .A4(new_n1104), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n883), .B1(new_n691), .B2(new_n791), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1088), .B1(new_n1106), .B2(new_n1097), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1107), .A2(KEYINPUT116), .ZN(new_n1108));
  INV_X1    g0908(.A(KEYINPUT116), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n1109), .B(new_n1088), .C1(new_n1106), .C2(new_n1097), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1105), .B1(new_n1108), .B2(new_n1110), .ZN(new_n1111));
  NAND4_X1  g0911(.A1(new_n440), .A2(G330), .A3(new_n441), .A4(new_n840), .ZN(new_n1112));
  INV_X1    g0912(.A(KEYINPUT115), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(new_n1112), .B(new_n1113), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1114), .A2(new_n603), .A3(new_n897), .ZN(new_n1115));
  OAI21_X1  g0915(.A(KEYINPUT117), .B1(new_n1111), .B2(new_n1115), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n1082), .A2(new_n789), .A3(new_n1083), .A4(new_n1104), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1110), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n1096), .B(new_n1094), .C1(new_n1081), .C2(new_n883), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1109), .B1(new_n1119), .B2(new_n1088), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1117), .B1(new_n1118), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(KEYINPUT117), .ZN(new_n1122));
  AND3_X1   g0922(.A1(new_n1114), .A2(new_n603), .A3(new_n897), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1121), .A2(new_n1122), .A3(new_n1123), .ZN(new_n1124));
  AND3_X1   g0924(.A1(new_n1116), .A2(KEYINPUT118), .A3(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(KEYINPUT118), .B1(new_n1116), .B2(new_n1124), .ZN(new_n1126));
  AND3_X1   g0926(.A1(new_n1080), .A2(new_n1082), .A3(new_n1086), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1098), .B1(new_n1080), .B2(new_n1086), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NOR3_X1   g0929(.A1(new_n1125), .A2(new_n1126), .A3(new_n1129), .ZN(new_n1130));
  NOR3_X1   g0930(.A1(new_n1111), .A2(KEYINPUT117), .A3(new_n1115), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1122), .B1(new_n1121), .B2(new_n1123), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1129), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1133), .A2(new_n696), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1102), .B1(new_n1130), .B2(new_n1134), .ZN(G378));
  NAND2_X1  g0935(.A1(new_n300), .A2(new_n849), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1136), .B1(new_n304), .B2(new_n309), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n304), .A2(new_n309), .A3(new_n1136), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1140));
  AND3_X1   g0940(.A1(new_n1138), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1140), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(KEYINPUT123), .ZN(new_n1144));
  INV_X1    g0944(.A(KEYINPUT123), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1145), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1144), .A2(new_n1146), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n865), .A2(G330), .A3(new_n1147), .A4(new_n872), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n872), .B(G330), .C1(KEYINPUT40), .C2(new_n864), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1149), .A2(new_n1143), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1148), .A2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n896), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1148), .A2(new_n1150), .A3(new_n896), .ZN(new_n1154));
  AND2_X1   g0954(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1144), .A2(new_n766), .A3(new_n1146), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n706), .B1(new_n201), .B2(new_n1056), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n743), .A2(G58), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(new_n1158), .B(KEYINPUT121), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n725), .A2(new_n529), .B1(new_n728), .B2(new_n208), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n262), .B1(new_n738), .B2(new_n203), .ZN(new_n1161));
  OAI22_X1  g0961(.A1(new_n734), .A2(new_n215), .B1(new_n739), .B2(new_n430), .ZN(new_n1162));
  NOR4_X1   g0962(.A1(new_n1159), .A2(new_n1160), .A3(new_n1161), .A4(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n377), .B1(new_n750), .B2(G97), .ZN(new_n1164));
  OAI211_X1 g0964(.A(new_n1163), .B(new_n1164), .C1(new_n719), .C2(new_n799), .ZN(new_n1165));
  XOR2_X1   g0965(.A(new_n1165), .B(KEYINPUT122), .Z(new_n1166));
  OR2_X1    g0966(.A1(new_n1166), .A2(KEYINPUT58), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1166), .A2(KEYINPUT58), .ZN(new_n1168));
  OAI211_X1 g0968(.A(new_n275), .B(new_n262), .C1(new_n742), .C2(new_n761), .ZN(new_n1169));
  AND2_X1   g0969(.A1(new_n716), .A2(G124), .ZN(new_n1170));
  INV_X1    g0970(.A(G128), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n1171), .A2(new_n734), .B1(new_n738), .B2(new_n1071), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1172), .B1(G137), .B2(new_n755), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(new_n724), .A2(G125), .B1(G150), .B2(new_n809), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n1173), .B(new_n1174), .C1(new_n749), .C2(new_n811), .ZN(new_n1175));
  AOI211_X1 g0975(.A(new_n1169), .B(new_n1170), .C1(KEYINPUT59), .C2(new_n1175), .ZN(new_n1176));
  OR2_X1    g0976(.A1(new_n1175), .A2(KEYINPUT59), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n262), .B1(new_n369), .B2(new_n275), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n1176), .A2(new_n1177), .B1(new_n290), .B2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1167), .A2(new_n1168), .A3(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1157), .B1(new_n1180), .B2(new_n708), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(new_n1155), .A2(new_n705), .B1(new_n1156), .B2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1133), .A2(new_n1123), .ZN(new_n1183));
  AOI21_X1  g0983(.A(KEYINPUT57), .B1(new_n1183), .B2(new_n1155), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1116), .A2(new_n1124), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1115), .B1(new_n1185), .B2(new_n1129), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1153), .A2(KEYINPUT57), .A3(new_n1154), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n696), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1182), .B1(new_n1184), .B2(new_n1188), .ZN(G375));
  INV_X1    g0989(.A(KEYINPUT118), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1185), .A2(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n955), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1116), .A2(KEYINPUT118), .A3(new_n1124), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1111), .A2(new_n1115), .ZN(new_n1194));
  NAND4_X1  g0994(.A1(new_n1191), .A2(new_n1192), .A3(new_n1193), .A4(new_n1194), .ZN(new_n1195));
  XOR2_X1   g0995(.A(new_n1195), .B(KEYINPUT124), .Z(new_n1196));
  OAI22_X1  g0996(.A1(new_n738), .A2(new_n506), .B1(new_n739), .B2(new_n215), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n251), .B1(new_n742), .B2(new_n203), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n1198), .A2(new_n1000), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1199), .B1(new_n727), .B2(new_n725), .ZN(new_n1200));
  AOI211_X1 g1000(.A(new_n1197), .B(new_n1200), .C1(G283), .C2(new_n1001), .ZN(new_n1201));
  OAI221_X1 g1001(.A(new_n1201), .B1(new_n529), .B2(new_n749), .C1(new_n719), .C2(new_n574), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n719), .A2(new_n1171), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1159), .B1(G137), .B2(new_n759), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n728), .A2(new_n290), .ZN(new_n1205));
  OAI22_X1  g1005(.A1(new_n738), .A2(new_n761), .B1(new_n739), .B2(new_n803), .ZN(new_n1206));
  AOI211_X1 g1006(.A(new_n1205), .B(new_n1206), .C1(G132), .C2(new_n724), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n369), .B1(new_n750), .B2(new_n1072), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1204), .A2(new_n1207), .A3(new_n1208), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1202), .B1(new_n1203), .B2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1210), .A2(new_n708), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n707), .B1(new_n208), .B2(new_n816), .ZN(new_n1212));
  OAI211_X1 g1012(.A(new_n1211), .B(new_n1212), .C1(new_n883), .C2(new_n767), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1213), .B1(new_n1111), .B2(new_n704), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1196), .A2(new_n1215), .ZN(G381));
  INV_X1    g1016(.A(G375), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n957), .A2(new_n987), .A3(new_n1053), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  XNOR2_X1  g1019(.A(new_n1099), .B(KEYINPUT119), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1078), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1087), .B1(new_n1092), .B2(new_n1098), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1191), .A2(new_n1223), .A3(new_n1193), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1223), .B1(new_n1116), .B2(new_n1124), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1225), .A2(new_n697), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1222), .B1(new_n1224), .B2(new_n1226), .ZN(new_n1227));
  NOR3_X1   g1027(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1217), .A2(new_n1219), .A3(new_n1227), .A4(new_n1228), .ZN(new_n1229));
  OR2_X1    g1029(.A1(new_n1229), .A2(G381), .ZN(G407));
  NAND3_X1  g1030(.A1(new_n1217), .A2(new_n642), .A3(new_n1227), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(G407), .A2(G213), .A3(new_n1231), .ZN(G409));
  OAI211_X1 g1032(.A(new_n1155), .B(new_n1192), .C1(new_n1225), .C2(new_n1115), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(new_n1182), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1224), .A2(new_n1226), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1234), .A2(new_n1235), .A3(new_n1102), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1236), .B1(G375), .B2(new_n1227), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT125), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  OAI211_X1 g1039(.A(new_n1155), .B(KEYINPUT57), .C1(new_n1225), .C2(new_n1115), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1241), .B1(new_n1133), .B2(new_n1123), .ZN(new_n1242));
  OAI211_X1 g1042(.A(new_n1240), .B(new_n696), .C1(new_n1242), .C2(KEYINPUT57), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1243), .A2(G378), .A3(new_n1182), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1244), .A2(KEYINPUT125), .A3(new_n1236), .ZN(new_n1245));
  INV_X1    g1045(.A(G213), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1246), .A2(G343), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1247), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1239), .A2(new_n1245), .A3(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT60), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n696), .B1(new_n1194), .B2(new_n1250), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1116), .A2(KEYINPUT60), .A3(new_n1124), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1251), .B1(new_n1252), .B2(new_n1194), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n819), .B1(new_n1253), .B2(new_n1214), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  NOR3_X1   g1055(.A1(new_n1253), .A2(new_n819), .A3(new_n1214), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  AND2_X1   g1057(.A1(new_n1247), .A2(G2897), .ZN(new_n1258));
  AND2_X1   g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1249), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1261));
  NAND4_X1  g1061(.A1(new_n1239), .A2(new_n1257), .A3(new_n1245), .A4(new_n1248), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT63), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1247), .B1(new_n1244), .B2(new_n1236), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1265), .A2(KEYINPUT63), .A3(new_n1257), .ZN(new_n1266));
  XNOR2_X1  g1066(.A(G393), .B(new_n781), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1218), .A2(KEYINPUT126), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1053), .B1(new_n957), .B2(new_n987), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1267), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1269), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1267), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1271), .A2(KEYINPUT126), .A3(new_n1218), .A4(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1270), .A2(new_n1273), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1274), .A2(KEYINPUT61), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1261), .A2(new_n1264), .A3(new_n1266), .A4(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT61), .ZN(new_n1277));
  NOR2_X1   g1077(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1277), .B1(new_n1278), .B2(new_n1265), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT62), .ZN(new_n1280));
  NOR3_X1   g1080(.A1(new_n1255), .A2(new_n1280), .A3(new_n1256), .ZN(new_n1281));
  AND4_X1   g1081(.A1(KEYINPUT127), .A2(new_n1237), .A3(new_n1248), .A4(new_n1281), .ZN(new_n1282));
  AOI21_X1  g1082(.A(KEYINPUT127), .B1(new_n1265), .B2(new_n1281), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1262), .A2(new_n1280), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1279), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1286));
  AND2_X1   g1086(.A1(new_n1270), .A2(new_n1273), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1276), .B1(new_n1286), .B2(new_n1287), .ZN(G405));
  NAND2_X1  g1088(.A1(G375), .A2(new_n1227), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1289), .A2(new_n1244), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1287), .A2(new_n1290), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1274), .A2(new_n1244), .A3(new_n1289), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1257), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1291), .A2(new_n1257), .A3(new_n1292), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1295), .A2(new_n1296), .ZN(G402));
endmodule


