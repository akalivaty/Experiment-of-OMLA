//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 1 1 1 0 1 1 0 1 1 0 0 0 0 1 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 1 1 0 1 1 0 0 1 1 1 0 1 1 1 0 0 0 0 1 0 0 0 0 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:39 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1195,
    new_n1196, new_n1197, new_n1198, new_n1199, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1253, new_n1254, new_n1255, new_n1256, new_n1257;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G116), .A2(G270), .ZN(new_n206));
  INV_X1    g0006(.A(G77), .ZN(new_n207));
  INV_X1    g0007(.A(G244), .ZN(new_n208));
  INV_X1    g0008(.A(G87), .ZN(new_n209));
  INV_X1    g0009(.A(G250), .ZN(new_n210));
  OAI221_X1 g0010(.A(new_n206), .B1(new_n207), .B2(new_n208), .C1(new_n209), .C2(new_n210), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G68), .A2(G238), .ZN(new_n213));
  INV_X1    g0013(.A(G226), .ZN(new_n214));
  OAI211_X1 g0014(.A(new_n212), .B(new_n213), .C1(new_n202), .C2(new_n214), .ZN(new_n215));
  AOI211_X1 g0015(.A(new_n211), .B(new_n215), .C1(G97), .C2(G257), .ZN(new_n216));
  AOI21_X1  g0016(.A(new_n216), .B1(G1), .B2(G20), .ZN(new_n217));
  XOR2_X1   g0017(.A(new_n217), .B(KEYINPUT1), .Z(new_n218));
  OR2_X1    g0018(.A1(KEYINPUT64), .A2(G20), .ZN(new_n219));
  NAND2_X1  g0019(.A1(KEYINPUT64), .A2(G20), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G13), .ZN(new_n222));
  OAI21_X1  g0022(.A(G50), .B1(G58), .B2(G68), .ZN(new_n223));
  NOR3_X1   g0023(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  INV_X1    g0024(.A(G1), .ZN(new_n225));
  INV_X1    g0025(.A(G20), .ZN(new_n226));
  NOR3_X1   g0026(.A1(new_n225), .A2(new_n226), .A3(G13), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n227), .B(G250), .C1(G257), .C2(G264), .ZN(new_n228));
  XOR2_X1   g0028(.A(new_n228), .B(KEYINPUT0), .Z(new_n229));
  NOR3_X1   g0029(.A1(new_n218), .A2(new_n224), .A3(new_n229), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT2), .B(G226), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G250), .B(G257), .Z(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XNOR2_X1  g0038(.A(G87), .B(G97), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT65), .ZN(new_n240));
  INV_X1    g0040(.A(G107), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  INV_X1    g0042(.A(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G68), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G58), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n244), .B(new_n247), .Z(G351));
  OAI21_X1  g0048(.A(new_n225), .B1(G41), .B2(G45), .ZN(new_n249));
  INV_X1    g0049(.A(G274), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  AND2_X1   g0051(.A1(G1), .A2(G13), .ZN(new_n252));
  NAND2_X1  g0052(.A1(G33), .A2(G41), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  AND2_X1   g0054(.A1(new_n254), .A2(new_n249), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n251), .B1(new_n255), .B2(G238), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n256), .B(KEYINPUT70), .ZN(new_n257));
  NAND2_X1  g0057(.A1(G33), .A2(G97), .ZN(new_n258));
  INV_X1    g0058(.A(G232), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G1698), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n260), .B1(G226), .B2(G1698), .ZN(new_n261));
  INV_X1    g0061(.A(G33), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(KEYINPUT3), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT3), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G33), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n258), .B1(new_n261), .B2(new_n266), .ZN(new_n267));
  AND2_X1   g0067(.A1(G33), .A2(G41), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT66), .ZN(new_n269));
  NOR3_X1   g0069(.A1(new_n268), .A2(new_n269), .A3(new_n222), .ZN(new_n270));
  AOI21_X1  g0070(.A(KEYINPUT66), .B1(new_n252), .B2(new_n253), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n267), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n257), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(KEYINPUT13), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT13), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n257), .A2(new_n276), .A3(new_n273), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G169), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(KEYINPUT14), .ZN(new_n280));
  INV_X1    g0080(.A(new_n278), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(G179), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT14), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n278), .A2(new_n283), .A3(G169), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n280), .A2(new_n282), .A3(new_n284), .ZN(new_n285));
  NAND3_X1  g0085(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(new_n222), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n221), .A2(G33), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n226), .A2(new_n262), .ZN(new_n289));
  OAI22_X1  g0089(.A1(new_n288), .A2(new_n207), .B1(new_n202), .B2(new_n289), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n226), .A2(G68), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n287), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT11), .ZN(new_n293));
  INV_X1    g0093(.A(G68), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n287), .B1(new_n225), .B2(G20), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  OAI22_X1  g0096(.A1(new_n292), .A2(new_n293), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  AND2_X1   g0097(.A1(new_n292), .A2(new_n293), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n291), .A2(new_n225), .A3(G13), .ZN(new_n299));
  XOR2_X1   g0099(.A(new_n299), .B(KEYINPUT12), .Z(new_n300));
  NOR3_X1   g0100(.A1(new_n297), .A2(new_n298), .A3(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n285), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G200), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n281), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(G190), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n301), .B1(new_n278), .B2(new_n306), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n303), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n203), .A2(G20), .ZN(new_n311));
  INV_X1    g0111(.A(G150), .ZN(new_n312));
  XNOR2_X1  g0112(.A(KEYINPUT8), .B(G58), .ZN(new_n313));
  OAI221_X1 g0113(.A(new_n311), .B1(new_n312), .B2(new_n289), .C1(new_n288), .C2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(G13), .ZN(new_n315));
  NOR3_X1   g0115(.A1(new_n315), .A2(new_n226), .A3(G1), .ZN(new_n316));
  AOI22_X1  g0116(.A1(new_n314), .A2(new_n287), .B1(new_n202), .B2(new_n316), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n317), .B1(new_n202), .B2(new_n296), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT9), .ZN(new_n319));
  OR2_X1    g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  XNOR2_X1  g0120(.A(KEYINPUT3), .B(G33), .ZN(new_n321));
  INV_X1    g0121(.A(G1698), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(G222), .ZN(new_n323));
  INV_X1    g0123(.A(G223), .ZN(new_n324));
  OAI211_X1 g0124(.A(new_n321), .B(new_n323), .C1(new_n324), .C2(new_n322), .ZN(new_n325));
  OAI211_X1 g0125(.A(new_n272), .B(new_n325), .C1(G77), .C2(new_n321), .ZN(new_n326));
  INV_X1    g0126(.A(new_n251), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n254), .A2(new_n249), .ZN(new_n328));
  OAI211_X1 g0128(.A(new_n326), .B(new_n327), .C1(new_n214), .C2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(G200), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n318), .A2(new_n319), .ZN(new_n331));
  OR2_X1    g0131(.A1(new_n329), .A2(new_n306), .ZN(new_n332));
  NAND4_X1  g0132(.A1(new_n320), .A2(new_n330), .A3(new_n331), .A4(new_n332), .ZN(new_n333));
  XNOR2_X1  g0133(.A(new_n333), .B(KEYINPUT10), .ZN(new_n334));
  INV_X1    g0134(.A(G169), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n329), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n318), .A2(new_n336), .ZN(new_n337));
  XOR2_X1   g0137(.A(new_n337), .B(KEYINPUT67), .Z(new_n338));
  OR2_X1    g0138(.A1(new_n329), .A2(G179), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n334), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT7), .ZN(new_n342));
  AND2_X1   g0142(.A1(KEYINPUT64), .A2(G20), .ZN(new_n343));
  NOR2_X1   g0143(.A1(KEYINPUT64), .A2(G20), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n342), .B1(new_n345), .B2(new_n321), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(KEYINPUT71), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n266), .A2(KEYINPUT7), .A3(new_n226), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT71), .ZN(new_n349));
  OAI211_X1 g0149(.A(new_n349), .B(new_n342), .C1(new_n345), .C2(new_n321), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n347), .A2(new_n348), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(G68), .ZN(new_n352));
  XNOR2_X1  g0152(.A(G58), .B(G68), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(G20), .ZN(new_n354));
  INV_X1    g0154(.A(G159), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n354), .B1(new_n355), .B2(new_n289), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n352), .A2(KEYINPUT16), .A3(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT16), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT72), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n360), .B1(new_n264), .B2(G33), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT73), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n362), .B1(new_n262), .B2(KEYINPUT3), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n262), .A2(KEYINPUT72), .A3(KEYINPUT3), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n264), .A2(KEYINPUT73), .A3(G33), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n361), .A2(new_n363), .A3(new_n364), .A4(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n366), .A2(KEYINPUT7), .A3(new_n221), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n342), .B1(new_n321), .B2(G20), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n294), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n359), .B1(new_n369), .B2(new_n356), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n358), .A2(new_n287), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n214), .A2(G1698), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n324), .A2(new_n322), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n321), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(G33), .A2(G87), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n251), .B1(new_n376), .B2(new_n272), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n328), .A2(new_n259), .ZN(new_n378));
  INV_X1    g0178(.A(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(new_n304), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n381), .B1(G190), .B2(new_n380), .ZN(new_n382));
  INV_X1    g0182(.A(new_n313), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n383), .A2(new_n316), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n384), .B1(new_n296), .B2(new_n383), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n371), .A2(new_n382), .A3(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT17), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(new_n287), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n356), .B1(new_n351), .B2(G68), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n390), .B1(new_n391), .B2(KEYINPUT16), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n385), .B1(new_n392), .B2(new_n370), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n393), .A2(KEYINPUT17), .A3(new_n382), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n389), .A2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT18), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n335), .B1(new_n377), .B2(new_n379), .ZN(new_n398));
  AND2_X1   g0198(.A1(new_n377), .A2(new_n379), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n398), .B1(G179), .B2(new_n399), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n397), .B1(new_n393), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n371), .A2(new_n386), .ZN(new_n402));
  INV_X1    g0202(.A(new_n400), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n402), .A2(KEYINPUT18), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n401), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n396), .A2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(new_n316), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n407), .A2(G77), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n296), .A2(new_n207), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n345), .A2(G77), .ZN(new_n410));
  XOR2_X1   g0210(.A(KEYINPUT15), .B(G87), .Z(new_n411));
  INV_X1    g0211(.A(KEYINPUT68), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  XNOR2_X1  g0213(.A(KEYINPUT15), .B(G87), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(KEYINPUT68), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  OAI221_X1 g0216(.A(new_n410), .B1(new_n289), .B2(new_n313), .C1(new_n416), .C2(new_n288), .ZN(new_n417));
  AOI211_X1 g0217(.A(new_n408), .B(new_n409), .C1(new_n417), .C2(new_n287), .ZN(new_n418));
  NAND2_X1  g0218(.A1(G238), .A2(G1698), .ZN(new_n419));
  OAI211_X1 g0219(.A(new_n321), .B(new_n419), .C1(new_n259), .C2(G1698), .ZN(new_n420));
  OAI211_X1 g0220(.A(new_n272), .B(new_n420), .C1(G107), .C2(new_n321), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n421), .B(new_n327), .C1(new_n208), .C2(new_n328), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(new_n335), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  OAI21_X1  g0224(.A(KEYINPUT69), .B1(new_n418), .B2(new_n424), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n408), .B1(new_n417), .B2(new_n287), .ZN(new_n426));
  INV_X1    g0226(.A(new_n409), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT69), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n428), .A2(new_n429), .A3(new_n423), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n425), .B(new_n430), .C1(G179), .C2(new_n422), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n422), .A2(G200), .ZN(new_n432));
  OAI211_X1 g0232(.A(new_n418), .B(new_n432), .C1(new_n306), .C2(new_n422), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  NOR4_X1   g0234(.A1(new_n310), .A2(new_n341), .A3(new_n406), .A4(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT23), .ZN(new_n436));
  NOR3_X1   g0236(.A1(new_n436), .A2(new_n226), .A3(G107), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n219), .A2(new_n241), .A3(new_n220), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n437), .B1(new_n438), .B2(new_n436), .ZN(new_n439));
  OAI211_X1 g0239(.A(new_n263), .B(new_n265), .C1(new_n343), .C2(new_n344), .ZN(new_n440));
  OAI21_X1  g0240(.A(KEYINPUT22), .B1(new_n440), .B2(new_n209), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT22), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n221), .A2(new_n321), .A3(new_n442), .A4(G87), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n439), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT24), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n262), .A2(new_n243), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(new_n226), .ZN(new_n447));
  XNOR2_X1  g0247(.A(new_n447), .B(KEYINPUT84), .ZN(new_n448));
  AND3_X1   g0248(.A1(new_n444), .A2(new_n445), .A3(new_n448), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n445), .B1(new_n444), .B2(new_n448), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n287), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(G41), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n452), .A2(KEYINPUT5), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n225), .A2(G45), .ZN(new_n454));
  OAI21_X1  g0254(.A(KEYINPUT76), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n452), .A2(KEYINPUT5), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT5), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(G41), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT76), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n458), .A2(new_n459), .A3(new_n225), .A4(G45), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n455), .A2(new_n456), .A3(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n461), .A2(G264), .A3(new_n254), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n210), .A2(new_n322), .ZN(new_n463));
  INV_X1    g0263(.A(G257), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(G1698), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n263), .A2(new_n463), .A3(new_n265), .A4(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(G33), .A2(G294), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(new_n272), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n462), .A2(new_n469), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n455), .A2(new_n460), .A3(G274), .A4(new_n456), .ZN(new_n471));
  INV_X1    g0271(.A(new_n254), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n304), .B1(new_n470), .B2(new_n473), .ZN(new_n474));
  OR2_X1    g0274(.A1(new_n471), .A2(new_n472), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n475), .A2(new_n306), .A3(new_n469), .A4(new_n462), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n316), .A2(KEYINPUT25), .A3(new_n241), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(KEYINPUT25), .B1(new_n316), .B2(new_n241), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n225), .A2(G33), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n407), .A2(new_n390), .A3(new_n481), .ZN(new_n482));
  OAI22_X1  g0282(.A1(new_n479), .A2(new_n480), .B1(new_n482), .B2(new_n241), .ZN(new_n483));
  INV_X1    g0283(.A(new_n483), .ZN(new_n484));
  AND3_X1   g0284(.A1(new_n451), .A2(new_n477), .A3(new_n484), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n335), .B1(new_n470), .B2(new_n473), .ZN(new_n486));
  INV_X1    g0286(.A(G179), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n475), .A2(new_n487), .A3(new_n469), .A4(new_n462), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n489), .B1(new_n451), .B2(new_n484), .ZN(new_n490));
  OAI21_X1  g0290(.A(KEYINPUT85), .B1(new_n485), .B2(new_n490), .ZN(new_n491));
  AND2_X1   g0291(.A1(new_n486), .A2(new_n488), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n441), .A2(new_n443), .ZN(new_n493));
  INV_X1    g0293(.A(new_n439), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n493), .A2(new_n448), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(KEYINPUT24), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n444), .A2(new_n445), .A3(new_n448), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n390), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n492), .B1(new_n498), .B2(new_n483), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT85), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n451), .A2(new_n477), .A3(new_n484), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n499), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n491), .A2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT82), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT81), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT78), .ZN(new_n506));
  INV_X1    g0306(.A(G45), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n506), .B(G250), .C1(new_n507), .C2(G1), .ZN(new_n508));
  AOI21_X1  g0308(.A(G274), .B1(KEYINPUT78), .B2(G250), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n508), .B1(new_n454), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(new_n254), .ZN(new_n511));
  NOR2_X1   g0311(.A1(G238), .A2(G1698), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n512), .B1(new_n208), .B2(G1698), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n446), .B1(new_n513), .B2(new_n321), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n269), .B1(new_n268), .B2(new_n222), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n252), .A2(KEYINPUT66), .A3(new_n253), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n511), .B1(new_n514), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(KEYINPUT79), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT79), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n511), .B(new_n520), .C1(new_n514), .C2(new_n517), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n505), .B1(new_n522), .B2(G190), .ZN(new_n523));
  AOI211_X1 g0323(.A(KEYINPUT81), .B(new_n306), .C1(new_n519), .C2(new_n521), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n504), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(new_n521), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n208), .A2(G1698), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n527), .B1(G238), .B2(G1698), .ZN(new_n528));
  OAI22_X1  g0328(.A1(new_n528), .A2(new_n266), .B1(new_n262), .B2(new_n243), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(new_n272), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n520), .B1(new_n530), .B2(new_n511), .ZN(new_n531));
  OAI21_X1  g0331(.A(G190), .B1(new_n526), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(KEYINPUT81), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n522), .A2(new_n505), .A3(G190), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n533), .A2(KEYINPUT82), .A3(new_n534), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n407), .B1(new_n413), .B2(new_n415), .ZN(new_n536));
  XNOR2_X1  g0336(.A(KEYINPUT80), .B(KEYINPUT19), .ZN(new_n537));
  INV_X1    g0337(.A(G97), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n537), .B1(new_n288), .B2(new_n538), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n221), .B1(new_n537), .B2(new_n258), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n209), .A2(new_n538), .A3(new_n241), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n539), .B(new_n542), .C1(new_n294), .C2(new_n440), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n536), .B1(new_n543), .B2(new_n287), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n544), .B1(new_n209), .B2(new_n482), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n522), .A2(new_n304), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n525), .A2(new_n535), .A3(new_n547), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n263), .A2(new_n265), .A3(G244), .A4(new_n322), .ZN(new_n549));
  XOR2_X1   g0349(.A(KEYINPUT75), .B(KEYINPUT4), .Z(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n210), .A2(new_n322), .ZN(new_n552));
  AOI22_X1  g0352(.A1(new_n321), .A2(new_n552), .B1(G33), .B2(G283), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT4), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(KEYINPUT75), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n321), .A2(G244), .A3(new_n322), .A4(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n551), .A2(new_n553), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(new_n272), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n461), .A2(G257), .A3(new_n254), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n558), .A2(new_n475), .A3(new_n559), .ZN(new_n560));
  AND2_X1   g0360(.A1(new_n560), .A2(G200), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n560), .A2(KEYINPUT77), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT77), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n558), .A2(new_n475), .A3(new_n563), .A4(new_n559), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n561), .B1(new_n565), .B2(G190), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n241), .B1(new_n367), .B2(new_n368), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT6), .ZN(new_n568));
  NOR3_X1   g0368(.A1(new_n568), .A2(new_n538), .A3(G107), .ZN(new_n569));
  XNOR2_X1  g0369(.A(G97), .B(G107), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n569), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  OAI22_X1  g0371(.A1(new_n571), .A2(new_n221), .B1(new_n207), .B2(new_n289), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n287), .B1(new_n567), .B2(new_n572), .ZN(new_n573));
  MUX2_X1   g0373(.A(new_n407), .B(new_n482), .S(G97), .Z(new_n574));
  NAND2_X1  g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(KEYINPUT74), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT74), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n573), .A2(new_n577), .A3(new_n574), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n566), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n562), .A2(new_n335), .A3(new_n564), .ZN(new_n581));
  OR2_X1    g0381(.A1(new_n560), .A2(G179), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n581), .A2(new_n582), .A3(new_n575), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n544), .B1(new_n416), .B2(new_n482), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n522), .A2(new_n487), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n584), .B(new_n585), .C1(G169), .C2(new_n522), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n548), .A2(new_n580), .A3(new_n583), .A4(new_n586), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n503), .B1(new_n587), .B2(KEYINPUT83), .ZN(new_n588));
  INV_X1    g0388(.A(new_n583), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n589), .B1(new_n579), .B2(new_n566), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT83), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n590), .A2(new_n591), .A3(new_n586), .A4(new_n548), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT21), .ZN(new_n593));
  AND3_X1   g0393(.A1(new_n461), .A2(G270), .A3(new_n254), .ZN(new_n594));
  INV_X1    g0394(.A(G303), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n264), .A2(G33), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n262), .A2(KEYINPUT3), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n595), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n322), .A2(G257), .ZN(new_n599));
  NAND2_X1  g0399(.A1(G264), .A2(G1698), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n263), .A2(new_n265), .A3(new_n599), .A4(new_n600), .ZN(new_n601));
  AND4_X1   g0401(.A1(new_n515), .A2(new_n598), .A3(new_n516), .A4(new_n601), .ZN(new_n602));
  NOR3_X1   g0402(.A1(new_n594), .A2(new_n473), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n316), .A2(new_n243), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n407), .A2(G116), .A3(new_n390), .A4(new_n481), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n262), .A2(G97), .ZN(new_n606));
  NAND2_X1  g0406(.A1(G33), .A2(G283), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n606), .B(new_n607), .C1(new_n343), .C2(new_n344), .ZN(new_n608));
  AOI22_X1  g0408(.A1(new_n286), .A2(new_n222), .B1(G20), .B2(new_n243), .ZN(new_n609));
  AND3_X1   g0409(.A1(new_n608), .A2(KEYINPUT20), .A3(new_n609), .ZN(new_n610));
  AOI21_X1  g0410(.A(KEYINPUT20), .B1(new_n608), .B2(new_n609), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n604), .B(new_n605), .C1(new_n610), .C2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(G169), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n593), .B1(new_n603), .B2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(new_n602), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n461), .A2(G270), .A3(new_n254), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n475), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n617), .A2(KEYINPUT21), .A3(G169), .A4(new_n612), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n603), .A2(G179), .A3(new_n612), .ZN(new_n619));
  AND3_X1   g0419(.A1(new_n614), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n617), .A2(G200), .ZN(new_n621));
  INV_X1    g0421(.A(new_n612), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n621), .B(new_n622), .C1(new_n306), .C2(new_n617), .ZN(new_n623));
  AND2_X1   g0423(.A1(new_n620), .A2(new_n623), .ZN(new_n624));
  AND4_X1   g0424(.A1(new_n435), .A2(new_n588), .A3(new_n592), .A4(new_n624), .ZN(G372));
  NAND2_X1  g0425(.A1(new_n303), .A2(new_n431), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n626), .A2(new_n309), .A3(new_n396), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(new_n405), .ZN(new_n628));
  AOI22_X1  g0428(.A1(new_n628), .A2(new_n334), .B1(new_n339), .B2(new_n338), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n548), .A2(new_n589), .A3(new_n586), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(KEYINPUT26), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n498), .A2(new_n483), .ZN(new_n632));
  AOI22_X1  g0432(.A1(new_n620), .A2(new_n499), .B1(new_n632), .B2(new_n477), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n545), .B1(new_n533), .B2(new_n534), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n518), .A2(G200), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n633), .A2(new_n583), .A3(new_n580), .A4(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT26), .ZN(new_n638));
  AND4_X1   g0438(.A1(new_n581), .A2(new_n576), .A3(new_n582), .A4(new_n578), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n636), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n518), .A2(new_n335), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n584), .A2(new_n585), .A3(new_n641), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n631), .A2(new_n637), .A3(new_n640), .A4(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n435), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n629), .A2(new_n644), .ZN(G369));
  INV_X1    g0445(.A(new_n503), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n221), .A2(new_n225), .A3(G13), .ZN(new_n647));
  OAI21_X1  g0447(.A(KEYINPUT86), .B1(new_n647), .B2(KEYINPUT27), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n345), .A2(new_n315), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT86), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT27), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n649), .A2(new_n650), .A3(new_n651), .A4(new_n225), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n648), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n647), .A2(KEYINPUT27), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n653), .A2(G213), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(KEYINPUT87), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT87), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n653), .A2(new_n657), .A3(G213), .A4(new_n654), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(G343), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n646), .B1(new_n632), .B2(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n662), .B1(new_n499), .B2(new_n661), .ZN(new_n663));
  INV_X1    g0463(.A(G343), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n659), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(new_n612), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n624), .A2(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n667), .B1(new_n620), .B2(new_n666), .ZN(new_n668));
  AND2_X1   g0468(.A1(new_n668), .A2(G330), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n663), .A2(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n499), .B1(new_n503), .B2(new_n620), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(new_n661), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n670), .A2(new_n672), .ZN(G399));
  INV_X1    g0473(.A(new_n227), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n674), .A2(G41), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n541), .A2(G116), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n676), .A2(G1), .A3(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n678), .B1(new_n223), .B2(new_n676), .ZN(new_n679));
  XNOR2_X1  g0479(.A(new_n679), .B(KEYINPUT28), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n643), .A2(new_n661), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT29), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(KEYINPUT88), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n636), .A2(new_n639), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(KEYINPUT26), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n686), .B1(KEYINPUT26), .B2(new_n630), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n637), .A2(new_n642), .ZN(new_n688));
  OAI211_X1 g0488(.A(KEYINPUT29), .B(new_n661), .C1(new_n687), .C2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT88), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n681), .A2(new_n690), .A3(new_n682), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n684), .A2(new_n689), .A3(new_n691), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n588), .A2(new_n592), .A3(new_n624), .A4(new_n661), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n617), .A2(new_n487), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n470), .B1(new_n519), .B2(new_n521), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n565), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT30), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n603), .A2(G179), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n475), .A2(new_n469), .A3(new_n462), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n699), .A2(new_n560), .A3(new_n518), .A4(new_n700), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n565), .A2(KEYINPUT30), .A3(new_n695), .A4(new_n694), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n698), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  AND3_X1   g0503(.A1(new_n703), .A2(KEYINPUT31), .A3(new_n665), .ZN(new_n704));
  AOI21_X1  g0504(.A(KEYINPUT31), .B1(new_n703), .B2(new_n665), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n693), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(G330), .ZN(new_n708));
  AND2_X1   g0508(.A1(new_n692), .A2(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n680), .B1(new_n709), .B2(G1), .ZN(G364));
  XOR2_X1   g0510(.A(new_n669), .B(KEYINPUT89), .Z(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n649), .A2(G45), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NOR3_X1   g0514(.A1(new_n714), .A2(new_n225), .A3(new_n675), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  OAI211_X1 g0516(.A(new_n712), .B(new_n716), .C1(G330), .C2(new_n668), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n222), .B1(G20), .B2(new_n335), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n304), .A2(G179), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n720), .A2(G20), .A3(G190), .ZN(new_n721));
  OR2_X1    g0521(.A1(new_n721), .A2(KEYINPUT95), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(KEYINPUT95), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n724), .A2(new_n209), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n345), .A2(new_n306), .A3(new_n720), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n221), .A2(new_n487), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(G190), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n728), .A2(new_n304), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  OAI221_X1 g0530(.A(new_n321), .B1(new_n241), .B2(new_n726), .C1(new_n730), .C2(new_n202), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n487), .A2(new_n304), .ZN(new_n732));
  XNOR2_X1  g0532(.A(new_n732), .B(KEYINPUT93), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n733), .A2(new_n306), .A3(new_n345), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  XOR2_X1   g0535(.A(KEYINPUT94), .B(KEYINPUT32), .Z(new_n736));
  NAND3_X1  g0536(.A1(new_n735), .A2(G159), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n727), .A2(new_n306), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n738), .A2(new_n304), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n737), .B1(new_n294), .B2(new_n740), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n736), .B1(new_n735), .B2(G159), .ZN(new_n742));
  OR4_X1    g0542(.A1(new_n725), .A2(new_n731), .A3(new_n741), .A4(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT92), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n728), .A2(G200), .ZN(new_n745));
  XNOR2_X1  g0545(.A(new_n745), .B(KEYINPUT91), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n738), .A2(G200), .ZN(new_n747));
  AOI22_X1  g0547(.A1(new_n746), .A2(G58), .B1(G77), .B2(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n743), .B1(new_n744), .B2(new_n748), .ZN(new_n749));
  AND2_X1   g0549(.A1(new_n733), .A2(G190), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(new_n221), .ZN(new_n751));
  OAI221_X1 g0551(.A(new_n749), .B1(new_n744), .B2(new_n748), .C1(new_n538), .C2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(G283), .ZN(new_n753));
  INV_X1    g0553(.A(G329), .ZN(new_n754));
  OAI221_X1 g0554(.A(new_n266), .B1(new_n753), .B2(new_n726), .C1(new_n734), .C2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(G317), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n739), .B1(KEYINPUT33), .B2(new_n756), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n757), .B1(KEYINPUT33), .B2(new_n756), .ZN(new_n758));
  AOI211_X1 g0558(.A(new_n755), .B(new_n758), .C1(G322), .C2(new_n746), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n729), .A2(G326), .ZN(new_n760));
  INV_X1    g0560(.A(new_n747), .ZN(new_n761));
  INV_X1    g0561(.A(G311), .ZN(new_n762));
  INV_X1    g0562(.A(G294), .ZN(new_n763));
  OAI221_X1 g0563(.A(new_n760), .B1(new_n761), .B2(new_n762), .C1(new_n763), .C2(new_n751), .ZN(new_n764));
  INV_X1    g0564(.A(KEYINPUT96), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  AND2_X1   g0566(.A1(new_n759), .A2(new_n766), .ZN(new_n767));
  OAI221_X1 g0567(.A(new_n767), .B1(new_n765), .B2(new_n764), .C1(new_n595), .C2(new_n724), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n719), .B1(new_n752), .B2(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(G13), .A2(G33), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(G20), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(new_n718), .ZN(new_n773));
  XOR2_X1   g0573(.A(new_n773), .B(KEYINPUT90), .Z(new_n774));
  NAND2_X1  g0574(.A1(new_n247), .A2(G45), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n674), .A2(new_n321), .ZN(new_n776));
  OAI211_X1 g0576(.A(new_n775), .B(new_n776), .C1(G45), .C2(new_n223), .ZN(new_n777));
  INV_X1    g0577(.A(G355), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n321), .A2(new_n227), .ZN(new_n779));
  OAI221_X1 g0579(.A(new_n777), .B1(G116), .B2(new_n227), .C1(new_n778), .C2(new_n779), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n769), .B1(new_n774), .B2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n772), .ZN(new_n782));
  OAI211_X1 g0582(.A(new_n781), .B(new_n715), .C1(new_n668), .C2(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n717), .A2(new_n783), .ZN(G396));
  NOR2_X1   g0584(.A1(new_n661), .A2(new_n418), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n785), .B1(new_n431), .B2(new_n433), .ZN(new_n786));
  AND2_X1   g0586(.A1(new_n431), .A2(new_n785), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n643), .A2(new_n661), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(KEYINPUT98), .ZN(new_n790));
  INV_X1    g0590(.A(new_n788), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n681), .A2(new_n791), .ZN(new_n792));
  XNOR2_X1  g0592(.A(new_n790), .B(new_n792), .ZN(new_n793));
  AND2_X1   g0593(.A1(new_n793), .A2(new_n708), .ZN(new_n794));
  OR2_X1    g0594(.A1(new_n794), .A2(KEYINPUT99), .ZN(new_n795));
  OR2_X1    g0595(.A1(new_n793), .A2(new_n708), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n794), .A2(KEYINPUT99), .ZN(new_n797));
  NAND4_X1  g0597(.A1(new_n795), .A2(new_n796), .A3(new_n716), .A4(new_n797), .ZN(new_n798));
  AND2_X1   g0598(.A1(new_n729), .A2(G137), .ZN(new_n799));
  OAI22_X1  g0599(.A1(new_n312), .A2(new_n740), .B1(new_n761), .B2(new_n355), .ZN(new_n800));
  AOI211_X1 g0600(.A(new_n799), .B(new_n800), .C1(G143), .C2(new_n746), .ZN(new_n801));
  XOR2_X1   g0601(.A(new_n801), .B(KEYINPUT34), .Z(new_n802));
  AOI21_X1  g0602(.A(new_n266), .B1(new_n735), .B2(G132), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n803), .B1(new_n202), .B2(new_n724), .ZN(new_n804));
  INV_X1    g0604(.A(new_n751), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n804), .B1(G58), .B2(new_n805), .ZN(new_n806));
  OAI211_X1 g0606(.A(new_n802), .B(new_n806), .C1(new_n294), .C2(new_n726), .ZN(new_n807));
  OAI22_X1  g0607(.A1(new_n730), .A2(new_n595), .B1(new_n209), .B2(new_n726), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n808), .B1(new_n746), .B2(G294), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n321), .B1(new_n735), .B2(G311), .ZN(new_n810));
  AOI22_X1  g0610(.A1(new_n805), .A2(G97), .B1(G116), .B2(new_n747), .ZN(new_n811));
  AND3_X1   g0611(.A1(new_n809), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  OR2_X1    g0612(.A1(new_n740), .A2(KEYINPUT97), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n740), .A2(KEYINPUT97), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  OAI221_X1 g0615(.A(new_n812), .B1(new_n241), .B2(new_n724), .C1(new_n753), .C2(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n719), .B1(new_n807), .B2(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n718), .A2(new_n770), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n817), .B1(new_n207), .B2(new_n818), .ZN(new_n819));
  OAI211_X1 g0619(.A(new_n819), .B(new_n715), .C1(new_n771), .C2(new_n788), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n798), .A2(new_n820), .ZN(G384));
  NOR2_X1   g0621(.A1(new_n431), .A2(new_n665), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n789), .A2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(KEYINPUT38), .ZN(new_n825));
  OR2_X1    g0625(.A1(new_n391), .A2(KEYINPUT16), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n826), .A2(new_n392), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n659), .B1(new_n827), .B2(new_n386), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n829), .B1(new_n396), .B2(new_n405), .ZN(new_n830));
  AOI22_X1  g0630(.A1(new_n827), .A2(new_n386), .B1(new_n400), .B2(new_n659), .ZN(new_n831));
  INV_X1    g0631(.A(new_n387), .ZN(new_n832));
  OAI21_X1  g0632(.A(KEYINPUT37), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  AOI22_X1  g0633(.A1(new_n371), .A2(new_n386), .B1(new_n659), .B2(new_n400), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT37), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n835), .A2(new_n836), .A3(new_n387), .ZN(new_n837));
  AND2_X1   g0637(.A1(new_n833), .A2(new_n837), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n825), .B1(new_n830), .B2(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(KEYINPUT18), .B1(new_n402), .B2(new_n403), .ZN(new_n840));
  AOI211_X1 g0640(.A(new_n397), .B(new_n400), .C1(new_n371), .C2(new_n386), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n828), .B1(new_n842), .B2(new_n395), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n833), .A2(new_n837), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n843), .A2(KEYINPUT38), .A3(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n839), .A2(new_n845), .ZN(new_n846));
  OAI211_X1 g0646(.A(new_n303), .B(new_n309), .C1(new_n301), .C2(new_n661), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n302), .B(new_n665), .C1(new_n285), .C2(new_n308), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  AND3_X1   g0649(.A1(new_n824), .A2(new_n846), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n402), .A2(new_n660), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n851), .B1(new_n396), .B2(new_n405), .ZN(new_n852));
  OAI21_X1  g0652(.A(KEYINPUT37), .B1(new_n832), .B2(new_n834), .ZN(new_n853));
  AND2_X1   g0653(.A1(new_n837), .A2(new_n853), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n825), .B1(new_n852), .B2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT39), .ZN(new_n856));
  AND3_X1   g0656(.A1(new_n855), .A2(new_n856), .A3(new_n845), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n856), .B1(new_n839), .B2(new_n845), .ZN(new_n858));
  OAI21_X1  g0658(.A(KEYINPUT101), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  AND3_X1   g0659(.A1(new_n843), .A2(KEYINPUT38), .A3(new_n844), .ZN(new_n860));
  AOI21_X1  g0660(.A(KEYINPUT38), .B1(new_n843), .B2(new_n844), .ZN(new_n861));
  OAI21_X1  g0661(.A(KEYINPUT39), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT101), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n859), .A2(new_n864), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n303), .A2(new_n665), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n850), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n842), .A2(new_n659), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND4_X1  g0669(.A1(new_n684), .A2(new_n435), .A3(new_n689), .A4(new_n691), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(new_n629), .ZN(new_n871));
  XOR2_X1   g0671(.A(new_n869), .B(new_n871), .Z(new_n872));
  AOI21_X1  g0672(.A(new_n791), .B1(new_n693), .B2(new_n706), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n873), .A2(new_n846), .A3(new_n849), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT40), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n855), .A2(new_n845), .ZN(new_n877));
  NAND4_X1  g0677(.A1(new_n873), .A2(KEYINPUT40), .A3(new_n877), .A4(new_n849), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n435), .A2(new_n707), .ZN(new_n880));
  XOR2_X1   g0680(.A(new_n879), .B(new_n880), .Z(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(G330), .ZN(new_n882));
  XNOR2_X1  g0682(.A(new_n872), .B(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n883), .B1(new_n225), .B2(new_n649), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT35), .ZN(new_n885));
  AOI211_X1 g0685(.A(new_n222), .B(new_n221), .C1(new_n571), .C2(new_n885), .ZN(new_n886));
  OAI211_X1 g0686(.A(new_n886), .B(G116), .C1(new_n885), .C2(new_n571), .ZN(new_n887));
  XNOR2_X1  g0687(.A(new_n887), .B(KEYINPUT36), .ZN(new_n888));
  INV_X1    g0688(.A(G58), .ZN(new_n889));
  OAI21_X1  g0689(.A(G77), .B1(new_n889), .B2(new_n294), .ZN(new_n890));
  OAI22_X1  g0690(.A1(new_n890), .A2(new_n223), .B1(G50), .B2(new_n294), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n891), .A2(G1), .A3(new_n315), .ZN(new_n892));
  XOR2_X1   g0692(.A(new_n892), .B(KEYINPUT100), .Z(new_n893));
  NAND3_X1  g0693(.A1(new_n884), .A2(new_n888), .A3(new_n893), .ZN(G367));
  OAI22_X1  g0694(.A1(new_n751), .A2(new_n294), .B1(new_n761), .B2(new_n202), .ZN(new_n895));
  AOI211_X1 g0695(.A(new_n266), .B(new_n895), .C1(G137), .C2(new_n735), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n729), .A2(G143), .ZN(new_n897));
  INV_X1    g0697(.A(new_n815), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(G159), .ZN(new_n899));
  OAI22_X1  g0699(.A1(new_n724), .A2(new_n889), .B1(new_n207), .B2(new_n726), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n900), .B1(new_n746), .B2(G150), .ZN(new_n901));
  NAND4_X1  g0701(.A1(new_n896), .A2(new_n897), .A3(new_n899), .A4(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n266), .B1(new_n730), .B2(new_n762), .ZN(new_n903));
  OAI22_X1  g0703(.A1(new_n751), .A2(new_n241), .B1(new_n761), .B2(new_n753), .ZN(new_n904));
  AOI211_X1 g0704(.A(new_n903), .B(new_n904), .C1(G317), .C2(new_n735), .ZN(new_n905));
  INV_X1    g0705(.A(new_n724), .ZN(new_n906));
  AOI21_X1  g0706(.A(KEYINPUT46), .B1(new_n906), .B2(G116), .ZN(new_n907));
  XOR2_X1   g0707(.A(new_n907), .B(KEYINPUT109), .Z(new_n908));
  NAND2_X1  g0708(.A1(new_n905), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n909), .B1(G294), .B2(new_n898), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n906), .A2(KEYINPUT46), .A3(G116), .ZN(new_n911));
  AOI22_X1  g0711(.A1(new_n746), .A2(G303), .B1(KEYINPUT108), .B2(new_n911), .ZN(new_n912));
  OAI211_X1 g0712(.A(new_n910), .B(new_n912), .C1(KEYINPUT108), .C2(new_n911), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n726), .A2(new_n538), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n902), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n915), .B(KEYINPUT110), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n916), .B(KEYINPUT47), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n716), .B1(new_n917), .B2(new_n718), .ZN(new_n918));
  INV_X1    g0718(.A(new_n776), .ZN(new_n919));
  OAI221_X1 g0719(.A(new_n773), .B1(new_n416), .B2(new_n227), .C1(new_n237), .C2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n665), .A2(new_n545), .ZN(new_n921));
  XOR2_X1   g0721(.A(new_n921), .B(KEYINPUT102), .Z(new_n922));
  INV_X1    g0722(.A(new_n636), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  MUX2_X1   g0724(.A(new_n922), .B(new_n924), .S(new_n642), .Z(new_n925));
  INV_X1    g0725(.A(KEYINPUT103), .ZN(new_n926));
  OR2_X1    g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n925), .A2(new_n926), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n927), .A2(new_n772), .A3(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n918), .A2(new_n920), .A3(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT43), .ZN(new_n931));
  AND3_X1   g0731(.A1(new_n927), .A2(new_n931), .A3(new_n928), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n931), .B1(new_n927), .B2(new_n928), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n590), .B1(new_n579), .B2(new_n661), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n639), .A2(new_n665), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n620), .A2(new_n665), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n646), .A2(new_n939), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n941), .B(KEYINPUT42), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n589), .B1(new_n937), .B2(new_n490), .ZN(new_n943));
  XOR2_X1   g0743(.A(new_n943), .B(KEYINPUT104), .Z(new_n944));
  OAI21_X1  g0744(.A(new_n942), .B1(new_n944), .B2(new_n665), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n934), .A2(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT105), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  OAI211_X1 g0748(.A(new_n932), .B(new_n942), .C1(new_n665), .C2(new_n944), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n934), .A2(KEYINPUT105), .A3(new_n945), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n948), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n670), .A2(new_n938), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n951), .B(new_n953), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n714), .A2(new_n225), .ZN(new_n955));
  INV_X1    g0755(.A(new_n955), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n672), .A2(new_n590), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n957), .B(KEYINPUT44), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n672), .A2(new_n937), .ZN(new_n959));
  XOR2_X1   g0759(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n960));
  XNOR2_X1  g0760(.A(new_n959), .B(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n958), .A2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(new_n670), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n962), .B(new_n963), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n940), .B1(new_n663), .B2(new_n939), .ZN(new_n965));
  INV_X1    g0765(.A(new_n669), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n967), .B1(new_n712), .B2(new_n965), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n968), .A2(new_n709), .ZN(new_n969));
  OR2_X1    g0769(.A1(new_n964), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n970), .A2(new_n709), .ZN(new_n971));
  XNOR2_X1  g0771(.A(KEYINPUT106), .B(KEYINPUT41), .ZN(new_n972));
  XOR2_X1   g0772(.A(new_n675), .B(new_n972), .Z(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n956), .B1(new_n971), .B2(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n930), .B1(new_n954), .B2(new_n975), .ZN(G387));
  NOR2_X1   g0776(.A1(new_n663), .A2(new_n782), .ZN(new_n977));
  AND2_X1   g0777(.A1(new_n735), .A2(G326), .ZN(new_n978));
  AOI22_X1  g0778(.A1(new_n746), .A2(G317), .B1(G322), .B2(new_n729), .ZN(new_n979));
  OAI221_X1 g0779(.A(new_n979), .B1(new_n595), .B2(new_n761), .C1(new_n815), .C2(new_n762), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(KEYINPUT48), .ZN(new_n981));
  OAI221_X1 g0781(.A(new_n981), .B1(new_n753), .B2(new_n751), .C1(new_n763), .C2(new_n724), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT49), .ZN(new_n983));
  AOI211_X1 g0783(.A(new_n321), .B(new_n978), .C1(new_n982), .C2(new_n983), .ZN(new_n984));
  OAI221_X1 g0784(.A(new_n984), .B1(new_n983), .B2(new_n982), .C1(new_n243), .C2(new_n726), .ZN(new_n985));
  OAI22_X1  g0785(.A1(new_n294), .A2(new_n761), .B1(new_n740), .B2(new_n313), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n321), .B1(new_n751), .B2(new_n416), .ZN(new_n987));
  NOR3_X1   g0787(.A1(new_n986), .A2(new_n987), .A3(new_n914), .ZN(new_n988));
  OAI22_X1  g0788(.A1(new_n730), .A2(new_n355), .B1(new_n734), .B2(new_n312), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n989), .B1(new_n746), .B2(G50), .ZN(new_n990));
  OAI211_X1 g0790(.A(new_n988), .B(new_n990), .C1(new_n207), .C2(new_n724), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n719), .B1(new_n985), .B2(new_n991), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n313), .A2(G50), .ZN(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n507), .B1(new_n994), .B2(KEYINPUT50), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n995), .B1(G68), .B2(G77), .ZN(new_n996));
  INV_X1    g0796(.A(new_n677), .ZN(new_n997));
  AOI22_X1  g0797(.A1(new_n994), .A2(KEYINPUT50), .B1(new_n997), .B2(KEYINPUT111), .ZN(new_n998));
  OAI211_X1 g0798(.A(new_n996), .B(new_n998), .C1(KEYINPUT111), .C2(new_n997), .ZN(new_n999));
  OAI211_X1 g0799(.A(new_n999), .B(new_n776), .C1(new_n234), .C2(new_n507), .ZN(new_n1000));
  OAI221_X1 g0800(.A(new_n1000), .B1(G107), .B2(new_n227), .C1(new_n677), .C2(new_n779), .ZN(new_n1001));
  AOI211_X1 g0801(.A(new_n977), .B(new_n992), .C1(new_n774), .C2(new_n1001), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(new_n1002), .A2(new_n715), .B1(new_n956), .B2(new_n968), .ZN(new_n1003));
  OR2_X1    g0803(.A1(new_n968), .A2(new_n709), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n1004), .A2(new_n675), .A3(new_n969), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1003), .A2(new_n1005), .ZN(G393));
  AOI21_X1  g0806(.A(new_n676), .B1(new_n964), .B2(new_n969), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n970), .A2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n321), .B1(new_n726), .B2(new_n209), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(new_n746), .A2(G159), .B1(G150), .B2(new_n729), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(KEYINPUT51), .ZN(new_n1011));
  AOI211_X1 g0811(.A(new_n1009), .B(new_n1011), .C1(G143), .C2(new_n735), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n751), .A2(new_n207), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1013), .B1(new_n898), .B2(G50), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1014), .B1(new_n313), .B2(new_n761), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1015), .B(KEYINPUT112), .ZN(new_n1016));
  OAI211_X1 g0816(.A(new_n1012), .B(new_n1016), .C1(new_n294), .C2(new_n724), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n746), .A2(G311), .B1(G317), .B2(new_n729), .ZN(new_n1018));
  XOR2_X1   g0818(.A(new_n1018), .B(KEYINPUT52), .Z(new_n1019));
  OAI21_X1  g0819(.A(new_n266), .B1(new_n726), .B2(new_n241), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1020), .B1(new_n735), .B2(G322), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n1021), .B1(new_n751), .B2(new_n243), .C1(new_n763), .C2(new_n761), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1022), .B1(new_n898), .B2(G303), .ZN(new_n1023));
  OAI211_X1 g0823(.A(new_n1019), .B(new_n1023), .C1(new_n753), .C2(new_n724), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1017), .A2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n716), .B1(new_n1025), .B2(new_n718), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n773), .B1(new_n538), .B2(new_n227), .C1(new_n244), .C2(new_n919), .ZN(new_n1027));
  OAI211_X1 g0827(.A(new_n1026), .B(new_n1027), .C1(new_n782), .C2(new_n937), .ZN(new_n1028));
  OAI211_X1 g0828(.A(new_n1008), .B(new_n1028), .C1(new_n955), .C2(new_n964), .ZN(new_n1029));
  XOR2_X1   g0829(.A(new_n1029), .B(KEYINPUT113), .Z(G390));
  NAND3_X1  g0830(.A1(new_n855), .A2(new_n856), .A3(new_n845), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n863), .B1(new_n862), .B2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n866), .B1(new_n824), .B2(new_n849), .ZN(new_n1033));
  AOI21_X1  g0833(.A(KEYINPUT101), .B1(new_n846), .B2(KEYINPUT39), .ZN(new_n1034));
  NOR3_X1   g0834(.A1(new_n1032), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n866), .ZN(new_n1036));
  OAI211_X1 g0836(.A(new_n788), .B(new_n661), .C1(new_n687), .C2(new_n688), .ZN(new_n1037));
  AND2_X1   g0837(.A1(new_n1037), .A2(new_n823), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n849), .ZN(new_n1039));
  OAI211_X1 g0839(.A(new_n1036), .B(new_n877), .C1(new_n1038), .C2(new_n1039), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n1040), .ZN(new_n1041));
  OAI21_X1  g0841(.A(KEYINPUT114), .B1(new_n1035), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT114), .ZN(new_n1043));
  OAI211_X1 g0843(.A(new_n1043), .B(new_n1040), .C1(new_n865), .C2(new_n1033), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n873), .A2(G330), .A3(new_n849), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1042), .A2(new_n1044), .A3(new_n1045), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n1035), .A2(new_n1041), .ZN(new_n1047));
  AND4_X1   g0847(.A1(G330), .A2(new_n707), .A3(new_n849), .A4(new_n788), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1047), .A2(new_n1043), .A3(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1046), .A2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n435), .A2(G330), .A3(new_n707), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n870), .A2(new_n629), .A3(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT115), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NAND4_X1  g0854(.A1(new_n870), .A2(KEYINPUT115), .A3(new_n629), .A4(new_n1051), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n707), .A2(G330), .A3(new_n788), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1057), .A2(new_n1039), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1058), .A2(new_n1045), .ZN(new_n1059));
  AOI21_X1  g0859(.A(KEYINPUT116), .B1(new_n1059), .B2(new_n824), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT116), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n824), .ZN(new_n1062));
  AOI211_X1 g0862(.A(new_n1061), .B(new_n1062), .C1(new_n1058), .C2(new_n1045), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n1060), .A2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1058), .A2(new_n1038), .A3(new_n1045), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1056), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1050), .A2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n849), .B1(new_n873), .B2(G330), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n824), .B1(new_n1048), .B2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1069), .A2(new_n1061), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1059), .A2(KEYINPUT116), .A3(new_n824), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1070), .A2(new_n1071), .A3(new_n1065), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1072), .A2(new_n1054), .A3(new_n1055), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1073), .A2(new_n1046), .A3(new_n1049), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1067), .A2(new_n1074), .A3(new_n675), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n859), .A2(new_n770), .A3(new_n864), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n734), .A2(new_n763), .B1(new_n294), .B2(new_n726), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n761), .A2(new_n538), .ZN(new_n1078));
  OR4_X1    g0878(.A1(new_n321), .A2(new_n1013), .A3(new_n1078), .A4(new_n725), .ZN(new_n1079));
  AOI211_X1 g0879(.A(new_n1077), .B(new_n1079), .C1(G116), .C2(new_n746), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n1080), .B1(new_n241), .B2(new_n815), .C1(new_n753), .C2(new_n730), .ZN(new_n1081));
  INV_X1    g0881(.A(G128), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n730), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n898), .A2(G137), .ZN(new_n1084));
  XOR2_X1   g0884(.A(KEYINPUT54), .B(G143), .Z(new_n1085));
  AOI22_X1  g0885(.A1(new_n805), .A2(G159), .B1(new_n747), .B2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n906), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1087));
  INV_X1    g0887(.A(KEYINPUT53), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1088), .B1(new_n724), .B2(new_n312), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n266), .B1(new_n735), .B2(G125), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1091), .B1(new_n202), .B2(new_n726), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(G132), .B2(new_n746), .ZN(new_n1093));
  NAND4_X1  g0893(.A1(new_n1084), .A2(new_n1086), .A3(new_n1090), .A4(new_n1093), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1081), .B1(new_n1083), .B2(new_n1094), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n1095), .A2(new_n718), .B1(new_n313), .B2(new_n818), .ZN(new_n1096));
  AND3_X1   g0896(.A1(new_n1076), .A2(new_n715), .A3(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1097), .B1(new_n1050), .B2(new_n956), .ZN(new_n1098));
  AND2_X1   g0898(.A1(new_n1075), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(G378));
  OAI211_X1 g0900(.A(new_n452), .B(new_n266), .C1(new_n724), .C2(new_n207), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n416), .A2(new_n761), .B1(new_n740), .B2(new_n538), .ZN(new_n1102));
  AOI211_X1 g0902(.A(new_n1101), .B(new_n1102), .C1(G68), .C2(new_n805), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n734), .A2(new_n753), .B1(new_n889), .B2(new_n726), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1104), .B1(new_n746), .B2(G107), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n1103), .B(new_n1105), .C1(new_n243), .C2(new_n730), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(new_n1106), .B(KEYINPUT58), .ZN(new_n1107));
  AOI21_X1  g0907(.A(G41), .B1(KEYINPUT3), .B2(G33), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1107), .B1(G50), .B2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n262), .B1(new_n726), .B2(new_n355), .ZN(new_n1110));
  AOI211_X1 g0910(.A(G41), .B(new_n1110), .C1(new_n735), .C2(G124), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n746), .A2(G128), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n906), .A2(new_n1085), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n805), .A2(G150), .B1(G137), .B2(new_n747), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(G125), .A2(new_n729), .B1(new_n739), .B2(G132), .ZN(new_n1115));
  NAND4_X1  g0915(.A1(new_n1112), .A2(new_n1113), .A3(new_n1114), .A4(new_n1115), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(KEYINPUT117), .B(KEYINPUT59), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(new_n1116), .B(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1109), .B1(new_n1111), .B2(new_n1118), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(new_n1119), .B(KEYINPUT118), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n716), .B1(new_n1120), .B2(new_n718), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n818), .A2(new_n202), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(new_n341), .B(KEYINPUT55), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n660), .A2(new_n318), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(new_n1124), .B(KEYINPUT56), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(new_n1123), .B(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1127), .A2(new_n770), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1121), .A2(new_n1122), .A3(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(G330), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1127), .B1(new_n879), .B2(new_n1130), .ZN(new_n1131));
  NAND4_X1  g0931(.A1(new_n1126), .A2(new_n876), .A3(G330), .A4(new_n878), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1133), .A2(new_n869), .ZN(new_n1134));
  NAND4_X1  g0934(.A1(new_n1131), .A2(new_n868), .A3(new_n867), .A4(new_n1132), .ZN(new_n1135));
  INV_X1    g0935(.A(KEYINPUT119), .ZN(new_n1136));
  INV_X1    g0936(.A(KEYINPUT120), .ZN(new_n1137));
  AND3_X1   g0937(.A1(new_n1135), .A2(new_n1136), .A3(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1137), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1134), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1141), .A2(KEYINPUT120), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1134), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1135), .A2(new_n1136), .A3(new_n1137), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1142), .A2(new_n1143), .A3(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1140), .A2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1129), .B1(new_n1146), .B2(new_n955), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1147), .ZN(new_n1148));
  AND2_X1   g0948(.A1(new_n1140), .A2(new_n1145), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1073), .B1(new_n1046), .B2(new_n1049), .ZN(new_n1150));
  OAI21_X1  g0950(.A(KEYINPUT121), .B1(new_n1150), .B2(new_n1056), .ZN(new_n1151));
  INV_X1    g0951(.A(KEYINPUT121), .ZN(new_n1152));
  AND2_X1   g0952(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1067), .A2(new_n1152), .A3(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1151), .A2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(KEYINPUT57), .B1(new_n1149), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT57), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1157), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1152), .B1(new_n1067), .B2(new_n1153), .ZN(new_n1159));
  AOI211_X1 g0959(.A(KEYINPUT121), .B(new_n1056), .C1(new_n1050), .C2(new_n1072), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1158), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1161), .A2(new_n675), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1148), .B1(new_n1156), .B2(new_n1162), .ZN(G375));
  NOR2_X1   g0963(.A1(new_n849), .A2(new_n771), .ZN(new_n1164));
  OAI22_X1  g0964(.A1(new_n751), .A2(new_n416), .B1(new_n207), .B2(new_n726), .ZN(new_n1165));
  AOI211_X1 g0965(.A(new_n321), .B(new_n1165), .C1(G107), .C2(new_n747), .ZN(new_n1166));
  OAI22_X1  g0966(.A1(new_n724), .A2(new_n538), .B1(new_n734), .B2(new_n595), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1167), .B1(new_n746), .B2(G283), .ZN(new_n1168));
  AND2_X1   g0968(.A1(new_n1166), .A2(new_n1168), .ZN(new_n1169));
  OAI221_X1 g0969(.A(new_n1169), .B1(new_n243), .B2(new_n815), .C1(new_n763), .C2(new_n730), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n761), .A2(new_n312), .B1(new_n889), .B2(new_n726), .ZN(new_n1171));
  AOI211_X1 g0971(.A(new_n266), .B(new_n1171), .C1(G50), .C2(new_n805), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n898), .A2(new_n1085), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n729), .A2(G132), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n724), .A2(new_n355), .B1(new_n734), .B2(new_n1082), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1175), .B1(new_n746), .B2(G137), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n1172), .A2(new_n1173), .A3(new_n1174), .A4(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n719), .B1(new_n1170), .B2(new_n1177), .ZN(new_n1178));
  NOR3_X1   g0978(.A1(new_n718), .A2(G68), .A3(new_n770), .ZN(new_n1179));
  NOR4_X1   g0979(.A1(new_n1164), .A2(new_n716), .A3(new_n1178), .A4(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1180), .B1(new_n1072), .B2(new_n956), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1073), .A2(new_n974), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n1153), .A2(new_n1072), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1181), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  XOR2_X1   g0984(.A(new_n1184), .B(KEYINPUT122), .Z(G381));
  AOI21_X1  g0985(.A(new_n676), .B1(new_n1155), .B2(new_n1158), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1157), .B1(new_n1187), .B2(new_n1146), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1147), .B1(new_n1186), .B2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1189), .A2(new_n1099), .ZN(new_n1190));
  OR3_X1    g0990(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(new_n1029), .B(KEYINPUT113), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n1192), .B(new_n930), .C1(new_n975), .C2(new_n954), .ZN(new_n1193));
  OR4_X1    g0993(.A1(G381), .A2(new_n1190), .A3(new_n1191), .A4(new_n1193), .ZN(G407));
  NAND2_X1  g0994(.A1(new_n664), .A2(G213), .ZN(new_n1195));
  XOR2_X1   g0995(.A(new_n1195), .B(KEYINPUT123), .Z(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n1190), .A2(new_n1197), .ZN(new_n1198));
  XOR2_X1   g0998(.A(new_n1198), .B(KEYINPUT124), .Z(new_n1199));
  NAND3_X1  g0999(.A1(new_n1199), .A2(G213), .A3(G407), .ZN(G409));
  NAND2_X1  g1000(.A1(new_n1196), .A2(G2897), .ZN(new_n1201));
  INV_X1    g1001(.A(KEYINPUT60), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1202), .B1(new_n1153), .B2(new_n1072), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1064), .A2(new_n1056), .A3(KEYINPUT60), .A4(new_n1065), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n1203), .A2(new_n675), .A3(new_n1204), .A4(new_n1073), .ZN(new_n1205));
  AND3_X1   g1005(.A1(new_n1205), .A2(G384), .A3(new_n1181), .ZN(new_n1206));
  AOI21_X1  g1006(.A(G384), .B1(new_n1205), .B2(new_n1181), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT125), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1201), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  OAI21_X1  g1010(.A(KEYINPUT125), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1205), .A2(new_n1181), .ZN(new_n1212));
  INV_X1    g1012(.A(G384), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1205), .A2(G384), .A3(new_n1181), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1214), .A2(new_n1209), .A3(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1211), .A2(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1210), .B1(new_n1201), .B2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1186), .A2(new_n1188), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1099), .B1(new_n1219), .B2(new_n1148), .ZN(new_n1220));
  AND3_X1   g1020(.A1(new_n1075), .A2(new_n1098), .A3(new_n1129), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1222), .A2(new_n956), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n1145), .B(new_n1140), .C1(new_n1159), .C2(new_n1160), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n1221), .B(new_n1223), .C1(new_n1224), .C2(new_n973), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1225), .A2(new_n1197), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1218), .B1(new_n1220), .B2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1227), .A2(KEYINPUT63), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(G375), .A2(G378), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1226), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1229), .A2(new_n1230), .A3(new_n1208), .ZN(new_n1231));
  AOI21_X1  g1031(.A(KEYINPUT61), .B1(new_n1228), .B2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(G390), .A2(G387), .ZN(new_n1233));
  XNOR2_X1  g1033(.A(G393), .B(G396), .ZN(new_n1234));
  AND3_X1   g1034(.A1(new_n1193), .A2(new_n1233), .A3(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1234), .B1(new_n1193), .B2(new_n1233), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1229), .A2(KEYINPUT63), .A3(new_n1230), .A4(new_n1208), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1232), .A2(new_n1237), .A3(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT62), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1240), .A2(KEYINPUT127), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1231), .A2(new_n1241), .ZN(new_n1242));
  XNOR2_X1  g1042(.A(KEYINPUT127), .B(KEYINPUT62), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1229), .A2(new_n1230), .A3(new_n1208), .A4(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1242), .A2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT126), .ZN(new_n1246));
  OAI211_X1 g1046(.A(new_n1197), .B(new_n1225), .C1(new_n1189), .C2(new_n1099), .ZN(new_n1247));
  AOI211_X1 g1047(.A(new_n1246), .B(KEYINPUT61), .C1(new_n1247), .C2(new_n1218), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT61), .ZN(new_n1249));
  AOI21_X1  g1049(.A(KEYINPUT126), .B1(new_n1227), .B2(new_n1249), .ZN(new_n1250));
  NOR3_X1   g1050(.A1(new_n1245), .A2(new_n1248), .A3(new_n1250), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1239), .B1(new_n1251), .B2(new_n1237), .ZN(G405));
  NAND2_X1  g1052(.A1(new_n1229), .A2(new_n1190), .ZN(new_n1253));
  OR2_X1    g1053(.A1(new_n1237), .A2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1237), .A2(new_n1253), .ZN(new_n1255));
  AND3_X1   g1055(.A1(new_n1254), .A2(new_n1208), .A3(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1208), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1256), .A2(new_n1257), .ZN(G402));
endmodule


