

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596;

  XNOR2_X1 U326 ( .A(n314), .B(n313), .ZN(n463) );
  NOR2_X1 U327 ( .A1(n401), .A2(n400), .ZN(n492) );
  XNOR2_X1 U328 ( .A(n458), .B(n457), .ZN(n508) );
  XOR2_X1 U329 ( .A(n416), .B(n322), .Z(n294) );
  INV_X1 U330 ( .A(KEYINPUT96), .ZN(n390) );
  XNOR2_X1 U331 ( .A(n301), .B(KEYINPUT79), .ZN(n302) );
  XNOR2_X1 U332 ( .A(n303), .B(n302), .ZN(n307) );
  INV_X1 U333 ( .A(G176GAT), .ZN(n326) );
  XNOR2_X1 U334 ( .A(n482), .B(KEYINPUT55), .ZN(n483) );
  XNOR2_X1 U335 ( .A(n312), .B(n311), .ZN(n313) );
  XNOR2_X1 U336 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U337 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U338 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U339 ( .A(n481), .B(KEYINPUT28), .Z(n543) );
  XNOR2_X1 U340 ( .A(n486), .B(KEYINPUT58), .ZN(n487) );
  XNOR2_X1 U341 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n459) );
  XNOR2_X1 U342 ( .A(n488), .B(n487), .ZN(G1351GAT) );
  XNOR2_X1 U343 ( .A(n460), .B(n459), .ZN(G1330GAT) );
  XNOR2_X1 U344 ( .A(KEYINPUT38), .B(KEYINPUT103), .ZN(n458) );
  XOR2_X1 U345 ( .A(G36GAT), .B(G190GAT), .Z(n355) );
  XOR2_X1 U346 ( .A(G92GAT), .B(KEYINPUT76), .Z(n296) );
  XNOR2_X1 U347 ( .A(G99GAT), .B(G85GAT), .ZN(n295) );
  XNOR2_X1 U348 ( .A(n296), .B(n295), .ZN(n447) );
  INV_X1 U349 ( .A(n447), .ZN(n298) );
  XOR2_X1 U350 ( .A(G50GAT), .B(G162GAT), .Z(n333) );
  INV_X1 U351 ( .A(n333), .ZN(n297) );
  NAND2_X1 U352 ( .A1(n298), .A2(n297), .ZN(n300) );
  NAND2_X1 U353 ( .A1(n333), .A2(n447), .ZN(n299) );
  NAND2_X1 U354 ( .A1(n300), .A2(n299), .ZN(n303) );
  AND2_X1 U355 ( .A1(G232GAT), .A2(G233GAT), .ZN(n301) );
  XOR2_X1 U356 ( .A(G29GAT), .B(G43GAT), .Z(n305) );
  XNOR2_X1 U357 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n304) );
  XNOR2_X1 U358 ( .A(n305), .B(n304), .ZN(n437) );
  XOR2_X1 U359 ( .A(n437), .B(KEYINPUT10), .Z(n306) );
  XNOR2_X1 U360 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U361 ( .A(n355), .B(n308), .Z(n314) );
  XOR2_X1 U362 ( .A(KEYINPUT9), .B(KEYINPUT11), .Z(n310) );
  XNOR2_X1 U363 ( .A(G106GAT), .B(KEYINPUT78), .ZN(n309) );
  XNOR2_X1 U364 ( .A(n310), .B(n309), .ZN(n312) );
  XNOR2_X1 U365 ( .A(G134GAT), .B(G218GAT), .ZN(n311) );
  XNOR2_X1 U366 ( .A(KEYINPUT36), .B(n463), .ZN(n594) );
  XOR2_X1 U367 ( .A(KEYINPUT81), .B(KEYINPUT19), .Z(n316) );
  XNOR2_X1 U368 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n315) );
  XNOR2_X1 U369 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U370 ( .A(n317), .B(KEYINPUT82), .Z(n319) );
  XNOR2_X1 U371 ( .A(G169GAT), .B(G183GAT), .ZN(n318) );
  XNOR2_X1 U372 ( .A(n319), .B(n318), .ZN(n360) );
  XOR2_X1 U373 ( .A(G15GAT), .B(G127GAT), .Z(n416) );
  XOR2_X1 U374 ( .A(G71GAT), .B(G190GAT), .Z(n321) );
  XNOR2_X1 U375 ( .A(G43GAT), .B(G99GAT), .ZN(n320) );
  XNOR2_X1 U376 ( .A(n321), .B(n320), .ZN(n322) );
  NAND2_X1 U377 ( .A1(G227GAT), .A2(G233GAT), .ZN(n323) );
  XNOR2_X1 U378 ( .A(n294), .B(n323), .ZN(n329) );
  XOR2_X1 U379 ( .A(G120GAT), .B(KEYINPUT0), .Z(n325) );
  XNOR2_X1 U380 ( .A(G113GAT), .B(G134GAT), .ZN(n324) );
  XNOR2_X1 U381 ( .A(n325), .B(n324), .ZN(n376) );
  XNOR2_X1 U382 ( .A(n376), .B(KEYINPUT20), .ZN(n327) );
  XOR2_X2 U383 ( .A(n360), .B(n330), .Z(n541) );
  XOR2_X1 U384 ( .A(G78GAT), .B(G148GAT), .Z(n332) );
  XNOR2_X1 U385 ( .A(G106GAT), .B(G204GAT), .ZN(n331) );
  XNOR2_X1 U386 ( .A(n332), .B(n331), .ZN(n448) );
  XNOR2_X1 U387 ( .A(n333), .B(n448), .ZN(n334) );
  XOR2_X1 U388 ( .A(G22GAT), .B(G155GAT), .Z(n415) );
  XNOR2_X1 U389 ( .A(n334), .B(n415), .ZN(n340) );
  XOR2_X1 U390 ( .A(KEYINPUT3), .B(KEYINPUT86), .Z(n336) );
  XNOR2_X1 U391 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n335) );
  XNOR2_X1 U392 ( .A(n336), .B(n335), .ZN(n373) );
  XOR2_X1 U393 ( .A(n373), .B(KEYINPUT84), .Z(n338) );
  NAND2_X1 U394 ( .A1(G228GAT), .A2(G233GAT), .ZN(n337) );
  XNOR2_X1 U395 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U396 ( .A(n340), .B(n339), .Z(n348) );
  XOR2_X1 U397 ( .A(KEYINPUT85), .B(G218GAT), .Z(n342) );
  XNOR2_X1 U398 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n341) );
  XNOR2_X1 U399 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U400 ( .A(G197GAT), .B(n343), .Z(n356) );
  XOR2_X1 U401 ( .A(KEYINPUT83), .B(KEYINPUT23), .Z(n345) );
  XNOR2_X1 U402 ( .A(KEYINPUT22), .B(KEYINPUT24), .ZN(n344) );
  XNOR2_X1 U403 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U404 ( .A(n356), .B(n346), .ZN(n347) );
  XNOR2_X1 U405 ( .A(n348), .B(n347), .ZN(n481) );
  XOR2_X1 U406 ( .A(G176GAT), .B(G64GAT), .Z(n451) );
  XOR2_X1 U407 ( .A(n451), .B(KEYINPUT91), .Z(n350) );
  NAND2_X1 U408 ( .A1(G226GAT), .A2(G233GAT), .ZN(n349) );
  XNOR2_X1 U409 ( .A(n350), .B(n349), .ZN(n354) );
  XOR2_X1 U410 ( .A(KEYINPUT92), .B(G92GAT), .Z(n352) );
  XNOR2_X1 U411 ( .A(G8GAT), .B(G204GAT), .ZN(n351) );
  XNOR2_X1 U412 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U413 ( .A(n354), .B(n353), .Z(n358) );
  XNOR2_X1 U414 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U415 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U416 ( .A(n360), .B(n359), .Z(n477) );
  XOR2_X1 U417 ( .A(n477), .B(KEYINPUT93), .Z(n361) );
  XNOR2_X1 U418 ( .A(KEYINPUT27), .B(n361), .ZN(n536) );
  NOR2_X1 U419 ( .A1(n543), .A2(n536), .ZN(n384) );
  INV_X1 U420 ( .A(n384), .ZN(n383) );
  XOR2_X1 U421 ( .A(KEYINPUT88), .B(KEYINPUT87), .Z(n363) );
  XNOR2_X1 U422 ( .A(KEYINPUT89), .B(KEYINPUT90), .ZN(n362) );
  XNOR2_X1 U423 ( .A(n363), .B(n362), .ZN(n367) );
  XOR2_X1 U424 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n365) );
  XNOR2_X1 U425 ( .A(G1GAT), .B(G57GAT), .ZN(n364) );
  XNOR2_X1 U426 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U427 ( .A(n367), .B(n366), .ZN(n371) );
  XOR2_X1 U428 ( .A(G155GAT), .B(G148GAT), .Z(n369) );
  XNOR2_X1 U429 ( .A(G127GAT), .B(G162GAT), .ZN(n368) );
  XNOR2_X1 U430 ( .A(n369), .B(n368), .ZN(n370) );
  XNOR2_X1 U431 ( .A(n371), .B(n370), .ZN(n372) );
  XOR2_X1 U432 ( .A(n372), .B(KEYINPUT5), .Z(n375) );
  XNOR2_X1 U433 ( .A(n373), .B(KEYINPUT4), .ZN(n374) );
  XNOR2_X1 U434 ( .A(n375), .B(n374), .ZN(n381) );
  XOR2_X1 U435 ( .A(G85GAT), .B(n376), .Z(n378) );
  NAND2_X1 U436 ( .A1(G225GAT), .A2(G233GAT), .ZN(n377) );
  XNOR2_X1 U437 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X1 U438 ( .A(G29GAT), .B(n379), .Z(n380) );
  XNOR2_X1 U439 ( .A(n381), .B(n380), .ZN(n539) );
  NAND2_X1 U440 ( .A1(KEYINPUT94), .A2(n539), .ZN(n382) );
  NOR2_X1 U441 ( .A1(n383), .A2(n382), .ZN(n386) );
  NOR2_X1 U442 ( .A1(KEYINPUT94), .A2(n384), .ZN(n385) );
  NOR2_X1 U443 ( .A1(n386), .A2(n385), .ZN(n387) );
  NOR2_X1 U444 ( .A1(n541), .A2(n387), .ZN(n401) );
  NOR2_X1 U445 ( .A1(n541), .A2(KEYINPUT94), .ZN(n398) );
  XNOR2_X1 U446 ( .A(KEYINPUT26), .B(KEYINPUT95), .ZN(n389) );
  NOR2_X1 U447 ( .A1(n541), .A2(n481), .ZN(n388) );
  XNOR2_X1 U448 ( .A(n389), .B(n388), .ZN(n557) );
  NOR2_X1 U449 ( .A1(n557), .A2(n536), .ZN(n391) );
  XNOR2_X1 U450 ( .A(n391), .B(n390), .ZN(n396) );
  INV_X1 U451 ( .A(n477), .ZN(n527) );
  NAND2_X1 U452 ( .A1(n527), .A2(n541), .ZN(n392) );
  NAND2_X1 U453 ( .A1(n392), .A2(n481), .ZN(n393) );
  XNOR2_X1 U454 ( .A(n393), .B(KEYINPUT25), .ZN(n394) );
  XNOR2_X1 U455 ( .A(KEYINPUT97), .B(n394), .ZN(n395) );
  NAND2_X1 U456 ( .A1(n396), .A2(n395), .ZN(n397) );
  NOR2_X1 U457 ( .A1(n398), .A2(n397), .ZN(n399) );
  NOR2_X1 U458 ( .A1(n539), .A2(n399), .ZN(n400) );
  XOR2_X1 U459 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n403) );
  NAND2_X1 U460 ( .A1(G231GAT), .A2(G233GAT), .ZN(n402) );
  XNOR2_X1 U461 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U462 ( .A(n404), .B(KEYINPUT15), .Z(n410) );
  XOR2_X1 U463 ( .A(G1GAT), .B(G8GAT), .Z(n406) );
  XNOR2_X1 U464 ( .A(KEYINPUT71), .B(KEYINPUT72), .ZN(n405) );
  XNOR2_X1 U465 ( .A(n406), .B(n405), .ZN(n436) );
  XOR2_X1 U466 ( .A(KEYINPUT13), .B(KEYINPUT75), .Z(n408) );
  XNOR2_X1 U467 ( .A(G71GAT), .B(G57GAT), .ZN(n407) );
  XNOR2_X1 U468 ( .A(n408), .B(n407), .ZN(n456) );
  XNOR2_X1 U469 ( .A(n436), .B(n456), .ZN(n409) );
  XNOR2_X1 U470 ( .A(n410), .B(n409), .ZN(n414) );
  XOR2_X1 U471 ( .A(G64GAT), .B(G78GAT), .Z(n412) );
  XNOR2_X1 U472 ( .A(G183GAT), .B(G211GAT), .ZN(n411) );
  XNOR2_X1 U473 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U474 ( .A(n414), .B(n413), .Z(n418) );
  XNOR2_X1 U475 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U476 ( .A(n418), .B(n417), .ZN(n577) );
  INV_X1 U477 ( .A(n577), .ZN(n590) );
  NOR2_X1 U478 ( .A1(n492), .A2(n590), .ZN(n419) );
  XOR2_X1 U479 ( .A(KEYINPUT102), .B(n419), .Z(n420) );
  NOR2_X1 U480 ( .A1(n594), .A2(n420), .ZN(n421) );
  XOR2_X1 U481 ( .A(KEYINPUT37), .B(n421), .Z(n523) );
  NAND2_X1 U482 ( .A1(G229GAT), .A2(G233GAT), .ZN(n427) );
  XOR2_X1 U483 ( .A(G22GAT), .B(G197GAT), .Z(n423) );
  XNOR2_X1 U484 ( .A(G169GAT), .B(G141GAT), .ZN(n422) );
  XNOR2_X1 U485 ( .A(n423), .B(n422), .ZN(n425) );
  XOR2_X1 U486 ( .A(G50GAT), .B(G36GAT), .Z(n424) );
  XNOR2_X1 U487 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U488 ( .A(n427), .B(n426), .ZN(n443) );
  XOR2_X1 U489 ( .A(KEYINPUT69), .B(KEYINPUT70), .Z(n429) );
  XNOR2_X1 U490 ( .A(KEYINPUT66), .B(KEYINPUT29), .ZN(n428) );
  XNOR2_X1 U491 ( .A(n429), .B(n428), .ZN(n441) );
  XOR2_X1 U492 ( .A(KEYINPUT73), .B(KEYINPUT74), .Z(n431) );
  XNOR2_X1 U493 ( .A(G15GAT), .B(G113GAT), .ZN(n430) );
  XNOR2_X1 U494 ( .A(n431), .B(n430), .ZN(n435) );
  XOR2_X1 U495 ( .A(KEYINPUT65), .B(KEYINPUT30), .Z(n433) );
  XNOR2_X1 U496 ( .A(KEYINPUT67), .B(KEYINPUT68), .ZN(n432) );
  XNOR2_X1 U497 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U498 ( .A(n435), .B(n434), .Z(n439) );
  XNOR2_X1 U499 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U500 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U501 ( .A(n441), .B(n440), .Z(n442) );
  XNOR2_X1 U502 ( .A(n443), .B(n442), .ZN(n581) );
  XOR2_X1 U503 ( .A(KEYINPUT31), .B(KEYINPUT32), .Z(n445) );
  NAND2_X1 U504 ( .A1(G230GAT), .A2(G233GAT), .ZN(n444) );
  XNOR2_X1 U505 ( .A(n445), .B(n444), .ZN(n446) );
  XOR2_X1 U506 ( .A(n446), .B(KEYINPUT33), .Z(n450) );
  XNOR2_X1 U507 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U508 ( .A(n450), .B(n449), .ZN(n452) );
  XOR2_X1 U509 ( .A(n452), .B(n451), .Z(n454) );
  XNOR2_X1 U510 ( .A(G120GAT), .B(KEYINPUT77), .ZN(n453) );
  XNOR2_X1 U511 ( .A(n454), .B(n453), .ZN(n455) );
  XOR2_X1 U512 ( .A(n456), .B(n455), .Z(n586) );
  NOR2_X1 U513 ( .A1(n581), .A2(n586), .ZN(n493) );
  NAND2_X1 U514 ( .A1(n523), .A2(n493), .ZN(n457) );
  NAND2_X1 U515 ( .A1(n508), .A2(n541), .ZN(n460) );
  XNOR2_X1 U516 ( .A(KEYINPUT113), .B(KEYINPUT47), .ZN(n467) );
  XNOR2_X1 U517 ( .A(KEYINPUT41), .B(n586), .ZN(n560) );
  NOR2_X1 U518 ( .A1(n581), .A2(n560), .ZN(n462) );
  XNOR2_X1 U519 ( .A(KEYINPUT112), .B(KEYINPUT46), .ZN(n461) );
  XNOR2_X1 U520 ( .A(n462), .B(n461), .ZN(n465) );
  NAND2_X1 U521 ( .A1(n577), .A2(n463), .ZN(n464) );
  NOR2_X1 U522 ( .A1(n465), .A2(n464), .ZN(n466) );
  XNOR2_X1 U523 ( .A(n467), .B(n466), .ZN(n475) );
  XNOR2_X1 U524 ( .A(KEYINPUT64), .B(KEYINPUT45), .ZN(n469) );
  NOR2_X1 U525 ( .A1(n577), .A2(n594), .ZN(n468) );
  XOR2_X1 U526 ( .A(n469), .B(n468), .Z(n470) );
  NOR2_X1 U527 ( .A1(n586), .A2(n470), .ZN(n472) );
  INV_X1 U528 ( .A(KEYINPUT114), .ZN(n471) );
  XNOR2_X1 U529 ( .A(n472), .B(n471), .ZN(n473) );
  INV_X1 U530 ( .A(n581), .ZN(n544) );
  NOR2_X1 U531 ( .A1(n473), .A2(n544), .ZN(n474) );
  NOR2_X1 U532 ( .A1(n475), .A2(n474), .ZN(n476) );
  XNOR2_X1 U533 ( .A(n476), .B(KEYINPUT48), .ZN(n537) );
  NOR2_X1 U534 ( .A1(n477), .A2(n537), .ZN(n479) );
  INV_X1 U535 ( .A(KEYINPUT54), .ZN(n478) );
  XNOR2_X1 U536 ( .A(n479), .B(n478), .ZN(n480) );
  NOR2_X1 U537 ( .A1(n480), .A2(n539), .ZN(n580) );
  NAND2_X1 U538 ( .A1(n580), .A2(n481), .ZN(n484) );
  XOR2_X1 U539 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n482) );
  NAND2_X1 U540 ( .A1(n485), .A2(n541), .ZN(n576) );
  NOR2_X1 U541 ( .A1(n576), .A2(n463), .ZN(n488) );
  INV_X1 U542 ( .A(G190GAT), .ZN(n486) );
  XOR2_X1 U543 ( .A(KEYINPUT34), .B(KEYINPUT98), .Z(n495) );
  NAND2_X1 U544 ( .A1(n590), .A2(n463), .ZN(n489) );
  XNOR2_X1 U545 ( .A(n489), .B(KEYINPUT80), .ZN(n490) );
  XNOR2_X1 U546 ( .A(n490), .B(KEYINPUT16), .ZN(n491) );
  NOR2_X1 U547 ( .A1(n492), .A2(n491), .ZN(n511) );
  AND2_X1 U548 ( .A1(n493), .A2(n511), .ZN(n501) );
  NAND2_X1 U549 ( .A1(n501), .A2(n539), .ZN(n494) );
  XNOR2_X1 U550 ( .A(n495), .B(n494), .ZN(n496) );
  XOR2_X1 U551 ( .A(G1GAT), .B(n496), .Z(G1324GAT) );
  NAND2_X1 U552 ( .A1(n527), .A2(n501), .ZN(n497) );
  XNOR2_X1 U553 ( .A(n497), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U554 ( .A(KEYINPUT35), .B(KEYINPUT99), .Z(n499) );
  NAND2_X1 U555 ( .A1(n501), .A2(n541), .ZN(n498) );
  XNOR2_X1 U556 ( .A(n499), .B(n498), .ZN(n500) );
  XOR2_X1 U557 ( .A(G15GAT), .B(n500), .Z(G1326GAT) );
  NAND2_X1 U558 ( .A1(n501), .A2(n543), .ZN(n502) );
  XNOR2_X1 U559 ( .A(n502), .B(KEYINPUT100), .ZN(n503) );
  XNOR2_X1 U560 ( .A(G22GAT), .B(n503), .ZN(G1327GAT) );
  NAND2_X1 U561 ( .A1(n508), .A2(n539), .ZN(n506) );
  XNOR2_X1 U562 ( .A(G29GAT), .B(KEYINPUT101), .ZN(n504) );
  XNOR2_X1 U563 ( .A(n504), .B(KEYINPUT39), .ZN(n505) );
  XNOR2_X1 U564 ( .A(n506), .B(n505), .ZN(G1328GAT) );
  NAND2_X1 U565 ( .A1(n508), .A2(n527), .ZN(n507) );
  XNOR2_X1 U566 ( .A(n507), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U567 ( .A1(n508), .A2(n543), .ZN(n509) );
  XNOR2_X1 U568 ( .A(n509), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U569 ( .A(KEYINPUT105), .B(n560), .Z(n571) );
  NOR2_X1 U570 ( .A1(n544), .A2(n571), .ZN(n510) );
  XOR2_X1 U571 ( .A(KEYINPUT106), .B(n510), .Z(n525) );
  INV_X1 U572 ( .A(n511), .ZN(n512) );
  NOR2_X1 U573 ( .A1(n525), .A2(n512), .ZN(n520) );
  NAND2_X1 U574 ( .A1(n539), .A2(n520), .ZN(n515) );
  XNOR2_X1 U575 ( .A(G57GAT), .B(KEYINPUT104), .ZN(n513) );
  XNOR2_X1 U576 ( .A(n513), .B(KEYINPUT42), .ZN(n514) );
  XNOR2_X1 U577 ( .A(n515), .B(n514), .ZN(G1332GAT) );
  XOR2_X1 U578 ( .A(G64GAT), .B(KEYINPUT107), .Z(n517) );
  NAND2_X1 U579 ( .A1(n520), .A2(n527), .ZN(n516) );
  XNOR2_X1 U580 ( .A(n517), .B(n516), .ZN(G1333GAT) );
  NAND2_X1 U581 ( .A1(n520), .A2(n541), .ZN(n518) );
  XNOR2_X1 U582 ( .A(n518), .B(KEYINPUT108), .ZN(n519) );
  XNOR2_X1 U583 ( .A(G71GAT), .B(n519), .ZN(G1334GAT) );
  XOR2_X1 U584 ( .A(G78GAT), .B(KEYINPUT43), .Z(n522) );
  NAND2_X1 U585 ( .A1(n520), .A2(n543), .ZN(n521) );
  XNOR2_X1 U586 ( .A(n522), .B(n521), .ZN(G1335GAT) );
  INV_X1 U587 ( .A(n523), .ZN(n524) );
  NOR2_X1 U588 ( .A1(n525), .A2(n524), .ZN(n532) );
  NAND2_X1 U589 ( .A1(n539), .A2(n532), .ZN(n526) );
  XNOR2_X1 U590 ( .A(n526), .B(G85GAT), .ZN(G1336GAT) );
  XOR2_X1 U591 ( .A(G92GAT), .B(KEYINPUT109), .Z(n529) );
  NAND2_X1 U592 ( .A1(n532), .A2(n527), .ZN(n528) );
  XNOR2_X1 U593 ( .A(n529), .B(n528), .ZN(G1337GAT) );
  NAND2_X1 U594 ( .A1(n532), .A2(n541), .ZN(n530) );
  XNOR2_X1 U595 ( .A(n530), .B(KEYINPUT110), .ZN(n531) );
  XNOR2_X1 U596 ( .A(G99GAT), .B(n531), .ZN(G1338GAT) );
  XOR2_X1 U597 ( .A(KEYINPUT111), .B(KEYINPUT44), .Z(n534) );
  NAND2_X1 U598 ( .A1(n532), .A2(n543), .ZN(n533) );
  XNOR2_X1 U599 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U600 ( .A(G106GAT), .B(n535), .ZN(G1339GAT) );
  NOR2_X1 U601 ( .A1(n537), .A2(n536), .ZN(n538) );
  NAND2_X1 U602 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U603 ( .A(n540), .B(KEYINPUT115), .ZN(n558) );
  NAND2_X1 U604 ( .A1(n541), .A2(n558), .ZN(n542) );
  NOR2_X1 U605 ( .A1(n543), .A2(n542), .ZN(n550) );
  NAND2_X1 U606 ( .A1(n544), .A2(n550), .ZN(n545) );
  XNOR2_X1 U607 ( .A(n545), .B(KEYINPUT116), .ZN(n546) );
  XNOR2_X1 U608 ( .A(G113GAT), .B(n546), .ZN(G1340GAT) );
  INV_X1 U609 ( .A(n550), .ZN(n554) );
  NOR2_X1 U610 ( .A1(n571), .A2(n554), .ZN(n548) );
  XNOR2_X1 U611 ( .A(KEYINPUT117), .B(KEYINPUT49), .ZN(n547) );
  XNOR2_X1 U612 ( .A(n548), .B(n547), .ZN(n549) );
  XOR2_X1 U613 ( .A(G120GAT), .B(n549), .Z(G1341GAT) );
  XOR2_X1 U614 ( .A(KEYINPUT50), .B(KEYINPUT118), .Z(n552) );
  NAND2_X1 U615 ( .A1(n550), .A2(n590), .ZN(n551) );
  XNOR2_X1 U616 ( .A(n552), .B(n551), .ZN(n553) );
  XOR2_X1 U617 ( .A(G127GAT), .B(n553), .Z(G1342GAT) );
  NOR2_X1 U618 ( .A1(n463), .A2(n554), .ZN(n556) );
  XNOR2_X1 U619 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n555) );
  XNOR2_X1 U620 ( .A(n556), .B(n555), .ZN(G1343GAT) );
  INV_X1 U621 ( .A(n557), .ZN(n579) );
  NAND2_X1 U622 ( .A1(n558), .A2(n579), .ZN(n566) );
  NOR2_X1 U623 ( .A1(n581), .A2(n566), .ZN(n559) );
  XOR2_X1 U624 ( .A(G141GAT), .B(n559), .Z(G1344GAT) );
  NOR2_X1 U625 ( .A1(n560), .A2(n566), .ZN(n562) );
  XNOR2_X1 U626 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n561) );
  XNOR2_X1 U627 ( .A(n562), .B(n561), .ZN(n563) );
  XNOR2_X1 U628 ( .A(G148GAT), .B(n563), .ZN(G1345GAT) );
  NOR2_X1 U629 ( .A1(n577), .A2(n566), .ZN(n565) );
  XNOR2_X1 U630 ( .A(G155GAT), .B(KEYINPUT119), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n565), .B(n564), .ZN(G1346GAT) );
  NOR2_X1 U632 ( .A1(n463), .A2(n566), .ZN(n567) );
  XOR2_X1 U633 ( .A(KEYINPUT120), .B(n567), .Z(n568) );
  XNOR2_X1 U634 ( .A(G162GAT), .B(n568), .ZN(G1347GAT) );
  NOR2_X1 U635 ( .A1(n581), .A2(n576), .ZN(n570) );
  XNOR2_X1 U636 ( .A(G169GAT), .B(KEYINPUT123), .ZN(n569) );
  XNOR2_X1 U637 ( .A(n570), .B(n569), .ZN(G1348GAT) );
  XNOR2_X1 U638 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n575) );
  NOR2_X1 U639 ( .A1(n576), .A2(n571), .ZN(n573) );
  XNOR2_X1 U640 ( .A(G176GAT), .B(KEYINPUT124), .ZN(n572) );
  XNOR2_X1 U641 ( .A(n573), .B(n572), .ZN(n574) );
  XNOR2_X1 U642 ( .A(n575), .B(n574), .ZN(G1349GAT) );
  NOR2_X1 U643 ( .A1(n577), .A2(n576), .ZN(n578) );
  XOR2_X1 U644 ( .A(G183GAT), .B(n578), .Z(G1350GAT) );
  NAND2_X1 U645 ( .A1(n580), .A2(n579), .ZN(n593) );
  NOR2_X1 U646 ( .A1(n581), .A2(n593), .ZN(n583) );
  XNOR2_X1 U647 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(n585) );
  XOR2_X1 U649 ( .A(KEYINPUT60), .B(KEYINPUT125), .Z(n584) );
  XNOR2_X1 U650 ( .A(n585), .B(n584), .ZN(G1352GAT) );
  XOR2_X1 U651 ( .A(G204GAT), .B(KEYINPUT61), .Z(n588) );
  INV_X1 U652 ( .A(n593), .ZN(n589) );
  NAND2_X1 U653 ( .A1(n589), .A2(n586), .ZN(n587) );
  XNOR2_X1 U654 ( .A(n588), .B(n587), .ZN(G1353GAT) );
  NAND2_X1 U655 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U656 ( .A(n591), .B(KEYINPUT126), .ZN(n592) );
  XNOR2_X1 U657 ( .A(G211GAT), .B(n592), .ZN(G1354GAT) );
  NOR2_X1 U658 ( .A1(n594), .A2(n593), .ZN(n595) );
  XOR2_X1 U659 ( .A(KEYINPUT62), .B(n595), .Z(n596) );
  XNOR2_X1 U660 ( .A(G218GAT), .B(n596), .ZN(G1355GAT) );
endmodule

