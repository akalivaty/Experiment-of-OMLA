//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 0 0 1 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 0 1 0 0 0 0 1 0 0 0 0 0 1 1 1 1 1 0 0 1 0 1 0 1 0 1 0 0 1 1 1 1 1 1 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:29 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n257, new_n258, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1273, new_n1274, new_n1275, new_n1277, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1351;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT64), .ZN(G353));
  INV_X1    g0005(.A(G97), .ZN(new_n206));
  INV_X1    g0006(.A(G107), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G87), .ZN(G355));
  NAND2_X1  g0009(.A1(G1), .A2(G20), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n211));
  INV_X1    g0011(.A(G68), .ZN(new_n212));
  INV_X1    g0012(.A(G238), .ZN(new_n213));
  INV_X1    g0013(.A(G87), .ZN(new_n214));
  INV_X1    g0014(.A(G250), .ZN(new_n215));
  OAI221_X1 g0015(.A(new_n211), .B1(new_n212), .B2(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n210), .B1(new_n216), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n220), .A2(KEYINPUT1), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n221), .B(KEYINPUT66), .ZN(new_n222));
  OR2_X1    g0022(.A1(new_n220), .A2(KEYINPUT1), .ZN(new_n223));
  INV_X1    g0023(.A(new_n223), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n210), .A2(G13), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n225), .B(G250), .C1(G257), .C2(G264), .ZN(new_n226));
  INV_X1    g0026(.A(new_n226), .ZN(new_n227));
  OR2_X1    g0027(.A1(new_n227), .A2(KEYINPUT0), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n227), .A2(KEYINPUT0), .ZN(new_n229));
  AND3_X1   g0029(.A1(KEYINPUT65), .A2(G1), .A3(G13), .ZN(new_n230));
  AOI21_X1  g0030(.A(KEYINPUT65), .B1(G1), .B2(G13), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  INV_X1    g0032(.A(G20), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  INV_X1    g0034(.A(new_n234), .ZN(new_n235));
  INV_X1    g0035(.A(new_n201), .ZN(new_n236));
  NAND2_X1  g0036(.A1(new_n236), .A2(G50), .ZN(new_n237));
  OAI211_X1 g0037(.A(new_n228), .B(new_n229), .C1(new_n235), .C2(new_n237), .ZN(new_n238));
  NOR3_X1   g0038(.A1(new_n222), .A2(new_n224), .A3(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT67), .ZN(G361));
  XOR2_X1   g0040(.A(G238), .B(G244), .Z(new_n241));
  XNOR2_X1  g0041(.A(KEYINPUT68), .B(G232), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(KEYINPUT2), .B(G226), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G250), .B(G257), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(KEYINPUT69), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G264), .B(G270), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n245), .B(new_n249), .ZN(G358));
  XOR2_X1   g0050(.A(G107), .B(G116), .Z(new_n251));
  XNOR2_X1  g0051(.A(G87), .B(G97), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n202), .A2(G68), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n212), .A2(G50), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  XNOR2_X1  g0056(.A(G58), .B(G77), .ZN(new_n257));
  XNOR2_X1  g0057(.A(new_n256), .B(new_n257), .ZN(new_n258));
  XNOR2_X1  g0058(.A(new_n253), .B(new_n258), .ZN(G351));
  NAND2_X1  g0059(.A1(KEYINPUT71), .A2(G58), .ZN(new_n260));
  XNOR2_X1  g0060(.A(new_n260), .B(KEYINPUT8), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n233), .A2(G33), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  NOR2_X1   g0064(.A1(G20), .A2(G33), .ZN(new_n265));
  AOI22_X1  g0065(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(G1), .A2(G13), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT65), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g0070(.A1(KEYINPUT65), .A2(G1), .A3(G13), .ZN(new_n271));
  NAND3_X1  g0071(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n270), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G1), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n274), .A2(G13), .A3(G20), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  AOI22_X1  g0076(.A1(new_n267), .A2(new_n273), .B1(new_n202), .B2(new_n276), .ZN(new_n277));
  NAND4_X1  g0077(.A1(new_n270), .A2(new_n275), .A3(new_n271), .A4(new_n272), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n274), .A2(G20), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n279), .A2(G50), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n277), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(G33), .A2(G41), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n283), .A2(G1), .A3(G13), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G41), .ZN(new_n286));
  INV_X1    g0086(.A(G45), .ZN(new_n287));
  AOI21_X1  g0087(.A(G1), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n285), .A2(new_n288), .ZN(new_n289));
  XOR2_X1   g0089(.A(KEYINPUT70), .B(G226), .Z(new_n290));
  AND2_X1   g0090(.A1(new_n284), .A2(G274), .ZN(new_n291));
  AOI22_X1  g0091(.A1(new_n289), .A2(new_n290), .B1(new_n291), .B2(new_n288), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n283), .B1(new_n230), .B2(new_n231), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  XNOR2_X1  g0094(.A(KEYINPUT3), .B(G33), .ZN(new_n295));
  NOR2_X1   g0095(.A1(G222), .A2(G1698), .ZN(new_n296));
  INV_X1    g0096(.A(G1698), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n297), .A2(G223), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n295), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n294), .B(new_n299), .C1(G77), .C2(new_n295), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n292), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G169), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G179), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n292), .A2(new_n300), .A3(new_n304), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n282), .A2(new_n303), .A3(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n282), .A2(KEYINPUT9), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT9), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n277), .A2(new_n309), .A3(new_n281), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(G190), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n301), .A2(new_n312), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n313), .B1(G200), .B2(new_n301), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n311), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(KEYINPUT10), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT10), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n311), .A2(new_n314), .A3(new_n317), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n307), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  XOR2_X1   g0119(.A(KEYINPUT75), .B(KEYINPUT13), .Z(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(G226), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(new_n297), .ZN(new_n323));
  OAI211_X1 g0123(.A(new_n295), .B(new_n323), .C1(G232), .C2(new_n297), .ZN(new_n324));
  NAND2_X1  g0124(.A1(G33), .A2(G97), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT74), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g0127(.A1(KEYINPUT74), .A2(G33), .A3(G97), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n293), .B1(new_n324), .B2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n288), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(new_n284), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n284), .A2(G274), .ZN(new_n334));
  OAI22_X1  g0134(.A1(new_n333), .A2(new_n213), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n321), .B1(new_n331), .B2(new_n336), .ZN(new_n337));
  NOR3_X1   g0137(.A1(new_n330), .A2(new_n335), .A3(new_n320), .ZN(new_n338));
  OAI21_X1  g0138(.A(G169), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(KEYINPUT14), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n330), .A2(new_n335), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT13), .ZN(new_n342));
  OAI21_X1  g0142(.A(KEYINPUT76), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT76), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n344), .B(KEYINPUT13), .C1(new_n330), .C2(new_n335), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n341), .A2(new_n321), .ZN(new_n346));
  NAND4_X1  g0146(.A1(new_n343), .A2(G179), .A3(new_n345), .A4(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT14), .ZN(new_n348));
  OAI211_X1 g0148(.A(new_n348), .B(G169), .C1(new_n337), .C2(new_n338), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n340), .A2(new_n347), .A3(new_n349), .ZN(new_n350));
  AOI22_X1  g0150(.A1(new_n265), .A2(G50), .B1(G20), .B2(new_n212), .ZN(new_n351));
  INV_X1    g0151(.A(G77), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n351), .B1(new_n352), .B2(new_n262), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(new_n273), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT11), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT77), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n276), .A2(new_n212), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n357), .B1(new_n358), .B2(KEYINPUT78), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n356), .B1(KEYINPUT12), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n279), .A2(KEYINPUT73), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT73), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n278), .A2(new_n362), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n361), .A2(G68), .A3(new_n280), .A4(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(new_n359), .ZN(new_n365));
  AOI21_X1  g0165(.A(KEYINPUT12), .B1(new_n358), .B2(new_n357), .ZN(new_n366));
  AOI22_X1  g0166(.A1(new_n365), .A2(new_n366), .B1(new_n354), .B2(new_n355), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n360), .A2(new_n364), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n350), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n368), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n343), .A2(G190), .A3(new_n345), .A4(new_n346), .ZN(new_n371));
  OAI21_X1  g0171(.A(G200), .B1(new_n337), .B2(new_n338), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n370), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n352), .B1(new_n274), .B2(G20), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n361), .A2(new_n363), .A3(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(new_n375), .ZN(new_n376));
  AND3_X1   g0176(.A1(new_n270), .A2(new_n271), .A3(new_n272), .ZN(new_n377));
  XNOR2_X1  g0177(.A(KEYINPUT8), .B(G58), .ZN(new_n378));
  OR2_X1    g0178(.A1(new_n378), .A2(KEYINPUT72), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(KEYINPUT72), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n379), .A2(new_n265), .A3(new_n380), .ZN(new_n381));
  XNOR2_X1  g0181(.A(KEYINPUT15), .B(G87), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  AOI22_X1  g0183(.A1(new_n383), .A2(new_n263), .B1(G20), .B2(G77), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n377), .B1(new_n381), .B2(new_n384), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n275), .A2(G77), .ZN(new_n386));
  OR3_X1    g0186(.A1(new_n376), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n295), .A2(G232), .A3(new_n297), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n388), .B1(new_n207), .B2(new_n295), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT3), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(G33), .ZN(new_n391));
  INV_X1    g0191(.A(G33), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(KEYINPUT3), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  NOR3_X1   g0194(.A1(new_n394), .A2(new_n213), .A3(new_n297), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n294), .B1(new_n389), .B2(new_n395), .ZN(new_n396));
  AOI22_X1  g0196(.A1(new_n289), .A2(G244), .B1(new_n291), .B2(new_n288), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(new_n302), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n396), .A2(new_n304), .A3(new_n397), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n387), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  NOR3_X1   g0201(.A1(new_n376), .A2(new_n385), .A3(new_n386), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n398), .A2(G200), .ZN(new_n403));
  OAI211_X1 g0203(.A(new_n402), .B(new_n403), .C1(new_n312), .C2(new_n398), .ZN(new_n404));
  AND2_X1   g0204(.A1(new_n401), .A2(new_n404), .ZN(new_n405));
  NAND4_X1  g0205(.A1(new_n319), .A2(new_n369), .A3(new_n373), .A4(new_n405), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n261), .A2(new_n275), .ZN(new_n407));
  AND2_X1   g0207(.A1(new_n261), .A2(new_n280), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n407), .B1(new_n408), .B2(new_n279), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT79), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n391), .A2(new_n393), .A3(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT80), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT7), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n413), .A2(G20), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n390), .A2(KEYINPUT79), .A3(G33), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n411), .A2(new_n412), .A3(new_n414), .A4(new_n415), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n413), .B1(new_n295), .B2(G20), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  AND2_X1   g0218(.A1(new_n415), .A2(new_n414), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n412), .B1(new_n419), .B2(new_n411), .ZN(new_n420));
  OAI21_X1  g0220(.A(G68), .B1(new_n418), .B2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(G58), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n422), .A2(new_n212), .ZN(new_n423));
  OAI21_X1  g0223(.A(G20), .B1(new_n423), .B2(new_n201), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n265), .A2(G159), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(KEYINPUT16), .B1(new_n421), .B2(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(KEYINPUT7), .B1(new_n394), .B2(new_n233), .ZN(new_n429));
  AOI211_X1 g0229(.A(new_n413), .B(G20), .C1(new_n391), .C2(new_n393), .ZN(new_n430));
  OAI21_X1  g0230(.A(G68), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(new_n427), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT16), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n273), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n409), .B1(new_n428), .B2(new_n434), .ZN(new_n435));
  AOI22_X1  g0235(.A1(new_n289), .A2(G232), .B1(new_n291), .B2(new_n288), .ZN(new_n436));
  OR2_X1    g0236(.A1(G223), .A2(G1698), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n322), .A2(G1698), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n391), .A2(new_n437), .A3(new_n393), .A4(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(G33), .A2(G87), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n439), .A2(KEYINPUT81), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(new_n294), .ZN(new_n442));
  AOI21_X1  g0242(.A(KEYINPUT81), .B1(new_n439), .B2(new_n440), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n436), .B(KEYINPUT82), .C1(new_n442), .C2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n439), .A2(new_n440), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT81), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n448), .A2(new_n294), .A3(new_n441), .ZN(new_n449));
  AOI21_X1  g0249(.A(KEYINPUT82), .B1(new_n449), .B2(new_n436), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n302), .B1(new_n445), .B2(new_n450), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n449), .A2(new_n304), .A3(new_n436), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n435), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(KEYINPUT18), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT17), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n449), .A2(new_n312), .A3(new_n436), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n436), .B1(new_n442), .B2(new_n443), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT82), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(new_n444), .ZN(new_n461));
  INV_X1    g0261(.A(G200), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n457), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n455), .B1(new_n463), .B2(new_n435), .ZN(new_n464));
  INV_X1    g0264(.A(new_n409), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n421), .A2(new_n427), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(new_n433), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n394), .A2(new_n414), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n417), .A2(new_n468), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n426), .B1(new_n469), .B2(G68), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n377), .B1(new_n470), .B2(KEYINPUT16), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n465), .B1(new_n467), .B2(new_n471), .ZN(new_n472));
  AOI21_X1  g0272(.A(G200), .B1(new_n460), .B2(new_n444), .ZN(new_n473));
  OAI211_X1 g0273(.A(new_n472), .B(KEYINPUT17), .C1(new_n473), .C2(new_n457), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT18), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n435), .A2(new_n451), .A3(new_n475), .A4(new_n452), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n454), .A2(new_n464), .A3(new_n474), .A4(new_n476), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n406), .A2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n274), .A2(G45), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT5), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(new_n286), .ZN(new_n482));
  NAND2_X1  g0282(.A1(KEYINPUT5), .A2(G41), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n480), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n484), .A2(new_n285), .ZN(new_n485));
  AOI22_X1  g0285(.A1(new_n485), .A2(G264), .B1(new_n291), .B2(new_n484), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n391), .A2(new_n393), .A3(G257), .A4(G1698), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n391), .A2(new_n393), .A3(G250), .A4(new_n297), .ZN(new_n488));
  INV_X1    g0288(.A(G294), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n487), .B(new_n488), .C1(new_n392), .C2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(new_n294), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n486), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(G169), .ZN(new_n493));
  AOI22_X1  g0293(.A1(new_n490), .A2(new_n294), .B1(new_n291), .B2(new_n484), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n287), .A2(G1), .ZN(new_n495));
  INV_X1    g0295(.A(new_n483), .ZN(new_n496));
  NOR2_X1   g0296(.A1(KEYINPUT5), .A2(G41), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n498), .A2(G264), .A3(new_n284), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT87), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n498), .A2(KEYINPUT87), .A3(G264), .A4(new_n284), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n494), .A2(new_n503), .A3(G179), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n493), .A2(new_n504), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n391), .A2(new_n393), .A3(new_n233), .A4(G87), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(KEYINPUT22), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT22), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n295), .A2(new_n508), .A3(new_n233), .A4(G87), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT23), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n511), .A2(new_n207), .A3(G20), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(KEYINPUT86), .ZN(new_n513));
  NAND2_X1  g0313(.A1(KEYINPUT23), .A2(G107), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n516));
  OAI22_X1  g0316(.A1(new_n512), .A2(KEYINPUT86), .B1(new_n516), .B2(G20), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n510), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(KEYINPUT24), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT24), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n510), .A2(new_n518), .A3(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n377), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT85), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n392), .A2(G1), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n377), .A2(new_n524), .A3(new_n275), .A4(new_n526), .ZN(new_n527));
  OAI21_X1  g0327(.A(KEYINPUT85), .B1(new_n278), .B2(new_n525), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n207), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n276), .A2(new_n207), .ZN(new_n530));
  XNOR2_X1  g0330(.A(new_n530), .B(KEYINPUT25), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(new_n532), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n505), .B1(new_n523), .B2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(G116), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n525), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n361), .A2(new_n363), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n535), .A2(G20), .ZN(new_n538));
  INV_X1    g0338(.A(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(G13), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n540), .A2(G1), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n206), .A2(KEYINPUT83), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT83), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(G97), .ZN(new_n545));
  AOI21_X1  g0345(.A(G33), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(G33), .A2(G283), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(new_n233), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n273), .B(new_n538), .C1(new_n546), .C2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT20), .ZN(new_n550));
  AND2_X1   g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n549), .A2(new_n550), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n537), .B(new_n542), .C1(new_n551), .C2(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n295), .A2(G264), .A3(G1698), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n295), .A2(G257), .A3(new_n297), .ZN(new_n555));
  INV_X1    g0355(.A(G303), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n554), .B(new_n555), .C1(new_n556), .C2(new_n295), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(new_n294), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n291), .A2(new_n484), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n498), .A2(G270), .A3(new_n284), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(new_n561), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n302), .B1(new_n558), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n553), .A2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT21), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n558), .A2(new_n562), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n567), .A2(new_n304), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(new_n553), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n553), .A2(new_n563), .A3(KEYINPUT21), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n534), .A2(new_n566), .A3(new_n569), .A4(new_n570), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n391), .A2(new_n393), .A3(G244), .A4(new_n297), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT4), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n295), .A2(KEYINPUT4), .A3(G244), .A4(new_n297), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n295), .A2(G250), .A3(G1698), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n574), .A2(new_n575), .A3(new_n547), .A4(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n294), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n485), .A2(G257), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n578), .A2(new_n559), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(new_n462), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n581), .B1(G190), .B2(new_n580), .ZN(new_n582));
  OAI21_X1  g0382(.A(G107), .B1(new_n418), .B2(new_n420), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(KEYINPUT84), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n419), .A2(new_n411), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(KEYINPUT80), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n586), .A2(new_n417), .A3(new_n416), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT84), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n587), .A2(new_n588), .A3(G107), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n265), .A2(G77), .ZN(new_n590));
  XNOR2_X1  g0390(.A(KEYINPUT83), .B(G97), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n207), .A2(KEYINPUT6), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(G97), .A2(G107), .ZN(new_n594));
  AOI21_X1  g0394(.A(KEYINPUT6), .B1(new_n208), .B2(new_n594), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n590), .B1(new_n596), .B2(new_n233), .ZN(new_n597));
  INV_X1    g0397(.A(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n584), .A2(new_n589), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(new_n273), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n275), .A2(G97), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n527), .A2(new_n528), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n601), .B1(new_n602), .B2(G97), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n582), .A2(new_n600), .A3(new_n603), .ZN(new_n604));
  AOI22_X1  g0404(.A1(new_n577), .A2(new_n294), .B1(G257), .B2(new_n485), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n605), .A2(new_n304), .A3(new_n559), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n580), .A2(new_n302), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n597), .B1(new_n583), .B2(KEYINPUT84), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n377), .B1(new_n608), .B2(new_n589), .ZN(new_n609));
  INV_X1    g0409(.A(new_n603), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n606), .B(new_n607), .C1(new_n609), .C2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n604), .A2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(new_n551), .ZN(new_n613));
  INV_X1    g0413(.A(new_n552), .ZN(new_n614));
  AOI22_X1  g0414(.A1(new_n613), .A2(new_n614), .B1(new_n541), .B2(new_n539), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n567), .A2(G200), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n561), .B1(new_n294), .B2(new_n557), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(G190), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n615), .A2(new_n616), .A3(new_n537), .A4(new_n618), .ZN(new_n619));
  AND3_X1   g0419(.A1(new_n510), .A2(new_n518), .A3(new_n521), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n521), .B1(new_n510), .B2(new_n518), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n273), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(G200), .B1(new_n494), .B2(new_n503), .ZN(new_n623));
  AND3_X1   g0423(.A1(new_n486), .A2(new_n312), .A3(new_n491), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n622), .B(new_n532), .C1(new_n623), .C2(new_n624), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n391), .A2(new_n393), .A3(G238), .A4(new_n297), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n391), .A2(new_n393), .A3(G244), .A4(G1698), .ZN(new_n627));
  OAI211_X1 g0427(.A(new_n626), .B(new_n627), .C1(new_n392), .C2(new_n535), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(new_n294), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n480), .A2(G250), .ZN(new_n630));
  OAI22_X1  g0430(.A1(new_n334), .A2(new_n480), .B1(new_n285), .B2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n629), .A2(new_n304), .A3(new_n632), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n631), .B1(new_n628), .B2(new_n294), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n295), .A2(new_n233), .A3(G68), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n591), .A2(new_n262), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n635), .B1(new_n636), .B2(KEYINPUT19), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n327), .A2(KEYINPUT19), .A3(new_n328), .ZN(new_n638));
  NOR2_X1   g0438(.A1(G87), .A2(G107), .ZN(new_n639));
  AOI22_X1  g0439(.A1(new_n638), .A2(new_n233), .B1(new_n591), .B2(new_n639), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n273), .B1(new_n637), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n382), .A2(new_n276), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n382), .B1(new_n527), .B2(new_n528), .ZN(new_n644));
  OAI221_X1 g0444(.A(new_n633), .B1(G169), .B2(new_n634), .C1(new_n643), .C2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n643), .ZN(new_n646));
  INV_X1    g0446(.A(new_n634), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(G200), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n602), .A2(G87), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n629), .A2(G190), .A3(new_n632), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n646), .A2(new_n648), .A3(new_n649), .A4(new_n650), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n619), .A2(new_n625), .A3(new_n645), .A4(new_n651), .ZN(new_n652));
  NOR4_X1   g0452(.A1(new_n479), .A2(new_n571), .A3(new_n612), .A4(new_n652), .ZN(G372));
  AND3_X1   g0453(.A1(new_n370), .A2(new_n371), .A3(new_n372), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n369), .B1(new_n654), .B2(new_n401), .ZN(new_n655));
  AND2_X1   g0455(.A1(new_n464), .A2(new_n474), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n454), .A2(new_n476), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n316), .A2(new_n318), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n307), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  AND3_X1   g0462(.A1(new_n625), .A2(new_n645), .A3(new_n651), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n663), .A2(new_n571), .A3(new_n611), .A4(new_n604), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n610), .B1(new_n599), .B2(new_n273), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n607), .A2(new_n606), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n643), .A2(new_n644), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n633), .B1(G169), .B2(new_n634), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n650), .B1(new_n462), .B2(new_n634), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n649), .A2(new_n641), .A3(new_n642), .ZN(new_n671));
  OAI22_X1  g0471(.A1(new_n668), .A2(new_n669), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  AOI21_X1  g0473(.A(KEYINPUT26), .B1(new_n667), .B2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT26), .ZN(new_n675));
  NOR4_X1   g0475(.A1(new_n665), .A2(new_n672), .A3(new_n675), .A4(new_n666), .ZN(new_n676));
  OAI211_X1 g0476(.A(new_n664), .B(new_n645), .C1(new_n674), .C2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n478), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n662), .A2(new_n678), .ZN(G369));
  INV_X1    g0479(.A(new_n619), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n566), .A2(new_n569), .A3(new_n570), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n541), .A2(new_n233), .ZN(new_n682));
  OR2_X1    g0482(.A1(new_n682), .A2(KEYINPUT27), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(KEYINPUT27), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n683), .A2(G213), .A3(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(G343), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n681), .A2(new_n553), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n553), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n566), .A2(new_n569), .A3(new_n570), .A4(new_n690), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n680), .B1(new_n689), .B2(new_n691), .ZN(new_n692));
  AOI21_X1  g0492(.A(KEYINPUT88), .B1(new_n692), .B2(G330), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n692), .A2(KEYINPUT88), .A3(G330), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n534), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n688), .B1(new_n523), .B2(new_n533), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n697), .B1(new_n625), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n697), .A2(new_n687), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n696), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n681), .A2(new_n687), .ZN(new_n704));
  OR2_X1    g0504(.A1(new_n704), .A2(KEYINPUT89), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(KEYINPUT89), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n701), .B1(new_n707), .B2(new_n702), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n703), .A2(new_n708), .ZN(G399));
  INV_X1    g0509(.A(new_n225), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n710), .A2(G41), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(G1), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n591), .A2(new_n535), .A3(new_n639), .ZN(new_n714));
  OAI22_X1  g0514(.A1(new_n713), .A2(new_n714), .B1(new_n237), .B2(new_n712), .ZN(new_n715));
  XOR2_X1   g0515(.A(KEYINPUT90), .B(KEYINPUT28), .Z(new_n716));
  XNOR2_X1  g0516(.A(new_n715), .B(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(G330), .ZN(new_n718));
  AND2_X1   g0518(.A1(new_n605), .A2(new_n634), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n494), .A2(new_n503), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n719), .A2(new_n568), .A3(KEYINPUT30), .A4(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT30), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n617), .A2(G179), .A3(new_n503), .A4(new_n494), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n605), .A2(new_n634), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n723), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NOR3_X1   g0526(.A1(new_n617), .A2(G179), .A3(new_n634), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n727), .A2(new_n720), .A3(new_n580), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n722), .A2(new_n726), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(new_n688), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT31), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n729), .A2(KEYINPUT31), .A3(new_n688), .ZN(new_n733));
  AND2_X1   g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n612), .A2(new_n652), .ZN(new_n735));
  INV_X1    g0535(.A(new_n571), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n735), .A2(new_n736), .A3(new_n687), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n718), .B1(new_n734), .B2(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n677), .A2(new_n687), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT29), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n739), .B1(KEYINPUT91), .B2(new_n740), .ZN(new_n741));
  AND2_X1   g0541(.A1(new_n740), .A2(KEYINPUT91), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n740), .A2(KEYINPUT91), .ZN(new_n743));
  OAI211_X1 g0543(.A(new_n677), .B(new_n687), .C1(new_n742), .C2(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n738), .B1(new_n741), .B2(new_n744), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n717), .B1(new_n745), .B2(G1), .ZN(G364));
  INV_X1    g0546(.A(new_n696), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n540), .A2(G20), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n274), .B1(new_n748), .B2(G45), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n711), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  OAI211_X1 g0552(.A(new_n747), .B(new_n752), .C1(G330), .C2(new_n692), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n232), .B1(G20), .B2(new_n302), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n233), .A2(G179), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n755), .A2(G190), .A3(G200), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n394), .B1(new_n756), .B2(new_n556), .ZN(new_n757));
  XNOR2_X1  g0557(.A(new_n757), .B(KEYINPUT93), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n233), .A2(new_n304), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NOR3_X1   g0560(.A1(new_n760), .A2(new_n312), .A3(G200), .ZN(new_n761));
  NOR2_X1   g0561(.A1(G190), .A2(G200), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n759), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  AOI22_X1  g0564(.A1(new_n761), .A2(G322), .B1(G311), .B2(new_n764), .ZN(new_n765));
  NOR3_X1   g0565(.A1(new_n760), .A2(new_n312), .A3(new_n462), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n755), .A2(new_n762), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  AOI22_X1  g0568(.A1(new_n766), .A2(G326), .B1(G329), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n765), .A2(new_n769), .ZN(new_n770));
  NOR3_X1   g0570(.A1(new_n312), .A2(G179), .A3(G200), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(new_n233), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n770), .B1(G294), .B2(new_n773), .ZN(new_n774));
  NOR3_X1   g0574(.A1(new_n760), .A2(new_n462), .A3(G190), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  XNOR2_X1  g0576(.A(KEYINPUT33), .B(G317), .ZN(new_n777));
  XNOR2_X1  g0577(.A(new_n777), .B(KEYINPUT94), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n774), .B1(new_n776), .B2(new_n778), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n755), .A2(new_n312), .A3(G200), .ZN(new_n780));
  INV_X1    g0580(.A(KEYINPUT92), .ZN(new_n781));
  OR2_X1    g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n780), .A2(new_n781), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  AOI211_X1 g0585(.A(new_n758), .B(new_n779), .C1(G283), .C2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(KEYINPUT32), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n768), .A2(new_n787), .A3(G159), .ZN(new_n788));
  OAI221_X1 g0588(.A(new_n788), .B1(new_n214), .B2(new_n756), .C1(new_n206), .C2(new_n772), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n787), .B1(new_n768), .B2(G159), .ZN(new_n790));
  AOI211_X1 g0590(.A(new_n394), .B(new_n790), .C1(G68), .C2(new_n775), .ZN(new_n791));
  AOI22_X1  g0591(.A1(new_n761), .A2(G58), .B1(new_n766), .B2(G50), .ZN(new_n792));
  OAI211_X1 g0592(.A(new_n791), .B(new_n792), .C1(new_n352), .C2(new_n763), .ZN(new_n793));
  AOI211_X1 g0593(.A(new_n789), .B(new_n793), .C1(G107), .C2(new_n785), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n754), .B1(new_n786), .B2(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n710), .A2(new_n394), .ZN(new_n796));
  AOI22_X1  g0596(.A1(new_n796), .A2(G355), .B1(new_n535), .B2(new_n710), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n258), .A2(new_n287), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n710), .A2(new_n295), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n799), .B1(G45), .B2(new_n237), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n797), .B1(new_n798), .B2(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(G13), .A2(G33), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n803), .A2(G20), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n754), .A2(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n752), .B1(new_n801), .B2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n804), .ZN(new_n807));
  OAI211_X1 g0607(.A(new_n795), .B(new_n806), .C1(new_n692), .C2(new_n807), .ZN(new_n808));
  AND2_X1   g0608(.A1(new_n753), .A2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(G396));
  INV_X1    g0610(.A(KEYINPUT99), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n387), .A2(new_n811), .A3(new_n688), .ZN(new_n812));
  OAI21_X1  g0612(.A(KEYINPUT99), .B1(new_n402), .B2(new_n687), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n401), .A2(KEYINPUT98), .ZN(new_n815));
  INV_X1    g0615(.A(KEYINPUT98), .ZN(new_n816));
  NAND4_X1  g0616(.A1(new_n387), .A2(new_n399), .A3(new_n816), .A4(new_n400), .ZN(new_n817));
  NAND4_X1  g0617(.A1(new_n814), .A2(new_n815), .A3(new_n404), .A4(new_n817), .ZN(new_n818));
  OR2_X1    g0618(.A1(new_n401), .A2(new_n687), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  MUX2_X1   g0620(.A(new_n818), .B(new_n820), .S(new_n739), .Z(new_n821));
  INV_X1    g0621(.A(new_n738), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n751), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n823), .B1(new_n822), .B2(new_n821), .ZN(new_n824));
  INV_X1    g0624(.A(G283), .ZN(new_n825));
  INV_X1    g0625(.A(new_n761), .ZN(new_n826));
  OAI22_X1  g0626(.A1(new_n825), .A2(new_n776), .B1(new_n826), .B2(new_n489), .ZN(new_n827));
  INV_X1    g0627(.A(new_n766), .ZN(new_n828));
  INV_X1    g0628(.A(G311), .ZN(new_n829));
  OAI22_X1  g0629(.A1(new_n828), .A2(new_n556), .B1(new_n767), .B2(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n827), .A2(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n394), .B1(new_n763), .B2(new_n535), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n832), .B1(G97), .B2(new_n773), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n785), .A2(G87), .ZN(new_n834));
  INV_X1    g0634(.A(new_n756), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n835), .A2(G107), .ZN(new_n836));
  NAND4_X1  g0636(.A1(new_n831), .A2(new_n833), .A3(new_n834), .A4(new_n836), .ZN(new_n837));
  XOR2_X1   g0637(.A(KEYINPUT96), .B(G143), .Z(new_n838));
  AOI22_X1  g0638(.A1(new_n838), .A2(new_n761), .B1(new_n766), .B2(G137), .ZN(new_n839));
  INV_X1    g0639(.A(G150), .ZN(new_n840));
  INV_X1    g0640(.A(G159), .ZN(new_n841));
  OAI221_X1 g0641(.A(new_n839), .B1(new_n840), .B2(new_n776), .C1(new_n841), .C2(new_n763), .ZN(new_n842));
  XNOR2_X1  g0642(.A(KEYINPUT97), .B(KEYINPUT34), .ZN(new_n843));
  XNOR2_X1  g0643(.A(new_n842), .B(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(G132), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n295), .B1(new_n767), .B2(new_n845), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n846), .B1(G50), .B2(new_n835), .ZN(new_n847));
  OAI221_X1 g0647(.A(new_n847), .B1(new_n422), .B2(new_n772), .C1(new_n784), .C2(new_n212), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n837), .B1(new_n844), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n849), .A2(new_n754), .ZN(new_n850));
  INV_X1    g0650(.A(new_n754), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n851), .A2(new_n803), .ZN(new_n852));
  XOR2_X1   g0652(.A(new_n852), .B(KEYINPUT95), .Z(new_n853));
  OAI221_X1 g0653(.A(new_n850), .B1(G77), .B2(new_n853), .C1(new_n820), .C2(new_n803), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(new_n751), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n824), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(KEYINPUT100), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT100), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n824), .A2(new_n858), .A3(new_n855), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(G384));
  NOR2_X1   g0661(.A1(new_n748), .A2(new_n274), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT40), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n426), .B1(new_n587), .B2(G68), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n471), .B1(new_n864), .B2(KEYINPUT16), .ZN(new_n865));
  OAI211_X1 g0665(.A(new_n865), .B(new_n409), .C1(new_n473), .C2(new_n457), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n435), .A2(new_n686), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n866), .A2(new_n453), .A3(new_n867), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n868), .A2(KEYINPUT37), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n461), .A2(new_n462), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n435), .B1(new_n870), .B2(new_n456), .ZN(new_n871));
  AOI21_X1  g0671(.A(G169), .B1(new_n460), .B2(new_n444), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n432), .A2(new_n433), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n465), .B1(new_n471), .B2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n452), .ZN(new_n875));
  NOR3_X1   g0675(.A1(new_n872), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  OAI21_X1  g0676(.A(KEYINPUT102), .B1(new_n871), .B2(new_n876), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n470), .A2(KEYINPUT16), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n409), .B1(new_n434), .B2(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n451), .A2(new_n879), .A3(new_n452), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT102), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n866), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n874), .A2(new_n685), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n877), .A2(new_n882), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n869), .B1(new_n885), .B2(KEYINPUT37), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n477), .A2(new_n883), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(KEYINPUT38), .ZN(new_n888));
  OAI21_X1  g0688(.A(KEYINPUT103), .B1(new_n886), .B2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT103), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT38), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n891), .B1(new_n477), .B2(new_n883), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT37), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n866), .A2(new_n880), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n883), .B1(new_n894), .B2(KEYINPUT102), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n893), .B1(new_n895), .B2(new_n882), .ZN(new_n896));
  OAI211_X1 g0696(.A(new_n890), .B(new_n892), .C1(new_n896), .C2(new_n869), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n887), .B1(new_n896), .B2(new_n869), .ZN(new_n898));
  AOI22_X1  g0698(.A1(new_n889), .A2(new_n897), .B1(new_n891), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n368), .A2(new_n688), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n369), .A2(new_n373), .A3(new_n900), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n368), .B(new_n688), .C1(new_n654), .C2(new_n350), .ZN(new_n902));
  AOI22_X1  g0702(.A1(new_n901), .A2(new_n902), .B1(new_n818), .B2(new_n819), .ZN(new_n903));
  NOR4_X1   g0703(.A1(new_n612), .A2(new_n571), .A3(new_n652), .A4(new_n688), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n732), .A2(new_n733), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n903), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT104), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n734), .A2(new_n737), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n909), .A2(KEYINPUT104), .A3(new_n903), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n863), .B1(new_n899), .B2(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n909), .A2(KEYINPUT40), .A3(new_n903), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n867), .B1(new_n659), .B2(new_n656), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n868), .B(new_n893), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n891), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n892), .B1(new_n896), .B2(new_n869), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n914), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n912), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n909), .A2(new_n478), .ZN(new_n922));
  AND2_X1   g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n921), .A2(new_n922), .ZN(new_n924));
  NOR3_X1   g0724(.A1(new_n923), .A2(new_n924), .A3(new_n718), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n889), .A2(new_n897), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n898), .A2(new_n891), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(new_n818), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n677), .A2(new_n687), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n815), .A2(new_n817), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(new_n687), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n901), .A2(new_n902), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(KEYINPUT101), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT101), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n934), .A2(new_n938), .A3(new_n935), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n929), .A2(new_n937), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n658), .A2(new_n685), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT39), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n917), .A2(new_n918), .A3(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(new_n943), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n944), .B1(new_n929), .B2(KEYINPUT39), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n369), .A2(new_n688), .ZN(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  OAI211_X1 g0747(.A(new_n940), .B(new_n941), .C1(new_n945), .C2(new_n947), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n741), .A2(new_n478), .A3(new_n744), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n949), .A2(new_n662), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n948), .B(new_n950), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n862), .B1(new_n926), .B2(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n952), .B1(new_n951), .B2(new_n926), .ZN(new_n953));
  INV_X1    g0753(.A(new_n596), .ZN(new_n954));
  AOI211_X1 g0754(.A(new_n535), .B(new_n235), .C1(new_n954), .C2(KEYINPUT35), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(KEYINPUT35), .B2(new_n954), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n956), .B(KEYINPUT36), .ZN(new_n957));
  OAI21_X1  g0757(.A(G77), .B1(new_n422), .B2(new_n212), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n254), .B1(new_n237), .B2(new_n958), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n959), .A2(G1), .A3(new_n540), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n953), .A2(new_n957), .A3(new_n960), .ZN(G367));
  INV_X1    g0761(.A(new_n799), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n249), .A2(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n805), .B1(new_n225), .B2(new_n382), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n751), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  OAI221_X1 g0765(.A(new_n394), .B1(new_n207), .B2(new_n772), .C1(new_n826), .C2(new_n556), .ZN(new_n966));
  OAI22_X1  g0766(.A1(new_n828), .A2(new_n829), .B1(new_n763), .B2(new_n825), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n768), .A2(G317), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n776), .B2(new_n489), .ZN(new_n969));
  NOR3_X1   g0769(.A1(new_n966), .A2(new_n967), .A3(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT109), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n971), .B1(new_n756), .B2(new_n535), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n970), .B1(KEYINPUT46), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(KEYINPUT46), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n974), .B1(new_n784), .B2(new_n591), .ZN(new_n975));
  AOI22_X1  g0775(.A1(new_n775), .A2(G159), .B1(G50), .B2(new_n764), .ZN(new_n976));
  XOR2_X1   g0776(.A(new_n976), .B(KEYINPUT110), .Z(new_n977));
  NAND2_X1  g0777(.A1(new_n785), .A2(G77), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n394), .B1(new_n768), .B2(G137), .ZN(new_n979));
  AOI22_X1  g0779(.A1(new_n838), .A2(new_n766), .B1(new_n761), .B2(G150), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n772), .A2(new_n212), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n981), .B1(G58), .B2(new_n835), .ZN(new_n982));
  NAND4_X1  g0782(.A1(new_n978), .A2(new_n979), .A3(new_n980), .A4(new_n982), .ZN(new_n983));
  OAI22_X1  g0783(.A1(new_n973), .A2(new_n975), .B1(new_n977), .B2(new_n983), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n984), .B(KEYINPUT47), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n965), .B1(new_n985), .B2(new_n754), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n671), .A2(new_n688), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT105), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n988), .A2(new_n645), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n989), .B1(new_n673), .B2(new_n988), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(new_n804), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n986), .A2(new_n991), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n749), .B(KEYINPUT108), .ZN(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT45), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n707), .A2(new_n702), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n996), .A2(new_n700), .ZN(new_n997));
  OAI211_X1 g0797(.A(new_n604), .B(new_n611), .C1(new_n665), .C2(new_n687), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n667), .A2(new_n688), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n1000), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n995), .B1(new_n997), .B2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n708), .A2(KEYINPUT45), .A3(new_n1000), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n997), .A2(KEYINPUT44), .A3(new_n1001), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT44), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1006), .B1(new_n708), .B2(new_n1000), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1004), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n703), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n702), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1012), .A2(new_n705), .A3(new_n706), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1013), .A2(new_n996), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n695), .ZN(new_n1016));
  OAI21_X1  g0816(.A(KEYINPUT106), .B1(new_n1016), .B2(new_n693), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT106), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n694), .A2(new_n1018), .A3(new_n695), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1015), .A2(new_n1017), .A3(new_n1019), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n696), .A2(new_n1014), .A3(KEYINPUT106), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1022), .A2(KEYINPUT107), .A3(new_n745), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1004), .A2(new_n1008), .A3(new_n703), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1011), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(KEYINPUT107), .B1(new_n1022), .B2(new_n745), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n745), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  XOR2_X1   g0827(.A(new_n711), .B(KEYINPUT41), .Z(new_n1028));
  INV_X1    g0828(.A(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n994), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT43), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n990), .A2(new_n1031), .ZN(new_n1032));
  OR2_X1    g0832(.A1(new_n998), .A2(new_n534), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n688), .B1(new_n1033), .B2(new_n611), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n707), .A2(new_n702), .A3(new_n1000), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1034), .B1(new_n1035), .B2(KEYINPUT42), .ZN(new_n1036));
  OR2_X1    g0836(.A1(new_n1035), .A2(KEYINPUT42), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1032), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n990), .A2(new_n1031), .ZN(new_n1039));
  OR2_X1    g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(new_n703), .B2(new_n1001), .ZN(new_n1043));
  NAND4_X1  g0843(.A1(new_n1040), .A2(new_n1010), .A3(new_n1000), .A4(new_n1041), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n992), .B1(new_n1030), .B2(new_n1045), .ZN(G387));
  NAND2_X1  g0846(.A1(new_n1022), .A2(new_n994), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n828), .A2(new_n841), .B1(new_n767), .B2(new_n840), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1048), .B1(G68), .B2(new_n764), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n295), .B1(new_n826), .B2(new_n202), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1050), .B1(G77), .B2(new_n835), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n785), .A2(G97), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n261), .A2(new_n775), .B1(new_n773), .B2(new_n383), .ZN(new_n1053));
  NAND4_X1  g0853(.A1(new_n1049), .A2(new_n1051), .A3(new_n1052), .A4(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n295), .B1(new_n768), .B2(G326), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n772), .A2(new_n825), .B1(new_n756), .B2(new_n489), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n761), .A2(G317), .B1(new_n766), .B2(G322), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n1057), .B1(new_n556), .B2(new_n763), .C1(new_n829), .C2(new_n776), .ZN(new_n1058));
  INV_X1    g0858(.A(KEYINPUT48), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1056), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1060), .B1(new_n1059), .B2(new_n1058), .ZN(new_n1061));
  INV_X1    g0861(.A(KEYINPUT49), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n1055), .B1(new_n535), .B2(new_n784), .C1(new_n1061), .C2(new_n1062), .ZN(new_n1063));
  AND2_X1   g0863(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1054), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1065), .A2(new_n754), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n796), .A2(new_n714), .B1(new_n207), .B2(new_n710), .ZN(new_n1067));
  AND2_X1   g0867(.A1(new_n379), .A2(new_n380), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1068), .A2(new_n202), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n1069), .B(KEYINPUT50), .ZN(new_n1070));
  AOI211_X1 g0870(.A(G45), .B(new_n714), .C1(G68), .C2(G77), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT111), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n1070), .A2(new_n1072), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n799), .B1(new_n245), .B2(new_n287), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1067), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n752), .B1(new_n1075), .B2(new_n805), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n1066), .B(new_n1076), .C1(new_n702), .C2(new_n807), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1022), .A2(new_n745), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1078), .A2(new_n711), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n1022), .A2(new_n745), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n1047), .B(new_n1077), .C1(new_n1079), .C2(new_n1080), .ZN(G393));
  INV_X1    g0881(.A(KEYINPUT107), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1078), .A2(new_n1082), .ZN(new_n1083));
  NAND4_X1  g0883(.A1(new_n1083), .A2(new_n1023), .A3(new_n1011), .A4(new_n1024), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1024), .A2(KEYINPUT112), .ZN(new_n1085));
  XOR2_X1   g0885(.A(new_n1085), .B(new_n1011), .Z(new_n1086));
  INV_X1    g0886(.A(new_n1078), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n711), .B(new_n1084), .C1(new_n1086), .C2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1001), .A2(new_n804), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n805), .B1(new_n225), .B2(new_n591), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n253), .A2(new_n962), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n751), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n761), .A2(G159), .B1(new_n766), .B2(G150), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(KEYINPUT113), .B(KEYINPUT51), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(new_n1093), .B(new_n1094), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1068), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1095), .B1(new_n1096), .B2(new_n763), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n768), .A2(new_n838), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n394), .B1(new_n775), .B2(G50), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n772), .A2(new_n352), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1100), .B1(G68), .B2(new_n835), .ZN(new_n1101));
  NAND4_X1  g0901(.A1(new_n834), .A2(new_n1098), .A3(new_n1099), .A4(new_n1101), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n761), .A2(G311), .B1(new_n766), .B2(G317), .ZN(new_n1103));
  XNOR2_X1  g0903(.A(new_n1103), .B(KEYINPUT52), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n785), .A2(G107), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n295), .B1(new_n764), .B2(G294), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n775), .A2(G303), .B1(G322), .B2(new_n768), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n773), .A2(G116), .B1(new_n835), .B2(G283), .ZN(new_n1108));
  NAND4_X1  g0908(.A1(new_n1105), .A2(new_n1106), .A3(new_n1107), .A4(new_n1108), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n1097), .A2(new_n1102), .B1(new_n1104), .B2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1092), .B1(new_n1110), .B2(new_n754), .ZN(new_n1111));
  XOR2_X1   g0911(.A(new_n1111), .B(KEYINPUT114), .Z(new_n1112));
  AOI22_X1  g0912(.A1(new_n1086), .A2(new_n994), .B1(new_n1089), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1088), .A2(new_n1113), .ZN(G390));
  NAND2_X1  g0914(.A1(new_n936), .A2(new_n947), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n1115), .B(new_n943), .C1(new_n942), .C2(new_n899), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n936), .A2(new_n947), .A3(new_n919), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n738), .A2(new_n820), .A3(new_n935), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1116), .A2(new_n1119), .A3(new_n1117), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n738), .A2(new_n478), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n949), .A2(new_n662), .A3(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n935), .B1(new_n738), .B2(new_n820), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n934), .B1(new_n1120), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n738), .A2(new_n820), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n935), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n1130), .A2(new_n931), .A3(new_n933), .A4(new_n1119), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1125), .B1(new_n1127), .B2(new_n1131), .ZN(new_n1132));
  OR2_X1    g0932(.A1(new_n1132), .A2(KEYINPUT115), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(KEYINPUT115), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1123), .A2(new_n1133), .A3(new_n1134), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1121), .A2(new_n1122), .A3(new_n1132), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1135), .A2(new_n711), .A3(new_n1136), .ZN(new_n1137));
  AND3_X1   g0937(.A1(new_n1116), .A2(new_n1119), .A3(new_n1117), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1119), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n945), .A2(new_n802), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n751), .B1(new_n853), .B2(new_n261), .ZN(new_n1142));
  OAI22_X1  g0942(.A1(new_n826), .A2(new_n535), .B1(new_n828), .B2(new_n825), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n776), .A2(new_n207), .B1(new_n591), .B2(new_n763), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n394), .B1(new_n767), .B2(new_n489), .ZN(new_n1146));
  AOI211_X1 g0946(.A(new_n1146), .B(new_n1100), .C1(G87), .C2(new_n835), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n1145), .B(new_n1147), .C1(new_n212), .C2(new_n784), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n756), .A2(new_n840), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(new_n1149), .B(KEYINPUT53), .ZN(new_n1150));
  AND2_X1   g0950(.A1(new_n775), .A2(G137), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(G125), .B2(new_n768), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(new_n761), .A2(G132), .B1(new_n766), .B2(G128), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(KEYINPUT54), .B(G143), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n295), .B1(new_n763), .B2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1155), .B1(G159), .B2(new_n773), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n1150), .A2(new_n1152), .A3(new_n1153), .A4(new_n1156), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n784), .A2(new_n202), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1148), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1142), .B1(new_n1159), .B2(new_n754), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(new_n1140), .A2(new_n994), .B1(new_n1141), .B2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1137), .A2(new_n1161), .ZN(G378));
  INV_X1    g0962(.A(KEYINPUT120), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n943), .B1(new_n899), .B2(new_n942), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(new_n1164), .A2(new_n946), .B1(new_n658), .B2(new_n685), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1163), .B1(new_n1165), .B2(new_n940), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n718), .B1(new_n914), .B2(new_n919), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n912), .A2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n282), .A2(new_n686), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(new_n1169), .B(KEYINPUT118), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(KEYINPUT117), .B1(new_n661), .B2(new_n306), .ZN(new_n1172));
  INV_X1    g0972(.A(KEYINPUT117), .ZN(new_n1173));
  AOI211_X1 g0973(.A(new_n1173), .B(new_n307), .C1(new_n316), .C2(new_n318), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1171), .B1(new_n1172), .B2(new_n1174), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n318), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n317), .B1(new_n311), .B2(new_n314), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n306), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1179), .A2(new_n1173), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n319), .A2(KEYINPUT117), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1180), .A2(new_n1181), .A3(new_n1170), .ZN(new_n1182));
  AND3_X1   g0982(.A1(new_n1175), .A2(new_n1176), .A3(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1176), .B1(new_n1175), .B2(new_n1182), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1168), .A2(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(KEYINPUT119), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1188), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1176), .ZN(new_n1190));
  NOR3_X1   g0990(.A1(new_n1172), .A2(new_n1174), .A3(new_n1171), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1170), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1190), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1175), .A2(new_n1182), .A3(new_n1176), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1193), .A2(KEYINPUT119), .A3(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1189), .A2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n912), .A2(new_n1167), .A3(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1187), .A2(new_n1197), .ZN(new_n1198));
  XNOR2_X1  g0998(.A(new_n1166), .B(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1199), .A2(new_n994), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1189), .A2(new_n802), .A3(new_n1195), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n751), .B1(new_n852), .B2(G50), .ZN(new_n1202));
  XNOR2_X1  g1002(.A(new_n1202), .B(KEYINPUT116), .ZN(new_n1203));
  OAI211_X1 g1003(.A(new_n286), .B(new_n394), .C1(new_n767), .C2(new_n825), .ZN(new_n1204));
  AOI211_X1 g1004(.A(new_n1204), .B(new_n981), .C1(G77), .C2(new_n835), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n785), .A2(G58), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(new_n761), .A2(G107), .B1(new_n383), .B2(new_n764), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n775), .A2(G97), .B1(new_n766), .B2(G116), .ZN(new_n1208));
  NAND4_X1  g1008(.A1(new_n1205), .A2(new_n1206), .A3(new_n1207), .A4(new_n1208), .ZN(new_n1209));
  XNOR2_X1  g1009(.A(new_n1209), .B(KEYINPUT58), .ZN(new_n1210));
  AOI21_X1  g1010(.A(G50), .B1(new_n392), .B2(new_n286), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1211), .B1(new_n295), .B2(G41), .ZN(new_n1212));
  AOI211_X1 g1012(.A(G33), .B(G41), .C1(new_n768), .C2(G124), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n775), .A2(G132), .B1(new_n766), .B2(G125), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n761), .A2(G128), .B1(G137), .B2(new_n764), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n772), .A2(new_n840), .B1(new_n756), .B2(new_n1154), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT59), .ZN(new_n1219));
  OAI221_X1 g1019(.A(new_n1213), .B1(new_n841), .B2(new_n784), .C1(new_n1218), .C2(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1218), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n1221), .A2(KEYINPUT59), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n1210), .B(new_n1212), .C1(new_n1220), .C2(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1203), .B1(new_n1223), .B2(new_n754), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1201), .A2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1200), .A2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1127), .A2(new_n1131), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1125), .B1(new_n1140), .B2(new_n1227), .ZN(new_n1228));
  AND3_X1   g1028(.A1(new_n912), .A2(new_n1167), .A3(new_n1196), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1185), .B1(new_n912), .B2(new_n1167), .ZN(new_n1230));
  OAI211_X1 g1030(.A(new_n940), .B(new_n1165), .C1(new_n1229), .C2(new_n1230), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n948), .A2(new_n1187), .A3(new_n1197), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1231), .A2(new_n1232), .A3(KEYINPUT57), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n711), .B1(new_n1228), .B2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT121), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1125), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1136), .A2(new_n1236), .ZN(new_n1237));
  AND2_X1   g1037(.A1(new_n1166), .A2(new_n1198), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1166), .A2(new_n1198), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1237), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT57), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(new_n1234), .A2(new_n1235), .B1(new_n1240), .B2(new_n1241), .ZN(new_n1242));
  OAI211_X1 g1042(.A(KEYINPUT121), .B(new_n711), .C1(new_n1228), .C2(new_n1233), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1226), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  XNOR2_X1  g1044(.A(new_n1244), .B(KEYINPUT122), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(G375));
  NAND3_X1  g1046(.A1(new_n1127), .A2(new_n1131), .A3(new_n1125), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(new_n1133), .A2(new_n1029), .A3(new_n1134), .A4(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1227), .A2(new_n994), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n751), .B1(new_n853), .B2(G68), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n756), .A2(new_n841), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n295), .B1(new_n763), .B2(new_n840), .ZN(new_n1252));
  AOI211_X1 g1052(.A(new_n1251), .B(new_n1252), .C1(G50), .C2(new_n773), .ZN(new_n1253));
  AOI22_X1  g1053(.A1(new_n766), .A2(G132), .B1(G128), .B2(new_n768), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1154), .ZN(new_n1255));
  AOI22_X1  g1055(.A1(new_n1255), .A2(new_n775), .B1(new_n761), .B2(G137), .ZN(new_n1256));
  NAND4_X1  g1056(.A1(new_n1206), .A2(new_n1253), .A3(new_n1254), .A4(new_n1256), .ZN(new_n1257));
  OAI22_X1  g1057(.A1(new_n776), .A2(new_n535), .B1(new_n828), .B2(new_n489), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1258), .B1(G283), .B2(new_n761), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n773), .A2(new_n383), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n295), .B1(new_n764), .B2(G107), .ZN(new_n1261));
  NAND4_X1  g1061(.A1(new_n1259), .A2(new_n978), .A3(new_n1260), .A4(new_n1261), .ZN(new_n1262));
  OAI22_X1  g1062(.A1(new_n756), .A2(new_n206), .B1(new_n767), .B2(new_n556), .ZN(new_n1263));
  XNOR2_X1  g1063(.A(new_n1263), .B(KEYINPUT123), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1257), .B1(new_n1262), .B2(new_n1264), .ZN(new_n1265));
  OR2_X1    g1065(.A1(new_n1265), .A2(KEYINPUT124), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n851), .B1(new_n1265), .B2(KEYINPUT124), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1250), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1268), .B1(new_n935), .B2(new_n803), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1249), .A2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1248), .A2(new_n1271), .ZN(G381));
  INV_X1    g1072(.A(G378), .ZN(new_n1273));
  OR3_X1    g1073(.A1(G384), .A2(G396), .A3(G393), .ZN(new_n1274));
  NOR4_X1   g1074(.A1(new_n1274), .A2(G390), .A3(G387), .A4(G381), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1245), .A2(new_n1273), .A3(new_n1275), .ZN(G407));
  NAND2_X1  g1076(.A1(new_n1245), .A2(new_n1273), .ZN(new_n1277));
  OAI211_X1 g1077(.A(G407), .B(G213), .C1(new_n1277), .C2(G343), .ZN(G409));
  INV_X1    g1078(.A(G390), .ZN(new_n1279));
  XNOR2_X1  g1079(.A(G393), .B(new_n809), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT126), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1280), .B1(G387), .B2(new_n1281), .ZN(new_n1282));
  XNOR2_X1  g1082(.A(G393), .B(G396), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1028), .B1(new_n1084), .B2(new_n745), .ZN(new_n1284));
  OAI211_X1 g1084(.A(new_n1044), .B(new_n1043), .C1(new_n1284), .C2(new_n994), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1283), .B1(new_n1285), .B2(new_n992), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1279), .B1(new_n1282), .B2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(G387), .A2(new_n1280), .ZN(new_n1288));
  AOI21_X1  g1088(.A(KEYINPUT126), .B1(new_n1285), .B2(new_n992), .ZN(new_n1289));
  OAI211_X1 g1089(.A(new_n1288), .B(G390), .C1(new_n1289), .C2(new_n1280), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1287), .A2(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(G213), .ZN(new_n1293));
  NOR2_X1   g1093(.A1(new_n1293), .A2(G343), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1294), .A2(G2897), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT60), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1247), .B1(new_n1132), .B2(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1297), .A2(new_n711), .ZN(new_n1298));
  NOR3_X1   g1098(.A1(new_n1227), .A2(new_n1236), .A3(new_n1296), .ZN(new_n1299));
  OAI21_X1  g1099(.A(KEYINPUT125), .B1(new_n1298), .B2(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1299), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT125), .ZN(new_n1302));
  NAND4_X1  g1102(.A1(new_n1301), .A2(new_n1302), .A3(new_n711), .A4(new_n1297), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1300), .A2(new_n1303), .ZN(new_n1304));
  AOI21_X1  g1104(.A(G384), .B1(new_n1304), .B2(new_n1271), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1305), .ZN(new_n1306));
  AOI211_X1 g1106(.A(new_n1270), .B(new_n860), .C1(new_n1300), .C2(new_n1303), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1307), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1295), .B1(new_n1306), .B2(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1295), .ZN(new_n1310));
  NOR3_X1   g1110(.A1(new_n1305), .A2(new_n1307), .A3(new_n1310), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1309), .A2(new_n1311), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1199), .A2(new_n1029), .A3(new_n1237), .ZN(new_n1313));
  AND2_X1   g1113(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1314));
  AOI22_X1  g1114(.A1(new_n1314), .A2(new_n994), .B1(new_n1201), .B2(new_n1224), .ZN(new_n1315));
  AOI21_X1  g1115(.A(G378), .B1(new_n1313), .B2(new_n1315), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n1316), .B1(new_n1244), .B2(G378), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1312), .B1(new_n1317), .B2(new_n1294), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1319), .A2(new_n1243), .A3(new_n1320), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1226), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1321), .A2(G378), .A3(new_n1322), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1316), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1323), .A2(new_n1324), .ZN(new_n1325));
  INV_X1    g1125(.A(KEYINPUT62), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1294), .ZN(new_n1327));
  NOR2_X1   g1127(.A1(new_n1305), .A2(new_n1307), .ZN(new_n1328));
  NAND4_X1  g1128(.A1(new_n1325), .A2(new_n1326), .A3(new_n1327), .A4(new_n1328), .ZN(new_n1329));
  INV_X1    g1129(.A(KEYINPUT61), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1318), .A2(new_n1329), .A3(new_n1330), .ZN(new_n1331));
  AOI21_X1  g1131(.A(new_n1294), .B1(new_n1323), .B2(new_n1324), .ZN(new_n1332));
  AOI21_X1  g1132(.A(new_n1326), .B1(new_n1332), .B2(new_n1328), .ZN(new_n1333));
  OAI21_X1  g1133(.A(new_n1292), .B1(new_n1331), .B2(new_n1333), .ZN(new_n1334));
  INV_X1    g1134(.A(KEYINPUT127), .ZN(new_n1335));
  AOI21_X1  g1135(.A(new_n1335), .B1(new_n1291), .B2(new_n1330), .ZN(new_n1336));
  AOI211_X1 g1136(.A(KEYINPUT127), .B(KEYINPUT61), .C1(new_n1287), .C2(new_n1290), .ZN(new_n1337));
  NOR2_X1   g1137(.A1(new_n1336), .A2(new_n1337), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1332), .A2(new_n1328), .ZN(new_n1339));
  INV_X1    g1139(.A(KEYINPUT63), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1339), .A2(new_n1340), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1332), .A2(KEYINPUT63), .A3(new_n1328), .ZN(new_n1342));
  NAND4_X1  g1142(.A1(new_n1338), .A2(new_n1341), .A3(new_n1318), .A4(new_n1342), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1334), .A2(new_n1343), .ZN(G405));
  XOR2_X1   g1144(.A(new_n1291), .B(new_n1328), .Z(new_n1345));
  NOR2_X1   g1145(.A1(new_n1244), .A2(new_n1273), .ZN(new_n1346));
  INV_X1    g1146(.A(new_n1346), .ZN(new_n1347));
  NAND3_X1  g1147(.A1(new_n1345), .A2(new_n1277), .A3(new_n1347), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1277), .A2(new_n1347), .ZN(new_n1349));
  XNOR2_X1  g1149(.A(new_n1291), .B(new_n1328), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1349), .A2(new_n1350), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1348), .A2(new_n1351), .ZN(G402));
endmodule


