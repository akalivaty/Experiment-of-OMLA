//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 0 1 0 0 0 0 0 1 1 0 1 1 1 1 1 1 1 0 1 1 1 0 0 1 0 1 1 0 1 0 0 1 0 1 0 0 1 0 0 0 0 1 0 1 1 1 0 1 0 0 0 0 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:30 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1252, new_n1253, new_n1254, new_n1255,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1330, new_n1331;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  XOR2_X1   g0006(.A(KEYINPUT64), .B(G68), .Z(new_n207));
  INV_X1    g0007(.A(G238), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G58), .A2(G232), .B1(G87), .B2(G250), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G97), .A2(G257), .B1(G116), .B2(G270), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G107), .A2(G264), .ZN(new_n213));
  NAND4_X1  g0013(.A1(new_n210), .A2(new_n211), .A3(new_n212), .A4(new_n213), .ZN(new_n214));
  OAI21_X1  g0014(.A(new_n206), .B1(new_n209), .B2(new_n214), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT65), .ZN(new_n216));
  INV_X1    g0016(.A(KEYINPUT1), .ZN(new_n217));
  AND2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n216), .A2(new_n217), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n206), .A2(G13), .ZN(new_n220));
  OAI211_X1 g0020(.A(new_n220), .B(G250), .C1(G257), .C2(G264), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT0), .Z(new_n222));
  OAI21_X1  g0022(.A(G50), .B1(G58), .B2(G68), .ZN(new_n223));
  INV_X1    g0023(.A(G20), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  NOR3_X1   g0025(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  NOR4_X1   g0026(.A1(new_n218), .A2(new_n219), .A3(new_n222), .A4(new_n226), .ZN(G361));
  XOR2_X1   g0027(.A(G238), .B(G244), .Z(new_n228));
  XNOR2_X1  g0028(.A(KEYINPUT66), .B(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT2), .B(G226), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n232), .B(new_n235), .Z(G358));
  XNOR2_X1  g0036(.A(G50), .B(G68), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT67), .ZN(new_n238));
  XOR2_X1   g0038(.A(G58), .B(G77), .Z(new_n239));
  XOR2_X1   g0039(.A(new_n238), .B(new_n239), .Z(new_n240));
  XNOR2_X1  g0040(.A(G87), .B(G97), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n240), .B(new_n243), .Z(G351));
  OR2_X1    g0044(.A1(KEYINPUT68), .A2(G1), .ZN(new_n245));
  NAND2_X1  g0045(.A1(KEYINPUT68), .A2(G1), .ZN(new_n246));
  NAND4_X1  g0046(.A1(new_n245), .A2(G13), .A3(G20), .A4(new_n246), .ZN(new_n247));
  INV_X1    g0047(.A(new_n247), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(new_n202), .ZN(new_n249));
  NAND3_X1  g0049(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(new_n225), .ZN(new_n251));
  AND2_X1   g0051(.A1(KEYINPUT68), .A2(G1), .ZN(new_n252));
  NOR2_X1   g0052(.A1(KEYINPUT68), .A2(G1), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n251), .B1(new_n254), .B2(G20), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n249), .B1(new_n256), .B2(new_n202), .ZN(new_n257));
  NOR2_X1   g0057(.A1(G20), .A2(G33), .ZN(new_n258));
  AOI22_X1  g0058(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G58), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n260), .A2(KEYINPUT8), .ZN(new_n261));
  XNOR2_X1  g0061(.A(KEYINPUT69), .B(G58), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n261), .B1(new_n262), .B2(KEYINPUT8), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n224), .A2(G33), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n259), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n257), .B1(new_n251), .B2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT3), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n267), .A2(G33), .ZN(new_n268));
  INV_X1    g0068(.A(G33), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n269), .A2(KEYINPUT3), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G1698), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n271), .A2(G222), .A3(new_n272), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n271), .A2(G223), .A3(G1698), .ZN(new_n274));
  INV_X1    g0074(.A(G77), .ZN(new_n275));
  OAI211_X1 g0075(.A(new_n273), .B(new_n274), .C1(new_n275), .C2(new_n271), .ZN(new_n276));
  AND2_X1   g0076(.A1(G33), .A2(G41), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n277), .A2(new_n225), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  NOR2_X1   g0079(.A1(G41), .A2(G45), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G1), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n281), .A2(new_n282), .A3(G274), .ZN(new_n283));
  INV_X1    g0083(.A(G226), .ZN(new_n284));
  INV_X1    g0084(.A(G41), .ZN(new_n285));
  OAI211_X1 g0085(.A(G1), .B(G13), .C1(new_n269), .C2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n245), .A2(new_n246), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n286), .B1(new_n287), .B2(new_n280), .ZN(new_n288));
  OAI211_X1 g0088(.A(new_n279), .B(new_n283), .C1(new_n284), .C2(new_n288), .ZN(new_n289));
  XOR2_X1   g0089(.A(KEYINPUT70), .B(G179), .Z(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G169), .ZN(new_n293));
  AOI211_X1 g0093(.A(new_n266), .B(new_n292), .C1(new_n293), .C2(new_n289), .ZN(new_n294));
  XNOR2_X1  g0094(.A(new_n266), .B(KEYINPUT9), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n289), .A2(G200), .ZN(new_n296));
  INV_X1    g0096(.A(G190), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n296), .B1(new_n297), .B2(new_n289), .ZN(new_n298));
  OR3_X1    g0098(.A1(new_n295), .A2(new_n298), .A3(KEYINPUT10), .ZN(new_n299));
  OAI21_X1  g0099(.A(KEYINPUT10), .B1(new_n298), .B2(new_n295), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n294), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  XNOR2_X1  g0101(.A(KEYINPUT64), .B(G68), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n302), .A2(new_n224), .ZN(new_n303));
  INV_X1    g0103(.A(new_n258), .ZN(new_n304));
  OAI22_X1  g0104(.A1(new_n304), .A2(new_n202), .B1(new_n264), .B2(new_n275), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n251), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT11), .ZN(new_n307));
  XNOR2_X1  g0107(.A(new_n306), .B(new_n307), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n248), .A2(KEYINPUT12), .A3(new_n207), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n309), .B1(KEYINPUT12), .B2(new_n248), .ZN(new_n310));
  INV_X1    g0110(.A(G68), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n311), .B1(new_n256), .B2(KEYINPUT12), .ZN(new_n312));
  NOR3_X1   g0112(.A1(new_n308), .A2(new_n310), .A3(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  OR2_X1    g0114(.A1(new_n293), .A2(KEYINPUT73), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n283), .B1(new_n288), .B2(new_n208), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n269), .A2(KEYINPUT3), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n284), .A2(new_n272), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n267), .A2(G33), .ZN(new_n319));
  INV_X1    g0119(.A(G232), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(G1698), .ZN(new_n321));
  NAND4_X1  g0121(.A1(new_n317), .A2(new_n318), .A3(new_n319), .A4(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(G33), .A2(G97), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n286), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  OAI21_X1  g0124(.A(KEYINPUT13), .B1(new_n316), .B2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n283), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n278), .B1(new_n254), .B2(new_n281), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n326), .B1(new_n327), .B2(G238), .ZN(new_n328));
  INV_X1    g0128(.A(new_n324), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT13), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n328), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n315), .B1(new_n325), .B2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT14), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n325), .A2(new_n331), .ZN(new_n334));
  INV_X1    g0134(.A(G179), .ZN(new_n335));
  OAI22_X1  g0135(.A1(new_n332), .A2(new_n333), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  AOI211_X1 g0136(.A(KEYINPUT14), .B(new_n315), .C1(new_n325), .C2(new_n331), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n314), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n325), .A2(new_n331), .A3(G190), .ZN(new_n339));
  AND2_X1   g0139(.A1(new_n313), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n334), .A2(G200), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NOR2_X1   g0142(.A1(G232), .A2(G1698), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n272), .A2(G238), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n271), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  OAI211_X1 g0145(.A(new_n345), .B(new_n278), .C1(G107), .C2(new_n271), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n326), .B1(new_n327), .B2(G244), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n348), .A2(new_n297), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT72), .ZN(new_n350));
  XNOR2_X1  g0150(.A(new_n258), .B(KEYINPUT71), .ZN(new_n351));
  XNOR2_X1  g0151(.A(KEYINPUT8), .B(G58), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  XNOR2_X1  g0153(.A(KEYINPUT15), .B(G87), .ZN(new_n354));
  OAI22_X1  g0154(.A1(new_n354), .A2(new_n264), .B1(new_n224), .B2(new_n275), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n251), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n255), .A2(G77), .ZN(new_n357));
  OAI211_X1 g0157(.A(new_n356), .B(new_n357), .C1(G77), .C2(new_n247), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n349), .B1(new_n350), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n348), .A2(G200), .ZN(new_n360));
  OAI211_X1 g0160(.A(new_n359), .B(new_n360), .C1(new_n350), .C2(new_n358), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n348), .A2(new_n293), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n346), .A2(new_n290), .A3(new_n347), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n362), .A2(new_n358), .A3(new_n363), .ZN(new_n364));
  AND2_X1   g0164(.A1(new_n361), .A2(new_n364), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n301), .A2(new_n338), .A3(new_n342), .A4(new_n365), .ZN(new_n366));
  OAI22_X1  g0166(.A1(new_n207), .A2(new_n262), .B1(G58), .B2(G68), .ZN(new_n367));
  AOI22_X1  g0167(.A1(new_n367), .A2(G20), .B1(G159), .B2(new_n258), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n267), .A2(KEYINPUT74), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT74), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(KEYINPUT3), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n369), .A2(new_n371), .A3(G33), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(new_n317), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT7), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n373), .A2(new_n374), .A3(new_n224), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(G68), .ZN(new_n376));
  AOI21_X1  g0176(.A(G20), .B1(new_n372), .B2(new_n317), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n377), .A2(new_n374), .ZN(new_n378));
  OAI211_X1 g0178(.A(new_n368), .B(KEYINPUT16), .C1(new_n376), .C2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT16), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n374), .B1(new_n271), .B2(G20), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n374), .A2(G20), .ZN(new_n382));
  AOI21_X1  g0182(.A(G33), .B1(new_n369), .B2(new_n371), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n382), .B1(new_n383), .B2(new_n270), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n207), .B1(new_n381), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n258), .A2(G159), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n260), .A2(KEYINPUT69), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT69), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(G58), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n201), .B1(new_n390), .B2(new_n302), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n386), .B1(new_n391), .B2(new_n224), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n380), .B1(new_n385), .B2(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n379), .A2(new_n393), .A3(new_n251), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n263), .A2(new_n248), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n395), .B1(new_n256), .B2(new_n263), .ZN(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(G200), .ZN(new_n398));
  NOR2_X1   g0198(.A1(G223), .A2(G1698), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n399), .B1(new_n284), .B2(G1698), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n400), .A2(new_n372), .A3(new_n317), .ZN(new_n401));
  NAND2_X1  g0201(.A1(G33), .A2(G87), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n286), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n283), .B1(new_n288), .B2(new_n320), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n398), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n326), .B1(new_n327), .B2(G232), .ZN(new_n406));
  AND2_X1   g0206(.A1(new_n401), .A2(new_n402), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n406), .B1(new_n407), .B2(new_n286), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n405), .B1(new_n408), .B2(G190), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n394), .A2(new_n397), .A3(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT17), .ZN(new_n411));
  OR2_X1    g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n394), .A2(new_n397), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n408), .A2(G169), .ZN(new_n414));
  OAI211_X1 g0214(.A(new_n406), .B(new_n291), .C1(new_n407), .C2(new_n286), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n413), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(KEYINPUT18), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT18), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n413), .A2(new_n419), .A3(new_n416), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n410), .A2(new_n411), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n412), .A2(new_n418), .A3(new_n420), .A4(new_n421), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n366), .A2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT85), .ZN(new_n424));
  MUX2_X1   g0224(.A(G250), .B(G257), .S(G1698), .Z(new_n425));
  NAND3_X1  g0225(.A1(new_n425), .A2(new_n372), .A3(new_n317), .ZN(new_n426));
  NAND2_X1  g0226(.A1(G33), .A2(G294), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n286), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  XOR2_X1   g0228(.A(KEYINPUT5), .B(G41), .Z(new_n429));
  NAND3_X1  g0229(.A1(new_n245), .A2(G45), .A3(new_n246), .ZN(new_n430));
  OAI211_X1 g0230(.A(G264), .B(new_n286), .C1(new_n429), .C2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n428), .A2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(G45), .ZN(new_n434));
  NOR3_X1   g0234(.A1(new_n252), .A2(new_n253), .A3(new_n434), .ZN(new_n435));
  XNOR2_X1  g0235(.A(KEYINPUT5), .B(G41), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n435), .A2(G274), .A3(new_n286), .A4(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n293), .B1(new_n433), .B2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n437), .ZN(new_n439));
  NOR4_X1   g0239(.A1(new_n428), .A2(new_n432), .A3(new_n439), .A4(new_n335), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n424), .B1(new_n438), .B2(new_n440), .ZN(new_n441));
  NOR3_X1   g0241(.A1(new_n428), .A2(new_n432), .A3(new_n439), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(G179), .ZN(new_n443));
  XNOR2_X1  g0243(.A(KEYINPUT74), .B(KEYINPUT3), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n268), .B1(new_n444), .B2(G33), .ZN(new_n445));
  AOI22_X1  g0245(.A1(new_n445), .A2(new_n425), .B1(G33), .B2(G294), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n431), .B(new_n437), .C1(new_n446), .C2(new_n286), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(G169), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n443), .A2(KEYINPUT85), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n441), .A2(new_n449), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n372), .A2(new_n224), .A3(G87), .A4(new_n317), .ZN(new_n451));
  AND3_X1   g0251(.A1(new_n451), .A2(KEYINPUT82), .A3(KEYINPUT22), .ZN(new_n452));
  AOI21_X1  g0252(.A(KEYINPUT82), .B1(new_n451), .B2(KEYINPUT22), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n317), .A2(new_n319), .ZN(new_n454));
  INV_X1    g0254(.A(G87), .ZN(new_n455));
  NOR4_X1   g0255(.A1(new_n454), .A2(KEYINPUT22), .A3(G20), .A4(new_n455), .ZN(new_n456));
  NOR3_X1   g0256(.A1(new_n452), .A2(new_n453), .A3(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT23), .ZN(new_n458));
  INV_X1    g0258(.A(G107), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n458), .B1(G20), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(KEYINPUT83), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n460), .A2(KEYINPUT83), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n458), .A2(new_n459), .A3(G20), .ZN(new_n464));
  INV_X1    g0264(.A(G116), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n464), .B1(new_n465), .B2(new_n264), .ZN(new_n466));
  NOR3_X1   g0266(.A1(new_n462), .A2(new_n463), .A3(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  NOR3_X1   g0268(.A1(new_n457), .A2(KEYINPUT24), .A3(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT24), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n451), .A2(KEYINPUT22), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT82), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n456), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n451), .A2(KEYINPUT82), .A3(KEYINPUT22), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n470), .B1(new_n475), .B2(new_n467), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n251), .B1(new_n469), .B2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(new_n251), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n245), .A2(G33), .A3(new_n246), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n247), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n480), .A2(new_n459), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n248), .A2(new_n459), .ZN(new_n482));
  XOR2_X1   g0282(.A(KEYINPUT84), .B(KEYINPUT25), .Z(new_n483));
  OR2_X1    g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n482), .A2(new_n483), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n481), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n450), .B1(new_n477), .B2(new_n486), .ZN(new_n487));
  OAI21_X1  g0287(.A(KEYINPUT24), .B1(new_n457), .B2(new_n468), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n475), .A2(new_n470), .A3(new_n467), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n478), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(new_n486), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n442), .A2(new_n297), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n447), .A2(new_n398), .ZN(new_n493));
  AND2_X1   g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NOR3_X1   g0294(.A1(new_n490), .A2(new_n491), .A3(new_n494), .ZN(new_n495));
  OAI21_X1  g0295(.A(KEYINPUT86), .B1(new_n487), .B2(new_n495), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n441), .B(new_n449), .C1(new_n490), .C2(new_n491), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n492), .A2(new_n493), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n477), .A2(new_n486), .A3(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT86), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n497), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n496), .A2(new_n501), .ZN(new_n502));
  OAI211_X1 g0302(.A(G270), .B(new_n286), .C1(new_n429), .C2(new_n430), .ZN(new_n503));
  MUX2_X1   g0303(.A(G257), .B(G264), .S(G1698), .Z(new_n504));
  XNOR2_X1  g0304(.A(KEYINPUT80), .B(G303), .ZN(new_n505));
  AOI22_X1  g0305(.A1(new_n445), .A2(new_n504), .B1(new_n454), .B2(new_n505), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n437), .B(new_n503), .C1(new_n506), .C2(new_n286), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n247), .A2(new_n478), .A3(new_n479), .A4(G116), .ZN(new_n508));
  AOI22_X1  g0308(.A1(new_n250), .A2(new_n225), .B1(G20), .B2(new_n465), .ZN(new_n509));
  NAND2_X1  g0309(.A1(G33), .A2(G283), .ZN(new_n510));
  INV_X1    g0310(.A(G97), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n510), .B(new_n224), .C1(G33), .C2(new_n511), .ZN(new_n512));
  AND3_X1   g0312(.A1(new_n509), .A2(KEYINPUT20), .A3(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(KEYINPUT20), .B1(new_n509), .B2(new_n512), .ZN(new_n514));
  OAI221_X1 g0314(.A(new_n508), .B1(G116), .B2(new_n247), .C1(new_n513), .C2(new_n514), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n507), .A2(G169), .A3(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT21), .ZN(new_n517));
  OR2_X1    g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n507), .A2(new_n335), .ZN(new_n519));
  AOI22_X1  g0319(.A1(new_n517), .A2(new_n516), .B1(new_n519), .B2(new_n515), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n507), .A2(G200), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT81), .ZN(new_n522));
  INV_X1    g0322(.A(new_n515), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n524), .B1(new_n297), .B2(new_n507), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n522), .B1(new_n521), .B2(new_n523), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n518), .B(new_n520), .C1(new_n525), .C2(new_n526), .ZN(new_n527));
  MUX2_X1   g0327(.A(G238), .B(G244), .S(G1698), .Z(new_n528));
  NAND3_X1  g0328(.A1(new_n528), .A2(new_n372), .A3(new_n317), .ZN(new_n529));
  NAND2_X1  g0329(.A1(G33), .A2(G116), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(new_n278), .ZN(new_n532));
  OAI21_X1  g0332(.A(G250), .B1(new_n277), .B2(new_n225), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT76), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n533), .B1(new_n534), .B2(new_n430), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n254), .A2(KEYINPUT76), .A3(G45), .ZN(new_n536));
  AND2_X1   g0336(.A1(new_n286), .A2(G274), .ZN(new_n537));
  AOI22_X1  g0337(.A1(new_n535), .A2(new_n536), .B1(new_n537), .B2(new_n435), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n532), .A2(new_n538), .A3(G190), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(KEYINPUT79), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT79), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n532), .A2(new_n538), .A3(new_n541), .A4(G190), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n480), .A2(new_n455), .ZN(new_n544));
  INV_X1    g0344(.A(new_n354), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n545), .A2(new_n247), .ZN(new_n546));
  NOR2_X1   g0346(.A1(G97), .A2(G107), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n547), .A2(new_n455), .B1(new_n323), .B2(new_n224), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT19), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(G97), .ZN(new_n550));
  OAI22_X1  g0350(.A1(new_n548), .A2(new_n549), .B1(new_n264), .B2(new_n550), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n372), .A2(new_n224), .A3(G68), .A4(new_n317), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT77), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n478), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n551), .A2(new_n552), .A3(KEYINPUT77), .ZN(new_n556));
  AOI211_X1 g0356(.A(new_n544), .B(new_n546), .C1(new_n555), .C2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n430), .A2(new_n534), .ZN(new_n558));
  INV_X1    g0358(.A(new_n533), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n558), .A2(new_n536), .A3(new_n559), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n254), .A2(new_n286), .A3(G45), .A4(G274), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n286), .B1(new_n529), .B2(new_n530), .ZN(new_n563));
  OAI21_X1  g0363(.A(G200), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n543), .A2(new_n557), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n546), .B1(new_n555), .B2(new_n556), .ZN(new_n566));
  XOR2_X1   g0366(.A(new_n354), .B(KEYINPUT78), .Z(new_n567));
  OR2_X1    g0367(.A1(new_n567), .A2(new_n480), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n293), .B1(new_n562), .B2(new_n563), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n532), .A2(new_n538), .A3(new_n290), .ZN(new_n571));
  AND2_X1   g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n565), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n459), .B1(new_n381), .B2(new_n384), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT6), .ZN(new_n576));
  NOR3_X1   g0376(.A1(new_n576), .A2(new_n511), .A3(G107), .ZN(new_n577));
  XNOR2_X1  g0377(.A(G97), .B(G107), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n577), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  OAI22_X1  g0379(.A1(new_n579), .A2(new_n224), .B1(new_n275), .B2(new_n304), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n251), .B1(new_n575), .B2(new_n580), .ZN(new_n581));
  MUX2_X1   g0381(.A(new_n247), .B(new_n480), .S(G97), .Z(new_n582));
  NAND2_X1  g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(new_n583), .ZN(new_n584));
  OAI211_X1 g0384(.A(G257), .B(new_n286), .C1(new_n429), .C2(new_n430), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(new_n437), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n372), .A2(G244), .A3(new_n272), .A4(new_n317), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT4), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n317), .A2(new_n319), .A3(G250), .A4(G1698), .ZN(new_n590));
  AND2_X1   g0390(.A1(KEYINPUT4), .A2(G244), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n317), .A2(new_n319), .A3(new_n591), .A4(new_n272), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n590), .A2(new_n592), .A3(new_n510), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n589), .A2(new_n594), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n586), .B1(new_n595), .B2(new_n278), .ZN(new_n596));
  OAI21_X1  g0396(.A(KEYINPUT75), .B1(new_n596), .B2(new_n398), .ZN(new_n597));
  AND2_X1   g0397(.A1(new_n585), .A2(new_n437), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n593), .B1(new_n588), .B2(new_n587), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n598), .B1(new_n599), .B2(new_n286), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT75), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n600), .A2(new_n601), .A3(G200), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n598), .B(G190), .C1(new_n599), .C2(new_n286), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n584), .A2(new_n597), .A3(new_n602), .A4(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n600), .A2(new_n293), .ZN(new_n605));
  OAI211_X1 g0405(.A(new_n598), .B(new_n290), .C1(new_n599), .C2(new_n286), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n605), .A2(new_n583), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n604), .A2(new_n607), .ZN(new_n608));
  NOR3_X1   g0408(.A1(new_n527), .A2(new_n574), .A3(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n423), .A2(new_n502), .A3(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(new_n610), .ZN(G372));
  INV_X1    g0411(.A(new_n420), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n419), .B1(new_n413), .B2(new_n416), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(new_n338), .ZN(new_n615));
  INV_X1    g0415(.A(new_n364), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n615), .B1(new_n342), .B2(new_n616), .ZN(new_n617));
  XNOR2_X1  g0417(.A(new_n410), .B(KEYINPUT17), .ZN(new_n618));
  INV_X1    g0418(.A(new_n618), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n614), .B1(new_n617), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n299), .A2(new_n300), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n294), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(new_n423), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n570), .A2(new_n571), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n624), .B1(new_n566), .B2(new_n568), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n555), .A2(new_n556), .ZN(new_n626));
  INV_X1    g0426(.A(new_n544), .ZN(new_n627));
  INV_X1    g0427(.A(new_n546), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n626), .A2(new_n564), .A3(new_n627), .A4(new_n628), .ZN(new_n629));
  AOI22_X1  g0429(.A1(new_n629), .A2(KEYINPUT87), .B1(new_n542), .B2(new_n540), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT87), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n557), .A2(new_n631), .A3(new_n564), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n625), .B1(new_n630), .B2(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT26), .ZN(new_n634));
  AND3_X1   g0434(.A1(new_n605), .A2(new_n583), .A3(new_n606), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n633), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n565), .A2(new_n635), .A3(new_n573), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n625), .B1(new_n637), .B2(KEYINPUT26), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n603), .A2(new_n581), .A3(new_n582), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n601), .B1(new_n600), .B2(G200), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n635), .B1(new_n641), .B2(new_n602), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n633), .A2(new_n642), .A3(new_n499), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n520), .A2(new_n518), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n477), .A2(new_n486), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n443), .A2(new_n448), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n644), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  OAI211_X1 g0447(.A(new_n636), .B(new_n638), .C1(new_n643), .C2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n622), .B1(new_n623), .B2(new_n649), .ZN(G369));
  INV_X1    g0450(.A(G13), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n651), .A2(G20), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  OAI21_X1  g0453(.A(KEYINPUT27), .B1(new_n287), .B2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT27), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n254), .A2(new_n655), .A3(new_n652), .ZN(new_n656));
  AND3_X1   g0456(.A1(new_n654), .A2(G213), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(G343), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n497), .A2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n658), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n645), .A2(new_n660), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n659), .B1(new_n502), .B2(new_n661), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n523), .A2(new_n658), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n644), .A2(new_n663), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n664), .B1(new_n527), .B2(new_n663), .ZN(new_n665));
  XOR2_X1   g0465(.A(KEYINPUT88), .B(G330), .Z(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n662), .A2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n645), .A2(new_n646), .A3(new_n658), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n644), .A2(new_n658), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  AND3_X1   g0473(.A1(new_n497), .A2(new_n500), .A3(new_n499), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n500), .B1(new_n497), .B2(new_n499), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n673), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n670), .A2(new_n671), .A3(new_n676), .ZN(G399));
  INV_X1    g0477(.A(new_n220), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n678), .A2(G41), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n547), .A2(new_n455), .A3(new_n465), .ZN(new_n680));
  NOR3_X1   g0480(.A1(new_n679), .A2(new_n680), .A3(new_n282), .ZN(new_n681));
  INV_X1    g0481(.A(new_n223), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n681), .B1(new_n682), .B2(new_n679), .ZN(new_n683));
  XOR2_X1   g0483(.A(new_n683), .B(KEYINPUT28), .Z(new_n684));
  INV_X1    g0484(.A(KEYINPUT89), .ZN(new_n685));
  INV_X1    g0485(.A(new_n450), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n644), .B1(new_n645), .B2(new_n686), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n685), .B1(new_n643), .B2(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n495), .A2(new_n608), .ZN(new_n689));
  AND2_X1   g0489(.A1(new_n520), .A2(new_n518), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n490), .A2(new_n491), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n690), .B1(new_n691), .B2(new_n450), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n689), .A2(new_n692), .A3(KEYINPUT89), .A4(new_n633), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n565), .A2(new_n635), .A3(new_n634), .A4(new_n573), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(new_n573), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n633), .A2(new_n635), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n695), .B1(new_n696), .B2(KEYINPUT26), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n688), .A2(new_n693), .A3(new_n697), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n698), .A2(KEYINPUT29), .A3(new_n658), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n648), .A2(new_n658), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT29), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  AND2_X1   g0502(.A1(new_n699), .A2(new_n702), .ZN(new_n703));
  OAI211_X1 g0503(.A(new_n609), .B(new_n658), .C1(new_n674), .C2(new_n675), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n562), .A2(new_n563), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n519), .A2(new_n433), .A3(new_n705), .A4(new_n596), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT30), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  AND2_X1   g0508(.A1(new_n705), .A2(new_n433), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n709), .A2(KEYINPUT30), .A3(new_n519), .A4(new_n596), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n705), .A2(new_n291), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n711), .A2(new_n447), .A3(new_n507), .A4(new_n600), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n708), .A2(new_n710), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(new_n660), .ZN(new_n714));
  XNOR2_X1  g0514(.A(new_n714), .B(KEYINPUT31), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n666), .B1(new_n704), .B2(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n703), .A2(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n684), .B1(new_n717), .B2(G1), .ZN(G364));
  INV_X1    g0518(.A(new_n668), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n282), .B1(new_n652), .B2(G45), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n679), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n719), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n723), .B1(new_n667), .B2(new_n665), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n225), .B1(G20), .B2(new_n293), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(G322), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n290), .A2(new_n224), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n297), .A2(G200), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n297), .A2(new_n398), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n728), .A2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(G326), .ZN(new_n733));
  OAI22_X1  g0533(.A1(new_n727), .A2(new_n730), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n731), .A2(G20), .A3(new_n335), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n224), .A2(G190), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n737), .A2(new_n335), .A3(new_n398), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  AOI22_X1  g0539(.A1(G303), .A2(new_n736), .B1(new_n739), .B2(G329), .ZN(new_n740));
  INV_X1    g0540(.A(G283), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n737), .A2(new_n335), .A3(G200), .ZN(new_n742));
  OAI211_X1 g0542(.A(new_n740), .B(new_n454), .C1(new_n741), .C2(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n729), .A2(new_n335), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(G20), .ZN(new_n745));
  AOI211_X1 g0545(.A(new_n734), .B(new_n743), .C1(G294), .C2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(G311), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n728), .A2(new_n297), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n749), .A2(KEYINPUT92), .A3(new_n398), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT92), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n751), .B1(new_n748), .B2(G200), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n749), .A2(G200), .ZN(new_n755));
  XOR2_X1   g0555(.A(KEYINPUT33), .B(G317), .Z(new_n756));
  OAI221_X1 g0556(.A(new_n746), .B1(new_n747), .B2(new_n754), .C1(new_n755), .C2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n745), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(new_n511), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n739), .A2(G159), .ZN(new_n760));
  XNOR2_X1  g0560(.A(new_n760), .B(KEYINPUT32), .ZN(new_n761));
  INV_X1    g0561(.A(new_n755), .ZN(new_n762));
  AOI211_X1 g0562(.A(new_n759), .B(new_n761), .C1(new_n762), .C2(G68), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n732), .A2(new_n202), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n736), .A2(G87), .ZN(new_n765));
  OAI211_X1 g0565(.A(new_n765), .B(new_n271), .C1(new_n459), .C2(new_n742), .ZN(new_n766));
  INV_X1    g0566(.A(new_n730), .ZN(new_n767));
  AOI211_X1 g0567(.A(new_n764), .B(new_n766), .C1(new_n390), .C2(new_n767), .ZN(new_n768));
  OAI211_X1 g0568(.A(new_n763), .B(new_n768), .C1(new_n275), .C2(new_n754), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n726), .B1(new_n757), .B2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n722), .ZN(new_n771));
  NOR2_X1   g0571(.A1(G13), .A2(G33), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(G20), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(new_n725), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n445), .A2(new_n678), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n777), .B1(G45), .B2(new_n223), .ZN(new_n778));
  XNOR2_X1  g0578(.A(new_n778), .B(KEYINPUT91), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n779), .B1(new_n434), .B2(new_n240), .ZN(new_n780));
  XOR2_X1   g0580(.A(G355), .B(KEYINPUT90), .Z(new_n781));
  NOR2_X1   g0581(.A1(new_n678), .A2(new_n454), .ZN(new_n782));
  AOI22_X1  g0582(.A1(new_n781), .A2(new_n782), .B1(new_n465), .B2(new_n678), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n776), .B1(new_n780), .B2(new_n783), .ZN(new_n784));
  NOR3_X1   g0584(.A1(new_n770), .A2(new_n771), .A3(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n774), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n785), .B1(new_n665), .B2(new_n786), .ZN(new_n787));
  AND2_X1   g0587(.A1(new_n724), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(G396));
  INV_X1    g0589(.A(G150), .ZN(new_n790));
  INV_X1    g0590(.A(G137), .ZN(new_n791));
  OAI22_X1  g0591(.A1(new_n755), .A2(new_n790), .B1(new_n791), .B2(new_n732), .ZN(new_n792));
  XNOR2_X1  g0592(.A(new_n792), .B(KEYINPUT93), .ZN(new_n793));
  INV_X1    g0593(.A(G143), .ZN(new_n794));
  INV_X1    g0594(.A(G159), .ZN(new_n795));
  OAI221_X1 g0595(.A(new_n793), .B1(new_n794), .B2(new_n730), .C1(new_n795), .C2(new_n754), .ZN(new_n796));
  XOR2_X1   g0596(.A(new_n796), .B(KEYINPUT34), .Z(new_n797));
  INV_X1    g0597(.A(new_n742), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(G68), .ZN(new_n799));
  INV_X1    g0599(.A(G132), .ZN(new_n800));
  OAI221_X1 g0600(.A(new_n799), .B1(new_n202), .B2(new_n735), .C1(new_n800), .C2(new_n738), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n445), .B1(new_n758), .B2(new_n262), .ZN(new_n802));
  NOR3_X1   g0602(.A1(new_n797), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  AOI22_X1  g0603(.A1(G107), .A2(new_n736), .B1(new_n739), .B2(G311), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n798), .A2(G87), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n804), .A2(new_n454), .A3(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n806), .A2(new_n759), .ZN(new_n807));
  INV_X1    g0607(.A(new_n732), .ZN(new_n808));
  AOI22_X1  g0608(.A1(G294), .A2(new_n767), .B1(new_n808), .B2(G303), .ZN(new_n809));
  OAI211_X1 g0609(.A(new_n807), .B(new_n809), .C1(new_n741), .C2(new_n755), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n810), .B1(G116), .B2(new_n753), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n725), .B1(new_n803), .B2(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n725), .A2(new_n772), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n771), .B1(new_n275), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n358), .A2(new_n660), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n361), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(new_n364), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n616), .A2(new_n658), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  OAI211_X1 g0620(.A(new_n812), .B(new_n814), .C1(new_n773), .C2(new_n820), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n821), .B(KEYINPUT94), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n648), .A2(new_n820), .A3(new_n658), .ZN(new_n823));
  XOR2_X1   g0623(.A(new_n819), .B(KEYINPUT95), .Z(new_n824));
  INV_X1    g0624(.A(new_n700), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n823), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n716), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n722), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n828), .B1(new_n827), .B2(new_n826), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n822), .A2(new_n829), .ZN(G384));
  NAND2_X1  g0630(.A1(new_n704), .A2(new_n715), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT97), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n338), .A2(new_n832), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n313), .A2(new_n658), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n834), .B1(new_n340), .B2(new_n341), .ZN(new_n835));
  OAI211_X1 g0635(.A(KEYINPUT97), .B(new_n314), .C1(new_n336), .C2(new_n337), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n833), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n834), .B1(new_n336), .B2(new_n337), .ZN(new_n838));
  AND2_X1   g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n839), .A2(new_n819), .ZN(new_n840));
  AND2_X1   g0640(.A1(new_n831), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n311), .B1(new_n377), .B2(new_n374), .ZN(new_n842));
  OAI21_X1  g0642(.A(KEYINPUT7), .B1(new_n445), .B2(G20), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n392), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n478), .B1(new_n844), .B2(KEYINPUT16), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n368), .B1(new_n376), .B2(new_n378), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n846), .A2(new_n380), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n396), .B1(new_n845), .B2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n657), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n410), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  AND2_X1   g0650(.A1(new_n414), .A2(new_n415), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n848), .A2(new_n851), .ZN(new_n852));
  OAI21_X1  g0652(.A(KEYINPUT37), .B1(new_n850), .B2(new_n852), .ZN(new_n853));
  XOR2_X1   g0653(.A(new_n657), .B(KEYINPUT98), .Z(new_n854));
  NAND2_X1  g0654(.A1(new_n413), .A2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT37), .ZN(new_n856));
  NAND4_X1  g0656(.A1(new_n417), .A2(new_n855), .A3(new_n856), .A4(new_n410), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n853), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(KEYINPUT99), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT99), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n853), .A2(new_n860), .A3(new_n857), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n848), .A2(new_n849), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n422), .A2(new_n862), .ZN(new_n863));
  NAND4_X1  g0663(.A1(new_n859), .A2(KEYINPUT38), .A3(new_n861), .A4(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT38), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n417), .A2(new_n855), .A3(new_n410), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(KEYINPUT37), .ZN(new_n867));
  AND2_X1   g0667(.A1(new_n867), .A2(new_n857), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n855), .B1(new_n614), .B2(new_n618), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n865), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n864), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n841), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(KEYINPUT40), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n859), .A2(new_n861), .A3(new_n863), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(new_n865), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(new_n864), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT40), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n841), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n873), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n423), .A2(new_n831), .ZN(new_n880));
  XOR2_X1   g0680(.A(new_n879), .B(new_n880), .Z(new_n881));
  NOR2_X1   g0681(.A1(new_n881), .A2(new_n666), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n660), .B1(new_n833), .B2(new_n836), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT100), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT39), .ZN(new_n886));
  NAND4_X1  g0686(.A1(new_n864), .A2(new_n870), .A3(new_n885), .A4(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n886), .B1(new_n875), .B2(new_n864), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n864), .A2(new_n886), .A3(new_n870), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(KEYINPUT100), .ZN(new_n890));
  OAI211_X1 g0690(.A(new_n884), .B(new_n887), .C1(new_n888), .C2(new_n890), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n614), .A2(new_n854), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n839), .B1(new_n823), .B2(new_n818), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n892), .B1(new_n876), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n891), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n699), .A2(new_n423), .A3(new_n702), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(new_n622), .ZN(new_n897));
  XNOR2_X1  g0697(.A(new_n895), .B(new_n897), .ZN(new_n898));
  AOI22_X1  g0698(.A1(new_n883), .A2(new_n898), .B1(new_n287), .B2(new_n653), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n899), .B1(new_n898), .B2(new_n883), .ZN(new_n900));
  NOR3_X1   g0700(.A1(new_n225), .A2(new_n224), .A3(new_n465), .ZN(new_n901));
  XNOR2_X1  g0701(.A(new_n579), .B(KEYINPUT96), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT35), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n901), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n905), .B1(new_n904), .B2(new_n903), .ZN(new_n906));
  XOR2_X1   g0706(.A(new_n906), .B(KEYINPUT36), .Z(new_n907));
  OAI211_X1 g0707(.A(G77), .B(new_n682), .C1(new_n207), .C2(new_n262), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n908), .B1(G50), .B2(new_n311), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n909), .A2(new_n651), .A3(new_n287), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n900), .A2(new_n907), .A3(new_n910), .ZN(new_n911));
  XOR2_X1   g0711(.A(new_n911), .B(KEYINPUT101), .Z(G367));
  OAI21_X1  g0712(.A(new_n642), .B1(new_n584), .B2(new_n658), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n607), .B1(new_n913), .B2(new_n497), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT102), .ZN(new_n915));
  OR2_X1    g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n914), .A2(new_n915), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n916), .A2(new_n658), .A3(new_n917), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n672), .B1(new_n496), .B2(new_n501), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT103), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT42), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n635), .A2(new_n660), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n913), .A2(new_n922), .ZN(new_n923));
  NAND4_X1  g0723(.A1(new_n919), .A2(new_n920), .A3(new_n921), .A4(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n919), .A2(new_n923), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(KEYINPUT42), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n918), .A2(new_n924), .A3(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT43), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n633), .B1(new_n557), .B2(new_n658), .ZN(new_n930));
  OR3_X1    g0730(.A1(new_n573), .A2(new_n557), .A3(new_n658), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(KEYINPUT103), .B1(new_n925), .B2(KEYINPUT42), .ZN(new_n934));
  NAND4_X1  g0734(.A1(new_n928), .A2(new_n929), .A3(new_n933), .A4(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n933), .A2(new_n929), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n932), .A2(KEYINPUT43), .ZN(new_n937));
  INV_X1    g0737(.A(new_n934), .ZN(new_n938));
  OAI211_X1 g0738(.A(new_n936), .B(new_n937), .C1(new_n927), .C2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n669), .A2(new_n923), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  AND3_X1   g0741(.A1(new_n935), .A2(new_n939), .A3(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n941), .B1(new_n935), .B2(new_n939), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  XOR2_X1   g0744(.A(new_n679), .B(KEYINPUT41), .Z(new_n945));
  INV_X1    g0745(.A(new_n923), .ZN(new_n946));
  INV_X1    g0746(.A(new_n671), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n946), .B1(new_n919), .B2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT44), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  OAI211_X1 g0750(.A(KEYINPUT44), .B(new_n946), .C1(new_n919), .C2(new_n947), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n676), .A2(new_n671), .A3(new_n923), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT45), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND4_X1  g0754(.A1(new_n676), .A2(KEYINPUT45), .A3(new_n671), .A4(new_n923), .ZN(new_n955));
  AOI22_X1  g0755(.A1(new_n950), .A2(new_n951), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n670), .B1(new_n956), .B2(KEYINPUT104), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n950), .A2(new_n951), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n954), .A2(new_n955), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT104), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n960), .A2(new_n961), .A3(new_n669), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n661), .B1(new_n674), .B2(new_n675), .ZN(new_n963));
  INV_X1    g0763(.A(new_n659), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n963), .A2(new_n964), .A3(new_n672), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT105), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n919), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  AOI211_X1 g0768(.A(KEYINPUT105), .B(new_n672), .C1(new_n496), .C2(new_n501), .ZN(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n668), .B1(new_n968), .B2(new_n970), .ZN(new_n971));
  AOI211_X1 g0771(.A(new_n719), .B(new_n969), .C1(new_n965), .C2(new_n967), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n957), .A2(new_n962), .A3(new_n717), .A4(new_n973), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n945), .B1(new_n974), .B2(new_n717), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n944), .B1(new_n975), .B2(new_n721), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n776), .B1(new_n678), .B2(new_n545), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n235), .A2(new_n777), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n771), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  OAI22_X1  g0779(.A1(new_n794), .A2(new_n732), .B1(new_n730), .B2(new_n790), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n758), .A2(new_n311), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n271), .B1(new_n735), .B2(new_n262), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n798), .A2(G77), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n983), .B1(new_n791), .B2(new_n738), .ZN(new_n984));
  NOR4_X1   g0784(.A1(new_n980), .A2(new_n981), .A3(new_n982), .A4(new_n984), .ZN(new_n985));
  OAI221_X1 g0785(.A(new_n985), .B1(new_n795), .B2(new_n755), .C1(new_n754), .C2(new_n202), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n798), .A2(G97), .ZN(new_n987));
  INV_X1    g0787(.A(G317), .ZN(new_n988));
  OAI211_X1 g0788(.A(new_n987), .B(new_n373), .C1(new_n988), .C2(new_n738), .ZN(new_n989));
  XNOR2_X1  g0789(.A(KEYINPUT106), .B(G311), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n732), .A2(new_n990), .ZN(new_n991));
  AOI211_X1 g0791(.A(new_n989), .B(new_n991), .C1(new_n505), .C2(new_n767), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n736), .A2(KEYINPUT46), .A3(G116), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT46), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n994), .B1(new_n735), .B2(new_n465), .ZN(new_n995));
  OAI211_X1 g0795(.A(new_n993), .B(new_n995), .C1(new_n459), .C2(new_n758), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n996), .B1(new_n762), .B2(G294), .ZN(new_n997));
  OAI211_X1 g0797(.A(new_n992), .B(new_n997), .C1(new_n741), .C2(new_n754), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n986), .A2(new_n998), .ZN(new_n999));
  XOR2_X1   g0799(.A(new_n999), .B(KEYINPUT47), .Z(new_n1000));
  OAI221_X1 g0800(.A(new_n979), .B1(new_n932), .B2(new_n786), .C1(new_n1000), .C2(new_n726), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n976), .A2(new_n1001), .ZN(G387));
  OAI22_X1  g0802(.A1(new_n971), .A2(new_n972), .B1(new_n703), .B2(new_n716), .ZN(new_n1003));
  OR2_X1    g0803(.A1(new_n1003), .A2(KEYINPUT108), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n973), .A2(new_n717), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1003), .A2(KEYINPUT108), .ZN(new_n1006));
  NAND4_X1  g0806(.A1(new_n1004), .A2(new_n679), .A3(new_n1005), .A4(new_n1006), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(new_n782), .A2(new_n680), .B1(new_n459), .B2(new_n678), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n232), .A2(new_n434), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n352), .A2(G50), .ZN(new_n1010));
  XOR2_X1   g0810(.A(new_n1010), .B(KEYINPUT50), .Z(new_n1011));
  INV_X1    g0811(.A(new_n680), .ZN(new_n1012));
  OAI211_X1 g0812(.A(new_n1012), .B(new_n434), .C1(new_n311), .C2(new_n275), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n777), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1008), .B1(new_n1009), .B2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n771), .B1(new_n1015), .B2(new_n775), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n754), .A2(new_n311), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n736), .A2(G77), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n739), .A2(G150), .ZN(new_n1019));
  NAND4_X1  g0819(.A1(new_n1018), .A2(new_n987), .A3(new_n1019), .A4(new_n445), .ZN(new_n1020));
  XOR2_X1   g0820(.A(new_n1020), .B(KEYINPUT107), .Z(new_n1021));
  OR2_X1    g0821(.A1(new_n567), .A2(new_n758), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n1022), .B1(new_n730), .B2(new_n202), .C1(new_n795), .C2(new_n732), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n755), .A2(new_n263), .ZN(new_n1024));
  NOR4_X1   g0824(.A1(new_n1017), .A2(new_n1021), .A3(new_n1023), .A4(new_n1024), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n742), .A2(new_n465), .B1(new_n738), .B2(new_n733), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(G317), .A2(new_n767), .B1(new_n808), .B2(G322), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1027), .B1(new_n755), .B2(new_n990), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1028), .B1(new_n505), .B2(new_n753), .ZN(new_n1029));
  OR2_X1    g0829(.A1(new_n1029), .A2(KEYINPUT48), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1029), .A2(KEYINPUT48), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(G294), .A2(new_n736), .B1(new_n745), .B2(G283), .ZN(new_n1032));
  AND3_X1   g0832(.A1(new_n1030), .A2(new_n1031), .A3(new_n1032), .ZN(new_n1033));
  AOI211_X1 g0833(.A(new_n445), .B(new_n1026), .C1(new_n1033), .C2(KEYINPUT49), .ZN(new_n1034));
  OR2_X1    g0834(.A1(new_n1033), .A2(KEYINPUT49), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1025), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1016), .B1(new_n1036), .B2(new_n726), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1037), .B1(new_n662), .B2(new_n774), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1038), .B1(new_n973), .B2(new_n721), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1007), .A2(new_n1039), .ZN(G393));
  NOR2_X1   g0840(.A1(new_n960), .A2(new_n669), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n956), .A2(new_n670), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1043), .A2(new_n721), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n776), .B1(G97), .B2(new_n678), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n243), .A2(new_n777), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n771), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n505), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n755), .A2(new_n1048), .B1(new_n465), .B2(new_n758), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n1049), .A2(KEYINPUT110), .B1(new_n753), .B2(G294), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1050), .B1(KEYINPUT110), .B2(new_n1049), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n747), .A2(new_n730), .B1(new_n732), .B2(new_n988), .ZN(new_n1052));
  XOR2_X1   g0852(.A(new_n1052), .B(KEYINPUT52), .Z(new_n1053));
  OAI21_X1  g0853(.A(new_n454), .B1(new_n742), .B2(new_n459), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n735), .A2(new_n741), .B1(new_n738), .B2(new_n727), .ZN(new_n1055));
  NOR4_X1   g0855(.A1(new_n1051), .A2(new_n1053), .A3(new_n1054), .A4(new_n1055), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1056), .B(KEYINPUT111), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n754), .A2(new_n352), .B1(new_n202), .B2(new_n755), .ZN(new_n1058));
  INV_X1    g0858(.A(KEYINPUT109), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n790), .A2(new_n732), .B1(new_n730), .B2(new_n795), .ZN(new_n1061));
  XOR2_X1   g0861(.A(new_n1061), .B(KEYINPUT51), .Z(new_n1062));
  OAI221_X1 g0862(.A(new_n805), .B1(new_n794), .B2(new_n738), .C1(new_n207), .C2(new_n735), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n445), .B1(new_n758), .B2(new_n275), .ZN(new_n1064));
  NOR3_X1   g0864(.A1(new_n1062), .A2(new_n1063), .A3(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n1058), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1065), .B1(KEYINPUT109), .B2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1057), .B1(new_n1060), .B2(new_n1067), .ZN(new_n1068));
  XOR2_X1   g0868(.A(new_n1068), .B(KEYINPUT112), .Z(new_n1069));
  OAI221_X1 g0869(.A(new_n1047), .B1(new_n786), .B2(new_n923), .C1(new_n1069), .C2(new_n726), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1005), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1071), .A2(new_n679), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n974), .ZN(new_n1073));
  OAI211_X1 g0873(.A(new_n1044), .B(new_n1070), .C1(new_n1072), .C2(new_n1073), .ZN(G390));
  NAND3_X1  g0874(.A1(new_n698), .A2(new_n658), .A3(new_n817), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1075), .A2(new_n818), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n839), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n884), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1078), .A2(new_n1079), .A3(new_n871), .ZN(new_n1080));
  AOI211_X1 g0880(.A(new_n666), .B(new_n819), .C1(new_n704), .C2(new_n715), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1081), .A2(new_n1077), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n887), .ZN(new_n1083));
  AND2_X1   g0883(.A1(new_n889), .A2(KEYINPUT100), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n864), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n858), .A2(KEYINPUT99), .B1(new_n422), .B2(new_n862), .ZN(new_n1086));
  AOI21_X1  g0886(.A(KEYINPUT38), .B1(new_n1086), .B2(new_n861), .ZN(new_n1087));
  OAI21_X1  g0887(.A(KEYINPUT39), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1083), .B1(new_n1084), .B2(new_n1088), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n893), .A2(new_n884), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n1080), .B(new_n1082), .C1(new_n1089), .C2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n871), .A2(new_n1079), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(new_n1077), .B2(new_n1076), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n887), .B1(new_n888), .B2(new_n890), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1090), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1093), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n831), .A2(G330), .A3(new_n840), .ZN(new_n1097));
  OAI211_X1 g0897(.A(new_n1091), .B(new_n721), .C1(new_n1096), .C2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n762), .A2(G137), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n735), .A2(new_n790), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(new_n1100), .B(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1102), .B1(G159), .B2(new_n745), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n767), .A2(G132), .ZN(new_n1104));
  INV_X1    g0904(.A(G125), .ZN(new_n1105));
  OAI221_X1 g0905(.A(new_n271), .B1(new_n738), .B2(new_n1105), .C1(new_n202), .C2(new_n742), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1106), .B1(new_n808), .B2(G128), .ZN(new_n1107));
  NAND4_X1  g0907(.A1(new_n1099), .A2(new_n1103), .A3(new_n1104), .A4(new_n1107), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(KEYINPUT54), .B(G143), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n754), .A2(new_n1109), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n754), .A2(new_n511), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n739), .A2(G294), .ZN(new_n1112));
  NAND4_X1  g0912(.A1(new_n765), .A2(new_n799), .A3(new_n1112), .A4(new_n454), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1113), .B1(G77), .B2(new_n745), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(G116), .A2(new_n767), .B1(new_n808), .B2(G283), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n1114), .B(new_n1115), .C1(new_n459), .C2(new_n755), .ZN(new_n1116));
  OAI22_X1  g0916(.A1(new_n1108), .A2(new_n1110), .B1(new_n1111), .B2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1117), .A2(new_n725), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n771), .B1(new_n263), .B2(new_n813), .ZN(new_n1119));
  OAI211_X1 g0919(.A(new_n1118), .B(new_n1119), .C1(new_n1089), .C2(new_n773), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1098), .A2(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n679), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1091), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1123));
  INV_X1    g0923(.A(G330), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1124), .B1(new_n704), .B2(new_n715), .ZN(new_n1125));
  INV_X1    g0925(.A(KEYINPUT114), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n824), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  AOI211_X1 g0927(.A(KEYINPUT114), .B(new_n1124), .C1(new_n704), .C2(new_n715), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n839), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1076), .B1(new_n1077), .B2(new_n1081), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(KEYINPUT113), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n823), .A2(new_n818), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1077), .B1(new_n716), .B2(new_n820), .ZN(new_n1134));
  AND3_X1   g0934(.A1(new_n831), .A2(G330), .A3(new_n840), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n1132), .B(new_n1133), .C1(new_n1134), .C2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1097), .B1(new_n1081), .B2(new_n1077), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1132), .B1(new_n1138), .B2(new_n1133), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1131), .B1(new_n1137), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n423), .A2(new_n1125), .ZN(new_n1141));
  AND3_X1   g0941(.A1(new_n896), .A2(new_n622), .A3(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1122), .B1(new_n1123), .B2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1088), .A2(KEYINPUT100), .A3(new_n889), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1090), .B1(new_n1145), .B2(new_n887), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1135), .B1(new_n1146), .B2(new_n1093), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n1147), .A2(new_n1140), .A3(new_n1091), .A4(new_n1142), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1121), .B1(new_n1144), .B2(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(G378));
  NOR2_X1   g0950(.A1(new_n266), .A2(new_n849), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n301), .B(new_n1151), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n1152), .B(new_n1153), .ZN(new_n1154));
  AND3_X1   g0954(.A1(new_n891), .A2(new_n894), .A3(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n879), .A2(G330), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1154), .B1(new_n891), .B2(new_n894), .ZN(new_n1157));
  NOR3_X1   g0957(.A1(new_n1155), .A2(new_n1156), .A3(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1124), .B1(new_n873), .B2(new_n878), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1154), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n895), .A2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n891), .A2(new_n894), .A3(new_n1154), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1159), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n721), .B1(new_n1158), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1160), .A2(new_n772), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n813), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n722), .B1(G50), .B2(new_n1166), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n202), .B1(G33), .B2(G41), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1168), .B1(new_n373), .B2(new_n285), .ZN(new_n1169));
  OAI221_X1 g0969(.A(new_n1018), .B1(new_n741), .B2(new_n738), .C1(new_n262), .C2(new_n742), .ZN(new_n1170));
  AOI211_X1 g0970(.A(new_n981), .B(new_n1170), .C1(new_n762), .C2(G97), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n459), .A2(new_n730), .B1(new_n732), .B2(new_n465), .ZN(new_n1172));
  NOR3_X1   g0972(.A1(new_n1172), .A2(G41), .A3(new_n445), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n1171), .B(new_n1173), .C1(new_n567), .C2(new_n754), .ZN(new_n1174));
  INV_X1    g0974(.A(KEYINPUT58), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1169), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1109), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n736), .A2(new_n1177), .B1(new_n745), .B2(G150), .ZN(new_n1178));
  INV_X1    g0978(.A(G128), .ZN(new_n1179));
  OAI221_X1 g0979(.A(new_n1178), .B1(new_n730), .B2(new_n1179), .C1(new_n1105), .C2(new_n732), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n755), .A2(new_n800), .ZN(new_n1181));
  AOI211_X1 g0981(.A(new_n1180), .B(new_n1181), .C1(G137), .C2(new_n753), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1183), .A2(KEYINPUT59), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n798), .A2(G159), .ZN(new_n1185));
  AOI211_X1 g0985(.A(G33), .B(G41), .C1(new_n739), .C2(G124), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1184), .A2(new_n1185), .A3(new_n1186), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n1183), .A2(KEYINPUT59), .ZN(new_n1188));
  OAI221_X1 g0988(.A(new_n1176), .B1(new_n1175), .B2(new_n1174), .C1(new_n1187), .C2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1167), .B1(new_n1189), .B2(new_n725), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1165), .A2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1164), .A2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1148), .A2(new_n1142), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1156), .B1(new_n1155), .B2(new_n1157), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1161), .A2(new_n1159), .A3(new_n1162), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1194), .A2(KEYINPUT57), .A3(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1198), .A2(new_n679), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n1148), .A2(new_n1142), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n1200), .A2(KEYINPUT57), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1193), .B1(new_n1199), .B2(new_n1201), .ZN(G375));
  INV_X1    g1002(.A(new_n945), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1133), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1204), .A2(KEYINPUT113), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1205), .A2(new_n1136), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1142), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1206), .A2(new_n1207), .A3(new_n1131), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1143), .A2(new_n1203), .A3(new_n1208), .ZN(new_n1209));
  XNOR2_X1  g1009(.A(new_n1209), .B(KEYINPUT116), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n839), .A2(new_n772), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n722), .B1(G68), .B2(new_n1166), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1022), .A2(new_n454), .A3(new_n983), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(G116), .B2(new_n762), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n753), .A2(G107), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(G97), .A2(new_n736), .B1(new_n739), .B2(G303), .ZN(new_n1216));
  XOR2_X1   g1016(.A(new_n1216), .B(KEYINPUT117), .Z(new_n1217));
  AOI22_X1  g1017(.A1(G283), .A2(new_n767), .B1(new_n808), .B2(G294), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1214), .A2(new_n1215), .A3(new_n1217), .A4(new_n1218), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n753), .A2(G150), .B1(G50), .B2(new_n745), .ZN(new_n1220));
  XNOR2_X1  g1020(.A(new_n1220), .B(KEYINPUT118), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n762), .A2(new_n1177), .ZN(new_n1222));
  OAI22_X1  g1022(.A1(new_n742), .A2(new_n262), .B1(new_n738), .B2(new_n1179), .ZN(new_n1223));
  AOI211_X1 g1023(.A(new_n373), .B(new_n1223), .C1(G159), .C2(new_n736), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(G132), .A2(new_n808), .B1(new_n767), .B2(G137), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1222), .A2(new_n1224), .A3(new_n1225), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1219), .B1(new_n1221), .B2(new_n1226), .ZN(new_n1227));
  OR2_X1    g1027(.A1(new_n1227), .A2(KEYINPUT119), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n726), .B1(new_n1227), .B2(KEYINPUT119), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1212), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(new_n1140), .A2(new_n721), .B1(new_n1211), .B2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1210), .A2(new_n1231), .ZN(G381));
  AOI21_X1  g1032(.A(new_n1122), .B1(new_n1200), .B2(KEYINPUT57), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT57), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1082), .ZN(new_n1235));
  AOI211_X1 g1035(.A(new_n1235), .B(new_n1093), .C1(new_n1094), .C2(new_n1095), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1097), .B1(new_n1237), .B2(new_n1080), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1236), .A2(new_n1238), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1207), .B1(new_n1206), .B2(new_n1131), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1207), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1158), .A2(new_n1163), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1234), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1192), .B1(new_n1233), .B2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1244), .A2(new_n1149), .ZN(new_n1245));
  INV_X1    g1045(.A(G390), .ZN(new_n1246));
  INV_X1    g1046(.A(G384), .ZN(new_n1247));
  AND3_X1   g1047(.A1(new_n1007), .A2(new_n788), .A3(new_n1039), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1246), .A2(new_n1247), .A3(new_n1248), .ZN(new_n1249));
  NOR4_X1   g1049(.A1(new_n1245), .A2(G387), .A3(G381), .A4(new_n1249), .ZN(new_n1250));
  XNOR2_X1  g1050(.A(new_n1250), .B(KEYINPUT120), .ZN(G407));
  INV_X1    g1051(.A(G343), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1252), .A2(G213), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1245), .A2(new_n1253), .ZN(new_n1254));
  XNOR2_X1  g1054(.A(new_n1254), .B(KEYINPUT121), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(G407), .A2(G213), .A3(new_n1255), .ZN(G409));
  NAND3_X1  g1056(.A1(new_n1164), .A2(KEYINPUT122), .A3(new_n1191), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT122), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n720), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1191), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1258), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1194), .A2(new_n1203), .A3(new_n1197), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1257), .A2(new_n1261), .A3(new_n1149), .A4(new_n1262), .ZN(new_n1263));
  AND2_X1   g1063(.A1(new_n1263), .A2(new_n1253), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(G375), .A2(G378), .ZN(new_n1265));
  AOI221_X4 g1065(.A(new_n1142), .B1(new_n1129), .B2(new_n1130), .C1(new_n1205), .C2(new_n1136), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1266), .B1(KEYINPUT60), .B2(new_n1143), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1206), .A2(KEYINPUT60), .A3(new_n1207), .A4(new_n1131), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(new_n679), .ZN(new_n1269));
  OAI211_X1 g1069(.A(G384), .B(new_n1231), .C1(new_n1267), .C2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT123), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT60), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1208), .B1(new_n1240), .B2(new_n1273), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1274), .A2(new_n679), .A3(new_n1268), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1275), .A2(KEYINPUT123), .A3(G384), .A4(new_n1231), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1143), .A2(KEYINPUT60), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1269), .B1(new_n1208), .B2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1231), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1247), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1280));
  AND3_X1   g1080(.A1(new_n1272), .A2(new_n1276), .A3(new_n1280), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1264), .A2(new_n1265), .A3(new_n1281), .ZN(new_n1282));
  OR2_X1    g1082(.A1(new_n1282), .A2(KEYINPUT62), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT61), .ZN(new_n1284));
  OAI211_X1 g1084(.A(new_n1253), .B(new_n1263), .C1(new_n1244), .C2(new_n1149), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1252), .A2(G213), .A3(G2897), .ZN(new_n1286));
  XOR2_X1   g1086(.A(new_n1286), .B(KEYINPUT125), .Z(new_n1287));
  INV_X1    g1087(.A(new_n1287), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1272), .A2(new_n1276), .A3(new_n1280), .A4(new_n1288), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1272), .A2(new_n1276), .A3(new_n1280), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1290), .A2(new_n1287), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1285), .A2(new_n1289), .A3(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1282), .A2(KEYINPUT62), .ZN(new_n1293));
  NAND4_X1  g1093(.A1(new_n1283), .A2(new_n1284), .A3(new_n1292), .A4(new_n1293), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n788), .B1(new_n1007), .B2(new_n1039), .ZN(new_n1295));
  OR2_X1    g1095(.A1(new_n1248), .A2(new_n1295), .ZN(new_n1296));
  AND3_X1   g1096(.A1(new_n976), .A2(G390), .A3(new_n1001), .ZN(new_n1297));
  AOI21_X1  g1097(.A(G390), .B1(new_n976), .B2(new_n1001), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1296), .B1(new_n1297), .B2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(G387), .A2(new_n1246), .ZN(new_n1300));
  NOR2_X1   g1100(.A1(new_n1248), .A2(new_n1295), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n976), .A2(G390), .A3(new_n1001), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1300), .A2(new_n1301), .A3(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1299), .A2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1294), .A2(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT127), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT63), .ZN(new_n1307));
  OAI211_X1 g1107(.A(KEYINPUT124), .B(new_n1307), .C1(new_n1285), .C2(new_n1290), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1308), .ZN(new_n1309));
  AOI21_X1  g1109(.A(KEYINPUT124), .B1(new_n1282), .B2(new_n1307), .ZN(new_n1310));
  NOR2_X1   g1110(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1299), .A2(new_n1303), .A3(new_n1284), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1312), .A2(KEYINPUT126), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT126), .ZN(new_n1314));
  NAND4_X1  g1114(.A1(new_n1299), .A2(new_n1303), .A3(new_n1314), .A4(new_n1284), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1313), .A2(new_n1315), .ZN(new_n1316));
  NAND4_X1  g1116(.A1(new_n1264), .A2(new_n1265), .A3(new_n1281), .A4(KEYINPUT63), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1316), .A2(new_n1292), .A3(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1318), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1306), .B1(new_n1311), .B2(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT124), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1243), .A2(new_n679), .A3(new_n1198), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1149), .B1(new_n1322), .B2(new_n1193), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1263), .A2(new_n1253), .ZN(new_n1324));
  NOR3_X1   g1124(.A1(new_n1323), .A2(new_n1324), .A3(new_n1290), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1321), .B1(new_n1325), .B2(KEYINPUT63), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1326), .A2(new_n1308), .ZN(new_n1327));
  NOR3_X1   g1127(.A1(new_n1327), .A2(KEYINPUT127), .A3(new_n1318), .ZN(new_n1328));
  OAI21_X1  g1128(.A(new_n1305), .B1(new_n1320), .B2(new_n1328), .ZN(G405));
  NAND2_X1  g1129(.A1(new_n1265), .A2(new_n1245), .ZN(new_n1330));
  XNOR2_X1  g1130(.A(new_n1330), .B(new_n1290), .ZN(new_n1331));
  XNOR2_X1  g1131(.A(new_n1331), .B(new_n1304), .ZN(G402));
endmodule


