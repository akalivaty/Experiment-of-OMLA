//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 0 1 1 1 0 0 0 0 1 1 0 0 0 0 1 1 1 1 1 1 1 0 1 0 1 0 1 0 1 1 0 0 0 1 1 1 1 0 0 1 0 0 1 1 1 1 1 1 1 0 0 0 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:24 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n535, new_n536, new_n537, new_n538, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n553, new_n554, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n564, new_n565, new_n567, new_n568, new_n569,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n603, new_n604, new_n605, new_n606, new_n607, new_n608, new_n611,
    new_n612, new_n613, new_n614, new_n616, new_n617, new_n618, new_n619,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n856, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1185, new_n1186, new_n1187, new_n1189;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT65), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n450));
  XNOR2_X1  g025(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(G2105), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G137), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n462), .A2(G2105), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G101), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n463), .A2(new_n464), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G125), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n470), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n469), .A2(new_n474), .ZN(G160));
  NAND2_X1  g050(.A1(new_n471), .A2(G2105), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n465), .A2(G136), .ZN(new_n479));
  OR2_X1    g054(.A1(G100), .A2(G2105), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n480), .B(G2104), .C1(G112), .C2(new_n470), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n478), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G162));
  OAI21_X1  g058(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(G114), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n484), .B1(new_n485), .B2(G2105), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n486), .B1(new_n477), .B2(G126), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT4), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n465), .A2(G138), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT68), .ZN(new_n490));
  OAI21_X1  g065(.A(new_n488), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n488), .A2(KEYINPUT67), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n465), .A2(KEYINPUT68), .A3(G138), .A4(new_n492), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n489), .A2(KEYINPUT67), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n487), .A2(new_n491), .A3(new_n493), .A4(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(G164));
  OAI21_X1  g071(.A(G543), .B1(KEYINPUT71), .B2(KEYINPUT5), .ZN(new_n497));
  AND2_X1   g072(.A1(KEYINPUT71), .A2(KEYINPUT5), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AND2_X1   g074(.A1(KEYINPUT69), .A2(G543), .ZN(new_n500));
  NOR2_X1   g075(.A1(KEYINPUT69), .A2(G543), .ZN(new_n501));
  OAI21_X1  g076(.A(KEYINPUT5), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(KEYINPUT70), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT70), .ZN(new_n504));
  OAI211_X1 g079(.A(new_n504), .B(KEYINPUT5), .C1(new_n500), .C2(new_n501), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n499), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  AND2_X1   g081(.A1(KEYINPUT6), .A2(G651), .ZN(new_n507));
  NOR2_X1   g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(new_n510));
  XNOR2_X1  g085(.A(KEYINPUT72), .B(G88), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n506), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  AND2_X1   g087(.A1(new_n510), .A2(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G50), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(KEYINPUT73), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT73), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n512), .A2(new_n517), .A3(new_n514), .ZN(new_n518));
  NAND2_X1  g093(.A1(G75), .A2(G543), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n503), .A2(new_n505), .ZN(new_n520));
  INV_X1    g095(.A(new_n499), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(G62), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n519), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n516), .A2(new_n518), .B1(G651), .B2(new_n524), .ZN(G166));
  AOI211_X1 g100(.A(new_n509), .B(new_n499), .C1(new_n503), .C2(new_n505), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G89), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n506), .A2(G63), .A3(G651), .ZN(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(KEYINPUT7), .ZN(new_n530));
  OR2_X1    g105(.A1(new_n529), .A2(KEYINPUT7), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n513), .A2(G51), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n527), .A2(new_n528), .A3(new_n532), .ZN(G286));
  INV_X1    g108(.A(G286), .ZN(G168));
  AOI22_X1  g109(.A1(new_n506), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n535));
  INV_X1    g110(.A(G651), .ZN(new_n536));
  OR2_X1    g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n526), .A2(G90), .B1(G52), .B2(new_n513), .ZN(new_n538));
  AND2_X1   g113(.A1(new_n537), .A2(new_n538), .ZN(G171));
  AOI22_X1  g114(.A1(new_n506), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT74), .ZN(new_n541));
  AND2_X1   g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  OAI21_X1  g117(.A(G651), .B1(new_n540), .B2(new_n541), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n506), .A2(G81), .A3(new_n510), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT75), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n513), .A2(G43), .ZN(new_n546));
  AND3_X1   g121(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n545), .B1(new_n544), .B2(new_n546), .ZN(new_n548));
  OAI22_X1  g123(.A1(new_n542), .A2(new_n543), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND4_X1  g129(.A1(G319), .A2(G483), .A3(G661), .A4(new_n554), .ZN(G188));
  NAND3_X1  g130(.A1(new_n506), .A2(G91), .A3(new_n510), .ZN(new_n556));
  INV_X1    g131(.A(G53), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n557), .A2(KEYINPUT76), .ZN(new_n558));
  OAI211_X1 g133(.A(new_n558), .B(G543), .C1(new_n508), .C2(new_n507), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT9), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n506), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n561));
  OAI211_X1 g136(.A(new_n556), .B(new_n560), .C1(new_n561), .C2(new_n536), .ZN(G299));
  INV_X1    g137(.A(G171), .ZN(G301));
  NAND2_X1  g138(.A1(new_n516), .A2(new_n518), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n524), .A2(G651), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n564), .A2(new_n565), .ZN(G303));
  NAND2_X1  g141(.A1(new_n526), .A2(G87), .ZN(new_n567));
  OAI21_X1  g142(.A(G651), .B1(new_n506), .B2(G74), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n513), .A2(G49), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(G288));
  AOI22_X1  g145(.A1(new_n506), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n571));
  NOR2_X1   g146(.A1(new_n571), .A2(new_n536), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n513), .A2(G48), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n506), .A2(new_n510), .ZN(new_n574));
  INV_X1    g149(.A(G86), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n573), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  OR2_X1    g151(.A1(new_n572), .A2(new_n576), .ZN(G305));
  NAND2_X1  g152(.A1(new_n513), .A2(G47), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n526), .A2(G85), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n506), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n580), .A2(KEYINPUT77), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(new_n582));
  OAI21_X1  g157(.A(G651), .B1(new_n580), .B2(KEYINPUT77), .ZN(new_n583));
  OAI211_X1 g158(.A(new_n578), .B(new_n579), .C1(new_n582), .C2(new_n583), .ZN(G290));
  XNOR2_X1  g159(.A(KEYINPUT69), .B(G543), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n504), .B1(new_n585), .B2(KEYINPUT5), .ZN(new_n586));
  INV_X1    g161(.A(new_n505), .ZN(new_n587));
  OAI211_X1 g162(.A(G66), .B(new_n521), .C1(new_n586), .C2(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(G79), .A2(G543), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n590), .A2(G651), .B1(G54), .B2(new_n513), .ZN(new_n591));
  NAND4_X1  g166(.A1(new_n520), .A2(G92), .A3(new_n521), .A4(new_n510), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT10), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND4_X1  g169(.A1(new_n506), .A2(KEYINPUT10), .A3(G92), .A4(new_n510), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  AND3_X1   g171(.A1(new_n591), .A2(KEYINPUT78), .A3(new_n596), .ZN(new_n597));
  AOI21_X1  g172(.A(KEYINPUT78), .B1(new_n591), .B2(new_n596), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(G868), .ZN(new_n600));
  MUX2_X1   g175(.A(G301), .B(new_n599), .S(new_n600), .Z(G284));
  MUX2_X1   g176(.A(G301), .B(new_n599), .S(new_n600), .Z(G321));
  NAND2_X1  g177(.A1(G286), .A2(G868), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n506), .A2(G65), .ZN(new_n604));
  NAND2_X1  g179(.A1(G78), .A2(G543), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n536), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n556), .A2(new_n560), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n603), .B1(new_n608), .B2(G868), .ZN(G297));
  OAI21_X1  g184(.A(new_n603), .B1(new_n608), .B2(G868), .ZN(G280));
  INV_X1    g185(.A(new_n598), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n591), .A2(new_n596), .A3(KEYINPUT78), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(G559), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n613), .B1(new_n614), .B2(G860), .ZN(G148));
  OAI21_X1  g190(.A(new_n614), .B1(new_n597), .B2(new_n598), .ZN(new_n616));
  INV_X1    g191(.A(new_n616), .ZN(new_n617));
  OR3_X1    g192(.A1(new_n617), .A2(KEYINPUT79), .A3(new_n600), .ZN(new_n618));
  OAI21_X1  g193(.A(KEYINPUT79), .B1(new_n617), .B2(new_n600), .ZN(new_n619));
  OAI211_X1 g194(.A(new_n618), .B(new_n619), .C1(G868), .C2(new_n550), .ZN(G323));
  XNOR2_X1  g195(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g196(.A1(new_n471), .A2(new_n467), .ZN(new_n622));
  XOR2_X1   g197(.A(KEYINPUT80), .B(KEYINPUT12), .Z(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  XOR2_X1   g199(.A(KEYINPUT81), .B(KEYINPUT13), .Z(new_n625));
  XNOR2_X1  g200(.A(new_n624), .B(new_n625), .ZN(new_n626));
  INV_X1    g201(.A(G2100), .ZN(new_n627));
  OR2_X1    g202(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n626), .A2(new_n627), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n465), .A2(G135), .ZN(new_n630));
  NOR2_X1   g205(.A1(new_n470), .A2(G111), .ZN(new_n631));
  OAI21_X1  g206(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n632));
  INV_X1    g207(.A(G123), .ZN(new_n633));
  OAI221_X1 g208(.A(new_n630), .B1(new_n631), .B2(new_n632), .C1(new_n633), .C2(new_n476), .ZN(new_n634));
  INV_X1    g209(.A(G2096), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n628), .A2(new_n629), .A3(new_n636), .ZN(G156));
  INV_X1    g212(.A(KEYINPUT14), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2427), .B(G2438), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2430), .ZN(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT15), .B(G2435), .ZN(new_n641));
  AOI21_X1  g216(.A(new_n638), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  OAI21_X1  g217(.A(new_n642), .B1(new_n641), .B2(new_n640), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2451), .B(G2454), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT16), .ZN(new_n645));
  XNOR2_X1  g220(.A(G1341), .B(G1348), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n643), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2443), .B(G2446), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n648), .A2(new_n649), .ZN(new_n651));
  AND3_X1   g226(.A1(new_n650), .A2(G14), .A3(new_n651), .ZN(G401));
  XNOR2_X1  g227(.A(G2072), .B(G2078), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n653), .B(KEYINPUT17), .Z(new_n654));
  XNOR2_X1  g229(.A(G2067), .B(G2678), .ZN(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(new_n656));
  NOR2_X1   g231(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G2084), .B(G2090), .Z(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  OAI21_X1  g234(.A(new_n659), .B1(new_n655), .B2(new_n653), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT82), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n658), .A2(new_n655), .A3(new_n653), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT18), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n659), .A2(new_n655), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n664), .B1(new_n654), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n662), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(new_n635), .ZN(new_n668));
  XNOR2_X1  g243(.A(KEYINPUT83), .B(G2100), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(G227));
  XNOR2_X1  g245(.A(G1956), .B(G2474), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT85), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1961), .B(G1966), .ZN(new_n673));
  OR2_X1    g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n672), .A2(new_n673), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1971), .B(G1976), .ZN(new_n676));
  XNOR2_X1  g251(.A(KEYINPUT84), .B(KEYINPUT19), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n674), .A2(new_n675), .A3(new_n678), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n674), .A2(new_n678), .ZN(new_n680));
  INV_X1    g255(.A(KEYINPUT20), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NOR3_X1   g257(.A1(new_n674), .A2(KEYINPUT20), .A3(new_n678), .ZN(new_n683));
  OAI221_X1 g258(.A(new_n679), .B1(new_n678), .B2(new_n675), .C1(new_n682), .C2(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT86), .ZN(new_n685));
  XOR2_X1   g260(.A(G1981), .B(G1986), .Z(new_n686));
  XNOR2_X1  g261(.A(G1991), .B(G1996), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XOR2_X1   g263(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n685), .B(new_n690), .ZN(G229));
  NOR2_X1   g266(.A1(KEYINPUT90), .A2(KEYINPUT36), .ZN(new_n692));
  XOR2_X1   g267(.A(new_n692), .B(KEYINPUT91), .Z(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n572), .A2(new_n576), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n695), .A2(G16), .ZN(new_n696));
  INV_X1    g271(.A(KEYINPUT32), .ZN(new_n697));
  OR2_X1    g272(.A1(G6), .A2(G16), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n696), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n697), .B1(new_n696), .B2(new_n698), .ZN(new_n701));
  OAI21_X1  g276(.A(G1981), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(new_n701), .ZN(new_n703));
  INV_X1    g278(.A(G1981), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n703), .A2(new_n704), .A3(new_n699), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n702), .A2(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(G166), .A2(G16), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(G16), .B2(G22), .ZN(new_n709));
  INV_X1    g284(.A(G1971), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  OAI211_X1 g286(.A(new_n708), .B(G1971), .C1(G16), .C2(G22), .ZN(new_n712));
  INV_X1    g287(.A(G16), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G23), .ZN(new_n714));
  INV_X1    g289(.A(G288), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n714), .B1(new_n715), .B2(new_n713), .ZN(new_n716));
  XNOR2_X1  g291(.A(KEYINPUT33), .B(G1976), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n711), .A2(new_n712), .A3(new_n718), .ZN(new_n719));
  OAI21_X1  g294(.A(KEYINPUT34), .B1(new_n707), .B2(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(new_n719), .ZN(new_n722));
  INV_X1    g297(.A(KEYINPUT34), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n722), .A2(new_n723), .A3(new_n706), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n713), .A2(G24), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n579), .A2(new_n578), .ZN(new_n726));
  NAND2_X1  g301(.A1(G72), .A2(G543), .ZN(new_n727));
  INV_X1    g302(.A(G60), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n727), .B1(new_n522), .B2(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(KEYINPUT77), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n536), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n726), .B1(new_n731), .B2(new_n581), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n725), .B1(new_n732), .B2(new_n713), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n733), .A2(KEYINPUT89), .ZN(new_n734));
  INV_X1    g309(.A(KEYINPUT89), .ZN(new_n735));
  OAI211_X1 g310(.A(new_n735), .B(new_n725), .C1(new_n732), .C2(new_n713), .ZN(new_n736));
  INV_X1    g311(.A(G1986), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n734), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(G29), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n739), .A2(G25), .ZN(new_n740));
  XOR2_X1   g315(.A(new_n740), .B(KEYINPUT87), .Z(new_n741));
  NAND2_X1  g316(.A1(new_n465), .A2(G131), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT88), .ZN(new_n743));
  OAI21_X1  g318(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n744));
  INV_X1    g319(.A(G107), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n744), .B1(new_n745), .B2(G2105), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(new_n477), .B2(G119), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n743), .A2(new_n747), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n741), .B1(new_n748), .B2(G29), .ZN(new_n749));
  XOR2_X1   g324(.A(KEYINPUT35), .B(G1991), .Z(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(KEYINPUT90), .B2(KEYINPUT36), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n738), .A2(new_n752), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n737), .B1(new_n734), .B2(new_n736), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n724), .A2(new_n755), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n694), .B1(new_n721), .B2(new_n756), .ZN(new_n757));
  NAND4_X1  g332(.A1(new_n720), .A2(new_n724), .A3(new_n755), .A4(new_n693), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n613), .A2(new_n713), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(G4), .B2(new_n713), .ZN(new_n760));
  XNOR2_X1  g335(.A(KEYINPUT92), .B(G1348), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n713), .A2(G20), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT23), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(new_n608), .B2(new_n713), .ZN(new_n765));
  INV_X1    g340(.A(G1956), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n739), .A2(G32), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n477), .A2(G129), .ZN(new_n769));
  AOI22_X1  g344(.A1(new_n465), .A2(G141), .B1(G105), .B2(new_n467), .ZN(new_n770));
  NAND3_X1  g345(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n771));
  XOR2_X1   g346(.A(new_n771), .B(KEYINPUT26), .Z(new_n772));
  AND3_X1   g347(.A1(new_n769), .A2(new_n770), .A3(new_n772), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n768), .B1(new_n773), .B2(new_n739), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT27), .ZN(new_n775));
  INV_X1    g350(.A(G1996), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n739), .A2(G27), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT96), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(new_n495), .B2(G29), .ZN(new_n780));
  INV_X1    g355(.A(G2078), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n482), .A2(G29), .ZN(new_n783));
  AND2_X1   g358(.A1(new_n739), .A2(G35), .ZN(new_n784));
  INV_X1    g359(.A(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n783), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n786), .A2(KEYINPUT29), .ZN(new_n787));
  INV_X1    g362(.A(G2090), .ZN(new_n788));
  INV_X1    g363(.A(KEYINPUT29), .ZN(new_n789));
  NAND3_X1  g364(.A1(new_n783), .A2(new_n789), .A3(new_n785), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n787), .A2(new_n788), .A3(new_n790), .ZN(new_n791));
  NAND3_X1  g366(.A1(new_n777), .A2(new_n782), .A3(new_n791), .ZN(new_n792));
  OR2_X1    g367(.A1(new_n469), .A2(new_n474), .ZN(new_n793));
  INV_X1    g368(.A(KEYINPUT24), .ZN(new_n794));
  AND2_X1   g369(.A1(new_n794), .A2(G34), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n739), .B1(new_n794), .B2(G34), .ZN(new_n796));
  OAI22_X1  g371(.A1(new_n793), .A2(new_n739), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(G2084), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  XOR2_X1   g374(.A(KEYINPUT94), .B(G2067), .Z(new_n800));
  NAND2_X1  g375(.A1(new_n465), .A2(G140), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n470), .A2(G116), .ZN(new_n802));
  OAI21_X1  g377(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n803));
  INV_X1    g378(.A(G128), .ZN(new_n804));
  OAI221_X1 g379(.A(new_n801), .B1(new_n802), .B2(new_n803), .C1(new_n804), .C2(new_n476), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n805), .A2(G29), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n739), .A2(G26), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT28), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n799), .B1(new_n800), .B2(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n739), .A2(G33), .ZN(new_n811));
  AND2_X1   g386(.A1(new_n471), .A2(G127), .ZN(new_n812));
  AND2_X1   g387(.A1(G115), .A2(G2104), .ZN(new_n813));
  OAI21_X1  g388(.A(G2105), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(KEYINPUT25), .ZN(new_n815));
  NAND2_X1  g390(.A1(G103), .A2(G2104), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n815), .B1(new_n816), .B2(G2105), .ZN(new_n817));
  NAND4_X1  g392(.A1(new_n470), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n818));
  AOI22_X1  g393(.A1(new_n465), .A2(G139), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  AND2_X1   g394(.A1(new_n814), .A2(new_n819), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n811), .B1(new_n820), .B2(new_n739), .ZN(new_n821));
  INV_X1    g396(.A(G2072), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n821), .B(new_n822), .ZN(new_n823));
  OR2_X1    g398(.A1(new_n809), .A2(new_n800), .ZN(new_n824));
  XNOR2_X1  g399(.A(KEYINPUT30), .B(G28), .ZN(new_n825));
  OR2_X1    g400(.A1(KEYINPUT31), .A2(G11), .ZN(new_n826));
  NAND2_X1  g401(.A1(KEYINPUT31), .A2(G11), .ZN(new_n827));
  AOI22_X1  g402(.A1(new_n825), .A2(new_n739), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n828), .B1(new_n634), .B2(new_n739), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n829), .B1(new_n797), .B2(new_n798), .ZN(new_n830));
  NAND4_X1  g405(.A1(new_n810), .A2(new_n823), .A3(new_n824), .A4(new_n830), .ZN(new_n831));
  OAI22_X1  g406(.A1(new_n775), .A2(new_n776), .B1(new_n781), .B2(new_n780), .ZN(new_n832));
  NOR3_X1   g407(.A1(new_n792), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n713), .A2(G5), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n834), .B1(G171), .B2(new_n713), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n835), .B(G1961), .Z(new_n836));
  NAND4_X1  g411(.A1(new_n762), .A2(new_n767), .A3(new_n833), .A4(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(G168), .A2(G16), .ZN(new_n838));
  OR2_X1    g413(.A1(G16), .A2(G21), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n838), .A2(KEYINPUT95), .A3(new_n839), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n840), .B1(KEYINPUT95), .B2(new_n838), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n841), .A2(G1966), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n788), .B1(new_n787), .B2(new_n790), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT97), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  NOR2_X1   g420(.A1(G16), .A2(G19), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n846), .B1(new_n550), .B2(G16), .ZN(new_n847));
  XNOR2_X1  g422(.A(KEYINPUT93), .B(G1341), .ZN(new_n848));
  OR2_X1    g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n847), .A2(new_n848), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n841), .A2(G1966), .ZN(new_n851));
  NAND4_X1  g426(.A1(new_n845), .A2(new_n849), .A3(new_n850), .A4(new_n851), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n760), .A2(new_n761), .ZN(new_n853));
  NOR3_X1   g428(.A1(new_n837), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n757), .A2(new_n758), .A3(new_n854), .ZN(G150));
  INV_X1    g430(.A(KEYINPUT98), .ZN(new_n856));
  XNOR2_X1  g431(.A(G150), .B(new_n856), .ZN(G311));
  INV_X1    g432(.A(KEYINPUT100), .ZN(new_n858));
  AOI22_X1  g433(.A1(new_n526), .A2(G93), .B1(G55), .B2(new_n513), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n520), .A2(G67), .A3(new_n521), .ZN(new_n860));
  NAND2_X1  g435(.A1(G80), .A2(G543), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n536), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT99), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n859), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  AOI22_X1  g439(.A1(new_n506), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n865));
  NOR3_X1   g440(.A1(new_n865), .A2(KEYINPUT99), .A3(new_n536), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n858), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n862), .A2(new_n863), .ZN(new_n868));
  OAI21_X1  g443(.A(KEYINPUT99), .B1(new_n865), .B2(new_n536), .ZN(new_n869));
  NAND4_X1  g444(.A1(new_n868), .A2(new_n869), .A3(KEYINPUT100), .A4(new_n859), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n867), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n871), .A2(G860), .ZN(new_n872));
  XOR2_X1   g447(.A(new_n872), .B(KEYINPUT37), .Z(new_n873));
  NAND2_X1  g448(.A1(new_n613), .A2(G559), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(KEYINPUT38), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n867), .A2(new_n549), .A3(new_n870), .ZN(new_n876));
  OR2_X1    g451(.A1(new_n542), .A2(new_n543), .ZN(new_n877));
  OR2_X1    g452(.A1(new_n547), .A2(new_n548), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n868), .A2(new_n869), .A3(new_n859), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n876), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n875), .B(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(KEYINPUT39), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(KEYINPUT101), .ZN(new_n884));
  INV_X1    g459(.A(G860), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n885), .B1(new_n882), .B2(KEYINPUT39), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n873), .B1(new_n884), .B2(new_n886), .ZN(G145));
  INV_X1    g462(.A(G37), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n805), .B(KEYINPUT103), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(new_n820), .ZN(new_n890));
  XOR2_X1   g465(.A(new_n748), .B(new_n624), .Z(new_n891));
  XNOR2_X1  g466(.A(new_n890), .B(new_n891), .ZN(new_n892));
  XOR2_X1   g467(.A(new_n495), .B(new_n773), .Z(new_n893));
  OAI21_X1  g468(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n894));
  INV_X1    g469(.A(G118), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n894), .B1(new_n895), .B2(G2105), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n465), .A2(G142), .ZN(new_n897));
  XOR2_X1   g472(.A(new_n897), .B(KEYINPUT104), .Z(new_n898));
  AOI211_X1 g473(.A(new_n896), .B(new_n898), .C1(G130), .C2(new_n477), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n893), .B(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n892), .B(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n793), .B(KEYINPUT102), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n902), .B(G162), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n903), .B(new_n634), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n888), .B1(new_n901), .B2(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n905), .B1(new_n904), .B2(new_n901), .ZN(new_n906));
  XOR2_X1   g481(.A(new_n906), .B(KEYINPUT40), .Z(G395));
  XNOR2_X1  g482(.A(new_n695), .B(G288), .ZN(new_n908));
  NOR2_X1   g483(.A1(G303), .A2(new_n732), .ZN(new_n909));
  NOR2_X1   g484(.A1(G290), .A2(G166), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n908), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n695), .B(new_n715), .ZN(new_n912));
  NAND2_X1  g487(.A1(G290), .A2(G166), .ZN(new_n913));
  NAND2_X1  g488(.A1(G303), .A2(new_n732), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n911), .A2(new_n915), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n916), .B1(KEYINPUT106), .B2(KEYINPUT42), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  AND2_X1   g493(.A1(new_n594), .A2(new_n595), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n513), .A2(G54), .ZN(new_n920));
  AOI22_X1  g495(.A1(new_n506), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n920), .B1(new_n921), .B2(new_n536), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n608), .B1(new_n919), .B2(new_n922), .ZN(new_n923));
  NAND3_X1  g498(.A1(G299), .A2(new_n591), .A3(new_n596), .ZN(new_n924));
  AND3_X1   g499(.A1(new_n923), .A2(KEYINPUT41), .A3(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT105), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n923), .A2(new_n926), .ZN(new_n927));
  OAI211_X1 g502(.A(new_n608), .B(KEYINPUT105), .C1(new_n919), .C2(new_n922), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n927), .A2(new_n924), .A3(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT41), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n925), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  AND3_X1   g506(.A1(new_n876), .A2(new_n616), .A3(new_n880), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n616), .B1(new_n876), .B2(new_n880), .ZN(new_n933));
  NOR3_X1   g508(.A1(new_n931), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n881), .A2(new_n617), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n876), .A2(new_n616), .A3(new_n880), .ZN(new_n936));
  AOI22_X1  g511(.A1(new_n935), .A2(new_n936), .B1(new_n924), .B2(new_n923), .ZN(new_n937));
  NOR2_X1   g512(.A1(KEYINPUT106), .A2(KEYINPUT42), .ZN(new_n938));
  NOR3_X1   g513(.A1(new_n934), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n938), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n929), .A2(new_n930), .ZN(new_n941));
  INV_X1    g516(.A(new_n925), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n943), .A2(new_n935), .A3(new_n936), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n923), .A2(new_n924), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n945), .B1(new_n932), .B2(new_n933), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n940), .B1(new_n944), .B2(new_n946), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n918), .B1(new_n939), .B2(new_n947), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n938), .B1(new_n934), .B2(new_n937), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n935), .A2(new_n936), .ZN(new_n950));
  OAI211_X1 g525(.A(new_n946), .B(new_n940), .C1(new_n950), .C2(new_n931), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n949), .A2(new_n917), .A3(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n600), .B1(new_n948), .B2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(new_n871), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n954), .A2(G868), .ZN(new_n955));
  NOR3_X1   g530(.A1(new_n953), .A2(KEYINPUT107), .A3(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT107), .ZN(new_n957));
  AND3_X1   g532(.A1(new_n949), .A2(new_n917), .A3(new_n951), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n917), .B1(new_n949), .B2(new_n951), .ZN(new_n959));
  OAI21_X1  g534(.A(G868), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(new_n955), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n957), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n956), .A2(new_n962), .ZN(G295));
  NAND2_X1  g538(.A1(new_n960), .A2(new_n961), .ZN(G331));
  AND3_X1   g539(.A1(new_n537), .A2(G286), .A3(new_n538), .ZN(new_n965));
  AOI21_X1  g540(.A(G286), .B1(new_n537), .B2(new_n538), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  AND3_X1   g542(.A1(new_n876), .A2(new_n880), .A3(new_n967), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n967), .B1(new_n876), .B2(new_n880), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  OAI21_X1  g545(.A(KEYINPUT109), .B1(new_n970), .B2(new_n931), .ZN(new_n971));
  INV_X1    g546(.A(new_n967), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n881), .A2(new_n972), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n876), .A2(new_n967), .A3(new_n880), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT109), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n975), .A2(new_n976), .A3(new_n943), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n973), .A2(new_n945), .A3(new_n974), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n971), .A2(new_n977), .A3(new_n916), .A4(new_n978), .ZN(new_n979));
  NAND4_X1  g554(.A1(new_n927), .A2(KEYINPUT41), .A3(new_n924), .A4(new_n928), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n945), .A2(new_n930), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n982), .B1(new_n968), .B2(new_n969), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n983), .A2(new_n978), .A3(KEYINPUT111), .ZN(new_n984));
  AND3_X1   g559(.A1(new_n911), .A2(new_n915), .A3(KEYINPUT110), .ZN(new_n985));
  AOI21_X1  g560(.A(KEYINPUT110), .B1(new_n911), .B2(new_n915), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT111), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n975), .A2(new_n988), .A3(new_n982), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n984), .A2(new_n987), .A3(new_n989), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n979), .A2(new_n990), .A3(new_n888), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(KEYINPUT43), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n971), .A2(new_n978), .A3(new_n977), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(new_n987), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n994), .A2(new_n888), .A3(new_n979), .ZN(new_n995));
  OAI211_X1 g570(.A(new_n992), .B(KEYINPUT44), .C1(new_n995), .C2(KEYINPUT43), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT43), .ZN(new_n997));
  AND4_X1   g572(.A1(new_n997), .A2(new_n979), .A3(new_n990), .A4(new_n888), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n998), .B1(new_n995), .B2(KEYINPUT43), .ZN(new_n999));
  XNOR2_X1  g574(.A(KEYINPUT108), .B(KEYINPUT44), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n996), .B1(new_n999), .B2(new_n1000), .ZN(G397));
  INV_X1    g576(.A(G1384), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n495), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT45), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  XOR2_X1   g580(.A(KEYINPUT112), .B(G40), .Z(new_n1006));
  INV_X1    g581(.A(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(G160), .A2(new_n1007), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n1005), .A2(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g584(.A(new_n773), .B(G1996), .ZN(new_n1010));
  INV_X1    g585(.A(G2067), .ZN(new_n1011));
  XNOR2_X1  g586(.A(new_n805), .B(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(new_n1009), .ZN(new_n1014));
  XNOR2_X1  g589(.A(new_n1014), .B(KEYINPUT113), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n743), .A2(new_n750), .A3(new_n747), .ZN(new_n1016));
  XOR2_X1   g591(.A(new_n1016), .B(KEYINPUT126), .Z(new_n1017));
  NAND2_X1  g592(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1018), .B1(G2067), .B2(new_n805), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1009), .B1(new_n1019), .B2(KEYINPUT127), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1020), .B1(KEYINPUT127), .B2(new_n1019), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1009), .ZN(new_n1022));
  OR3_X1    g597(.A1(new_n1022), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1023));
  OAI21_X1  g598(.A(KEYINPUT46), .B1(new_n1022), .B2(G1996), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1012), .A2(new_n773), .ZN(new_n1025));
  AOI22_X1  g600(.A1(new_n1023), .A2(new_n1024), .B1(new_n1009), .B2(new_n1025), .ZN(new_n1026));
  XNOR2_X1  g601(.A(new_n1026), .B(KEYINPUT47), .ZN(new_n1027));
  XNOR2_X1  g602(.A(new_n748), .B(new_n750), .ZN(new_n1028));
  XOR2_X1   g603(.A(new_n1028), .B(KEYINPUT114), .Z(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(new_n1009), .ZN(new_n1030));
  AND2_X1   g605(.A1(new_n1030), .A2(new_n1015), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1009), .A2(new_n732), .A3(new_n737), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT48), .ZN(new_n1033));
  OR2_X1    g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1035));
  AND3_X1   g610(.A1(new_n1031), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  NOR3_X1   g611(.A1(new_n1021), .A2(new_n1027), .A3(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(G305), .A2(G1981), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n695), .A2(new_n704), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT49), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1038), .A2(KEYINPUT49), .A3(new_n1039), .ZN(new_n1043));
  AND2_X1   g618(.A1(new_n495), .A2(new_n1002), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1008), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(G8), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1042), .A2(new_n1043), .A3(new_n1048), .ZN(new_n1049));
  NOR2_X1   g624(.A1(G288), .A2(G1976), .ZN(new_n1050));
  AOI22_X1  g625(.A1(new_n1049), .A2(new_n1050), .B1(new_n704), .B2(new_n695), .ZN(new_n1051));
  OR2_X1    g626(.A1(new_n1051), .A2(KEYINPUT117), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1051), .A2(KEYINPUT117), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1052), .A2(new_n1048), .A3(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n495), .A2(KEYINPUT45), .A3(new_n1002), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1005), .A2(new_n1045), .A3(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(new_n710), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT115), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1003), .A2(KEYINPUT50), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT50), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n495), .A2(new_n1060), .A3(new_n1002), .ZN(new_n1061));
  AND3_X1   g636(.A1(new_n1059), .A2(new_n1045), .A3(new_n1061), .ZN(new_n1062));
  AOI22_X1  g637(.A1(new_n1057), .A2(new_n1058), .B1(new_n1062), .B2(new_n788), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1063), .B1(new_n1058), .B2(new_n1057), .ZN(new_n1064));
  INV_X1    g639(.A(G8), .ZN(new_n1065));
  NOR2_X1   g640(.A1(G166), .A2(new_n1065), .ZN(new_n1066));
  XNOR2_X1  g641(.A(new_n1066), .B(KEYINPUT55), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1064), .A2(G8), .A3(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(G1976), .ZN(new_n1069));
  OAI211_X1 g644(.A(new_n1046), .B(G8), .C1(new_n1069), .C2(G288), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT52), .ZN(new_n1072));
  OAI21_X1  g647(.A(KEYINPUT116), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT116), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1070), .A2(new_n1074), .A3(KEYINPUT52), .ZN(new_n1075));
  AOI21_X1  g650(.A(KEYINPUT52), .B1(G288), .B2(new_n1069), .ZN(new_n1076));
  AOI22_X1  g651(.A1(new_n1073), .A2(new_n1075), .B1(new_n1071), .B2(new_n1076), .ZN(new_n1077));
  AND3_X1   g652(.A1(new_n1005), .A2(new_n1045), .A3(new_n1055), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1008), .B1(new_n1003), .B2(KEYINPUT50), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(new_n1061), .ZN(new_n1080));
  OAI22_X1  g655(.A1(new_n1078), .A2(G1966), .B1(new_n1080), .B2(G2084), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(G8), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT63), .ZN(new_n1083));
  NOR3_X1   g658(.A1(new_n1082), .A2(new_n1083), .A3(G286), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1068), .A2(new_n1049), .A3(new_n1077), .A4(new_n1084), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1067), .B1(new_n1064), .B2(G8), .ZN(new_n1086));
  OAI21_X1  g661(.A(KEYINPUT63), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  AND2_X1   g662(.A1(new_n1077), .A2(new_n1049), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1068), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1054), .A2(new_n1087), .A3(new_n1090), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1045), .A2(new_n1002), .A3(new_n1011), .A4(new_n495), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(KEYINPUT121), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT121), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1044), .A2(new_n1094), .A3(new_n1011), .A4(new_n1045), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1096), .B1(G1348), .B2(new_n1062), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT60), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n599), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(G1348), .ZN(new_n1100));
  AOI22_X1  g675(.A1(new_n1080), .A2(new_n1100), .B1(new_n1093), .B2(new_n1095), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1101), .A2(KEYINPUT60), .A3(new_n613), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1099), .A2(new_n1102), .A3(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT61), .ZN(new_n1105));
  AOI21_X1  g680(.A(KEYINPUT57), .B1(new_n560), .B2(KEYINPUT119), .ZN(new_n1106));
  XNOR2_X1  g681(.A(G299), .B(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT118), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1061), .A2(new_n1108), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n495), .A2(KEYINPUT118), .A3(new_n1060), .A4(new_n1002), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1111), .A2(new_n1079), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1112), .A2(new_n766), .ZN(new_n1113));
  XNOR2_X1  g688(.A(KEYINPUT120), .B(KEYINPUT56), .ZN(new_n1114));
  XNOR2_X1  g689(.A(new_n1114), .B(new_n822), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1078), .A2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1107), .B1(new_n1113), .B2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g692(.A(G1956), .B1(new_n1111), .B2(new_n1079), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1115), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1056), .A2(new_n1119), .ZN(new_n1120));
  XNOR2_X1  g695(.A(new_n608), .B(new_n1106), .ZN(new_n1121));
  NOR3_X1   g696(.A1(new_n1118), .A2(new_n1120), .A3(new_n1121), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1105), .B1(new_n1117), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT59), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(KEYINPUT122), .ZN(new_n1125));
  XOR2_X1   g700(.A(KEYINPUT58), .B(G1341), .Z(new_n1126));
  NAND2_X1  g701(.A1(new_n1046), .A2(new_n1126), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1127), .B1(new_n1056), .B2(G1996), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1125), .B1(new_n1128), .B2(new_n550), .ZN(new_n1129));
  AND2_X1   g704(.A1(new_n1128), .A2(new_n550), .ZN(new_n1130));
  XNOR2_X1  g705(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1129), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1113), .A2(new_n1116), .A3(new_n1107), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1121), .B1(new_n1118), .B2(new_n1120), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1133), .A2(KEYINPUT61), .A3(new_n1134), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1104), .A2(new_n1123), .A3(new_n1132), .A4(new_n1135), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1101), .A2(new_n599), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1133), .B1(new_n1117), .B2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(G1966), .ZN(new_n1140));
  AOI22_X1  g715(.A1(new_n1062), .A2(new_n798), .B1(new_n1056), .B2(new_n1140), .ZN(new_n1141));
  NOR2_X1   g716(.A1(G168), .A2(new_n1065), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1142), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1144));
  OAI21_X1  g719(.A(KEYINPUT51), .B1(new_n1142), .B2(KEYINPUT123), .ZN(new_n1145));
  OAI211_X1 g720(.A(new_n1143), .B(new_n1145), .C1(new_n1141), .C2(new_n1065), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1145), .ZN(new_n1147));
  OAI211_X1 g722(.A(G8), .B(new_n1147), .C1(new_n1081), .C2(G286), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1144), .B1(new_n1146), .B2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT53), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1150), .A2(G2078), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1078), .A2(new_n1151), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1150), .B1(new_n1056), .B2(G2078), .ZN(new_n1153));
  XNOR2_X1  g728(.A(KEYINPUT124), .B(G1961), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1080), .A2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1152), .A2(new_n1153), .A3(new_n1155), .ZN(new_n1156));
  XOR2_X1   g731(.A(G171), .B(KEYINPUT54), .Z(new_n1157));
  AND2_X1   g732(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1153), .A2(new_n1155), .ZN(new_n1159));
  AND3_X1   g734(.A1(G160), .A2(G40), .A3(new_n1151), .ZN(new_n1160));
  AND3_X1   g735(.A1(new_n1005), .A2(new_n1055), .A3(new_n1160), .ZN(new_n1161));
  NOR3_X1   g736(.A1(new_n1157), .A2(new_n1159), .A3(new_n1161), .ZN(new_n1162));
  NOR3_X1   g737(.A1(new_n1149), .A2(new_n1158), .A3(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1139), .A2(new_n1163), .ZN(new_n1164));
  AND2_X1   g739(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1165));
  OAI211_X1 g740(.A(KEYINPUT125), .B(KEYINPUT62), .C1(new_n1165), .C2(new_n1144), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT125), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT62), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1167), .B1(new_n1149), .B2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1156), .A2(G171), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1170), .B1(new_n1149), .B2(new_n1168), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1166), .A2(new_n1169), .A3(new_n1171), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1082), .A2(G286), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1173), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1164), .A2(new_n1172), .A3(new_n1174), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1111), .A2(new_n788), .A3(new_n1079), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1065), .B1(new_n1176), .B2(new_n1057), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1088), .B1(new_n1067), .B2(new_n1177), .ZN(new_n1178));
  NOR2_X1   g753(.A1(new_n1178), .A2(new_n1089), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1091), .B1(new_n1175), .B2(new_n1179), .ZN(new_n1180));
  XNOR2_X1  g755(.A(new_n732), .B(G1986), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1031), .B1(new_n1022), .B2(new_n1181), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n1037), .B1(new_n1180), .B2(new_n1182), .ZN(G329));
  assign    G231 = 1'b0;
  OR4_X1    g758(.A1(new_n459), .A2(G227), .A3(G229), .A4(G401), .ZN(new_n1185));
  NOR2_X1   g759(.A1(new_n1185), .A2(new_n906), .ZN(new_n1186));
  INV_X1    g760(.A(new_n1186), .ZN(new_n1187));
  NOR2_X1   g761(.A1(new_n1187), .A2(new_n999), .ZN(G308));
  AND2_X1   g762(.A1(new_n995), .A2(KEYINPUT43), .ZN(new_n1189));
  OAI21_X1  g763(.A(new_n1186), .B1(new_n1189), .B2(new_n998), .ZN(G225));
endmodule


