

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823;

  NAND2_X1 U376 ( .A1(n489), .A2(n487), .ZN(n486) );
  BUF_X1 U377 ( .A(n652), .Z(n355) );
  XNOR2_X1 U378 ( .A(n649), .B(KEYINPUT33), .ZN(n792) );
  XNOR2_X1 U379 ( .A(n529), .B(n528), .ZN(n640) );
  BUF_X1 U380 ( .A(G116), .Z(n709) );
  INV_X1 U381 ( .A(G210), .ZN(n557) );
  NAND2_X1 U382 ( .A1(G237), .A2(G234), .ZN(n533) );
  XNOR2_X1 U383 ( .A(G113), .B(KEYINPUT75), .ZN(n495) );
  XNOR2_X1 U384 ( .A(n435), .B(n475), .ZN(n683) );
  NAND2_X1 U385 ( .A1(n683), .A2(n631), .ZN(n456) );
  NAND2_X4 U386 ( .A1(n693), .A2(G953), .ZN(n736) );
  XNOR2_X2 U387 ( .A(n429), .B(n670), .ZN(n671) );
  XOR2_X2 U388 ( .A(n719), .B(KEYINPUT59), .Z(n720) );
  XNOR2_X2 U389 ( .A(n688), .B(n690), .ZN(n691) );
  XNOR2_X2 U390 ( .A(n432), .B(n712), .ZN(n714) );
  XNOR2_X2 U391 ( .A(n356), .B(n555), .ZN(n687) );
  XNOR2_X2 U392 ( .A(n389), .B(n807), .ZN(n356) );
  NAND2_X2 U393 ( .A1(n464), .A2(n462), .ZN(n732) );
  XNOR2_X2 U394 ( .A(n357), .B(n493), .ZN(n425) );
  NAND2_X2 U395 ( .A1(n671), .A2(n672), .ZN(n357) );
  AND2_X2 U396 ( .A1(n411), .A2(n414), .ZN(n412) );
  XNOR2_X1 U397 ( .A(G137), .B(KEYINPUT5), .ZN(n497) );
  INV_X1 U398 ( .A(KEYINPUT15), .ZN(n522) );
  INV_X1 U399 ( .A(G902), .ZN(n520) );
  BUF_X1 U400 ( .A(G107), .Z(n450) );
  INV_X1 U401 ( .A(G953), .ZN(n504) );
  BUF_X1 U402 ( .A(G146), .Z(n360) );
  XNOR2_X1 U403 ( .A(KEYINPUT114), .B(KEYINPUT41), .ZN(n358) );
  NAND2_X2 U404 ( .A1(n421), .A2(n676), .ZN(n420) );
  NAND2_X2 U405 ( .A1(n380), .A2(n377), .ZN(n794) );
  AND2_X2 U406 ( .A1(n382), .A2(n381), .ZN(n380) );
  AND2_X2 U407 ( .A1(n539), .A2(n593), .ZN(n540) );
  XNOR2_X2 U408 ( .A(n477), .B(G119), .ZN(n496) );
  XNOR2_X1 U409 ( .A(n430), .B(KEYINPUT45), .ZN(n677) );
  NAND2_X1 U410 ( .A1(n379), .A2(n378), .ZN(n377) );
  NOR2_X1 U411 ( .A1(n763), .A2(n358), .ZN(n378) );
  OR2_X1 U412 ( .A1(n687), .A2(n669), .ZN(n388) );
  INV_X1 U413 ( .A(KEYINPUT109), .ZN(n457) );
  INV_X1 U414 ( .A(KEYINPUT6), .ZN(n458) );
  NOR2_X1 U415 ( .A1(n399), .A2(n398), .ZN(n409) );
  AND2_X1 U416 ( .A1(n466), .A2(n403), .ZN(n464) );
  NAND2_X1 U417 ( .A1(n763), .A2(n358), .ZN(n381) );
  NAND2_X1 U418 ( .A1(n639), .A2(n638), .ZN(n439) );
  BUF_X1 U419 ( .A(n772), .Z(n451) );
  AND2_X1 U420 ( .A1(n373), .A2(n387), .ZN(n386) );
  INV_X1 U421 ( .A(n560), .ZN(n359) );
  INV_X1 U422 ( .A(n669), .ZN(n385) );
  NOR2_X1 U423 ( .A1(n510), .A2(G953), .ZN(n513) );
  INV_X1 U424 ( .A(G234), .ZN(n510) );
  NOR2_X2 U425 ( .A1(G902), .A2(G237), .ZN(n502) );
  XNOR2_X1 U426 ( .A(G137), .B(G140), .ZN(n516) );
  INV_X2 U427 ( .A(G104), .ZN(n695) );
  XNOR2_X1 U428 ( .A(G128), .B(G143), .ZN(n547) );
  NOR2_X1 U429 ( .A1(n772), .A2(n361), .ZN(n649) );
  NAND2_X1 U430 ( .A1(n362), .A2(n659), .ZN(n361) );
  INV_X1 U431 ( .A(n652), .ZN(n362) );
  NAND2_X1 U432 ( .A1(n363), .A2(n407), .ZN(n413) );
  NAND2_X1 U433 ( .A1(n444), .A2(n443), .ZN(n363) );
  XNOR2_X1 U434 ( .A(n549), .B(n548), .ZN(n552) );
  XNOR2_X1 U435 ( .A(n449), .B(n507), .ZN(n739) );
  NAND2_X1 U436 ( .A1(n364), .A2(G472), .ZN(n715) );
  NAND2_X1 U437 ( .A1(n364), .A2(G478), .ZN(n735) );
  XNOR2_X1 U438 ( .A(n392), .B(KEYINPUT65), .ZN(n364) );
  NAND2_X1 U439 ( .A1(n365), .A2(G475), .ZN(n721) );
  NAND2_X1 U440 ( .A1(n365), .A2(G210), .ZN(n692) );
  XNOR2_X1 U441 ( .A(n686), .B(KEYINPUT65), .ZN(n365) );
  XNOR2_X1 U442 ( .A(n366), .B(KEYINPUT100), .ZN(n367) );
  XNOR2_X2 U443 ( .A(G110), .B(KEYINPUT24), .ZN(n366) );
  XNOR2_X1 U444 ( .A(n368), .B(n367), .ZN(n509) );
  XNOR2_X1 U445 ( .A(n370), .B(n369), .ZN(n368) );
  XNOR2_X2 U446 ( .A(G119), .B(KEYINPUT23), .ZN(n369) );
  XNOR2_X2 U447 ( .A(G128), .B(KEYINPUT86), .ZN(n370) );
  XNOR2_X2 U448 ( .A(n371), .B(n522), .ZN(n673) );
  XNOR2_X2 U449 ( .A(G902), .B(KEYINPUT93), .ZN(n371) );
  NAND2_X1 U450 ( .A1(n687), .A2(n560), .ZN(n373) );
  XNOR2_X2 U451 ( .A(KEYINPUT70), .B(KEYINPUT71), .ZN(n499) );
  XNOR2_X2 U452 ( .A(n375), .B(n564), .ZN(n815) );
  XNOR2_X2 U453 ( .A(n374), .B(G134), .ZN(n564) );
  XNOR2_X2 U454 ( .A(G128), .B(G143), .ZN(n374) );
  XNOR2_X1 U455 ( .A(n583), .B(n408), .ZN(n375) );
  XNOR2_X2 U456 ( .A(KEYINPUT64), .B(KEYINPUT4), .ZN(n408) );
  XNOR2_X2 U457 ( .A(KEYINPUT73), .B(G131), .ZN(n583) );
  AND2_X1 U458 ( .A1(n376), .A2(n650), .ZN(n603) );
  XNOR2_X2 U459 ( .A(n376), .B(n561), .ZN(n590) );
  NAND2_X1 U460 ( .A1(n626), .A2(n376), .ZN(n610) );
  NOR2_X1 U461 ( .A1(n629), .A2(n376), .ZN(n630) );
  NAND2_X2 U462 ( .A1(n397), .A2(n396), .ZN(n376) );
  NAND2_X1 U463 ( .A1(n794), .A2(n616), .ZN(n600) );
  INV_X1 U464 ( .A(n767), .ZN(n379) );
  NAND2_X1 U465 ( .A1(n767), .A2(n358), .ZN(n382) );
  XNOR2_X2 U466 ( .A(n461), .B(n591), .ZN(n767) );
  NAND2_X1 U467 ( .A1(n386), .A2(n383), .ZN(n628) );
  OR2_X1 U468 ( .A1(n687), .A2(n384), .ZN(n383) );
  NAND2_X1 U469 ( .A1(n359), .A2(n385), .ZN(n384) );
  NAND2_X1 U470 ( .A1(n560), .A2(n669), .ZN(n387) );
  INV_X1 U471 ( .A(n388), .ZN(n395) );
  NAND2_X1 U472 ( .A1(n388), .A2(n560), .ZN(n396) );
  XNOR2_X1 U473 ( .A(n552), .B(n551), .ZN(n389) );
  XNOR2_X2 U474 ( .A(n544), .B(n543), .ZN(n807) );
  NAND2_X1 U475 ( .A1(n732), .A2(n710), .ZN(n399) );
  BUF_X1 U476 ( .A(n739), .Z(n390) );
  XNOR2_X1 U477 ( .A(n439), .B(KEYINPUT0), .ZN(n391) );
  XNOR2_X1 U478 ( .A(n439), .B(KEYINPUT0), .ZN(n442) );
  NAND2_X1 U479 ( .A1(n436), .A2(n401), .ZN(n435) );
  NAND2_X1 U480 ( .A1(n422), .A2(n420), .ZN(n392) );
  NAND2_X1 U481 ( .A1(n422), .A2(n420), .ZN(n393) );
  BUF_X1 U482 ( .A(n710), .Z(n394) );
  NAND2_X1 U483 ( .A1(n422), .A2(n420), .ZN(n686) );
  XNOR2_X2 U484 ( .A(n456), .B(n455), .ZN(n672) );
  NAND2_X2 U485 ( .A1(n589), .A2(n750), .ZN(n453) );
  XNOR2_X2 U486 ( .A(n454), .B(n406), .ZN(n589) );
  NAND2_X1 U487 ( .A1(n412), .A2(n413), .ZN(n430) );
  XNOR2_X2 U488 ( .A(n453), .B(KEYINPUT40), .ZN(n733) );
  NAND2_X1 U489 ( .A1(n395), .A2(n359), .ZN(n397) );
  AND2_X1 U490 ( .A1(KEYINPUT44), .A2(n668), .ZN(n398) );
  XNOR2_X1 U491 ( .A(n660), .B(n458), .ZN(n652) );
  XNOR2_X2 U492 ( .A(n452), .B(KEYINPUT22), .ZN(n441) );
  INV_X1 U493 ( .A(KEYINPUT80), .ZN(n501) );
  XNOR2_X1 U494 ( .A(n415), .B(n667), .ZN(n414) );
  NAND2_X1 U495 ( .A1(n445), .A2(n698), .ZN(n415) );
  NAND2_X1 U496 ( .A1(n666), .A2(n765), .ZN(n445) );
  NOR2_X1 U497 ( .A1(n731), .A2(n416), .ZN(n444) );
  XNOR2_X1 U498 ( .A(n601), .B(n476), .ZN(n436) );
  INV_X1 U499 ( .A(KEYINPUT46), .ZN(n476) );
  INV_X1 U500 ( .A(KEYINPUT90), .ZN(n455) );
  INV_X1 U501 ( .A(n425), .ZN(n421) );
  AND2_X1 U502 ( .A1(n488), .A2(n494), .ZN(n487) );
  XNOR2_X1 U503 ( .A(n438), .B(n405), .ZN(n437) );
  NOR2_X1 U504 ( .A1(n643), .A2(n760), .ZN(n438) );
  NAND2_X1 U505 ( .A1(n659), .A2(n459), .ZN(n656) );
  OR2_X1 U506 ( .A1(n643), .A2(n644), .ZN(n465) );
  AND2_X1 U507 ( .A1(n451), .A2(n467), .ZN(n446) );
  XNOR2_X1 U508 ( .A(n391), .B(KEYINPUT98), .ZN(n665) );
  NOR2_X2 U509 ( .A1(G953), .A2(G237), .ZN(n577) );
  NOR2_X1 U510 ( .A1(n777), .A2(n459), .ZN(n778) );
  XOR2_X1 U511 ( .A(KEYINPUT20), .B(KEYINPUT101), .Z(n523) );
  XOR2_X1 U512 ( .A(KEYINPUT102), .B(KEYINPUT11), .Z(n579) );
  XNOR2_X1 U513 ( .A(G140), .B(G122), .ZN(n575) );
  XNOR2_X1 U514 ( .A(n408), .B(n545), .ZN(n549) );
  INV_X1 U515 ( .A(KEYINPUT48), .ZN(n475) );
  XNOR2_X1 U516 ( .A(n661), .B(n605), .ZN(n772) );
  XNOR2_X1 U517 ( .A(n559), .B(KEYINPUT95), .ZN(n560) );
  XNOR2_X1 U518 ( .A(KEYINPUT16), .B(G122), .ZN(n543) );
  XOR2_X1 U519 ( .A(KEYINPUT7), .B(G122), .Z(n563) );
  XNOR2_X1 U520 ( .A(n542), .B(n541), .ZN(n604) );
  NAND2_X1 U521 ( .A1(n540), .A2(n437), .ZN(n542) );
  INV_X1 U522 ( .A(G472), .ZN(n460) );
  NAND2_X1 U523 ( .A1(n480), .A2(n400), .ZN(n478) );
  NAND2_X1 U524 ( .A1(n463), .A2(KEYINPUT68), .ZN(n462) );
  INV_X1 U525 ( .A(KEYINPUT56), .ZN(n447) );
  AND2_X1 U526 ( .A1(n485), .A2(n479), .ZN(n400) );
  AND2_X1 U527 ( .A1(n624), .A2(n623), .ZN(n401) );
  XOR2_X1 U528 ( .A(n813), .B(n505), .Z(n402) );
  AND2_X1 U529 ( .A1(n465), .A2(n595), .ZN(n403) );
  XOR2_X1 U530 ( .A(n675), .B(KEYINPUT69), .Z(n404) );
  XOR2_X1 U531 ( .A(n503), .B(KEYINPUT30), .Z(n405) );
  NOR2_X1 U532 ( .A1(n404), .A2(KEYINPUT66), .ZN(n423) );
  XOR2_X1 U533 ( .A(KEYINPUT77), .B(KEYINPUT39), .Z(n406) );
  INV_X1 U534 ( .A(KEYINPUT68), .ZN(n644) );
  INV_X1 U535 ( .A(KEYINPUT44), .ZN(n416) );
  OR2_X1 U536 ( .A1(KEYINPUT67), .A2(KEYINPUT44), .ZN(n407) );
  INV_X1 U537 ( .A(KEYINPUT66), .ZN(n676) );
  NAND2_X1 U538 ( .A1(n409), .A2(n410), .ZN(n411) );
  NAND2_X1 U539 ( .A1(n731), .A2(n668), .ZN(n410) );
  AND2_X2 U540 ( .A1(n419), .A2(n417), .ZN(n422) );
  NOR2_X1 U541 ( .A1(n418), .A2(n423), .ZN(n417) );
  INV_X1 U542 ( .A(n758), .ZN(n418) );
  NAND2_X1 U543 ( .A1(n425), .A2(n424), .ZN(n419) );
  AND2_X1 U544 ( .A1(n404), .A2(KEYINPUT66), .ZN(n424) );
  XNOR2_X1 U545 ( .A(n426), .B(n553), .ZN(n427) );
  XNOR2_X2 U546 ( .A(n499), .B(G101), .ZN(n553) );
  XNOR2_X1 U547 ( .A(n498), .B(n497), .ZN(n426) );
  XNOR2_X1 U548 ( .A(n544), .B(n427), .ZN(n428) );
  XNOR2_X1 U549 ( .A(n507), .B(n428), .ZN(n713) );
  XNOR2_X2 U550 ( .A(n815), .B(n360), .ZN(n507) );
  NAND2_X1 U551 ( .A1(n677), .A2(n669), .ZN(n429) );
  NAND2_X1 U552 ( .A1(n604), .A2(n590), .ZN(n454) );
  NAND2_X1 U553 ( .A1(n792), .A2(KEYINPUT34), .ZN(n488) );
  BUF_X1 U554 ( .A(n792), .Z(n431) );
  BUF_X1 U555 ( .A(n713), .Z(n432) );
  XNOR2_X1 U556 ( .A(n393), .B(KEYINPUT65), .ZN(n433) );
  XOR2_X1 U557 ( .A(KEYINPUT12), .B(G143), .Z(n576) );
  BUF_X1 U558 ( .A(n807), .Z(n434) );
  XNOR2_X2 U559 ( .A(n660), .B(n457), .ZN(n643) );
  NAND2_X1 U560 ( .A1(n399), .A2(n668), .ZN(n443) );
  XNOR2_X2 U561 ( .A(n440), .B(KEYINPUT19), .ZN(n639) );
  NAND2_X1 U562 ( .A1(n628), .A2(n615), .ZN(n440) );
  NAND2_X1 U563 ( .A1(n441), .A2(n648), .ZN(n468) );
  NAND2_X1 U564 ( .A1(n441), .A2(n451), .ZN(n463) );
  NAND2_X1 U565 ( .A1(n441), .A2(n446), .ZN(n466) );
  NOR2_X2 U566 ( .A1(n442), .A2(n642), .ZN(n452) );
  OR2_X1 U567 ( .A1(n391), .A2(n780), .ZN(n658) );
  INV_X1 U568 ( .A(n463), .ZN(n654) );
  XNOR2_X1 U569 ( .A(n448), .B(n447), .ZN(G51) );
  NAND2_X1 U570 ( .A1(n694), .A2(n736), .ZN(n448) );
  XNOR2_X1 U571 ( .A(n509), .B(n812), .ZN(n519) );
  XNOR2_X1 U572 ( .A(n506), .B(n402), .ZN(n449) );
  INV_X1 U573 ( .A(n431), .ZN(n491) );
  INV_X1 U574 ( .A(n485), .ZN(n483) );
  INV_X1 U575 ( .A(n672), .ZN(n755) );
  INV_X1 U576 ( .A(n660), .ZN(n459) );
  XNOR2_X2 U577 ( .A(n500), .B(n460), .ZN(n660) );
  INV_X1 U578 ( .A(n590), .ZN(n761) );
  NAND2_X1 U579 ( .A1(n590), .A2(n615), .ZN(n461) );
  AND2_X1 U580 ( .A1(n643), .A2(n644), .ZN(n467) );
  XNOR2_X2 U581 ( .A(n468), .B(KEYINPUT32), .ZN(n710) );
  NAND2_X1 U582 ( .A1(n472), .A2(n640), .ZN(n531) );
  XNOR2_X2 U583 ( .A(n471), .B(n470), .ZN(n472) );
  INV_X1 U584 ( .A(n526), .ZN(n470) );
  INV_X1 U585 ( .A(n472), .ZN(n595) );
  OR2_X2 U586 ( .A1(n725), .A2(G902), .ZN(n471) );
  INV_X1 U587 ( .A(n725), .ZN(n521) );
  XNOR2_X2 U588 ( .A(n805), .B(KEYINPUT76), .ZN(n554) );
  XNOR2_X2 U589 ( .A(n474), .B(n473), .ZN(n805) );
  XNOR2_X2 U590 ( .A(G110), .B(KEYINPUT81), .ZN(n473) );
  XNOR2_X2 U591 ( .A(G104), .B(G107), .ZN(n474) );
  OR2_X2 U592 ( .A1(n713), .A2(G902), .ZN(n500) );
  INV_X1 U593 ( .A(n589), .ZN(n625) );
  XNOR2_X2 U594 ( .A(G116), .B(KEYINPUT3), .ZN(n477) );
  NAND2_X2 U595 ( .A1(n481), .A2(n478), .ZN(n731) );
  INV_X1 U596 ( .A(KEYINPUT35), .ZN(n479) );
  INV_X1 U597 ( .A(n486), .ZN(n480) );
  AND2_X2 U598 ( .A1(n484), .A2(n482), .ZN(n481) );
  NAND2_X1 U599 ( .A1(n483), .A2(KEYINPUT35), .ZN(n482) );
  NAND2_X1 U600 ( .A1(n486), .A2(KEYINPUT35), .ZN(n484) );
  NAND2_X1 U601 ( .A1(n665), .A2(KEYINPUT34), .ZN(n485) );
  OR2_X2 U602 ( .A1(n665), .A2(n490), .ZN(n489) );
  NAND2_X1 U603 ( .A1(n793), .A2(n492), .ZN(n490) );
  INV_X1 U604 ( .A(KEYINPUT34), .ZN(n492) );
  INV_X1 U605 ( .A(KEYINPUT87), .ZN(n493) );
  XNOR2_X1 U606 ( .A(n519), .B(n518), .ZN(n725) );
  XOR2_X1 U607 ( .A(n650), .B(KEYINPUT83), .Z(n494) );
  INV_X1 U608 ( .A(KEYINPUT88), .ZN(n670) );
  XNOR2_X2 U609 ( .A(n496), .B(n495), .ZN(n544) );
  AND2_X1 U610 ( .A1(n577), .A2(G210), .ZN(n498) );
  XNOR2_X1 U611 ( .A(n502), .B(n501), .ZN(n556) );
  AND2_X1 U612 ( .A1(n556), .A2(G214), .ZN(n760) );
  INV_X1 U613 ( .A(KEYINPUT112), .ZN(n503) );
  XNOR2_X1 U614 ( .A(n554), .B(n553), .ZN(n506) );
  XNOR2_X1 U615 ( .A(n516), .B(KEYINPUT99), .ZN(n813) );
  NAND2_X1 U616 ( .A1(G227), .A2(n504), .ZN(n505) );
  OR2_X2 U617 ( .A1(n739), .A2(G902), .ZN(n508) );
  XNOR2_X2 U618 ( .A(n508), .B(G469), .ZN(n661) );
  XNOR2_X2 U619 ( .A(G125), .B(G146), .ZN(n545) );
  XNOR2_X1 U620 ( .A(n545), .B(KEYINPUT10), .ZN(n812) );
  INV_X1 U621 ( .A(KEYINPUT8), .ZN(n512) );
  INV_X1 U622 ( .A(n513), .ZN(n511) );
  NAND2_X1 U623 ( .A1(n512), .A2(n511), .ZN(n515) );
  NAND2_X1 U624 ( .A1(KEYINPUT8), .A2(n513), .ZN(n514) );
  NAND2_X1 U625 ( .A1(n515), .A2(n514), .ZN(n566) );
  NAND2_X1 U626 ( .A1(n566), .A2(G221), .ZN(n517) );
  XNOR2_X1 U627 ( .A(n517), .B(n516), .ZN(n518) );
  NAND2_X1 U628 ( .A1(n673), .A2(G234), .ZN(n524) );
  XNOR2_X1 U629 ( .A(n524), .B(n523), .ZN(n527) );
  NAND2_X1 U630 ( .A1(n527), .A2(G217), .ZN(n525) );
  XNOR2_X1 U631 ( .A(n525), .B(KEYINPUT25), .ZN(n526) );
  NAND2_X1 U632 ( .A1(n527), .A2(G221), .ZN(n529) );
  INV_X1 U633 ( .A(KEYINPUT21), .ZN(n528) );
  INV_X1 U634 ( .A(n640), .ZN(n774) );
  INV_X1 U635 ( .A(KEYINPUT72), .ZN(n530) );
  XNOR2_X2 U636 ( .A(n531), .B(n530), .ZN(n655) );
  NAND2_X1 U637 ( .A1(n661), .A2(n655), .ZN(n532) );
  XNOR2_X1 U638 ( .A(n532), .B(KEYINPUT111), .ZN(n539) );
  XNOR2_X1 U639 ( .A(n533), .B(KEYINPUT14), .ZN(n535) );
  NAND2_X1 U640 ( .A1(G952), .A2(n535), .ZN(n534) );
  XOR2_X1 U641 ( .A(KEYINPUT96), .B(n534), .Z(n788) );
  NAND2_X1 U642 ( .A1(n504), .A2(n788), .ZN(n635) );
  NAND2_X1 U643 ( .A1(G902), .A2(n535), .ZN(n632) );
  NOR2_X1 U644 ( .A1(G900), .A2(n632), .ZN(n536) );
  NAND2_X1 U645 ( .A1(G953), .A2(n536), .ZN(n537) );
  NAND2_X1 U646 ( .A1(n635), .A2(n537), .ZN(n538) );
  XNOR2_X1 U647 ( .A(n538), .B(KEYINPUT84), .ZN(n593) );
  INV_X1 U648 ( .A(KEYINPUT82), .ZN(n541) );
  XNOR2_X1 U649 ( .A(KEYINPUT94), .B(KEYINPUT17), .ZN(n546) );
  XNOR2_X1 U650 ( .A(n547), .B(n546), .ZN(n548) );
  NAND2_X1 U651 ( .A1(n504), .A2(G224), .ZN(n550) );
  XNOR2_X1 U652 ( .A(n550), .B(KEYINPUT18), .ZN(n551) );
  XOR2_X1 U653 ( .A(n554), .B(n553), .Z(n555) );
  INV_X1 U654 ( .A(n673), .ZN(n669) );
  INV_X1 U655 ( .A(n556), .ZN(n558) );
  OR2_X1 U656 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U657 ( .A(KEYINPUT79), .B(KEYINPUT38), .ZN(n561) );
  XNOR2_X1 U658 ( .A(n450), .B(n709), .ZN(n562) );
  XNOR2_X1 U659 ( .A(n563), .B(n562), .ZN(n565) );
  XNOR2_X1 U660 ( .A(n564), .B(n565), .ZN(n570) );
  XOR2_X1 U661 ( .A(KEYINPUT9), .B(KEYINPUT103), .Z(n568) );
  NAND2_X1 U662 ( .A1(G217), .A2(n566), .ZN(n567) );
  XNOR2_X1 U663 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U664 ( .A(n570), .B(n569), .ZN(n734) );
  NAND2_X1 U665 ( .A1(n734), .A2(n520), .ZN(n574) );
  XNOR2_X1 U666 ( .A(KEYINPUT104), .B(KEYINPUT105), .ZN(n572) );
  INV_X1 U667 ( .A(G478), .ZN(n571) );
  XNOR2_X1 U668 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U669 ( .A(n574), .B(n573), .ZN(n602) );
  XNOR2_X1 U670 ( .A(n576), .B(n575), .ZN(n581) );
  NAND2_X1 U671 ( .A1(n577), .A2(G214), .ZN(n578) );
  XNOR2_X1 U672 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U673 ( .A(n581), .B(n580), .ZN(n586) );
  XNOR2_X1 U674 ( .A(n695), .B(G113), .ZN(n582) );
  XNOR2_X1 U675 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U676 ( .A(n812), .B(n584), .ZN(n585) );
  XNOR2_X1 U677 ( .A(n586), .B(n585), .ZN(n719) );
  NAND2_X1 U678 ( .A1(n719), .A2(n520), .ZN(n588) );
  XOR2_X1 U679 ( .A(KEYINPUT13), .B(G475), .Z(n587) );
  XNOR2_X1 U680 ( .A(n588), .B(n587), .ZN(n617) );
  INV_X1 U681 ( .A(n617), .ZN(n592) );
  OR2_X1 U682 ( .A1(n602), .A2(n592), .ZN(n705) );
  INV_X1 U683 ( .A(KEYINPUT113), .ZN(n591) );
  INV_X1 U684 ( .A(n602), .ZN(n618) );
  AND2_X1 U685 ( .A1(n618), .A2(n592), .ZN(n641) );
  INV_X1 U686 ( .A(n641), .ZN(n763) );
  AND2_X1 U687 ( .A1(n640), .A2(n593), .ZN(n594) );
  XNOR2_X1 U688 ( .A(KEYINPUT74), .B(n594), .ZN(n606) );
  NAND2_X1 U689 ( .A1(n606), .A2(n595), .ZN(n596) );
  OR2_X1 U690 ( .A1(n643), .A2(n596), .ZN(n598) );
  INV_X1 U691 ( .A(KEYINPUT28), .ZN(n597) );
  XNOR2_X1 U692 ( .A(n598), .B(n597), .ZN(n599) );
  AND2_X1 U693 ( .A1(n661), .A2(n599), .ZN(n616) );
  XNOR2_X1 U694 ( .A(n600), .B(KEYINPUT42), .ZN(n729) );
  NAND2_X1 U695 ( .A1(n733), .A2(n729), .ZN(n601) );
  AND2_X1 U696 ( .A1(n602), .A2(n617), .ZN(n650) );
  AND2_X1 U697 ( .A1(n604), .A2(n603), .ZN(n749) );
  INV_X1 U698 ( .A(KEYINPUT78), .ZN(n620) );
  NAND2_X1 U699 ( .A1(n620), .A2(KEYINPUT47), .ZN(n613) );
  INV_X1 U700 ( .A(KEYINPUT1), .ZN(n605) );
  INV_X1 U701 ( .A(n760), .ZN(n615) );
  NAND2_X1 U702 ( .A1(n606), .A2(n615), .ZN(n607) );
  INV_X1 U703 ( .A(n595), .ZN(n645) );
  NOR2_X1 U704 ( .A1(n607), .A2(n645), .ZN(n608) );
  INV_X1 U705 ( .A(n705), .ZN(n750) );
  NAND2_X1 U706 ( .A1(n608), .A2(n750), .ZN(n609) );
  NOR2_X1 U707 ( .A1(n355), .A2(n609), .ZN(n626) );
  XNOR2_X1 U708 ( .A(KEYINPUT36), .B(n610), .ZN(n611) );
  NOR2_X1 U709 ( .A1(n451), .A2(n611), .ZN(n753) );
  INV_X1 U710 ( .A(n753), .ZN(n612) );
  NAND2_X1 U711 ( .A1(n613), .A2(n612), .ZN(n614) );
  NOR2_X1 U712 ( .A1(n749), .A2(n614), .ZN(n624) );
  AND2_X1 U713 ( .A1(n639), .A2(n616), .ZN(n751) );
  OR2_X1 U714 ( .A1(n618), .A2(n617), .ZN(n619) );
  XNOR2_X1 U715 ( .A(n619), .B(KEYINPUT106), .ZN(n744) );
  NAND2_X1 U716 ( .A1(n744), .A2(n705), .ZN(n765) );
  NAND2_X1 U717 ( .A1(n751), .A2(n765), .ZN(n622) );
  NOR2_X1 U718 ( .A1(n620), .A2(KEYINPUT47), .ZN(n621) );
  XNOR2_X1 U719 ( .A(n622), .B(n621), .ZN(n623) );
  NOR2_X1 U720 ( .A1(n625), .A2(n744), .ZN(n711) );
  NAND2_X1 U721 ( .A1(n451), .A2(n626), .ZN(n627) );
  XOR2_X1 U722 ( .A(KEYINPUT43), .B(n627), .Z(n629) );
  XNOR2_X1 U723 ( .A(n630), .B(KEYINPUT110), .ZN(n823) );
  NOR2_X1 U724 ( .A1(n711), .A2(n823), .ZN(n631) );
  INV_X1 U725 ( .A(n632), .ZN(n633) );
  NOR2_X1 U726 ( .A1(G898), .A2(n504), .ZN(n808) );
  NAND2_X1 U727 ( .A1(n633), .A2(n808), .ZN(n634) );
  NAND2_X1 U728 ( .A1(n635), .A2(n634), .ZN(n637) );
  INV_X1 U729 ( .A(KEYINPUT97), .ZN(n636) );
  XNOR2_X1 U730 ( .A(n637), .B(n636), .ZN(n638) );
  NAND2_X1 U731 ( .A1(n641), .A2(n640), .ZN(n642) );
  INV_X1 U732 ( .A(KEYINPUT107), .ZN(n646) );
  XNOR2_X1 U733 ( .A(n595), .B(n646), .ZN(n775) );
  NAND2_X1 U734 ( .A1(n355), .A2(n775), .ZN(n647) );
  NOR2_X1 U735 ( .A1(n647), .A2(n451), .ZN(n648) );
  INV_X1 U736 ( .A(KEYINPUT67), .ZN(n668) );
  INV_X1 U737 ( .A(n655), .ZN(n771) );
  INV_X1 U738 ( .A(n775), .ZN(n651) );
  AND2_X1 U739 ( .A1(n355), .A2(n651), .ZN(n653) );
  NAND2_X1 U740 ( .A1(n654), .A2(n653), .ZN(n698) );
  BUF_X2 U741 ( .A(n655), .Z(n659) );
  OR2_X1 U742 ( .A1(n772), .A2(n656), .ZN(n780) );
  INV_X1 U743 ( .A(KEYINPUT31), .ZN(n657) );
  XNOR2_X1 U744 ( .A(n658), .B(n657), .ZN(n707) );
  NAND2_X1 U745 ( .A1(n660), .A2(n659), .ZN(n663) );
  INV_X1 U746 ( .A(n661), .ZN(n662) );
  OR2_X1 U747 ( .A1(n663), .A2(n662), .ZN(n664) );
  OR2_X1 U748 ( .A1(n665), .A2(n664), .ZN(n702) );
  NAND2_X1 U749 ( .A1(n707), .A2(n702), .ZN(n666) );
  INV_X1 U750 ( .A(KEYINPUT108), .ZN(n667) );
  XNOR2_X1 U751 ( .A(n673), .B(KEYINPUT89), .ZN(n674) );
  NAND2_X1 U752 ( .A1(n674), .A2(KEYINPUT2), .ZN(n675) );
  BUF_X1 U753 ( .A(n677), .Z(n678) );
  INV_X1 U754 ( .A(n711), .ZN(n679) );
  NAND2_X1 U755 ( .A1(n679), .A2(KEYINPUT2), .ZN(n680) );
  XOR2_X1 U756 ( .A(KEYINPUT85), .B(n680), .Z(n681) );
  NOR2_X1 U757 ( .A1(n681), .A2(n823), .ZN(n682) );
  NAND2_X1 U758 ( .A1(n678), .A2(n682), .ZN(n685) );
  INV_X1 U759 ( .A(n683), .ZN(n684) );
  OR2_X1 U760 ( .A1(n685), .A2(n684), .ZN(n758) );
  BUF_X1 U761 ( .A(n687), .Z(n688) );
  XNOR2_X1 U762 ( .A(KEYINPUT123), .B(KEYINPUT54), .ZN(n689) );
  XOR2_X1 U763 ( .A(n689), .B(KEYINPUT55), .Z(n690) );
  XNOR2_X1 U764 ( .A(n692), .B(n691), .ZN(n694) );
  INV_X1 U765 ( .A(G952), .ZN(n693) );
  NOR2_X1 U766 ( .A1(n702), .A2(n705), .ZN(n696) );
  XNOR2_X1 U767 ( .A(n696), .B(n695), .ZN(G6) );
  XOR2_X1 U768 ( .A(G101), .B(KEYINPUT115), .Z(n697) );
  XNOR2_X1 U769 ( .A(n698), .B(n697), .ZN(G3) );
  XOR2_X1 U770 ( .A(KEYINPUT117), .B(KEYINPUT27), .Z(n700) );
  XNOR2_X1 U771 ( .A(n450), .B(KEYINPUT26), .ZN(n699) );
  XNOR2_X1 U772 ( .A(n700), .B(n699), .ZN(n701) );
  XOR2_X1 U773 ( .A(KEYINPUT116), .B(n701), .Z(n704) );
  NOR2_X1 U774 ( .A1(n702), .A2(n744), .ZN(n703) );
  XOR2_X1 U775 ( .A(n704), .B(n703), .Z(G9) );
  NOR2_X1 U776 ( .A1(n707), .A2(n705), .ZN(n706) );
  XOR2_X1 U777 ( .A(G113), .B(n706), .Z(G15) );
  NOR2_X1 U778 ( .A1(n707), .A2(n744), .ZN(n708) );
  XOR2_X1 U779 ( .A(n709), .B(n708), .Z(G18) );
  XNOR2_X1 U780 ( .A(n394), .B(G119), .ZN(G21) );
  XOR2_X1 U781 ( .A(G134), .B(n711), .Z(G36) );
  XOR2_X1 U782 ( .A(KEYINPUT92), .B(KEYINPUT62), .Z(n712) );
  XNOR2_X1 U783 ( .A(n715), .B(n714), .ZN(n716) );
  NAND2_X1 U784 ( .A1(n716), .A2(n736), .ZN(n718) );
  XOR2_X1 U785 ( .A(KEYINPUT91), .B(KEYINPUT63), .Z(n717) );
  XNOR2_X1 U786 ( .A(n718), .B(n717), .ZN(G57) );
  XNOR2_X1 U787 ( .A(n721), .B(n720), .ZN(n722) );
  NAND2_X1 U788 ( .A1(n722), .A2(n736), .ZN(n724) );
  XOR2_X1 U789 ( .A(KEYINPUT124), .B(KEYINPUT60), .Z(n723) );
  XNOR2_X1 U790 ( .A(n724), .B(n723), .ZN(G60) );
  NAND2_X1 U791 ( .A1(n433), .A2(G217), .ZN(n726) );
  XNOR2_X1 U792 ( .A(n726), .B(n521), .ZN(n727) );
  NAND2_X1 U793 ( .A1(n727), .A2(n736), .ZN(n728) );
  XNOR2_X1 U794 ( .A(n728), .B(KEYINPUT125), .ZN(G66) );
  XNOR2_X1 U795 ( .A(n729), .B(G137), .ZN(G39) );
  XNOR2_X1 U796 ( .A(G122), .B(KEYINPUT127), .ZN(n730) );
  XNOR2_X1 U797 ( .A(n731), .B(n730), .ZN(G24) );
  XNOR2_X1 U798 ( .A(n732), .B(G110), .ZN(G12) );
  XNOR2_X1 U799 ( .A(n733), .B(G131), .ZN(G33) );
  XOR2_X1 U800 ( .A(n735), .B(n734), .Z(n737) );
  INV_X1 U801 ( .A(n736), .ZN(n742) );
  NOR2_X1 U802 ( .A1(n737), .A2(n742), .ZN(G63) );
  NAND2_X1 U803 ( .A1(n433), .A2(G469), .ZN(n741) );
  XOR2_X1 U804 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n738) );
  XNOR2_X1 U805 ( .A(n390), .B(n738), .ZN(n740) );
  XNOR2_X1 U806 ( .A(n741), .B(n740), .ZN(n743) );
  NOR2_X1 U807 ( .A1(n743), .A2(n742), .ZN(G54) );
  XOR2_X1 U808 ( .A(KEYINPUT29), .B(KEYINPUT118), .Z(n747) );
  INV_X1 U809 ( .A(n744), .ZN(n745) );
  NAND2_X1 U810 ( .A1(n751), .A2(n745), .ZN(n746) );
  XNOR2_X1 U811 ( .A(n747), .B(n746), .ZN(n748) );
  XNOR2_X1 U812 ( .A(G128), .B(n748), .ZN(G30) );
  XOR2_X1 U813 ( .A(G143), .B(n749), .Z(G45) );
  NAND2_X1 U814 ( .A1(n751), .A2(n750), .ZN(n752) );
  XNOR2_X1 U815 ( .A(n752), .B(n360), .ZN(G48) );
  XNOR2_X1 U816 ( .A(G125), .B(n753), .ZN(n754) );
  XNOR2_X1 U817 ( .A(n754), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U818 ( .A(KEYINPUT53), .B(KEYINPUT122), .Z(n800) );
  INV_X1 U819 ( .A(n678), .ZN(n756) );
  NOR2_X1 U820 ( .A1(n755), .A2(n756), .ZN(n757) );
  OR2_X1 U821 ( .A1(n757), .A2(KEYINPUT2), .ZN(n759) );
  NAND2_X1 U822 ( .A1(n759), .A2(n758), .ZN(n791) );
  NAND2_X1 U823 ( .A1(n761), .A2(n760), .ZN(n762) );
  XOR2_X1 U824 ( .A(KEYINPUT120), .B(n762), .Z(n764) );
  NOR2_X1 U825 ( .A1(n764), .A2(n763), .ZN(n769) );
  INV_X1 U826 ( .A(n765), .ZN(n766) );
  NOR2_X1 U827 ( .A1(n767), .A2(n766), .ZN(n768) );
  NOR2_X1 U828 ( .A1(n769), .A2(n768), .ZN(n770) );
  NOR2_X1 U829 ( .A1(n770), .A2(n431), .ZN(n786) );
  NAND2_X1 U830 ( .A1(n451), .A2(n771), .ZN(n773) );
  XNOR2_X1 U831 ( .A(n773), .B(KEYINPUT50), .ZN(n779) );
  NAND2_X1 U832 ( .A1(n775), .A2(n774), .ZN(n776) );
  XNOR2_X1 U833 ( .A(n776), .B(KEYINPUT49), .ZN(n777) );
  NAND2_X1 U834 ( .A1(n779), .A2(n778), .ZN(n781) );
  NAND2_X1 U835 ( .A1(n781), .A2(n780), .ZN(n782) );
  XOR2_X1 U836 ( .A(KEYINPUT51), .B(n782), .Z(n783) );
  NAND2_X1 U837 ( .A1(n783), .A2(n794), .ZN(n784) );
  XNOR2_X1 U838 ( .A(n784), .B(KEYINPUT119), .ZN(n785) );
  NOR2_X1 U839 ( .A1(n786), .A2(n785), .ZN(n787) );
  XOR2_X1 U840 ( .A(KEYINPUT52), .B(n787), .Z(n789) );
  NAND2_X1 U841 ( .A1(n789), .A2(n788), .ZN(n790) );
  NAND2_X1 U842 ( .A1(n791), .A2(n790), .ZN(n797) );
  INV_X1 U843 ( .A(n792), .ZN(n793) );
  NAND2_X1 U844 ( .A1(n794), .A2(n491), .ZN(n795) );
  XNOR2_X1 U845 ( .A(n795), .B(KEYINPUT121), .ZN(n796) );
  NOR2_X1 U846 ( .A1(n797), .A2(n796), .ZN(n798) );
  NAND2_X1 U847 ( .A1(n798), .A2(n504), .ZN(n799) );
  XNOR2_X1 U848 ( .A(n800), .B(n799), .ZN(G75) );
  NAND2_X1 U849 ( .A1(n678), .A2(n504), .ZN(n804) );
  NAND2_X1 U850 ( .A1(G953), .A2(G224), .ZN(n801) );
  XNOR2_X1 U851 ( .A(KEYINPUT61), .B(n801), .ZN(n802) );
  NAND2_X1 U852 ( .A1(n802), .A2(G898), .ZN(n803) );
  NAND2_X1 U853 ( .A1(n804), .A2(n803), .ZN(n811) );
  XNOR2_X1 U854 ( .A(n805), .B(G101), .ZN(n806) );
  XNOR2_X1 U855 ( .A(n434), .B(n806), .ZN(n809) );
  NOR2_X1 U856 ( .A1(n809), .A2(n808), .ZN(n810) );
  XNOR2_X1 U857 ( .A(n811), .B(n810), .ZN(G69) );
  XOR2_X1 U858 ( .A(n813), .B(n812), .Z(n814) );
  XNOR2_X1 U859 ( .A(n815), .B(n814), .ZN(n817) );
  XNOR2_X1 U860 ( .A(n755), .B(n817), .ZN(n816) );
  NAND2_X1 U861 ( .A1(n816), .A2(n504), .ZN(n822) );
  XNOR2_X1 U862 ( .A(n817), .B(G227), .ZN(n818) );
  NAND2_X1 U863 ( .A1(n818), .A2(G900), .ZN(n819) );
  XNOR2_X1 U864 ( .A(KEYINPUT126), .B(n819), .ZN(n820) );
  NAND2_X1 U865 ( .A1(n820), .A2(G953), .ZN(n821) );
  NAND2_X1 U866 ( .A1(n822), .A2(n821), .ZN(G72) );
  XOR2_X1 U867 ( .A(G140), .B(n823), .Z(G42) );
endmodule

