

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732;

  NOR2_X1 U374 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U375 ( .A(G110), .B(KEYINPUT76), .ZN(n441) );
  INV_X1 U376 ( .A(G953), .ZN(n719) );
  XOR2_X1 U377 ( .A(KEYINPUT72), .B(G469), .Z(n352) );
  XNOR2_X1 U378 ( .A(n691), .B(n690), .ZN(n353) );
  NOR2_X2 U379 ( .A1(n635), .A2(n636), .ZN(n489) );
  XNOR2_X2 U380 ( .A(n420), .B(n454), .ZN(n517) );
  NOR2_X2 U381 ( .A1(n562), .A2(n453), .ZN(n420) );
  NOR2_X2 U382 ( .A1(n731), .A2(n730), .ZN(n589) );
  XNOR2_X2 U383 ( .A(n387), .B(n360), .ZN(n636) );
  NOR2_X2 U384 ( .A1(n652), .A2(n523), .ZN(n406) );
  AND2_X2 U385 ( .A1(n413), .A2(n412), .ZN(n695) );
  OR2_X1 U386 ( .A1(n629), .A2(n630), .ZN(n412) );
  XNOR2_X1 U387 ( .A(n421), .B(n368), .ZN(n562) );
  XNOR2_X1 U388 ( .A(n716), .B(G146), .ZN(n361) );
  XNOR2_X1 U389 ( .A(n701), .B(n443), .ZN(n486) );
  XNOR2_X1 U390 ( .A(n455), .B(n407), .ZN(n716) );
  XNOR2_X1 U391 ( .A(n496), .B(n411), .ZN(n455) );
  XNOR2_X1 U392 ( .A(n444), .B(G143), .ZN(n496) );
  XOR2_X1 U393 ( .A(G146), .B(G125), .Z(n469) );
  INV_X1 U394 ( .A(KEYINPUT1), .ZN(n360) );
  XNOR2_X1 U395 ( .A(n356), .B(n355), .ZN(G60) );
  XNOR2_X1 U396 ( .A(n358), .B(n353), .ZN(n357) );
  NAND2_X1 U397 ( .A1(n695), .A2(G475), .ZN(n358) );
  AND2_X1 U398 ( .A1(n602), .A2(n601), .ZN(n717) );
  NOR2_X1 U399 ( .A1(n594), .A2(n585), .ZN(n586) );
  NAND2_X1 U400 ( .A1(n359), .A2(n387), .ZN(n522) );
  NOR2_X1 U401 ( .A1(n658), .A2(n657), .ZN(n424) );
  AND2_X1 U402 ( .A1(n555), .A2(n653), .ZN(n421) );
  XNOR2_X1 U403 ( .A(n361), .B(n487), .ZN(n682) );
  XNOR2_X1 U404 ( .A(n469), .B(G140), .ZN(n470) );
  INV_X1 U405 ( .A(n374), .ZN(n442) );
  INV_X1 U406 ( .A(n699), .ZN(n354) );
  XNOR2_X1 U407 ( .A(G116), .B(G113), .ZN(n416) );
  XNOR2_X1 U408 ( .A(G104), .B(G107), .ZN(n374) );
  XNOR2_X1 U409 ( .A(G128), .B(KEYINPUT65), .ZN(n444) );
  INV_X1 U410 ( .A(KEYINPUT60), .ZN(n355) );
  NAND2_X1 U411 ( .A1(n357), .A2(n354), .ZN(n356) );
  INV_X1 U412 ( .A(n635), .ZN(n359) );
  XNOR2_X2 U413 ( .A(n488), .B(n352), .ZN(n387) );
  XNOR2_X1 U414 ( .A(n361), .B(n462), .ZN(n606) );
  XNOR2_X1 U415 ( .A(n379), .B(n378), .ZN(n633) );
  XOR2_X1 U416 ( .A(KEYINPUT68), .B(G101), .Z(n456) );
  XNOR2_X1 U417 ( .A(n503), .B(n408), .ZN(n407) );
  XNOR2_X1 U418 ( .A(n409), .B(G137), .ZN(n408) );
  INV_X1 U419 ( .A(G134), .ZN(n409) );
  XNOR2_X1 U420 ( .A(n439), .B(n438), .ZN(n457) );
  XNOR2_X1 U421 ( .A(n416), .B(n437), .ZN(n439) );
  XOR2_X1 U422 ( .A(KEYINPUT70), .B(KEYINPUT10), .Z(n471) );
  NOR2_X1 U423 ( .A1(n606), .A2(G902), .ZN(n464) );
  NAND2_X1 U424 ( .A1(n695), .A2(G472), .ZN(n403) );
  NOR2_X1 U425 ( .A1(n627), .A2(n600), .ZN(n601) );
  AND2_X1 U426 ( .A1(n591), .A2(n366), .ZN(n383) );
  AND2_X1 U427 ( .A1(n601), .A2(n465), .ZN(n426) );
  XOR2_X1 U428 ( .A(KEYINPUT79), .B(G140), .Z(n484) );
  XNOR2_X1 U429 ( .A(n514), .B(n513), .ZN(n526) );
  NOR2_X1 U430 ( .A1(n559), .A2(n394), .ZN(n567) );
  NAND2_X1 U431 ( .A1(n396), .A2(n395), .ZN(n394) );
  INV_X1 U432 ( .A(n560), .ZN(n395) );
  INV_X1 U433 ( .A(n639), .ZN(n396) );
  INV_X1 U434 ( .A(n517), .ZN(n523) );
  XNOR2_X1 U435 ( .A(n551), .B(n373), .ZN(n568) );
  INV_X1 U436 ( .A(KEYINPUT6), .ZN(n373) );
  XNOR2_X1 U437 ( .A(n510), .B(n431), .ZN(n511) );
  XOR2_X1 U438 ( .A(KEYINPUT12), .B(G122), .Z(n505) );
  XNOR2_X1 U439 ( .A(n584), .B(n583), .ZN(n594) );
  XNOR2_X1 U440 ( .A(n518), .B(KEYINPUT22), .ZN(n534) );
  INV_X1 U441 ( .A(KEYINPUT69), .ZN(n378) );
  NOR2_X1 U442 ( .A1(n640), .A2(n639), .ZN(n379) );
  XNOR2_X1 U443 ( .A(G478), .B(n502), .ZN(n528) );
  NOR2_X2 U444 ( .A1(n534), .A2(n573), .ZN(n537) );
  XNOR2_X1 U445 ( .A(n457), .B(n388), .ZN(n461) );
  XNOR2_X1 U446 ( .A(n377), .B(n477), .ZN(n697) );
  XNOR2_X1 U447 ( .A(n715), .B(n474), .ZN(n377) );
  NAND2_X1 U448 ( .A1(n414), .A2(n604), .ZN(n413) );
  NAND2_X1 U449 ( .A1(n617), .A2(n566), .ZN(n576) );
  XNOR2_X1 U450 ( .A(n659), .B(n397), .ZN(n419) );
  INV_X1 U451 ( .A(KEYINPUT82), .ZN(n397) );
  NAND2_X1 U452 ( .A1(n576), .A2(KEYINPUT47), .ZN(n575) );
  INV_X1 U453 ( .A(KEYINPUT103), .ZN(n381) );
  XNOR2_X1 U454 ( .A(KEYINPUT4), .B(KEYINPUT64), .ZN(n411) );
  AND2_X1 U455 ( .A1(n398), .A2(n585), .ZN(n659) );
  OR2_X1 U456 ( .A1(G237), .A2(G902), .ZN(n452) );
  XNOR2_X1 U457 ( .A(KEYINPUT100), .B(KEYINPUT102), .ZN(n429) );
  XNOR2_X1 U458 ( .A(n410), .B(G131), .ZN(n503) );
  INV_X1 U459 ( .A(KEYINPUT71), .ZN(n410) );
  NAND2_X1 U460 ( .A1(G234), .A2(G237), .ZN(n432) );
  XNOR2_X1 U461 ( .A(n515), .B(KEYINPUT104), .ZN(n657) );
  XNOR2_X1 U462 ( .A(n458), .B(n456), .ZN(n388) );
  NOR2_X1 U463 ( .A1(G953), .A2(G237), .ZN(n459) );
  XNOR2_X1 U464 ( .A(KEYINPUT16), .B(G122), .ZN(n440) );
  XNOR2_X1 U465 ( .A(G128), .B(G137), .ZN(n472) );
  XOR2_X1 U466 ( .A(G110), .B(G119), .Z(n473) );
  XNOR2_X1 U467 ( .A(n430), .B(n428), .ZN(n498) );
  XNOR2_X1 U468 ( .A(n495), .B(n429), .ZN(n428) );
  XNOR2_X1 U469 ( .A(n494), .B(n493), .ZN(n430) );
  XNOR2_X1 U470 ( .A(G134), .B(G107), .ZN(n495) );
  XNOR2_X1 U471 ( .A(n392), .B(n391), .ZN(n499) );
  INV_X1 U472 ( .A(KEYINPUT8), .ZN(n391) );
  NAND2_X1 U473 ( .A1(n719), .A2(G234), .ZN(n392) );
  INV_X1 U474 ( .A(KEYINPUT83), .ZN(n427) );
  BUF_X1 U475 ( .A(n652), .Z(n670) );
  AND2_X1 U476 ( .A1(n554), .A2(n386), .ZN(n582) );
  AND2_X1 U477 ( .A1(n422), .A2(n387), .ZN(n587) );
  XNOR2_X1 U478 ( .A(n393), .B(n561), .ZN(n422) );
  NAND2_X1 U479 ( .A1(n551), .A2(n567), .ZN(n393) );
  XNOR2_X1 U480 ( .A(n400), .B(n399), .ZN(n691) );
  XNOR2_X1 U481 ( .A(n506), .B(n364), .ZN(n399) );
  XNOR2_X1 U482 ( .A(n715), .B(n511), .ZN(n400) );
  NOR2_X1 U483 ( .A1(n598), .A2(n595), .ZN(n572) );
  XNOR2_X1 U484 ( .A(n406), .B(n367), .ZN(n405) );
  XNOR2_X1 U485 ( .A(n535), .B(n376), .ZN(n729) );
  XNOR2_X1 U486 ( .A(KEYINPUT32), .B(KEYINPUT66), .ZN(n376) );
  OR2_X1 U487 ( .A1(n534), .A2(n533), .ZN(n535) );
  AND2_X1 U488 ( .A1(n587), .A2(n390), .ZN(n617) );
  INV_X1 U489 ( .A(n562), .ZN(n390) );
  XNOR2_X1 U490 ( .A(KEYINPUT106), .B(n538), .ZN(n732) );
  INV_X1 U491 ( .A(n585), .ZN(n619) );
  XNOR2_X1 U492 ( .A(n401), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U493 ( .A1(n402), .A2(n354), .ZN(n401) );
  XNOR2_X1 U494 ( .A(n403), .B(n369), .ZN(n402) );
  XNOR2_X1 U495 ( .A(n696), .B(n380), .ZN(n698) );
  XNOR2_X1 U496 ( .A(n697), .B(KEYINPUT122), .ZN(n380) );
  INV_X1 U497 ( .A(KEYINPUT56), .ZN(n384) );
  XOR2_X1 U498 ( .A(n556), .B(KEYINPUT80), .Z(n362) );
  XOR2_X1 U499 ( .A(n531), .B(KEYINPUT105), .Z(n363) );
  XOR2_X1 U500 ( .A(G143), .B(G104), .Z(n364) );
  NOR2_X1 U501 ( .A1(n527), .A2(n528), .ZN(n622) );
  INV_X1 U502 ( .A(n622), .ZN(n398) );
  AND2_X1 U503 ( .A1(n419), .A2(n645), .ZN(n365) );
  AND2_X1 U504 ( .A1(n616), .A2(n565), .ZN(n366) );
  XOR2_X1 U505 ( .A(KEYINPUT34), .B(KEYINPUT81), .Z(n367) );
  XOR2_X1 U506 ( .A(KEYINPUT19), .B(KEYINPUT67), .Z(n368) );
  XOR2_X1 U507 ( .A(n606), .B(n605), .Z(n369) );
  XNOR2_X1 U508 ( .A(n457), .B(n440), .ZN(n700) );
  XOR2_X1 U509 ( .A(n679), .B(n678), .Z(n370) );
  XOR2_X1 U510 ( .A(G902), .B(KEYINPUT15), .Z(n465) );
  NOR2_X1 U511 ( .A1(G952), .A2(n719), .ZN(n699) );
  XNOR2_X1 U512 ( .A(n371), .B(KEYINPUT85), .ZN(n545) );
  NAND2_X1 U513 ( .A1(n529), .A2(n530), .ZN(n371) );
  NAND2_X1 U514 ( .A1(n372), .A2(n545), .ZN(n546) );
  NAND2_X1 U515 ( .A1(n544), .A2(n543), .ZN(n372) );
  NAND2_X1 U516 ( .A1(n537), .A2(n536), .ZN(n538) );
  AND2_X1 U517 ( .A1(n590), .A2(n383), .ZN(n593) );
  AND2_X1 U518 ( .A1(n517), .A2(n633), .ZN(n520) );
  XNOR2_X1 U519 ( .A(n415), .B(n427), .ZN(n414) );
  XNOR2_X1 U520 ( .A(n382), .B(n381), .ZN(n375) );
  NOR2_X1 U521 ( .A1(n375), .A2(n607), .ZN(n529) );
  XNOR2_X2 U522 ( .A(n442), .B(n441), .ZN(n701) );
  NAND2_X1 U523 ( .A1(n418), .A2(n417), .ZN(n382) );
  NAND2_X1 U524 ( .A1(n654), .A2(n653), .ZN(n658) );
  XNOR2_X1 U525 ( .A(n486), .B(n455), .ZN(n389) );
  XNOR2_X1 U526 ( .A(n389), .B(n700), .ZN(n449) );
  XNOR2_X1 U527 ( .A(n385), .B(n384), .ZN(G51) );
  NAND2_X1 U528 ( .A1(n681), .A2(n354), .ZN(n385) );
  AND2_X1 U529 ( .A1(n633), .A2(n387), .ZN(n386) );
  XNOR2_X2 U530 ( .A(n470), .B(n471), .ZN(n715) );
  XNOR2_X2 U531 ( .A(n404), .B(KEYINPUT35), .ZN(n728) );
  NAND2_X1 U532 ( .A1(n405), .A2(n362), .ZN(n404) );
  NAND2_X1 U533 ( .A1(n717), .A2(n706), .ZN(n629) );
  NAND2_X1 U534 ( .A1(n425), .A2(n706), .ZN(n415) );
  AND2_X1 U535 ( .A1(n525), .A2(n645), .ZN(n609) );
  NAND2_X1 U536 ( .A1(n525), .A2(n365), .ZN(n417) );
  NAND2_X1 U537 ( .A1(n621), .A2(n419), .ZN(n418) );
  XNOR2_X2 U538 ( .A(n521), .B(KEYINPUT31), .ZN(n621) );
  NAND2_X1 U539 ( .A1(n631), .A2(n587), .ZN(n588) );
  XNOR2_X1 U540 ( .A(n424), .B(n423), .ZN(n631) );
  INV_X1 U541 ( .A(KEYINPUT41), .ZN(n423) );
  AND2_X1 U542 ( .A1(n602), .A2(n426), .ZN(n425) );
  XNOR2_X2 U543 ( .A(n546), .B(KEYINPUT45), .ZN(n706) );
  XNOR2_X1 U544 ( .A(n451), .B(n450), .ZN(n555) );
  XNOR2_X2 U545 ( .A(n482), .B(n481), .ZN(n640) );
  INV_X1 U546 ( .A(n555), .ZN(n598) );
  XOR2_X1 U547 ( .A(n509), .B(n508), .Z(n431) );
  XNOR2_X1 U548 ( .A(n542), .B(n539), .ZN(n540) );
  XNOR2_X1 U549 ( .A(n541), .B(n540), .ZN(n544) );
  INV_X1 U550 ( .A(KEYINPUT88), .ZN(n490) );
  INV_X1 U551 ( .A(n628), .ZN(n600) );
  XNOR2_X1 U552 ( .A(n490), .B(KEYINPUT33), .ZN(n491) );
  XNOR2_X1 U553 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U554 ( .A(n492), .B(n491), .ZN(n652) );
  XNOR2_X1 U555 ( .A(n512), .B(G475), .ZN(n513) );
  INV_X1 U556 ( .A(KEYINPUT39), .ZN(n583) );
  XNOR2_X1 U557 ( .A(n432), .B(KEYINPUT14), .ZN(n433) );
  NAND2_X1 U558 ( .A1(G952), .A2(n433), .ZN(n668) );
  NOR2_X1 U559 ( .A1(G953), .A2(n668), .ZN(n550) );
  NAND2_X1 U560 ( .A1(n433), .A2(G902), .ZN(n434) );
  XNOR2_X1 U561 ( .A(n434), .B(KEYINPUT91), .ZN(n547) );
  NOR2_X1 U562 ( .A1(G898), .A2(n719), .ZN(n705) );
  NAND2_X1 U563 ( .A1(n547), .A2(n705), .ZN(n435) );
  XOR2_X1 U564 ( .A(KEYINPUT92), .B(n435), .Z(n436) );
  NOR2_X1 U565 ( .A1(n550), .A2(n436), .ZN(n453) );
  INV_X1 U566 ( .A(KEYINPUT3), .ZN(n437) );
  XOR2_X1 U567 ( .A(KEYINPUT73), .B(G119), .Z(n438) );
  INV_X1 U568 ( .A(n456), .ZN(n443) );
  XOR2_X1 U569 ( .A(KEYINPUT18), .B(n469), .Z(n446) );
  NAND2_X1 U570 ( .A1(G224), .A2(n719), .ZN(n445) );
  XNOR2_X1 U571 ( .A(n446), .B(n445), .ZN(n447) );
  XOR2_X1 U572 ( .A(n447), .B(KEYINPUT17), .Z(n448) );
  XNOR2_X1 U573 ( .A(n449), .B(n448), .ZN(n679) );
  NOR2_X1 U574 ( .A1(n679), .A2(n465), .ZN(n451) );
  NAND2_X1 U575 ( .A1(G210), .A2(n452), .ZN(n450) );
  NAND2_X1 U576 ( .A1(G214), .A2(n452), .ZN(n653) );
  XOR2_X1 U577 ( .A(KEYINPUT87), .B(KEYINPUT0), .Z(n454) );
  XOR2_X1 U578 ( .A(KEYINPUT75), .B(KEYINPUT5), .Z(n458) );
  XOR2_X1 U579 ( .A(KEYINPUT77), .B(n459), .Z(n507) );
  NAND2_X1 U580 ( .A1(n507), .A2(G210), .ZN(n460) );
  XNOR2_X1 U581 ( .A(G472), .B(KEYINPUT95), .ZN(n463) );
  XNOR2_X2 U582 ( .A(n464), .B(n463), .ZN(n551) );
  XOR2_X1 U583 ( .A(KEYINPUT21), .B(KEYINPUT93), .Z(n468) );
  INV_X1 U584 ( .A(n465), .ZN(n603) );
  NAND2_X1 U585 ( .A1(n603), .A2(G234), .ZN(n466) );
  XNOR2_X1 U586 ( .A(n466), .B(KEYINPUT20), .ZN(n478) );
  NAND2_X1 U587 ( .A1(G221), .A2(n478), .ZN(n467) );
  XNOR2_X1 U588 ( .A(n468), .B(n467), .ZN(n639) );
  XNOR2_X1 U589 ( .A(n473), .B(n472), .ZN(n474) );
  XOR2_X1 U590 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n476) );
  NAND2_X1 U591 ( .A1(G221), .A2(n499), .ZN(n475) );
  XNOR2_X1 U592 ( .A(n476), .B(n475), .ZN(n477) );
  NOR2_X1 U593 ( .A1(n697), .A2(G902), .ZN(n482) );
  XOR2_X1 U594 ( .A(KEYINPUT25), .B(KEYINPUT78), .Z(n480) );
  NAND2_X1 U595 ( .A1(G217), .A2(n478), .ZN(n479) );
  XNOR2_X1 U596 ( .A(n480), .B(n479), .ZN(n481) );
  INV_X1 U597 ( .A(n633), .ZN(n635) );
  NAND2_X1 U598 ( .A1(G227), .A2(n719), .ZN(n483) );
  XNOR2_X1 U599 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U600 ( .A(n486), .B(n485), .ZN(n487) );
  NOR2_X1 U601 ( .A1(n682), .A2(G902), .ZN(n488) );
  NAND2_X1 U602 ( .A1(n568), .A2(n489), .ZN(n492) );
  XOR2_X1 U603 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n494) );
  XNOR2_X1 U604 ( .A(G116), .B(G122), .ZN(n493) );
  XNOR2_X1 U605 ( .A(n496), .B(KEYINPUT101), .ZN(n497) );
  XNOR2_X1 U606 ( .A(n498), .B(n497), .ZN(n501) );
  NAND2_X1 U607 ( .A1(n499), .A2(G217), .ZN(n500) );
  XOR2_X1 U608 ( .A(n501), .B(n500), .Z(n693) );
  NOR2_X1 U609 ( .A1(G902), .A2(n693), .ZN(n502) );
  XNOR2_X1 U610 ( .A(n503), .B(G113), .ZN(n504) );
  XNOR2_X1 U611 ( .A(n505), .B(n504), .ZN(n506) );
  NAND2_X1 U612 ( .A1(G214), .A2(n507), .ZN(n510) );
  XOR2_X1 U613 ( .A(KEYINPUT98), .B(KEYINPUT96), .Z(n509) );
  XNOR2_X1 U614 ( .A(KEYINPUT97), .B(KEYINPUT11), .ZN(n508) );
  NOR2_X1 U615 ( .A1(G902), .A2(n691), .ZN(n514) );
  XNOR2_X1 U616 ( .A(KEYINPUT99), .B(KEYINPUT13), .ZN(n512) );
  OR2_X1 U617 ( .A1(n528), .A2(n526), .ZN(n556) );
  NAND2_X1 U618 ( .A1(n728), .A2(KEYINPUT44), .ZN(n530) );
  INV_X1 U619 ( .A(n636), .ZN(n573) );
  NAND2_X1 U620 ( .A1(n526), .A2(n528), .ZN(n515) );
  NOR2_X1 U621 ( .A1(n639), .A2(n657), .ZN(n516) );
  NAND2_X1 U622 ( .A1(n517), .A2(n516), .ZN(n518) );
  INV_X1 U623 ( .A(n568), .ZN(n532) );
  NAND2_X1 U624 ( .A1(n537), .A2(n532), .ZN(n519) );
  NOR2_X1 U625 ( .A1(n640), .A2(n519), .ZN(n607) );
  INV_X1 U626 ( .A(n551), .ZN(n645) );
  NOR2_X1 U627 ( .A1(n645), .A2(n636), .ZN(n634) );
  NAND2_X1 U628 ( .A1(n520), .A2(n634), .ZN(n521) );
  XNOR2_X1 U629 ( .A(n524), .B(KEYINPUT94), .ZN(n525) );
  INV_X1 U630 ( .A(n526), .ZN(n527) );
  NAND2_X1 U631 ( .A1(n528), .A2(n527), .ZN(n585) );
  INV_X1 U632 ( .A(n640), .ZN(n559) );
  NOR2_X1 U633 ( .A1(n559), .A2(n636), .ZN(n531) );
  NAND2_X1 U634 ( .A1(n532), .A2(n363), .ZN(n533) );
  NOR2_X1 U635 ( .A1(n551), .A2(n559), .ZN(n536) );
  NAND2_X1 U636 ( .A1(n729), .A2(n732), .ZN(n541) );
  INV_X1 U637 ( .A(KEYINPUT44), .ZN(n542) );
  INV_X1 U638 ( .A(KEYINPUT86), .ZN(n539) );
  NAND2_X1 U639 ( .A1(n542), .A2(n728), .ZN(n543) );
  NAND2_X1 U640 ( .A1(G953), .A2(n547), .ZN(n548) );
  NOR2_X1 U641 ( .A1(G900), .A2(n548), .ZN(n549) );
  NOR2_X1 U642 ( .A1(n550), .A2(n549), .ZN(n560) );
  NAND2_X1 U643 ( .A1(n551), .A2(n653), .ZN(n552) );
  XNOR2_X1 U644 ( .A(KEYINPUT30), .B(n552), .ZN(n553) );
  NOR2_X1 U645 ( .A1(n560), .A2(n553), .ZN(n554) );
  NOR2_X1 U646 ( .A1(n598), .A2(n556), .ZN(n557) );
  NAND2_X1 U647 ( .A1(n582), .A2(n557), .ZN(n616) );
  XNOR2_X1 U648 ( .A(KEYINPUT28), .B(KEYINPUT109), .ZN(n558) );
  XNOR2_X1 U649 ( .A(n558), .B(KEYINPUT108), .ZN(n561) );
  INV_X1 U650 ( .A(n617), .ZN(n563) );
  NOR2_X1 U651 ( .A1(KEYINPUT82), .A2(n563), .ZN(n564) );
  NAND2_X1 U652 ( .A1(n659), .A2(n564), .ZN(n565) );
  INV_X1 U653 ( .A(n659), .ZN(n566) );
  INV_X1 U654 ( .A(n567), .ZN(n570) );
  NAND2_X1 U655 ( .A1(n619), .A2(n568), .ZN(n569) );
  NOR2_X1 U656 ( .A1(n570), .A2(n569), .ZN(n571) );
  NAND2_X1 U657 ( .A1(n571), .A2(n653), .ZN(n595) );
  XNOR2_X1 U658 ( .A(KEYINPUT36), .B(n572), .ZN(n574) );
  NAND2_X1 U659 ( .A1(n574), .A2(n573), .ZN(n624) );
  NAND2_X1 U660 ( .A1(n575), .A2(n624), .ZN(n580) );
  INV_X1 U661 ( .A(n576), .ZN(n577) );
  NAND2_X1 U662 ( .A1(KEYINPUT82), .A2(n577), .ZN(n578) );
  NOR2_X1 U663 ( .A1(KEYINPUT47), .A2(n578), .ZN(n579) );
  NOR2_X1 U664 ( .A1(n580), .A2(n579), .ZN(n591) );
  XNOR2_X1 U665 ( .A(KEYINPUT38), .B(KEYINPUT74), .ZN(n581) );
  XNOR2_X1 U666 ( .A(n581), .B(n598), .ZN(n654) );
  NAND2_X1 U667 ( .A1(n582), .A2(n654), .ZN(n584) );
  XNOR2_X1 U668 ( .A(n586), .B(KEYINPUT40), .ZN(n731) );
  XOR2_X1 U669 ( .A(KEYINPUT42), .B(n588), .Z(n730) );
  XNOR2_X1 U670 ( .A(n589), .B(KEYINPUT46), .ZN(n590) );
  XNOR2_X1 U671 ( .A(KEYINPUT48), .B(KEYINPUT84), .ZN(n592) );
  XNOR2_X1 U672 ( .A(n593), .B(n592), .ZN(n602) );
  NOR2_X1 U673 ( .A1(n594), .A2(n398), .ZN(n627) );
  XNOR2_X1 U674 ( .A(KEYINPUT107), .B(n595), .ZN(n596) );
  NAND2_X1 U675 ( .A1(n596), .A2(n636), .ZN(n597) );
  XNOR2_X1 U676 ( .A(n597), .B(KEYINPUT43), .ZN(n599) );
  NAND2_X1 U677 ( .A1(n599), .A2(n598), .ZN(n628) );
  INV_X1 U678 ( .A(KEYINPUT2), .ZN(n630) );
  OR2_X1 U679 ( .A1(n603), .A2(n630), .ZN(n604) );
  XOR2_X1 U680 ( .A(KEYINPUT62), .B(KEYINPUT89), .Z(n605) );
  XOR2_X1 U681 ( .A(G101), .B(n607), .Z(G3) );
  NAND2_X1 U682 ( .A1(n609), .A2(n619), .ZN(n608) );
  XNOR2_X1 U683 ( .A(n608), .B(G104), .ZN(G6) );
  XNOR2_X1 U684 ( .A(G107), .B(KEYINPUT110), .ZN(n613) );
  XOR2_X1 U685 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n611) );
  NAND2_X1 U686 ( .A1(n609), .A2(n622), .ZN(n610) );
  XNOR2_X1 U687 ( .A(n611), .B(n610), .ZN(n612) );
  XNOR2_X1 U688 ( .A(n613), .B(n612), .ZN(G9) );
  XOR2_X1 U689 ( .A(G128), .B(KEYINPUT29), .Z(n615) );
  NAND2_X1 U690 ( .A1(n617), .A2(n622), .ZN(n614) );
  XNOR2_X1 U691 ( .A(n615), .B(n614), .ZN(G30) );
  XNOR2_X1 U692 ( .A(G143), .B(n616), .ZN(G45) );
  NAND2_X1 U693 ( .A1(n617), .A2(n619), .ZN(n618) );
  XNOR2_X1 U694 ( .A(n618), .B(G146), .ZN(G48) );
  NAND2_X1 U695 ( .A1(n621), .A2(n619), .ZN(n620) );
  XNOR2_X1 U696 ( .A(n620), .B(G113), .ZN(G15) );
  NAND2_X1 U697 ( .A1(n621), .A2(n622), .ZN(n623) );
  XNOR2_X1 U698 ( .A(n623), .B(G116), .ZN(G18) );
  XNOR2_X1 U699 ( .A(KEYINPUT111), .B(KEYINPUT37), .ZN(n625) );
  XNOR2_X1 U700 ( .A(n625), .B(n624), .ZN(n626) );
  XNOR2_X1 U701 ( .A(G125), .B(n626), .ZN(G27) );
  XOR2_X1 U702 ( .A(G134), .B(n627), .Z(G36) );
  XNOR2_X1 U703 ( .A(G140), .B(n628), .ZN(G42) );
  XNOR2_X1 U704 ( .A(n630), .B(n629), .ZN(n675) );
  INV_X1 U705 ( .A(n631), .ZN(n671) );
  XNOR2_X1 U706 ( .A(KEYINPUT51), .B(KEYINPUT115), .ZN(n632) );
  XNOR2_X1 U707 ( .A(n632), .B(KEYINPUT114), .ZN(n650) );
  NAND2_X1 U708 ( .A1(n634), .A2(n633), .ZN(n648) );
  NAND2_X1 U709 ( .A1(n636), .A2(n635), .ZN(n637) );
  XNOR2_X1 U710 ( .A(n637), .B(KEYINPUT113), .ZN(n638) );
  XNOR2_X1 U711 ( .A(KEYINPUT50), .B(n638), .ZN(n644) );
  NAND2_X1 U712 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U713 ( .A(n641), .B(KEYINPUT49), .ZN(n642) );
  XNOR2_X1 U714 ( .A(KEYINPUT112), .B(n642), .ZN(n643) );
  NOR2_X1 U715 ( .A1(n644), .A2(n643), .ZN(n646) );
  NAND2_X1 U716 ( .A1(n646), .A2(n645), .ZN(n647) );
  NAND2_X1 U717 ( .A1(n648), .A2(n647), .ZN(n649) );
  XOR2_X1 U718 ( .A(n650), .B(n649), .Z(n651) );
  NOR2_X1 U719 ( .A1(n671), .A2(n651), .ZN(n665) );
  NOR2_X1 U720 ( .A1(n654), .A2(n653), .ZN(n655) );
  XNOR2_X1 U721 ( .A(n655), .B(KEYINPUT116), .ZN(n656) );
  NOR2_X1 U722 ( .A1(n657), .A2(n656), .ZN(n662) );
  NOR2_X1 U723 ( .A1(n659), .A2(n658), .ZN(n660) );
  XOR2_X1 U724 ( .A(KEYINPUT117), .B(n660), .Z(n661) );
  NOR2_X1 U725 ( .A1(n662), .A2(n661), .ZN(n663) );
  NOR2_X1 U726 ( .A1(n670), .A2(n663), .ZN(n664) );
  NOR2_X1 U727 ( .A1(n665), .A2(n664), .ZN(n666) );
  XNOR2_X1 U728 ( .A(n666), .B(KEYINPUT52), .ZN(n667) );
  NOR2_X1 U729 ( .A1(n668), .A2(n667), .ZN(n669) );
  XNOR2_X1 U730 ( .A(n669), .B(KEYINPUT118), .ZN(n673) );
  NOR2_X1 U731 ( .A1(n671), .A2(n670), .ZN(n672) );
  NOR2_X1 U732 ( .A1(n673), .A2(n672), .ZN(n674) );
  NAND2_X1 U733 ( .A1(n675), .A2(n674), .ZN(n676) );
  NOR2_X1 U734 ( .A1(n676), .A2(G953), .ZN(n677) );
  XNOR2_X1 U735 ( .A(n677), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U736 ( .A1(n695), .A2(G210), .ZN(n680) );
  XOR2_X1 U737 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n678) );
  XNOR2_X1 U738 ( .A(n680), .B(n370), .ZN(n681) );
  XNOR2_X1 U739 ( .A(KEYINPUT58), .B(KEYINPUT119), .ZN(n684) );
  XNOR2_X1 U740 ( .A(n682), .B(KEYINPUT57), .ZN(n683) );
  XNOR2_X1 U741 ( .A(n684), .B(n683), .ZN(n686) );
  NAND2_X1 U742 ( .A1(n695), .A2(G469), .ZN(n685) );
  XNOR2_X1 U743 ( .A(n686), .B(n685), .ZN(n687) );
  NOR2_X1 U744 ( .A1(n699), .A2(n687), .ZN(G54) );
  XOR2_X1 U745 ( .A(KEYINPUT121), .B(KEYINPUT90), .Z(n689) );
  XNOR2_X1 U746 ( .A(KEYINPUT59), .B(KEYINPUT120), .ZN(n688) );
  XNOR2_X1 U747 ( .A(n689), .B(n688), .ZN(n690) );
  NAND2_X1 U748 ( .A1(G478), .A2(n695), .ZN(n692) );
  XNOR2_X1 U749 ( .A(n693), .B(n692), .ZN(n694) );
  NOR2_X1 U750 ( .A1(n699), .A2(n694), .ZN(G63) );
  NAND2_X1 U751 ( .A1(n695), .A2(G217), .ZN(n696) );
  NOR2_X1 U752 ( .A1(n699), .A2(n698), .ZN(G66) );
  XOR2_X1 U753 ( .A(KEYINPUT125), .B(n700), .Z(n703) );
  XNOR2_X1 U754 ( .A(n701), .B(G101), .ZN(n702) );
  XNOR2_X1 U755 ( .A(n703), .B(n702), .ZN(n704) );
  NOR2_X1 U756 ( .A1(n705), .A2(n704), .ZN(n713) );
  NAND2_X1 U757 ( .A1(n706), .A2(n719), .ZN(n707) );
  XOR2_X1 U758 ( .A(KEYINPUT123), .B(n707), .Z(n711) );
  NAND2_X1 U759 ( .A1(G953), .A2(G224), .ZN(n708) );
  XNOR2_X1 U760 ( .A(KEYINPUT61), .B(n708), .ZN(n709) );
  NAND2_X1 U761 ( .A1(n709), .A2(G898), .ZN(n710) );
  NAND2_X1 U762 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U763 ( .A(n713), .B(n712), .ZN(n714) );
  XNOR2_X1 U764 ( .A(KEYINPUT124), .B(n714), .ZN(G69) );
  XOR2_X1 U765 ( .A(n716), .B(n715), .Z(n722) );
  INV_X1 U766 ( .A(n722), .ZN(n718) );
  XNOR2_X1 U767 ( .A(n718), .B(n717), .ZN(n720) );
  NAND2_X1 U768 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U769 ( .A(KEYINPUT126), .B(n721), .ZN(n727) );
  XNOR2_X1 U770 ( .A(G227), .B(n722), .ZN(n723) );
  NAND2_X1 U771 ( .A1(n723), .A2(G900), .ZN(n724) );
  NAND2_X1 U772 ( .A1(n724), .A2(G953), .ZN(n725) );
  XOR2_X1 U773 ( .A(KEYINPUT127), .B(n725), .Z(n726) );
  NAND2_X1 U774 ( .A1(n727), .A2(n726), .ZN(G72) );
  XOR2_X1 U775 ( .A(n728), .B(G122), .Z(G24) );
  XNOR2_X1 U776 ( .A(n729), .B(G119), .ZN(G21) );
  XOR2_X1 U777 ( .A(n730), .B(G137), .Z(G39) );
  XOR2_X1 U778 ( .A(n731), .B(G131), .Z(G33) );
  XNOR2_X1 U779 ( .A(n732), .B(G110), .ZN(G12) );
endmodule

