//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 1 1 1 0 0 1 0 0 0 1 0 0 0 0 0 1 1 0 1 1 0 0 1 1 0 0 0 1 0 0 0 0 1 0 0 0 1 0 1 1 1 1 1 1 1 0 0 1 1 1 0 0 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:20 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1285, new_n1286, new_n1287,
    new_n1288, new_n1289;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n211));
  INV_X1    g0011(.A(G77), .ZN(new_n212));
  INV_X1    g0012(.A(G244), .ZN(new_n213));
  INV_X1    g0013(.A(G87), .ZN(new_n214));
  INV_X1    g0014(.A(G250), .ZN(new_n215));
  OAI221_X1 g0015(.A(new_n211), .B1(new_n212), .B2(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n217));
  INV_X1    g0017(.A(G232), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n217), .B1(new_n202), .B2(new_n218), .C1(new_n203), .C2(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n210), .B1(new_n216), .B2(new_n220), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT64), .Z(new_n222));
  NAND2_X1  g0022(.A1(new_n222), .A2(KEYINPUT1), .ZN(new_n223));
  XOR2_X1   g0023(.A(new_n223), .B(KEYINPUT65), .Z(new_n224));
  OAI21_X1  g0024(.A(G50), .B1(G58), .B2(G68), .ZN(new_n225));
  INV_X1    g0025(.A(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n227), .A2(new_n208), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n210), .A2(G13), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n230), .B(G250), .C1(G257), .C2(G264), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT0), .ZN(new_n232));
  OAI211_X1 g0032(.A(new_n229), .B(new_n232), .C1(new_n222), .C2(KEYINPUT1), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n224), .A2(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT2), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(new_n218), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XOR2_X1   g0042(.A(G68), .B(G77), .Z(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G58), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  NAND2_X1  g0049(.A1(new_n202), .A2(KEYINPUT8), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT8), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G58), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  NOR2_X1   g0053(.A1(G20), .A2(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n208), .A2(G33), .ZN(new_n256));
  XNOR2_X1  g0056(.A(KEYINPUT15), .B(G87), .ZN(new_n257));
  OAI221_X1 g0057(.A(new_n255), .B1(new_n208), .B2(new_n212), .C1(new_n256), .C2(new_n257), .ZN(new_n258));
  NAND3_X1  g0058(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(new_n227), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n207), .A2(G13), .A3(G20), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n263), .A2(new_n260), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n212), .B1(new_n207), .B2(G20), .ZN(new_n265));
  AOI22_X1  g0065(.A1(new_n264), .A2(new_n265), .B1(new_n212), .B2(new_n263), .ZN(new_n266));
  AND2_X1   g0066(.A1(new_n261), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  OR2_X1    g0068(.A1(KEYINPUT3), .A2(G33), .ZN(new_n269));
  NAND2_X1  g0069(.A1(KEYINPUT3), .A2(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(G238), .A2(G1698), .ZN(new_n272));
  OAI211_X1 g0072(.A(new_n271), .B(new_n272), .C1(new_n218), .C2(G1698), .ZN(new_n273));
  NAND2_X1  g0073(.A1(G33), .A2(G41), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n274), .A2(G1), .A3(G13), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  OAI211_X1 g0076(.A(new_n273), .B(new_n276), .C1(G107), .C2(new_n271), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT66), .ZN(new_n278));
  AND2_X1   g0078(.A1(G33), .A2(G41), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n278), .B1(new_n279), .B2(new_n227), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NAND4_X1  g0082(.A1(new_n274), .A2(KEYINPUT66), .A3(G1), .A4(G13), .ZN(new_n283));
  NAND4_X1  g0083(.A1(new_n280), .A2(new_n282), .A3(G274), .A4(new_n283), .ZN(new_n284));
  AND2_X1   g0084(.A1(new_n280), .A2(new_n283), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n285), .A2(G244), .A3(new_n281), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n277), .A2(new_n284), .A3(new_n286), .ZN(new_n287));
  XOR2_X1   g0087(.A(KEYINPUT68), .B(G200), .Z(new_n288));
  AOI21_X1  g0088(.A(new_n268), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G190), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n289), .B1(new_n290), .B2(new_n287), .ZN(new_n291));
  INV_X1    g0091(.A(G169), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n267), .B1(new_n292), .B2(new_n287), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT69), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n294), .B1(new_n287), .B2(G179), .ZN(new_n295));
  OR3_X1    g0095(.A1(new_n287), .A2(new_n294), .A3(G179), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n293), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  AND2_X1   g0097(.A1(new_n291), .A2(new_n297), .ZN(new_n298));
  NAND4_X1  g0098(.A1(new_n280), .A2(G238), .A3(new_n281), .A4(new_n283), .ZN(new_n299));
  INV_X1    g0099(.A(G33), .ZN(new_n300));
  INV_X1    g0100(.A(G97), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NOR2_X1   g0102(.A1(G226), .A2(G1698), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n303), .B1(new_n218), .B2(G1698), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n302), .B1(new_n304), .B2(new_n271), .ZN(new_n305));
  OAI211_X1 g0105(.A(new_n284), .B(new_n299), .C1(new_n305), .C2(new_n275), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(KEYINPUT13), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n218), .A2(G1698), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n308), .B1(G226), .B2(G1698), .ZN(new_n309));
  AND2_X1   g0109(.A1(KEYINPUT3), .A2(G33), .ZN(new_n310));
  NOR2_X1   g0110(.A1(KEYINPUT3), .A2(G33), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  OAI22_X1  g0112(.A1(new_n309), .A2(new_n312), .B1(new_n300), .B2(new_n301), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(new_n276), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT13), .ZN(new_n315));
  NAND4_X1  g0115(.A1(new_n314), .A2(new_n315), .A3(new_n284), .A4(new_n299), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n307), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(G200), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT70), .ZN(new_n319));
  XNOR2_X1  g0119(.A(new_n318), .B(new_n319), .ZN(new_n320));
  AND3_X1   g0120(.A1(new_n306), .A2(KEYINPUT71), .A3(KEYINPUT13), .ZN(new_n321));
  AOI21_X1  g0121(.A(KEYINPUT71), .B1(new_n306), .B2(KEYINPUT13), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n323), .A2(G190), .A3(new_n316), .ZN(new_n324));
  INV_X1    g0124(.A(new_n260), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT67), .ZN(new_n326));
  XNOR2_X1  g0126(.A(new_n256), .B(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(G77), .ZN(new_n328));
  AOI22_X1  g0128(.A1(new_n254), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n325), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  OR2_X1    g0130(.A1(new_n330), .A2(KEYINPUT11), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(KEYINPUT11), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT72), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n333), .B1(new_n262), .B2(G68), .ZN(new_n334));
  XNOR2_X1  g0134(.A(new_n334), .B(KEYINPUT12), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n203), .B1(new_n207), .B2(G20), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n335), .B1(new_n264), .B2(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n331), .A2(new_n332), .A3(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n324), .A2(new_n339), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n320), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n285), .A2(G226), .A3(new_n281), .ZN(new_n343));
  INV_X1    g0143(.A(G1698), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(G222), .ZN(new_n345));
  NAND2_X1  g0145(.A1(G223), .A2(G1698), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n271), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  OAI211_X1 g0147(.A(new_n347), .B(new_n276), .C1(G77), .C2(new_n271), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n343), .A2(new_n348), .A3(new_n284), .ZN(new_n349));
  OR2_X1    g0149(.A1(new_n349), .A2(new_n290), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n288), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n327), .A2(new_n253), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n204), .A2(G20), .B1(G150), .B2(new_n254), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n325), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n207), .A2(G20), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n264), .A2(G50), .A3(new_n355), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n356), .B1(G50), .B2(new_n262), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n354), .A2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT9), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NOR3_X1   g0160(.A1(new_n354), .A2(new_n357), .A3(KEYINPUT9), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n350), .B(new_n351), .C1(new_n360), .C2(new_n361), .ZN(new_n362));
  XNOR2_X1  g0162(.A(new_n362), .B(KEYINPUT10), .ZN(new_n363));
  OR2_X1    g0163(.A1(new_n349), .A2(G179), .ZN(new_n364));
  INV_X1    g0164(.A(new_n358), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n349), .A2(new_n292), .ZN(new_n366));
  AND3_X1   g0166(.A1(new_n364), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(new_n367), .ZN(new_n368));
  NAND4_X1  g0168(.A1(new_n298), .A2(new_n342), .A3(new_n363), .A4(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n317), .A2(G169), .ZN(new_n370));
  AOI21_X1  g0170(.A(KEYINPUT73), .B1(new_n370), .B2(KEYINPUT14), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n292), .B1(new_n307), .B2(new_n316), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT73), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT14), .ZN(new_n374));
  NOR3_X1   g0174(.A1(new_n372), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  OAI22_X1  g0175(.A1(new_n371), .A2(new_n375), .B1(KEYINPUT14), .B2(new_n370), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT74), .ZN(new_n377));
  AND2_X1   g0177(.A1(new_n316), .A2(G179), .ZN(new_n378));
  INV_X1    g0178(.A(new_n322), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n306), .A2(KEYINPUT71), .A3(KEYINPUT13), .ZN(new_n380));
  AND4_X1   g0180(.A1(new_n377), .A2(new_n378), .A3(new_n379), .A4(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n377), .B1(new_n323), .B2(new_n378), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n338), .B1(new_n376), .B2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n280), .A2(G232), .A3(new_n281), .A4(new_n283), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n300), .A2(new_n214), .ZN(new_n387));
  NOR2_X1   g0187(.A1(G223), .A2(G1698), .ZN(new_n388));
  INV_X1    g0188(.A(G226), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n388), .B1(new_n389), .B2(G1698), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n387), .B1(new_n390), .B2(new_n271), .ZN(new_n391));
  OAI211_X1 g0191(.A(new_n386), .B(new_n284), .C1(new_n391), .C2(new_n275), .ZN(new_n392));
  INV_X1    g0192(.A(G179), .ZN(new_n393));
  OR2_X1    g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n392), .A2(G169), .ZN(new_n395));
  AOI21_X1  g0195(.A(KEYINPUT7), .B1(new_n312), .B2(new_n208), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT7), .ZN(new_n397));
  NOR4_X1   g0197(.A1(new_n310), .A2(new_n311), .A3(new_n397), .A4(G20), .ZN(new_n398));
  OAI21_X1  g0198(.A(G68), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n202), .A2(new_n203), .ZN(new_n400));
  NOR2_X1   g0200(.A1(G58), .A2(G68), .ZN(new_n401));
  OAI21_X1  g0201(.A(G20), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n254), .A2(G159), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n399), .A2(KEYINPUT16), .A3(new_n405), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n269), .A2(KEYINPUT7), .A3(new_n208), .A4(new_n270), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(KEYINPUT75), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n397), .B1(new_n271), .B2(G20), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT75), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n312), .A2(new_n410), .A3(KEYINPUT7), .A4(new_n208), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n408), .A2(new_n409), .A3(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n404), .B1(new_n412), .B2(G68), .ZN(new_n413));
  OAI211_X1 g0213(.A(new_n260), .B(new_n406), .C1(new_n413), .C2(KEYINPUT16), .ZN(new_n414));
  AND2_X1   g0214(.A1(new_n253), .A2(new_n355), .ZN(new_n415));
  INV_X1    g0215(.A(new_n253), .ZN(new_n416));
  AOI22_X1  g0216(.A1(new_n415), .A2(new_n264), .B1(new_n263), .B2(new_n416), .ZN(new_n417));
  AOI221_X4 g0217(.A(KEYINPUT18), .B1(new_n394), .B2(new_n395), .C1(new_n414), .C2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT18), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n414), .A2(new_n417), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n394), .A2(new_n395), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n419), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n418), .A2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(G200), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n392), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n389), .A2(G1698), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n426), .B1(G223), .B2(G1698), .ZN(new_n427));
  OAI22_X1  g0227(.A1(new_n427), .A2(new_n312), .B1(new_n300), .B2(new_n214), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(new_n276), .ZN(new_n429));
  AND2_X1   g0229(.A1(new_n290), .A2(KEYINPUT76), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n290), .A2(KEYINPUT76), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n429), .A2(new_n386), .A3(new_n284), .A4(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n425), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n412), .A2(G68), .ZN(new_n435));
  AOI21_X1  g0235(.A(KEYINPUT16), .B1(new_n435), .B2(new_n405), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n406), .A2(new_n260), .ZN(new_n437));
  OAI211_X1 g0237(.A(new_n417), .B(new_n434), .C1(new_n436), .C2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(KEYINPUT17), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT17), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n414), .A2(new_n440), .A3(new_n417), .A4(new_n434), .ZN(new_n441));
  AND3_X1   g0241(.A1(new_n439), .A2(KEYINPUT77), .A3(new_n441), .ZN(new_n442));
  AOI21_X1  g0242(.A(KEYINPUT77), .B1(new_n439), .B2(new_n441), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n423), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NOR3_X1   g0244(.A1(new_n369), .A2(new_n385), .A3(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT85), .ZN(new_n447));
  OAI21_X1  g0247(.A(KEYINPUT23), .B1(new_n208), .B2(G107), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT23), .ZN(new_n449));
  INV_X1    g0249(.A(G107), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n449), .A2(new_n450), .A3(G20), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n208), .A2(G33), .A3(G116), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n448), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(KEYINPUT83), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT83), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n448), .A2(new_n451), .A3(new_n452), .A4(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT81), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT22), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n208), .B1(new_n310), .B2(new_n311), .ZN(new_n460));
  OAI211_X1 g0260(.A(new_n458), .B(new_n459), .C1(new_n460), .C2(new_n214), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n214), .B1(KEYINPUT81), .B2(KEYINPUT22), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n458), .A2(new_n459), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n271), .A2(new_n462), .A3(new_n208), .A4(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n457), .A2(new_n461), .A3(new_n464), .ZN(new_n465));
  XNOR2_X1  g0265(.A(KEYINPUT82), .B(KEYINPUT24), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n457), .A2(new_n466), .A3(new_n461), .A4(new_n464), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n325), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT84), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT25), .ZN(new_n472));
  AOI211_X1 g0272(.A(G107), .B(new_n262), .C1(new_n471), .C2(new_n472), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n471), .A2(new_n472), .ZN(new_n474));
  OR2_X1    g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n473), .A2(new_n474), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n207), .A2(G33), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n325), .A2(new_n262), .A3(new_n478), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n477), .B1(new_n450), .B2(new_n479), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n447), .B1(new_n470), .B2(new_n480), .ZN(new_n481));
  AND2_X1   g0281(.A1(new_n461), .A2(new_n464), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n466), .B1(new_n482), .B2(new_n457), .ZN(new_n483));
  INV_X1    g0283(.A(new_n469), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n260), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  AND3_X1   g0285(.A1(new_n325), .A2(new_n262), .A3(new_n478), .ZN(new_n486));
  AOI22_X1  g0286(.A1(new_n475), .A2(new_n476), .B1(G107), .B2(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n485), .A2(KEYINPUT85), .A3(new_n487), .ZN(new_n488));
  OAI211_X1 g0288(.A(G250), .B(new_n344), .C1(new_n310), .C2(new_n311), .ZN(new_n489));
  OAI211_X1 g0289(.A(G257), .B(G1698), .C1(new_n310), .C2(new_n311), .ZN(new_n490));
  INV_X1    g0290(.A(G294), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n489), .B(new_n490), .C1(new_n300), .C2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(new_n276), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(KEYINPUT86), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT86), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n492), .A2(new_n495), .A3(new_n276), .ZN(new_n496));
  INV_X1    g0296(.A(G45), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n497), .A2(G1), .ZN(new_n498));
  INV_X1    g0298(.A(G41), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(KEYINPUT5), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT5), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(G41), .ZN(new_n502));
  AND3_X1   g0302(.A1(new_n498), .A2(new_n500), .A3(new_n502), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n503), .A2(G274), .A3(new_n280), .A4(new_n283), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n498), .A2(new_n500), .A3(new_n502), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n505), .A2(new_n280), .A3(G264), .A4(new_n283), .ZN(new_n506));
  AND2_X1   g0306(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n494), .A2(new_n496), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(G169), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n493), .A2(new_n504), .A3(new_n506), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n509), .B1(new_n393), .B2(new_n510), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n481), .A2(new_n488), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n510), .A2(new_n424), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n513), .B1(new_n508), .B2(G190), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n514), .A2(new_n485), .A3(new_n487), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n512), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n344), .A2(G257), .ZN(new_n517));
  NAND2_X1  g0317(.A1(G264), .A2(G1698), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n271), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n519), .B(new_n276), .C1(G303), .C2(new_n271), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n505), .A2(new_n280), .A3(G270), .A4(new_n283), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n520), .A2(new_n504), .A3(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n264), .A2(G116), .A3(new_n478), .ZN(new_n523));
  INV_X1    g0323(.A(G116), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n263), .A2(new_n524), .ZN(new_n525));
  AOI22_X1  g0325(.A1(new_n259), .A2(new_n227), .B1(G20), .B2(new_n524), .ZN(new_n526));
  NAND2_X1  g0326(.A1(G33), .A2(G283), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n527), .B(new_n208), .C1(G33), .C2(new_n301), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n526), .A2(KEYINPUT20), .A3(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(new_n529), .ZN(new_n530));
  AOI21_X1  g0330(.A(KEYINPUT20), .B1(new_n526), .B2(new_n528), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n523), .B(new_n525), .C1(new_n530), .C2(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n522), .A2(new_n532), .A3(G169), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT21), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n522), .A2(G200), .ZN(new_n536));
  INV_X1    g0336(.A(new_n532), .ZN(new_n537));
  INV_X1    g0337(.A(new_n432), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n520), .A2(new_n504), .A3(new_n538), .A4(new_n521), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n536), .A2(new_n537), .A3(new_n539), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n522), .A2(new_n393), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(new_n532), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n522), .A2(new_n532), .A3(KEYINPUT21), .A4(G169), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n535), .A2(new_n540), .A3(new_n542), .A4(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n214), .A2(new_n301), .A3(new_n450), .ZN(new_n545));
  OAI211_X1 g0345(.A(KEYINPUT19), .B(new_n545), .C1(new_n302), .C2(G20), .ZN(new_n546));
  OAI211_X1 g0346(.A(new_n208), .B(G68), .C1(new_n310), .C2(new_n311), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT19), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n548), .B1(new_n256), .B2(new_n301), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n546), .A2(new_n547), .A3(new_n549), .ZN(new_n550));
  AOI22_X1  g0350(.A1(new_n550), .A2(new_n260), .B1(new_n263), .B2(new_n257), .ZN(new_n551));
  INV_X1    g0351(.A(new_n257), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(KEYINPUT80), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT80), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n257), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n486), .A2(new_n553), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n551), .A2(new_n556), .ZN(new_n557));
  OR3_X1    g0357(.A1(new_n497), .A2(G1), .A3(G274), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n215), .B1(new_n497), .B2(G1), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n280), .A2(new_n558), .A3(new_n283), .A4(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n219), .A2(new_n344), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n213), .A2(G1698), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n562), .B(new_n563), .C1(new_n310), .C2(new_n311), .ZN(new_n564));
  NAND2_X1  g0364(.A1(G33), .A2(G116), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n275), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n561), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(new_n393), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n292), .B1(new_n561), .B2(new_n566), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n557), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  AND2_X1   g0370(.A1(new_n564), .A2(new_n565), .ZN(new_n571));
  OAI211_X1 g0371(.A(G190), .B(new_n560), .C1(new_n571), .C2(new_n275), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n288), .B1(new_n561), .B2(new_n566), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n486), .A2(G87), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n572), .A2(new_n573), .A3(new_n551), .A4(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n570), .A2(new_n575), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n544), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n263), .A2(new_n301), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n578), .B1(new_n479), .B2(new_n301), .ZN(new_n579));
  INV_X1    g0379(.A(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT78), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n412), .A2(G107), .ZN(new_n582));
  XNOR2_X1  g0382(.A(G97), .B(G107), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT6), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NOR3_X1   g0385(.A1(new_n584), .A2(new_n301), .A3(G107), .ZN(new_n586));
  INV_X1    g0386(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  AOI22_X1  g0388(.A1(new_n588), .A2(G20), .B1(G77), .B2(new_n254), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n582), .A2(new_n589), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n581), .B1(new_n590), .B2(new_n260), .ZN(new_n591));
  AOI211_X1 g0391(.A(KEYINPUT78), .B(new_n325), .C1(new_n582), .C2(new_n589), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n580), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n271), .A2(G250), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n344), .B1(new_n594), .B2(KEYINPUT4), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT4), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n596), .A2(G1698), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n597), .B(G244), .C1(new_n311), .C2(new_n310), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n213), .B1(new_n269), .B2(new_n270), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n598), .B(new_n527), .C1(new_n599), .C2(KEYINPUT4), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n276), .B1(new_n595), .B2(new_n600), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n505), .A2(new_n280), .A3(G257), .A4(new_n283), .ZN(new_n602));
  AND2_X1   g0402(.A1(new_n504), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(new_n292), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n601), .A2(new_n603), .A3(new_n393), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n593), .A2(new_n608), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n424), .B1(new_n601), .B2(new_n603), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n601), .A2(new_n603), .A3(G190), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT79), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n601), .A2(new_n603), .A3(KEYINPUT79), .A4(G190), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n610), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n254), .A2(G77), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n586), .B1(new_n584), .B2(new_n583), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n616), .B1(new_n617), .B2(new_n208), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n618), .B1(G107), .B2(new_n412), .ZN(new_n619));
  OAI21_X1  g0419(.A(KEYINPUT78), .B1(new_n619), .B2(new_n325), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n590), .A2(new_n581), .A3(new_n260), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n579), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n615), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n577), .A2(new_n609), .A3(new_n623), .ZN(new_n624));
  NOR3_X1   g0424(.A1(new_n446), .A2(new_n516), .A3(new_n624), .ZN(G372));
  NOR2_X1   g0425(.A1(new_n341), .A2(new_n297), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n385), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n442), .A2(new_n443), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n423), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n367), .B1(new_n629), .B2(new_n363), .ZN(new_n630));
  INV_X1    g0430(.A(new_n570), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT87), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n573), .A2(new_n551), .A3(new_n632), .A4(new_n574), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(new_n572), .ZN(new_n634));
  INV_X1    g0434(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n550), .A2(new_n260), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n257), .A2(new_n263), .ZN(new_n637));
  AND3_X1   g0437(.A1(new_n636), .A2(new_n574), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(new_n573), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(KEYINPUT87), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n631), .B1(new_n635), .B2(new_n640), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n609), .A2(new_n623), .A3(new_n515), .A4(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n485), .A2(new_n487), .ZN(new_n643));
  AND2_X1   g0443(.A1(new_n511), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n535), .A2(new_n542), .A3(new_n543), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n642), .A2(new_n646), .ZN(new_n647));
  OAI21_X1  g0447(.A(KEYINPUT26), .B1(new_n609), .B2(new_n576), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n620), .A2(new_n621), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n607), .B1(new_n649), .B2(new_n580), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT26), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n650), .A2(new_n641), .A3(new_n651), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n648), .A2(new_n652), .A3(new_n570), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n445), .B1(new_n647), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n630), .A2(new_n654), .ZN(G369));
  NAND3_X1  g0455(.A1(new_n207), .A2(new_n208), .A3(G13), .ZN(new_n656));
  OR2_X1    g0456(.A1(new_n656), .A2(KEYINPUT27), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(KEYINPUT27), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n657), .A2(G213), .A3(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(G343), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n537), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g0462(.A(new_n662), .B(KEYINPUT88), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(new_n645), .ZN(new_n664));
  OR2_X1    g0464(.A1(new_n664), .A2(KEYINPUT89), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(KEYINPUT89), .ZN(new_n666));
  OAI211_X1 g0466(.A(new_n665), .B(new_n666), .C1(new_n544), .C2(new_n663), .ZN(new_n667));
  XNOR2_X1  g0467(.A(KEYINPUT90), .B(G330), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT91), .ZN(new_n671));
  XNOR2_X1  g0471(.A(new_n670), .B(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n661), .ZN(new_n673));
  AND3_X1   g0473(.A1(new_n481), .A2(new_n488), .A3(new_n673), .ZN(new_n674));
  OAI22_X1  g0474(.A1(new_n516), .A2(new_n674), .B1(new_n512), .B2(new_n661), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n645), .A2(new_n661), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n516), .A2(new_n677), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n678), .B1(new_n644), .B2(new_n661), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n676), .A2(new_n679), .ZN(G399));
  INV_X1    g0480(.A(new_n230), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n681), .A2(G41), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n545), .A2(G116), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n683), .A2(G1), .A3(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n685), .B1(new_n225), .B2(new_n683), .ZN(new_n686));
  XNOR2_X1  g0486(.A(new_n686), .B(KEYINPUT28), .ZN(new_n687));
  AND2_X1   g0487(.A1(new_n601), .A2(new_n603), .ZN(new_n688));
  AND2_X1   g0488(.A1(new_n493), .A2(new_n506), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n688), .A2(new_n541), .A3(new_n689), .A4(new_n567), .ZN(new_n690));
  XNOR2_X1  g0490(.A(new_n690), .B(KEYINPUT30), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n567), .A2(G179), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n604), .A2(new_n692), .A3(new_n510), .A4(new_n522), .ZN(new_n693));
  XNOR2_X1  g0493(.A(new_n693), .B(KEYINPUT92), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n661), .B1(new_n691), .B2(new_n694), .ZN(new_n695));
  AND2_X1   g0495(.A1(new_n512), .A2(new_n515), .ZN(new_n696));
  AND2_X1   g0496(.A1(new_n609), .A2(new_n623), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n696), .A2(new_n697), .A3(new_n577), .A4(new_n661), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n695), .B1(new_n698), .B2(KEYINPUT31), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT31), .ZN(new_n700));
  AOI211_X1 g0500(.A(new_n700), .B(new_n661), .C1(new_n691), .C2(new_n693), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n669), .B1(new_n699), .B2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n645), .ZN(new_n704));
  AND2_X1   g0504(.A1(new_n512), .A2(new_n704), .ZN(new_n705));
  OAI21_X1  g0505(.A(KEYINPUT94), .B1(new_n705), .B2(new_n642), .ZN(new_n706));
  AND2_X1   g0506(.A1(new_n641), .A2(new_n515), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n512), .A2(new_n704), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT94), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n697), .A2(new_n707), .A3(new_n708), .A4(new_n709), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n651), .B1(new_n650), .B2(new_n641), .ZN(new_n711));
  NOR4_X1   g0511(.A1(new_n622), .A2(new_n576), .A3(new_n607), .A4(KEYINPUT26), .ZN(new_n712));
  NOR3_X1   g0512(.A1(new_n711), .A2(new_n712), .A3(new_n631), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n706), .A2(new_n710), .A3(new_n713), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n714), .A2(KEYINPUT29), .A3(new_n661), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n661), .B1(new_n647), .B2(new_n653), .ZN(new_n716));
  XNOR2_X1  g0516(.A(KEYINPUT93), .B(KEYINPUT29), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n703), .B1(new_n715), .B2(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n687), .B1(new_n719), .B2(G1), .ZN(G364));
  AND2_X1   g0520(.A1(new_n208), .A2(G13), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(G45), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n683), .A2(G1), .A3(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n681), .A2(new_n312), .ZN(new_n725));
  AOI22_X1  g0525(.A1(new_n725), .A2(G355), .B1(new_n524), .B2(new_n681), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n681), .A2(new_n271), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n727), .B1(G45), .B2(new_n225), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n245), .A2(new_n497), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n726), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  AND2_X1   g0530(.A1(new_n730), .A2(KEYINPUT95), .ZN(new_n731));
  NOR2_X1   g0531(.A1(G13), .A2(G33), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n733), .A2(G20), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n227), .B1(G20), .B2(new_n292), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n736), .B1(new_n730), .B2(KEYINPUT95), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n724), .B1(new_n731), .B2(new_n737), .ZN(new_n738));
  NOR4_X1   g0538(.A1(new_n208), .A2(G179), .A3(G190), .A4(G200), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n271), .B1(new_n739), .B2(G329), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n208), .A2(new_n393), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(new_n424), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n742), .A2(G190), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(G311), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n740), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n288), .A2(G20), .A3(new_n393), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(G190), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n746), .B1(G283), .B2(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n432), .A2(new_n742), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n741), .A2(G200), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n432), .A2(new_n751), .ZN(new_n752));
  AOI22_X1  g0552(.A1(G322), .A2(new_n750), .B1(new_n752), .B2(G326), .ZN(new_n753));
  NOR3_X1   g0553(.A1(new_n290), .A2(G179), .A3(G200), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(new_n208), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n751), .A2(G190), .ZN(new_n757));
  XNOR2_X1  g0557(.A(KEYINPUT33), .B(G317), .ZN(new_n758));
  AOI22_X1  g0558(.A1(G294), .A2(new_n756), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n747), .A2(new_n290), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(G303), .ZN(new_n761));
  NAND4_X1  g0561(.A1(new_n749), .A2(new_n753), .A3(new_n759), .A4(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n760), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(new_n214), .ZN(new_n764));
  INV_X1    g0564(.A(new_n748), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(new_n450), .ZN(new_n766));
  NOR3_X1   g0566(.A1(new_n764), .A2(new_n766), .A3(new_n312), .ZN(new_n767));
  XOR2_X1   g0567(.A(new_n767), .B(KEYINPUT96), .Z(new_n768));
  NAND2_X1  g0568(.A1(new_n739), .A2(G159), .ZN(new_n769));
  XOR2_X1   g0569(.A(new_n769), .B(KEYINPUT32), .Z(new_n770));
  NAND2_X1  g0570(.A1(new_n757), .A2(G68), .ZN(new_n771));
  AOI22_X1  g0571(.A1(new_n750), .A2(G58), .B1(new_n756), .B2(G97), .ZN(new_n772));
  AOI22_X1  g0572(.A1(new_n752), .A2(G50), .B1(new_n743), .B2(G77), .ZN(new_n773));
  NAND4_X1  g0573(.A1(new_n770), .A2(new_n771), .A3(new_n772), .A4(new_n773), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n762), .B1(new_n768), .B2(new_n774), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n738), .B1(new_n775), .B2(new_n735), .ZN(new_n776));
  INV_X1    g0576(.A(new_n734), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n776), .B1(new_n667), .B2(new_n777), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n723), .B1(new_n667), .B2(new_n669), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n778), .B1(new_n672), .B2(new_n779), .ZN(G396));
  NAND2_X1  g0580(.A1(new_n297), .A2(KEYINPUT99), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n268), .A2(new_n673), .ZN(new_n782));
  INV_X1    g0582(.A(KEYINPUT99), .ZN(new_n783));
  NAND4_X1  g0583(.A1(new_n293), .A2(new_n783), .A3(new_n295), .A4(new_n296), .ZN(new_n784));
  NAND4_X1  g0584(.A1(new_n781), .A2(new_n291), .A3(new_n782), .A4(new_n784), .ZN(new_n785));
  OR2_X1    g0585(.A1(new_n297), .A2(new_n782), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  XNOR2_X1  g0587(.A(new_n716), .B(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(new_n702), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n724), .B1(new_n789), .B2(new_n702), .ZN(new_n792));
  INV_X1    g0592(.A(new_n787), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(new_n732), .ZN(new_n794));
  INV_X1    g0594(.A(new_n735), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(new_n733), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n724), .B1(G77), .B2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n739), .ZN(new_n798));
  OAI221_X1 g0598(.A(new_n312), .B1(new_n755), .B2(new_n301), .C1(new_n745), .C2(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n799), .B1(G87), .B2(new_n748), .ZN(new_n800));
  AOI22_X1  g0600(.A1(new_n750), .A2(G294), .B1(new_n743), .B2(G116), .ZN(new_n801));
  AOI22_X1  g0601(.A1(new_n752), .A2(G303), .B1(new_n757), .B2(G283), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n760), .A2(G107), .ZN(new_n803));
  NAND4_X1  g0603(.A1(new_n800), .A2(new_n801), .A3(new_n802), .A4(new_n803), .ZN(new_n804));
  AOI22_X1  g0604(.A1(new_n752), .A2(G137), .B1(new_n743), .B2(G159), .ZN(new_n805));
  INV_X1    g0605(.A(G150), .ZN(new_n806));
  INV_X1    g0606(.A(new_n757), .ZN(new_n807));
  INV_X1    g0607(.A(new_n750), .ZN(new_n808));
  XNOR2_X1  g0608(.A(KEYINPUT97), .B(G143), .ZN(new_n809));
  OAI221_X1 g0609(.A(new_n805), .B1(new_n806), .B2(new_n807), .C1(new_n808), .C2(new_n809), .ZN(new_n810));
  XNOR2_X1  g0610(.A(new_n810), .B(KEYINPUT98), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(KEYINPUT34), .ZN(new_n812));
  INV_X1    g0612(.A(G132), .ZN(new_n813));
  OAI221_X1 g0613(.A(new_n271), .B1(new_n755), .B2(new_n202), .C1(new_n813), .C2(new_n798), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n814), .B1(G68), .B2(new_n748), .ZN(new_n815));
  OAI211_X1 g0615(.A(new_n812), .B(new_n815), .C1(new_n201), .C2(new_n763), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n811), .A2(KEYINPUT34), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n804), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n797), .B1(new_n818), .B2(new_n735), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n791), .A2(new_n792), .B1(new_n794), .B2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(G384));
  OR2_X1    g0621(.A1(new_n588), .A2(KEYINPUT35), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n588), .A2(KEYINPUT35), .ZN(new_n823));
  NAND4_X1  g0623(.A1(new_n822), .A2(G116), .A3(new_n228), .A4(new_n823), .ZN(new_n824));
  XOR2_X1   g0624(.A(new_n824), .B(KEYINPUT36), .Z(new_n825));
  OAI211_X1 g0625(.A(new_n226), .B(G77), .C1(new_n202), .C2(new_n203), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n201), .A2(G68), .ZN(new_n827));
  AOI211_X1 g0627(.A(new_n207), .B(G13), .C1(new_n826), .C2(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n825), .A2(new_n828), .ZN(new_n829));
  OAI211_X1 g0629(.A(new_n787), .B(new_n661), .C1(new_n647), .C2(new_n653), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n781), .A2(new_n784), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n831), .A2(new_n661), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n384), .A2(KEYINPUT100), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n370), .A2(KEYINPUT73), .A3(KEYINPUT14), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n373), .B1(new_n372), .B2(new_n374), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n834), .A2(new_n835), .B1(new_n374), .B2(new_n372), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n378), .A2(new_n379), .A3(new_n380), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n837), .A2(KEYINPUT74), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n323), .A2(new_n377), .A3(new_n378), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n836), .A2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT100), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n841), .A2(new_n842), .A3(new_n338), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n338), .A2(new_n673), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT101), .ZN(new_n845));
  XNOR2_X1  g0645(.A(new_n844), .B(new_n845), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n846), .A2(new_n341), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n833), .A2(new_n843), .A3(new_n847), .ZN(new_n848));
  OAI211_X1 g0648(.A(new_n338), .B(new_n673), .C1(new_n841), .C2(new_n341), .ZN(new_n849));
  AOI22_X1  g0649(.A1(new_n830), .A2(new_n832), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n437), .ZN(new_n851));
  AND2_X1   g0651(.A1(new_n399), .A2(new_n405), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n851), .B1(KEYINPUT16), .B2(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n659), .B1(new_n853), .B2(new_n417), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n444), .A2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n421), .ZN(new_n856));
  AOI22_X1  g0656(.A1(new_n853), .A2(new_n417), .B1(new_n856), .B2(new_n659), .ZN(new_n857));
  INV_X1    g0657(.A(new_n438), .ZN(new_n858));
  OAI21_X1  g0658(.A(KEYINPUT37), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n420), .A2(new_n421), .ZN(new_n860));
  XNOR2_X1  g0660(.A(new_n659), .B(KEYINPUT102), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n420), .A2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT37), .ZN(new_n863));
  NAND4_X1  g0663(.A1(new_n860), .A2(new_n862), .A3(new_n863), .A4(new_n438), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n859), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n855), .A2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT38), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n855), .A2(KEYINPUT38), .A3(new_n865), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n850), .A2(new_n870), .ZN(new_n871));
  OR2_X1    g0671(.A1(new_n423), .A2(new_n861), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n842), .B1(new_n841), .B2(new_n338), .ZN(new_n874));
  AOI211_X1 g0674(.A(KEYINPUT100), .B(new_n339), .C1(new_n836), .C2(new_n840), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n661), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(new_n877));
  AOI221_X4 g0677(.A(new_n867), .B1(new_n859), .B2(new_n864), .C1(new_n444), .C2(new_n854), .ZN(new_n878));
  AOI21_X1  g0678(.A(KEYINPUT38), .B1(new_n855), .B2(new_n865), .ZN(new_n879));
  OAI21_X1  g0679(.A(KEYINPUT39), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n860), .A2(new_n862), .A3(new_n438), .ZN(new_n881));
  XNOR2_X1  g0681(.A(new_n881), .B(new_n863), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n439), .A2(new_n441), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n862), .B1(new_n423), .B2(new_n883), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n867), .B1(new_n882), .B2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT39), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n869), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n880), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n873), .B1(new_n877), .B2(new_n888), .ZN(new_n889));
  XNOR2_X1  g0689(.A(new_n889), .B(KEYINPUT103), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n715), .A2(new_n445), .A3(new_n718), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n630), .A2(new_n891), .ZN(new_n892));
  XNOR2_X1  g0692(.A(new_n890), .B(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT40), .ZN(new_n894));
  INV_X1    g0694(.A(new_n695), .ZN(new_n895));
  NOR3_X1   g0695(.A1(new_n624), .A2(new_n516), .A3(new_n673), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n895), .B1(new_n896), .B2(new_n700), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n695), .A2(KEYINPUT31), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n793), .B1(new_n848), .B2(new_n849), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n870), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  AND2_X1   g0701(.A1(new_n900), .A2(new_n899), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n894), .B1(new_n869), .B2(new_n885), .ZN(new_n903));
  AOI22_X1  g0703(.A1(new_n894), .A2(new_n901), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  AND3_X1   g0704(.A1(new_n904), .A2(new_n445), .A3(new_n899), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n904), .B1(new_n445), .B2(new_n899), .ZN(new_n906));
  OR3_X1    g0706(.A1(new_n905), .A2(new_n906), .A3(new_n668), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n893), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n908), .B1(new_n207), .B2(new_n721), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n893), .A2(new_n907), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n829), .B1(new_n909), .B2(new_n910), .ZN(G367));
  NAND2_X1  g0711(.A1(new_n727), .A2(new_n241), .ZN(new_n912));
  INV_X1    g0712(.A(new_n736), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n913), .B1(new_n681), .B2(new_n552), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n723), .B1(new_n912), .B2(new_n914), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n638), .A2(new_n661), .ZN(new_n916));
  MUX2_X1   g0716(.A(new_n641), .B(new_n631), .S(new_n916), .Z(new_n917));
  INV_X1    g0717(.A(G317), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n312), .B1(new_n798), .B2(new_n918), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n765), .A2(new_n301), .ZN(new_n920));
  AOI211_X1 g0720(.A(new_n919), .B(new_n920), .C1(G303), .C2(new_n750), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n760), .A2(G116), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n922), .B(KEYINPUT46), .ZN(new_n923));
  AOI22_X1  g0723(.A1(new_n752), .A2(G311), .B1(new_n756), .B2(G107), .ZN(new_n924));
  AOI22_X1  g0724(.A1(G283), .A2(new_n743), .B1(new_n757), .B2(G294), .ZN(new_n925));
  NAND4_X1  g0725(.A1(new_n921), .A2(new_n923), .A3(new_n924), .A4(new_n925), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n926), .B(KEYINPUT108), .ZN(new_n927));
  INV_X1    g0727(.A(new_n809), .ZN(new_n928));
  AOI22_X1  g0728(.A1(new_n752), .A2(new_n928), .B1(new_n743), .B2(G50), .ZN(new_n929));
  INV_X1    g0729(.A(G159), .ZN(new_n930));
  OAI221_X1 g0730(.A(new_n929), .B1(new_n806), .B2(new_n808), .C1(new_n930), .C2(new_n807), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n760), .A2(G58), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n748), .A2(G77), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n755), .A2(new_n203), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n312), .B1(new_n739), .B2(G137), .ZN(new_n936));
  NAND4_X1  g0736(.A1(new_n932), .A2(new_n933), .A3(new_n935), .A4(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n927), .B1(new_n931), .B2(new_n937), .ZN(new_n938));
  XOR2_X1   g0738(.A(new_n938), .B(KEYINPUT47), .Z(new_n939));
  OAI221_X1 g0739(.A(new_n915), .B1(new_n777), .B2(new_n917), .C1(new_n939), .C2(new_n795), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n697), .B1(new_n622), .B2(new_n661), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n650), .A2(new_n673), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(new_n678), .ZN(new_n944));
  OR2_X1    g0744(.A1(new_n944), .A2(KEYINPUT42), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n609), .B1(new_n941), .B2(new_n512), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(new_n661), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n944), .A2(KEYINPUT42), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n945), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n949), .B(KEYINPUT105), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n917), .A2(KEYINPUT43), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n672), .A2(new_n675), .A3(new_n943), .ZN(new_n953));
  OR2_X1    g0753(.A1(new_n953), .A2(KEYINPUT104), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n953), .A2(KEYINPUT104), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  OR2_X1    g0756(.A1(new_n952), .A2(new_n956), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n917), .A2(KEYINPUT43), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n952), .A2(new_n956), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n957), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n952), .A2(new_n956), .ZN(new_n961));
  AOI22_X1  g0761(.A1(new_n950), .A2(new_n951), .B1(new_n954), .B2(new_n955), .ZN(new_n962));
  OAI22_X1  g0762(.A1(new_n961), .A2(new_n962), .B1(KEYINPUT43), .B2(new_n917), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n960), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n722), .A2(G1), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n965), .B(KEYINPUT107), .Z(new_n966));
  INV_X1    g0766(.A(new_n966), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n679), .A2(new_n943), .ZN(new_n968));
  XOR2_X1   g0768(.A(new_n968), .B(KEYINPUT44), .Z(new_n969));
  NAND2_X1  g0769(.A1(new_n679), .A2(new_n943), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(KEYINPUT45), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n972), .B(new_n676), .ZN(new_n973));
  INV_X1    g0773(.A(new_n678), .ZN(new_n974));
  INV_X1    g0774(.A(new_n677), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n974), .B1(new_n675), .B2(new_n975), .ZN(new_n976));
  AND2_X1   g0776(.A1(new_n672), .A2(KEYINPUT106), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n672), .A2(KEYINPUT106), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n976), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  OR2_X1    g0779(.A1(new_n978), .A2(new_n976), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n979), .A2(new_n980), .A3(new_n719), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n719), .B1(new_n973), .B2(new_n981), .ZN(new_n982));
  XOR2_X1   g0782(.A(new_n682), .B(KEYINPUT41), .Z(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n967), .B1(new_n982), .B2(new_n984), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n940), .B1(new_n964), .B2(new_n985), .ZN(G387));
  OAI21_X1  g0786(.A(new_n271), .B1(new_n798), .B2(new_n806), .ZN(new_n987));
  AOI211_X1 g0787(.A(new_n987), .B(new_n920), .C1(G50), .C2(new_n750), .ZN(new_n988));
  INV_X1    g0788(.A(new_n752), .ZN(new_n989));
  OAI22_X1  g0789(.A1(new_n989), .A2(new_n930), .B1(new_n807), .B2(new_n416), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n990), .B1(G68), .B2(new_n743), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n763), .A2(new_n212), .ZN(new_n992));
  INV_X1    g0792(.A(new_n992), .ZN(new_n993));
  AND2_X1   g0793(.A1(new_n553), .A2(new_n555), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(new_n756), .ZN(new_n995));
  NAND4_X1  g0795(.A1(new_n988), .A2(new_n991), .A3(new_n993), .A4(new_n995), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n271), .B1(new_n739), .B2(G326), .ZN(new_n997));
  INV_X1    g0797(.A(G283), .ZN(new_n998));
  OAI22_X1  g0798(.A1(new_n763), .A2(new_n491), .B1(new_n998), .B2(new_n755), .ZN(new_n999));
  AOI22_X1  g0799(.A1(new_n752), .A2(G322), .B1(new_n757), .B2(G311), .ZN(new_n1000));
  INV_X1    g0800(.A(G303), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n1000), .B1(new_n1001), .B2(new_n744), .C1(new_n918), .C2(new_n808), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT48), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n999), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1004), .B1(new_n1003), .B2(new_n1002), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT49), .ZN(new_n1006));
  OAI221_X1 g0806(.A(new_n997), .B1(new_n524), .B2(new_n765), .C1(new_n1005), .C2(new_n1006), .ZN(new_n1007));
  AND2_X1   g0807(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n996), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n723), .B1(new_n1009), .B2(new_n735), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n684), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n725), .A2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(G107), .B2(new_n230), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n238), .A2(G45), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n727), .ZN(new_n1015));
  AOI211_X1 g0815(.A(G45), .B(new_n1011), .C1(G68), .C2(G77), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n253), .A2(new_n201), .ZN(new_n1017));
  XOR2_X1   g0817(.A(new_n1017), .B(KEYINPUT50), .Z(new_n1018));
  AOI21_X1  g0818(.A(new_n1015), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1013), .B1(new_n1014), .B2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n913), .B1(new_n1020), .B2(KEYINPUT109), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1021), .B1(KEYINPUT109), .B2(new_n1020), .ZN(new_n1022));
  OAI211_X1 g0822(.A(new_n1010), .B(new_n1022), .C1(new_n675), .C2(new_n777), .ZN(new_n1023));
  XOR2_X1   g0823(.A(new_n1023), .B(KEYINPUT110), .Z(new_n1024));
  AND2_X1   g0824(.A1(new_n979), .A2(new_n980), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1024), .B1(new_n1025), .B2(new_n967), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n1025), .A2(new_n719), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n981), .A2(new_n682), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1026), .B1(new_n1027), .B2(new_n1028), .ZN(G393));
  OR2_X1    g0829(.A1(new_n972), .A2(new_n676), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n972), .A2(new_n676), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1030), .A2(new_n1031), .A3(new_n967), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n312), .B1(new_n928), .B2(new_n739), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n1033), .B1(new_n763), .B2(new_n203), .C1(new_n214), .C2(new_n765), .ZN(new_n1034));
  XOR2_X1   g0834(.A(new_n1034), .B(KEYINPUT111), .Z(new_n1035));
  AOI22_X1  g0835(.A1(G150), .A2(new_n752), .B1(new_n750), .B2(G159), .ZN(new_n1036));
  XOR2_X1   g0836(.A(new_n1036), .B(KEYINPUT51), .Z(new_n1037));
  NAND2_X1  g0837(.A1(new_n757), .A2(G50), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(G77), .A2(new_n756), .B1(new_n743), .B2(new_n253), .ZN(new_n1039));
  NAND4_X1  g0839(.A1(new_n1035), .A2(new_n1037), .A3(new_n1038), .A4(new_n1039), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(G294), .A2(new_n743), .B1(new_n757), .B2(G303), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1041), .B1(new_n524), .B2(new_n755), .ZN(new_n1042));
  XOR2_X1   g0842(.A(new_n1042), .B(KEYINPUT112), .Z(new_n1043));
  AOI22_X1  g0843(.A1(G311), .A2(new_n750), .B1(new_n752), .B2(G317), .ZN(new_n1044));
  XOR2_X1   g0844(.A(new_n1044), .B(KEYINPUT52), .Z(new_n1045));
  INV_X1    g0845(.A(G322), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n312), .B1(new_n798), .B2(new_n1046), .ZN(new_n1047));
  AOI211_X1 g0847(.A(new_n1047), .B(new_n766), .C1(G283), .C2(new_n760), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1043), .A2(new_n1045), .A3(new_n1048), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n795), .B1(new_n1040), .B2(new_n1049), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n1015), .A2(new_n248), .ZN(new_n1051));
  AOI211_X1 g0851(.A(new_n913), .B(new_n1051), .C1(G97), .C2(new_n681), .ZN(new_n1052));
  NOR3_X1   g0852(.A1(new_n1050), .A2(new_n723), .A3(new_n1052), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(new_n943), .B2(new_n777), .ZN(new_n1054));
  AND2_X1   g0854(.A1(new_n1032), .A2(new_n1054), .ZN(new_n1055));
  AND2_X1   g0855(.A1(new_n973), .A2(new_n981), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n682), .B1(new_n973), .B2(new_n981), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1055), .B1(new_n1056), .B2(new_n1057), .ZN(G390));
  INV_X1    g0858(.A(KEYINPUT113), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n830), .A2(new_n832), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n848), .A2(new_n849), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n877), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n841), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n844), .B1(new_n1063), .B2(new_n342), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n874), .A2(new_n875), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1064), .B1(new_n1065), .B2(new_n847), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n714), .A2(new_n661), .A3(new_n787), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1066), .B1(new_n1067), .B2(new_n832), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n869), .A2(new_n885), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1069), .A2(new_n876), .ZN(new_n1070));
  OAI22_X1  g0870(.A1(new_n888), .A2(new_n1062), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n669), .B(new_n787), .C1(new_n699), .C2(new_n701), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n1072), .A2(new_n1066), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1059), .B1(new_n1071), .B2(new_n1073), .ZN(new_n1074));
  OR2_X1    g0874(.A1(new_n1068), .A2(new_n1070), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n880), .B(new_n887), .C1(new_n850), .C2(new_n877), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n1073), .ZN(new_n1077));
  NAND4_X1  g0877(.A1(new_n1075), .A2(KEYINPUT113), .A3(new_n1076), .A4(new_n1077), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1071), .A2(G330), .A3(new_n902), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1074), .A2(new_n1078), .A3(new_n1079), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n899), .A2(G330), .A3(new_n445), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n630), .A2(new_n891), .A3(new_n1081), .ZN(new_n1082));
  INV_X1    g0882(.A(KEYINPUT114), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NAND4_X1  g0884(.A1(new_n630), .A2(new_n891), .A3(new_n1081), .A4(KEYINPUT114), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n832), .B(new_n1067), .C1(new_n1072), .C2(new_n1066), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n898), .ZN(new_n1087));
  OAI21_X1  g0887(.A(G330), .B1(new_n699), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(KEYINPUT115), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n899), .A2(KEYINPUT115), .A3(G330), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1090), .A2(new_n787), .A3(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1086), .B1(new_n1092), .B2(new_n1066), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1072), .A2(new_n1066), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n900), .A2(new_n899), .A3(G330), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n1094), .A2(new_n1095), .B1(new_n830), .B2(new_n832), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n1084), .B(new_n1085), .C1(new_n1093), .C2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n682), .B1(new_n1080), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(KEYINPUT116), .ZN(new_n1099));
  INV_X1    g0899(.A(KEYINPUT116), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n1100), .B(new_n682), .C1(new_n1080), .C2(new_n1097), .ZN(new_n1101));
  INV_X1    g0901(.A(KEYINPUT117), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1080), .A2(new_n1102), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n1074), .A2(new_n1078), .A3(new_n1079), .A4(KEYINPUT117), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1103), .A2(new_n1097), .A3(new_n1104), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1099), .A2(new_n1101), .A3(new_n1105), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n1080), .A2(new_n966), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n880), .A2(new_n732), .A3(new_n887), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n312), .B1(new_n739), .B2(G125), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(KEYINPUT54), .B(G143), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1109), .B1(new_n744), .B2(new_n1110), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n752), .A2(G128), .B1(new_n757), .B2(G137), .ZN(new_n1112));
  OAI221_X1 g0912(.A(new_n1112), .B1(new_n813), .B2(new_n808), .C1(new_n930), .C2(new_n755), .ZN(new_n1113));
  AOI211_X1 g0913(.A(new_n1111), .B(new_n1113), .C1(G50), .C2(new_n748), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n760), .A2(G150), .ZN(new_n1115));
  XOR2_X1   g0915(.A(new_n1115), .B(KEYINPUT53), .Z(new_n1116));
  OAI22_X1  g0916(.A1(new_n524), .A2(new_n808), .B1(new_n989), .B2(new_n998), .ZN(new_n1117));
  OAI22_X1  g0917(.A1(new_n807), .A2(new_n450), .B1(new_n744), .B2(new_n301), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  OAI221_X1 g0919(.A(new_n312), .B1(new_n755), .B2(new_n212), .C1(new_n491), .C2(new_n798), .ZN(new_n1120));
  AOI211_X1 g0920(.A(new_n1120), .B(new_n764), .C1(G68), .C2(new_n748), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(new_n1114), .A2(new_n1116), .B1(new_n1119), .B2(new_n1121), .ZN(new_n1122));
  OAI221_X1 g0922(.A(new_n724), .B1(new_n253), .B2(new_n796), .C1(new_n1122), .C2(new_n795), .ZN(new_n1123));
  XOR2_X1   g0923(.A(new_n1123), .B(KEYINPUT118), .Z(new_n1124));
  AOI21_X1  g0924(.A(new_n1107), .B1(new_n1108), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1106), .A2(new_n1125), .ZN(G378));
  NAND2_X1  g0926(.A1(new_n900), .A2(new_n899), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n878), .A2(new_n879), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n894), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n903), .A2(new_n899), .A3(new_n900), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1129), .A2(G330), .A3(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n363), .A2(new_n368), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1133));
  XNOR2_X1  g0933(.A(new_n1132), .B(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n365), .A2(new_n660), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(new_n1134), .B(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1131), .A2(new_n1137), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n1129), .A2(G330), .A3(new_n1130), .A4(new_n1136), .ZN(new_n1139));
  AND3_X1   g0939(.A1(new_n1138), .A2(new_n889), .A3(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n889), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1141));
  INV_X1    g0941(.A(KEYINPUT121), .ZN(new_n1142));
  NOR3_X1   g0942(.A1(new_n1140), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n889), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1136), .B1(new_n904), .B2(G330), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1139), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1144), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1138), .A2(new_n889), .A3(new_n1139), .ZN(new_n1148));
  AOI21_X1  g0948(.A(KEYINPUT121), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n1143), .A2(new_n1149), .ZN(new_n1150));
  OR2_X1    g0950(.A1(new_n1080), .A2(new_n1097), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1152), .A2(KEYINPUT122), .ZN(new_n1153));
  INV_X1    g0953(.A(KEYINPUT122), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1084), .A2(new_n1154), .A3(new_n1085), .ZN(new_n1155));
  AND2_X1   g0955(.A1(new_n1153), .A2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(KEYINPUT57), .B1(new_n1151), .B2(new_n1156), .ZN(new_n1157));
  OAI211_X1 g0957(.A(new_n1153), .B(new_n1155), .C1(new_n1080), .C2(new_n1097), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(new_n1150), .A2(new_n1157), .B1(KEYINPUT57), .B2(new_n1160), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n1161), .A2(new_n683), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n724), .B1(G50), .B2(new_n796), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n765), .A2(new_n202), .ZN(new_n1164));
  AOI211_X1 g0964(.A(new_n992), .B(new_n1164), .C1(new_n994), .C2(new_n743), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n750), .A2(G107), .ZN(new_n1166));
  XOR2_X1   g0966(.A(new_n1166), .B(KEYINPUT119), .Z(new_n1167));
  NAND2_X1  g0967(.A1(new_n312), .A2(new_n499), .ZN(new_n1168));
  AOI211_X1 g0968(.A(new_n1168), .B(new_n934), .C1(G283), .C2(new_n739), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(new_n752), .A2(G116), .B1(new_n757), .B2(G97), .ZN(new_n1170));
  NAND4_X1  g0970(.A1(new_n1165), .A2(new_n1167), .A3(new_n1169), .A4(new_n1170), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(new_n1171), .B(KEYINPUT58), .ZN(new_n1172));
  INV_X1    g0972(.A(G137), .ZN(new_n1173));
  OAI22_X1  g0973(.A1(new_n807), .A2(new_n813), .B1(new_n744), .B2(new_n1173), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(G125), .A2(new_n752), .B1(new_n750), .B2(G128), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1175), .B1(new_n806), .B2(new_n755), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1110), .ZN(new_n1177));
  AOI211_X1 g0977(.A(new_n1174), .B(new_n1176), .C1(new_n760), .C2(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT59), .ZN(new_n1179));
  OR2_X1    g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n748), .A2(G159), .ZN(new_n1182));
  AOI211_X1 g0982(.A(G33), .B(G41), .C1(new_n739), .C2(G124), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n1180), .A2(new_n1181), .A3(new_n1182), .A4(new_n1183), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n1168), .B(new_n201), .C1(G33), .C2(G41), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1172), .A2(new_n1184), .A3(new_n1185), .ZN(new_n1186));
  OR2_X1    g0986(.A1(new_n1186), .A2(KEYINPUT120), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n795), .B1(new_n1186), .B2(KEYINPUT120), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1163), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1189), .B1(new_n1136), .B2(new_n733), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1191), .B1(new_n1150), .B2(new_n967), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n1162), .A2(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1194), .ZN(G375));
  NOR2_X1   g0995(.A1(new_n1093), .A2(new_n1096), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1066), .A2(new_n732), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n724), .B1(G68), .B2(new_n796), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n755), .A2(new_n201), .ZN(new_n1200));
  AOI211_X1 g1000(.A(new_n312), .B(new_n1200), .C1(G128), .C2(new_n739), .ZN(new_n1201));
  OAI221_X1 g1001(.A(new_n1201), .B1(new_n763), .B2(new_n930), .C1(new_n202), .C2(new_n765), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n752), .A2(G132), .B1(new_n757), .B2(new_n1177), .ZN(new_n1203));
  OAI221_X1 g1003(.A(new_n1203), .B1(new_n1173), .B2(new_n808), .C1(new_n806), .C2(new_n744), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n752), .A2(G294), .B1(new_n757), .B2(G116), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1205), .B1(new_n450), .B2(new_n744), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n312), .B1(new_n798), .B2(new_n1001), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1207), .B1(new_n750), .B2(G283), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n760), .A2(G97), .ZN(new_n1209));
  NAND4_X1  g1009(.A1(new_n1208), .A2(new_n995), .A3(new_n933), .A4(new_n1209), .ZN(new_n1210));
  OAI22_X1  g1010(.A1(new_n1202), .A2(new_n1204), .B1(new_n1206), .B2(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1199), .B1(new_n1211), .B2(new_n735), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n1197), .A2(new_n967), .B1(new_n1198), .B2(new_n1212), .ZN(new_n1213));
  AND2_X1   g1013(.A1(new_n1196), .A2(new_n1152), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1097), .A2(new_n984), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1213), .B1(new_n1214), .B2(new_n1215), .ZN(G381));
  INV_X1    g1016(.A(G390), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1217), .A2(new_n820), .ZN(new_n1218));
  OR2_X1    g1018(.A1(G393), .A2(G396), .ZN(new_n1219));
  NOR4_X1   g1019(.A1(new_n1218), .A2(G387), .A3(G381), .A4(new_n1219), .ZN(new_n1220));
  XOR2_X1   g1020(.A(new_n1220), .B(KEYINPUT123), .Z(new_n1221));
  INV_X1    g1021(.A(KEYINPUT124), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(G378), .A2(new_n1222), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1106), .A2(KEYINPUT124), .A3(new_n1125), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(G375), .A2(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1226), .ZN(new_n1227));
  OR2_X1    g1027(.A1(new_n1221), .A2(new_n1227), .ZN(G407));
  OAI211_X1 g1028(.A(G407), .B(G213), .C1(G343), .C2(new_n1227), .ZN(G409));
  INV_X1    g1029(.A(KEYINPUT61), .ZN(new_n1230));
  INV_X1    g1030(.A(G343), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1231), .A2(G213), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n983), .B1(new_n1151), .B2(new_n1156), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1150), .A2(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1191), .B1(new_n1159), .B2(new_n967), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1223), .A2(new_n1224), .A3(new_n1237), .ZN(new_n1238));
  OAI211_X1 g1038(.A(G378), .B(new_n1192), .C1(new_n1161), .C2(new_n683), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1233), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1214), .A2(KEYINPUT60), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1196), .A2(new_n1152), .A3(KEYINPUT60), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1242), .A2(new_n682), .A3(new_n1097), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1213), .B1(new_n1241), .B2(new_n1243), .ZN(new_n1244));
  OR2_X1    g1044(.A1(new_n1244), .A2(new_n820), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1244), .A2(new_n820), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(G2897), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1232), .A2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1247), .A2(new_n1249), .ZN(new_n1250));
  OAI211_X1 g1050(.A(new_n1245), .B(new_n1246), .C1(new_n1248), .C2(new_n1232), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1230), .B1(new_n1240), .B2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1247), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1254), .A2(new_n1232), .A3(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1253), .B1(KEYINPUT62), .B2(new_n1256), .ZN(new_n1257));
  OR2_X1    g1057(.A1(new_n1256), .A2(KEYINPUT62), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  OAI211_X1 g1059(.A(G390), .B(new_n940), .C1(new_n964), .C2(new_n985), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT126), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1262));
  XNOR2_X1  g1062(.A(G393), .B(G396), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(G387), .A2(new_n1217), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(new_n1260), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1264), .A2(new_n1266), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1265), .A2(KEYINPUT126), .A3(new_n1260), .A4(new_n1263), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1259), .A2(new_n1270), .ZN(new_n1271));
  AOI211_X1 g1071(.A(new_n1233), .B(new_n1247), .C1(new_n1238), .C2(new_n1239), .ZN(new_n1272));
  OAI21_X1  g1072(.A(KEYINPUT125), .B1(new_n1272), .B2(KEYINPUT63), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT125), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT63), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1256), .A2(new_n1274), .A3(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1273), .A2(new_n1276), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1254), .A2(KEYINPUT63), .A3(new_n1232), .A4(new_n1255), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1278), .A2(new_n1269), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1279), .A2(new_n1253), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT127), .ZN(new_n1281));
  AND3_X1   g1081(.A1(new_n1277), .A2(new_n1280), .A3(new_n1281), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1281), .B1(new_n1277), .B2(new_n1280), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1271), .B1(new_n1282), .B2(new_n1283), .ZN(G405));
  OR2_X1    g1084(.A1(new_n1194), .A2(new_n1225), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1285), .A2(new_n1239), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1286), .A2(new_n1255), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1285), .A2(new_n1247), .A3(new_n1239), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  XNOR2_X1  g1089(.A(new_n1289), .B(new_n1270), .ZN(G402));
endmodule


