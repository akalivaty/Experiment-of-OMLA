//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0 0 0 0 1 1 0 1 1 1 0 0 0 0 0 1 1 1 0 1 0 0 0 0 0 0 0 0 1 1 0 0 0 0 1 0 1 0 0 1 0 1 1 1 0 0 0 0 0 0 0 1 1 1 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:51 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1214, new_n1215, new_n1216, new_n1218, new_n1219,
    new_n1220, new_n1221, new_n1222, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1269,
    new_n1270, new_n1271, new_n1272, new_n1273, new_n1274;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(new_n207), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(new_n201), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(G50), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n218));
  INV_X1    g0018(.A(G77), .ZN(new_n219));
  INV_X1    g0019(.A(G244), .ZN(new_n220));
  INV_X1    g0020(.A(G107), .ZN(new_n221));
  INV_X1    g0021(.A(G264), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n218), .B1(new_n219), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n209), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n212), .B1(new_n215), .B2(new_n217), .C1(KEYINPUT1), .C2(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT2), .B(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XOR2_X1   g0037(.A(G87), .B(G97), .Z(new_n238));
  XNOR2_X1  g0038(.A(G107), .B(G116), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  NAND2_X1  g0040(.A1(new_n202), .A2(G68), .ZN(new_n241));
  INV_X1    g0041(.A(G68), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n242), .A2(G50), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G58), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n240), .B(new_n246), .ZN(G351));
  INV_X1    g0047(.A(G274), .ZN(new_n248));
  INV_X1    g0048(.A(new_n213), .ZN(new_n249));
  NAND2_X1  g0049(.A1(G33), .A2(G41), .ZN(new_n250));
  AOI21_X1  g0050(.A(new_n248), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n213), .B1(G33), .B2(G41), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n256), .A2(new_n253), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n255), .B1(G226), .B2(new_n257), .ZN(new_n258));
  XNOR2_X1  g0058(.A(KEYINPUT3), .B(G33), .ZN(new_n259));
  INV_X1    g0059(.A(G1698), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G222), .ZN(new_n262));
  OAI22_X1  g0062(.A1(new_n261), .A2(new_n262), .B1(new_n219), .B2(new_n259), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n259), .A2(G1698), .ZN(new_n264));
  XNOR2_X1  g0064(.A(new_n264), .B(KEYINPUT64), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n263), .B1(new_n265), .B2(G223), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n249), .A2(new_n250), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n258), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G179), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G13), .ZN(new_n272));
  NOR3_X1   g0072(.A1(new_n272), .A2(new_n207), .A3(G1), .ZN(new_n273));
  NAND3_X1  g0073(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(new_n213), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n206), .A2(G20), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n276), .A2(G50), .A3(new_n277), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n272), .A2(G1), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(G20), .ZN(new_n280));
  XNOR2_X1  g0080(.A(KEYINPUT8), .B(G58), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n207), .A2(G33), .ZN(new_n282));
  INV_X1    g0082(.A(G150), .ZN(new_n283));
  NOR2_X1   g0083(.A1(G20), .A2(G33), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  OAI22_X1  g0085(.A1(new_n281), .A2(new_n282), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n286), .B1(G20), .B2(new_n203), .ZN(new_n287));
  INV_X1    g0087(.A(new_n275), .ZN(new_n288));
  OAI221_X1 g0088(.A(new_n278), .B1(G50), .B2(new_n280), .C1(new_n287), .C2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G169), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n268), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n271), .A2(new_n289), .A3(new_n291), .ZN(new_n292));
  XOR2_X1   g0092(.A(new_n289), .B(KEYINPUT9), .Z(new_n293));
  INV_X1    g0093(.A(G200), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n269), .A2(new_n294), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT10), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n269), .A2(G190), .ZN(new_n298));
  AND3_X1   g0098(.A1(new_n296), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n297), .B1(new_n296), .B2(new_n298), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n292), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G223), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(new_n260), .ZN(new_n303));
  INV_X1    g0103(.A(G226), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(G1698), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(G33), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(KEYINPUT3), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT3), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(G33), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT68), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n308), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n307), .A2(KEYINPUT68), .A3(KEYINPUT3), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n306), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(G87), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n307), .A2(new_n315), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n256), .B1(new_n314), .B2(new_n316), .ZN(new_n317));
  AOI22_X1  g0117(.A1(new_n257), .A2(G232), .B1(new_n251), .B2(new_n253), .ZN(new_n318));
  AND3_X1   g0118(.A1(new_n317), .A2(new_n270), .A3(new_n318), .ZN(new_n319));
  AOI21_X1  g0119(.A(G169), .B1(new_n317), .B2(new_n318), .ZN(new_n320));
  OAI21_X1  g0120(.A(KEYINPUT71), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT72), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT71), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n317), .A2(new_n270), .A3(new_n318), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n267), .A2(new_n252), .ZN(new_n325));
  INV_X1    g0125(.A(G232), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n254), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n316), .ZN(new_n328));
  INV_X1    g0128(.A(new_n313), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n329), .B1(new_n311), .B2(new_n259), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n328), .B1(new_n330), .B2(new_n306), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n327), .B1(new_n331), .B2(new_n256), .ZN(new_n332));
  OAI211_X1 g0132(.A(new_n323), .B(new_n324), .C1(new_n332), .C2(G169), .ZN(new_n333));
  AND3_X1   g0133(.A1(new_n321), .A2(new_n322), .A3(new_n333), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n322), .B1(new_n321), .B2(new_n333), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT16), .ZN(new_n336));
  AND2_X1   g0136(.A1(G58), .A2(G68), .ZN(new_n337));
  OAI21_X1  g0137(.A(G20), .B1(new_n337), .B2(new_n201), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n284), .A2(G159), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT69), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n338), .A2(KEYINPUT69), .A3(new_n339), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT7), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n345), .B1(new_n259), .B2(G20), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n308), .A2(new_n310), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n347), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n242), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n336), .B1(new_n344), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(new_n275), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n312), .A2(new_n313), .A3(new_n207), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(KEYINPUT7), .ZN(new_n353));
  NAND4_X1  g0153(.A1(new_n312), .A2(new_n313), .A3(new_n345), .A4(new_n207), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n353), .A2(G68), .A3(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(new_n343), .ZN(new_n356));
  AOI21_X1  g0156(.A(KEYINPUT69), .B1(new_n338), .B2(new_n339), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n355), .A2(KEYINPUT16), .A3(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT70), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n355), .A2(new_n358), .A3(KEYINPUT70), .A4(KEYINPUT16), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n351), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n276), .ZN(new_n364));
  INV_X1    g0164(.A(new_n281), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(new_n277), .ZN(new_n366));
  OAI22_X1  g0166(.A1(new_n364), .A2(new_n366), .B1(new_n280), .B2(new_n365), .ZN(new_n367));
  OAI22_X1  g0167(.A1(new_n334), .A2(new_n335), .B1(new_n363), .B2(new_n367), .ZN(new_n368));
  XNOR2_X1  g0168(.A(KEYINPUT73), .B(KEYINPUT18), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(new_n351), .ZN(new_n371));
  AND2_X1   g0171(.A1(new_n354), .A2(G68), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n344), .B1(new_n372), .B2(new_n353), .ZN(new_n373));
  AOI21_X1  g0173(.A(KEYINPUT70), .B1(new_n373), .B2(KEYINPUT16), .ZN(new_n374));
  INV_X1    g0174(.A(new_n362), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n371), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n367), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n317), .A2(new_n318), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n378), .A2(G190), .ZN(new_n379));
  AOI21_X1  g0179(.A(G200), .B1(new_n317), .B2(new_n318), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  XOR2_X1   g0182(.A(KEYINPUT74), .B(KEYINPUT17), .Z(new_n383));
  INV_X1    g0183(.A(new_n383), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n376), .A2(new_n377), .A3(new_n382), .A4(new_n384), .ZN(new_n385));
  NOR3_X1   g0185(.A1(new_n363), .A2(new_n367), .A3(new_n381), .ZN(new_n386));
  NOR2_X1   g0186(.A1(KEYINPUT74), .A2(KEYINPUT17), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n385), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NOR3_X1   g0188(.A1(new_n319), .A2(new_n320), .A3(KEYINPUT71), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n378), .A2(new_n290), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n323), .B1(new_n390), .B2(new_n324), .ZN(new_n391));
  OAI21_X1  g0191(.A(KEYINPUT72), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n321), .A2(new_n333), .A3(new_n322), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n376), .A2(new_n377), .ZN(new_n395));
  INV_X1    g0195(.A(new_n369), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n394), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n370), .A2(new_n388), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n284), .A2(G50), .ZN(new_n399));
  XNOR2_X1  g0199(.A(new_n399), .B(KEYINPUT67), .ZN(new_n400));
  OAI22_X1  g0200(.A1(new_n282), .A2(new_n219), .B1(new_n207), .B2(G68), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n275), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT11), .ZN(new_n403));
  OR2_X1    g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n288), .A2(new_n280), .A3(KEYINPUT66), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT66), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n406), .B1(new_n273), .B2(new_n275), .ZN(new_n407));
  AND2_X1   g0207(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n408), .A2(G68), .A3(new_n277), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n402), .A2(new_n403), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n273), .A2(new_n242), .ZN(new_n411));
  XNOR2_X1  g0211(.A(new_n411), .B(KEYINPUT12), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n404), .A2(new_n409), .A3(new_n410), .A4(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT14), .ZN(new_n414));
  NAND2_X1  g0214(.A1(G33), .A2(G97), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n326), .A2(G1698), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n416), .B1(G226), .B2(G1698), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n415), .B1(new_n417), .B2(new_n347), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(new_n256), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n255), .B1(G238), .B2(new_n257), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT13), .ZN(new_n421));
  AND3_X1   g0221(.A1(new_n419), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n421), .B1(new_n420), .B2(new_n419), .ZN(new_n423));
  OAI211_X1 g0223(.A(new_n414), .B(G169), .C1(new_n422), .C2(new_n423), .ZN(new_n424));
  OR2_X1    g0224(.A1(new_n422), .A2(new_n423), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n424), .B1(new_n425), .B2(new_n270), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n414), .B1(new_n425), .B2(G169), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n413), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(new_n413), .ZN(new_n429));
  OAI21_X1  g0229(.A(G200), .B1(new_n422), .B2(new_n423), .ZN(new_n430));
  INV_X1    g0230(.A(G190), .ZN(new_n431));
  OAI211_X1 g0231(.A(new_n429), .B(new_n430), .C1(new_n425), .C2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n428), .A2(new_n432), .ZN(new_n433));
  XNOR2_X1  g0233(.A(KEYINPUT15), .B(G87), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n434), .A2(new_n282), .ZN(new_n435));
  AOI22_X1  g0235(.A1(new_n365), .A2(new_n284), .B1(G20), .B2(G77), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n435), .B1(new_n436), .B2(KEYINPUT65), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n437), .B1(KEYINPUT65), .B2(new_n436), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(new_n275), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n408), .A2(G77), .A3(new_n277), .ZN(new_n440));
  OAI211_X1 g0240(.A(new_n439), .B(new_n440), .C1(G77), .C2(new_n280), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n255), .B1(G244), .B2(new_n257), .ZN(new_n442));
  OAI22_X1  g0242(.A1(new_n261), .A2(new_n326), .B1(new_n221), .B2(new_n259), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n443), .B1(new_n265), .B2(G238), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n442), .B1(new_n444), .B2(new_n267), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n441), .B1(new_n446), .B2(G190), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n447), .B1(new_n294), .B2(new_n446), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n445), .A2(new_n290), .ZN(new_n449));
  AND2_X1   g0249(.A1(new_n441), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n446), .A2(new_n270), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n448), .A2(new_n452), .ZN(new_n453));
  NOR4_X1   g0253(.A1(new_n301), .A2(new_n398), .A3(new_n433), .A4(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(G250), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(new_n260), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n457), .B1(G257), .B2(new_n260), .ZN(new_n458));
  INV_X1    g0258(.A(G294), .ZN(new_n459));
  OAI22_X1  g0259(.A1(new_n330), .A2(new_n458), .B1(new_n307), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(new_n256), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT76), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT5), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n462), .B1(new_n463), .B2(G41), .ZN(new_n464));
  INV_X1    g0264(.A(G41), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n465), .A2(KEYINPUT76), .A3(KEYINPUT5), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n206), .B(G45), .C1(new_n465), .C2(KEYINPUT5), .ZN(new_n468));
  OAI211_X1 g0268(.A(G264), .B(new_n267), .C1(new_n467), .C2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(new_n467), .ZN(new_n470));
  INV_X1    g0270(.A(G45), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n471), .A2(G1), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT75), .ZN(new_n473));
  OAI211_X1 g0273(.A(new_n472), .B(new_n473), .C1(KEYINPUT5), .C2(new_n465), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n468), .A2(KEYINPUT75), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n470), .A2(new_n251), .A3(new_n474), .A4(new_n475), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n461), .A2(new_n469), .A3(new_n476), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n477), .A2(G179), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n478), .B1(new_n290), .B2(new_n477), .ZN(new_n479));
  AOI21_X1  g0279(.A(KEYINPUT23), .B1(new_n221), .B2(G20), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n221), .A2(KEYINPUT23), .A3(G20), .ZN(new_n482));
  INV_X1    g0282(.A(G116), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n307), .A2(new_n483), .ZN(new_n484));
  AOI22_X1  g0284(.A1(new_n481), .A2(new_n482), .B1(new_n484), .B2(new_n207), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n312), .A2(new_n313), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT22), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n487), .A2(new_n315), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n486), .A2(new_n207), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n207), .A2(G87), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n487), .B1(new_n347), .B2(new_n490), .ZN(new_n491));
  AND3_X1   g0291(.A1(new_n489), .A2(KEYINPUT83), .A3(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(KEYINPUT83), .B1(new_n489), .B2(new_n491), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n485), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(KEYINPUT24), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT24), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n496), .B(new_n485), .C1(new_n492), .C2(new_n493), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n288), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n206), .A2(G33), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n276), .A2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(new_n500), .ZN(new_n501));
  AOI21_X1  g0301(.A(KEYINPUT25), .B1(new_n273), .B2(new_n221), .ZN(new_n502));
  INV_X1    g0302(.A(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n273), .A2(KEYINPUT25), .A3(new_n221), .ZN(new_n504));
  AOI22_X1  g0304(.A1(new_n501), .A2(G107), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(new_n505), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n479), .B1(new_n498), .B2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT84), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n479), .B(KEYINPUT84), .C1(new_n498), .C2(new_n506), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n498), .A2(new_n506), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n477), .A2(new_n431), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n512), .B1(G200), .B2(new_n477), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n509), .A2(new_n510), .A3(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT21), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n405), .A2(new_n407), .A3(G116), .A4(new_n499), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n279), .A2(G20), .A3(new_n483), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(G33), .A2(G283), .ZN(new_n520));
  INV_X1    g0320(.A(G97), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n520), .B(new_n207), .C1(G33), .C2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT82), .ZN(new_n523));
  XNOR2_X1  g0323(.A(new_n522), .B(new_n523), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n288), .B1(G20), .B2(new_n483), .ZN(new_n525));
  AOI21_X1  g0325(.A(KEYINPUT20), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n524), .A2(KEYINPUT20), .A3(new_n525), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n519), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(G303), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n259), .A2(new_n530), .ZN(new_n531));
  NOR2_X1   g0331(.A1(G257), .A2(G1698), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n532), .B1(new_n222), .B2(G1698), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n531), .B1(new_n486), .B2(new_n533), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n534), .A2(new_n267), .ZN(new_n535));
  OAI211_X1 g0335(.A(G270), .B(new_n267), .C1(new_n467), .C2(new_n468), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n476), .A2(new_n536), .ZN(new_n537));
  OAI21_X1  g0337(.A(G169), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n516), .B1(new_n529), .B2(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(new_n528), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n518), .B(new_n517), .C1(new_n540), .C2(new_n526), .ZN(new_n541));
  INV_X1    g0341(.A(new_n537), .ZN(new_n542));
  AND2_X1   g0342(.A1(new_n486), .A2(new_n533), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n256), .B1(new_n543), .B2(new_n531), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n541), .A2(KEYINPUT21), .A3(G169), .A4(new_n545), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n535), .A2(new_n537), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n541), .A2(G179), .A3(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n542), .A2(new_n544), .A3(G190), .ZN(new_n549));
  OAI21_X1  g0349(.A(G200), .B1(new_n535), .B2(new_n537), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n529), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  AND4_X1   g0351(.A1(new_n539), .A2(new_n546), .A3(new_n548), .A4(new_n551), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n259), .A2(KEYINPUT4), .A3(G244), .A4(new_n260), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n553), .B(new_n520), .C1(new_n456), .C2(new_n264), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n220), .A2(G1698), .ZN(new_n555));
  AOI21_X1  g0355(.A(KEYINPUT4), .B1(new_n486), .B2(new_n555), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n256), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  OAI211_X1 g0357(.A(G257), .B(new_n267), .C1(new_n467), .C2(new_n468), .ZN(new_n558));
  AND2_X1   g0358(.A1(new_n476), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  OAI21_X1  g0360(.A(KEYINPUT77), .B1(new_n560), .B2(new_n431), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT77), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n557), .A2(new_n559), .A3(new_n562), .A4(G190), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT6), .ZN(new_n565));
  NOR3_X1   g0365(.A1(new_n565), .A2(new_n521), .A3(G107), .ZN(new_n566));
  XNOR2_X1  g0366(.A(G97), .B(G107), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n566), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  OAI22_X1  g0368(.A1(new_n568), .A2(new_n207), .B1(new_n219), .B2(new_n285), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n221), .B1(new_n346), .B2(new_n348), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n275), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n280), .A2(G97), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n572), .B1(new_n501), .B2(G97), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n574), .B1(G200), .B2(new_n560), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n557), .A2(new_n270), .A3(new_n559), .ZN(new_n576));
  AOI22_X1  g0376(.A1(new_n560), .A2(new_n290), .B1(new_n573), .B2(new_n571), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n564), .A2(new_n575), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT81), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n220), .A2(G1698), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n580), .B1(G238), .B2(G1698), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n330), .A2(new_n581), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n256), .B1(new_n582), .B2(new_n484), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n472), .A2(new_n248), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n584), .B(new_n267), .C1(G250), .C2(new_n472), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n579), .B1(new_n586), .B2(new_n431), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n583), .A2(KEYINPUT81), .A3(G190), .A4(new_n585), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n486), .A2(new_n207), .A3(G68), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT19), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n591), .B1(new_n415), .B2(new_n207), .ZN(new_n592));
  NOR2_X1   g0392(.A1(G87), .A2(G97), .ZN(new_n593));
  AND3_X1   g0393(.A1(new_n593), .A2(KEYINPUT78), .A3(new_n221), .ZN(new_n594));
  AOI21_X1  g0394(.A(KEYINPUT78), .B1(new_n593), .B2(new_n221), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n592), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n591), .B1(new_n282), .B2(new_n521), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n590), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(KEYINPUT79), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT79), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n590), .A2(new_n600), .A3(new_n596), .A4(new_n597), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n599), .A2(new_n275), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n434), .A2(new_n273), .ZN(new_n603));
  AND2_X1   g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n501), .A2(G87), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n586), .A2(G200), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n589), .A2(new_n604), .A3(new_n605), .A4(new_n606), .ZN(new_n607));
  OR2_X1    g0407(.A1(new_n500), .A2(new_n434), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n602), .A2(new_n603), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(KEYINPUT80), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT80), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n602), .A2(new_n611), .A3(new_n603), .A4(new_n608), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n586), .A2(G169), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n613), .B1(new_n270), .B2(new_n586), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n610), .A2(new_n612), .A3(new_n614), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n552), .A2(new_n578), .A3(new_n607), .A4(new_n615), .ZN(new_n616));
  NOR3_X1   g0416(.A1(new_n455), .A2(new_n515), .A3(new_n616), .ZN(G372));
  INV_X1    g0417(.A(new_n292), .ZN(new_n618));
  OAI22_X1  g0418(.A1(new_n363), .A2(new_n367), .B1(new_n391), .B2(new_n389), .ZN(new_n619));
  XNOR2_X1  g0419(.A(new_n619), .B(KEYINPUT18), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n432), .A2(new_n450), .A3(new_n451), .ZN(new_n622));
  AND2_X1   g0422(.A1(new_n428), .A2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n388), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n621), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT85), .ZN(new_n626));
  OR2_X1    g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n299), .A2(new_n300), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n628), .B1(new_n625), .B2(new_n626), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n618), .B1(new_n627), .B2(new_n629), .ZN(new_n630));
  AND2_X1   g0430(.A1(new_n577), .A2(new_n576), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n614), .A2(new_n609), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n607), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT26), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n615), .A2(new_n607), .A3(KEYINPUT26), .A4(new_n631), .ZN(new_n636));
  AND2_X1   g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n514), .A2(new_n607), .A3(new_n578), .A4(new_n632), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n546), .A2(new_n548), .ZN(new_n639));
  AND3_X1   g0439(.A1(new_n507), .A2(new_n539), .A3(new_n639), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n632), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n454), .B1(new_n637), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n630), .A2(new_n642), .ZN(G369));
  NAND2_X1  g0443(.A1(new_n639), .A2(new_n539), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n279), .A2(new_n207), .ZN(new_n645));
  OR2_X1    g0445(.A1(new_n645), .A2(KEYINPUT27), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(KEYINPUT27), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n646), .A2(G213), .A3(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(G343), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n644), .A2(new_n541), .A3(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n650), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n552), .B1(new_n529), .B2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT86), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n651), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n655), .B1(new_n654), .B2(new_n651), .ZN(new_n656));
  INV_X1    g0456(.A(G330), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n511), .A2(new_n652), .ZN(new_n659));
  OAI22_X1  g0459(.A1(new_n515), .A2(new_n659), .B1(new_n507), .B2(new_n652), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g0461(.A(new_n661), .B(KEYINPUT87), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n644), .A2(new_n652), .ZN(new_n663));
  XNOR2_X1  g0463(.A(new_n663), .B(KEYINPUT88), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(new_n660), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n665), .B1(new_n507), .B2(new_n650), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n662), .A2(new_n667), .ZN(G399));
  INV_X1    g0468(.A(KEYINPUT89), .ZN(new_n669));
  INV_X1    g0469(.A(new_n210), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n669), .B1(new_n670), .B2(G41), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n210), .A2(KEYINPUT89), .A3(new_n465), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  OR3_X1    g0473(.A1(new_n594), .A2(new_n595), .A3(G116), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n673), .A2(G1), .A3(new_n675), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n676), .B1(new_n217), .B2(new_n673), .ZN(new_n677));
  XNOR2_X1  g0477(.A(new_n677), .B(KEYINPUT28), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT90), .ZN(new_n679));
  AND2_X1   g0479(.A1(new_n509), .A2(new_n510), .ZN(new_n680));
  INV_X1    g0480(.A(new_n616), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n680), .A2(new_n681), .A3(new_n514), .A4(new_n652), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n583), .A2(new_n461), .A3(new_n469), .A4(new_n585), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n542), .A2(new_n544), .A3(G179), .ZN(new_n684));
  NOR3_X1   g0484(.A1(new_n683), .A2(new_n684), .A3(new_n560), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(KEYINPUT30), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n547), .A2(G179), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n688), .A2(new_n477), .A3(new_n586), .A4(new_n560), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n689), .B1(new_n685), .B2(KEYINPUT30), .ZN(new_n690));
  OAI211_X1 g0490(.A(KEYINPUT31), .B(new_n650), .C1(new_n687), .C2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT30), .ZN(new_n693));
  OR2_X1    g0493(.A1(new_n683), .A2(new_n684), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n693), .B1(new_n694), .B2(new_n560), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n695), .A2(new_n686), .A3(new_n689), .ZN(new_n696));
  AOI21_X1  g0496(.A(KEYINPUT31), .B1(new_n696), .B2(new_n650), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n692), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n682), .A2(new_n698), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n679), .B1(new_n699), .B2(G330), .ZN(new_n700));
  AOI211_X1 g0500(.A(KEYINPUT90), .B(new_n657), .C1(new_n682), .C2(new_n698), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n652), .B1(new_n641), .B2(new_n637), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT29), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n644), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n638), .B1(new_n680), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n633), .A2(KEYINPUT26), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n615), .A2(new_n607), .A3(new_n634), .A4(new_n631), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n708), .A2(new_n632), .A3(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n652), .B1(new_n707), .B2(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n705), .B1(new_n704), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n702), .A2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n678), .B1(new_n714), .B2(G1), .ZN(G364));
  INV_X1    g0515(.A(new_n673), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n272), .A2(G20), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n206), .B1(new_n717), .B2(G45), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n716), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n658), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n656), .A2(new_n657), .ZN(new_n722));
  NOR2_X1   g0522(.A1(G13), .A2(G33), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n724), .A2(G20), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n656), .A2(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n290), .A2(KEYINPUT92), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n207), .B1(KEYINPUT92), .B2(new_n290), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n213), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(G179), .A2(G200), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n207), .B1(new_n731), .B2(G190), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n732), .A2(new_n459), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n207), .A2(G190), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n294), .A2(G179), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(G283), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n347), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NAND3_X1  g0538(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n739), .A2(new_n431), .ZN(new_n740));
  AOI211_X1 g0540(.A(new_n733), .B(new_n738), .C1(G326), .C2(new_n740), .ZN(new_n741));
  XNOR2_X1  g0541(.A(KEYINPUT33), .B(G317), .ZN(new_n742));
  OR2_X1    g0542(.A1(new_n742), .A2(KEYINPUT95), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n739), .A2(G190), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n742), .A2(KEYINPUT95), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n743), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n207), .A2(new_n431), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n270), .A2(G200), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n748), .A2(new_n734), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  AOI22_X1  g0552(.A1(G322), .A2(new_n750), .B1(new_n752), .B2(G311), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n747), .A2(new_n735), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n734), .A2(new_n731), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  AOI22_X1  g0557(.A1(G303), .A2(new_n755), .B1(new_n757), .B2(G329), .ZN(new_n758));
  NAND4_X1  g0558(.A1(new_n741), .A2(new_n746), .A3(new_n753), .A4(new_n758), .ZN(new_n759));
  XOR2_X1   g0559(.A(new_n759), .B(KEYINPUT96), .Z(new_n760));
  AND2_X1   g0560(.A1(new_n751), .A2(KEYINPUT93), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n751), .A2(KEYINPUT93), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  AOI22_X1  g0564(.A1(new_n764), .A2(G77), .B1(G58), .B2(new_n750), .ZN(new_n765));
  AND2_X1   g0565(.A1(new_n765), .A2(KEYINPUT94), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n765), .A2(KEYINPUT94), .ZN(new_n767));
  INV_X1    g0567(.A(G159), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n756), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(KEYINPUT32), .ZN(new_n770));
  INV_X1    g0570(.A(new_n732), .ZN(new_n771));
  AOI22_X1  g0571(.A1(new_n769), .A2(new_n770), .B1(new_n771), .B2(G97), .ZN(new_n772));
  INV_X1    g0572(.A(new_n744), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n772), .B1(new_n242), .B2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n740), .ZN(new_n775));
  OAI22_X1  g0575(.A1(new_n769), .A2(new_n770), .B1(new_n202), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n755), .A2(G87), .ZN(new_n777));
  OAI211_X1 g0577(.A(new_n777), .B(new_n259), .C1(new_n221), .C2(new_n736), .ZN(new_n778));
  OR3_X1    g0578(.A1(new_n774), .A2(new_n776), .A3(new_n778), .ZN(new_n779));
  NOR3_X1   g0579(.A1(new_n766), .A2(new_n767), .A3(new_n779), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n730), .B1(new_n760), .B2(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n730), .A2(new_n725), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n670), .A2(new_n347), .ZN(new_n784));
  AOI22_X1  g0584(.A1(new_n784), .A2(G355), .B1(new_n483), .B2(new_n670), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n670), .A2(new_n486), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n786), .B1(G45), .B2(new_n217), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n246), .A2(new_n471), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n785), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n783), .B1(new_n789), .B2(KEYINPUT91), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n790), .B1(KEYINPUT91), .B2(new_n789), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n781), .A2(new_n720), .A3(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  AOI22_X1  g0593(.A1(new_n721), .A2(new_n722), .B1(new_n726), .B2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(G396));
  NOR2_X1   g0595(.A1(new_n452), .A2(new_n650), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n441), .A2(new_n650), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n448), .A2(new_n797), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n796), .B1(new_n798), .B2(new_n452), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n703), .A2(new_n800), .ZN(new_n801));
  OAI211_X1 g0601(.A(new_n652), .B(new_n799), .C1(new_n641), .C2(new_n637), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n720), .B1(new_n702), .B2(new_n803), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n804), .B1(new_n702), .B2(new_n803), .ZN(new_n805));
  INV_X1    g0605(.A(new_n730), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n806), .A2(new_n724), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n720), .B1(G77), .B2(new_n807), .ZN(new_n808));
  AOI22_X1  g0608(.A1(new_n750), .A2(G143), .B1(G137), .B2(new_n740), .ZN(new_n809));
  OAI221_X1 g0609(.A(new_n809), .B1(new_n283), .B2(new_n773), .C1(new_n763), .C2(new_n768), .ZN(new_n810));
  XNOR2_X1  g0610(.A(new_n810), .B(KEYINPUT34), .ZN(new_n811));
  INV_X1    g0611(.A(new_n736), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(G68), .ZN(new_n813));
  INV_X1    g0613(.A(G132), .ZN(new_n814));
  OAI221_X1 g0614(.A(new_n813), .B1(new_n202), .B2(new_n754), .C1(new_n814), .C2(new_n756), .ZN(new_n815));
  AOI211_X1 g0615(.A(new_n330), .B(new_n815), .C1(G58), .C2(new_n771), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n811), .A2(new_n816), .ZN(new_n817));
  OAI22_X1  g0617(.A1(new_n749), .A2(new_n459), .B1(new_n732), .B2(new_n521), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n818), .B(KEYINPUT97), .ZN(new_n819));
  OAI22_X1  g0619(.A1(new_n773), .A2(new_n737), .B1(new_n775), .B2(new_n530), .ZN(new_n820));
  INV_X1    g0620(.A(G311), .ZN(new_n821));
  OAI22_X1  g0621(.A1(new_n754), .A2(new_n221), .B1(new_n756), .B2(new_n821), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n347), .B1(new_n736), .B2(new_n315), .ZN(new_n823));
  NOR3_X1   g0623(.A1(new_n820), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n824), .B1(new_n483), .B2(new_n763), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n817), .B1(new_n819), .B2(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n808), .B1(new_n826), .B2(new_n730), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n827), .B1(new_n799), .B2(new_n724), .ZN(new_n828));
  AND2_X1   g0628(.A1(new_n805), .A2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(G384));
  INV_X1    g0630(.A(new_n568), .ZN(new_n831));
  AOI211_X1 g0631(.A(new_n483), .B(new_n215), .C1(new_n831), .C2(KEYINPUT35), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n832), .B1(KEYINPUT35), .B2(new_n831), .ZN(new_n833));
  XNOR2_X1  g0633(.A(KEYINPUT98), .B(KEYINPUT36), .ZN(new_n834));
  XNOR2_X1  g0634(.A(new_n833), .B(new_n834), .ZN(new_n835));
  OR3_X1    g0635(.A1(new_n217), .A2(new_n219), .A3(new_n337), .ZN(new_n836));
  AOI211_X1 g0636(.A(new_n206), .B(G13), .C1(new_n836), .C2(new_n241), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT102), .ZN(new_n839));
  INV_X1    g0639(.A(new_n648), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n840), .B1(new_n363), .B2(new_n367), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n841), .B1(new_n621), .B2(new_n388), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n376), .A2(new_n377), .A3(new_n382), .ZN(new_n843));
  AND2_X1   g0643(.A1(new_n843), .A2(new_n841), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(new_n619), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n845), .A2(KEYINPUT37), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT37), .ZN(new_n847));
  NAND4_X1  g0647(.A1(new_n368), .A2(new_n847), .A3(new_n843), .A4(new_n841), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT100), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(KEYINPUT37), .B1(new_n394), .B2(new_n395), .ZN(new_n851));
  AOI21_X1  g0651(.A(KEYINPUT100), .B1(new_n851), .B2(new_n844), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n846), .B1(new_n850), .B2(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n842), .B1(new_n853), .B2(KEYINPUT101), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n848), .A2(new_n849), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n851), .A2(new_n844), .A3(KEYINPUT100), .ZN(new_n856));
  AOI22_X1  g0656(.A1(new_n855), .A2(new_n856), .B1(KEYINPUT37), .B2(new_n845), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT101), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  AOI21_X1  g0659(.A(KEYINPUT38), .B1(new_n854), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n355), .A2(new_n358), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n288), .B1(new_n861), .B2(new_n336), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n862), .B1(new_n374), .B2(new_n375), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n648), .B1(new_n863), .B2(new_n377), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n398), .A2(new_n864), .ZN(new_n865));
  AOI22_X1  g0665(.A1(new_n863), .A2(new_n377), .B1(new_n321), .B2(new_n333), .ZN(new_n866));
  NOR3_X1   g0666(.A1(new_n866), .A2(new_n864), .A3(new_n386), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n848), .B1(new_n867), .B2(new_n847), .ZN(new_n868));
  AND3_X1   g0668(.A1(new_n865), .A2(KEYINPUT38), .A3(new_n868), .ZN(new_n869));
  OR2_X1    g0669(.A1(new_n869), .A2(KEYINPUT39), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n839), .B1(new_n860), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(KEYINPUT38), .B1(new_n865), .B2(new_n868), .ZN(new_n872));
  OAI21_X1  g0672(.A(KEYINPUT39), .B1(new_n869), .B2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT99), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  OAI211_X1 g0675(.A(KEYINPUT99), .B(KEYINPUT39), .C1(new_n869), .C2(new_n872), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT38), .ZN(new_n878));
  OAI211_X1 g0678(.A(new_n395), .B(new_n840), .C1(new_n620), .C2(new_n624), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n879), .B1(new_n857), .B2(new_n858), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n853), .A2(KEYINPUT101), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n878), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n869), .A2(KEYINPUT39), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n882), .A2(KEYINPUT102), .A3(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n871), .A2(new_n877), .A3(new_n884), .ZN(new_n885));
  OR2_X1    g0685(.A1(new_n428), .A2(new_n650), .ZN(new_n886));
  INV_X1    g0686(.A(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n796), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n802), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n413), .A2(new_n650), .ZN(new_n891));
  XNOR2_X1  g0691(.A(new_n433), .B(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n890), .A2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  OR2_X1    g0695(.A1(new_n869), .A2(new_n872), .ZN(new_n896));
  AOI22_X1  g0696(.A1(new_n895), .A2(new_n896), .B1(new_n620), .B2(new_n648), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n888), .A2(new_n897), .ZN(new_n898));
  OAI211_X1 g0698(.A(new_n705), .B(new_n454), .C1(new_n704), .C2(new_n711), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(new_n630), .ZN(new_n900));
  XOR2_X1   g0700(.A(new_n900), .B(KEYINPUT103), .Z(new_n901));
  XNOR2_X1  g0701(.A(new_n898), .B(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT105), .ZN(new_n903));
  XNOR2_X1  g0703(.A(new_n691), .B(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n696), .A2(new_n650), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT31), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n907), .A2(KEYINPUT104), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT104), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n697), .A2(new_n909), .ZN(new_n910));
  OAI211_X1 g0710(.A(new_n904), .B(new_n682), .C1(new_n908), .C2(new_n910), .ZN(new_n911));
  AND3_X1   g0711(.A1(new_n911), .A2(new_n799), .A3(new_n893), .ZN(new_n912));
  AOI21_X1  g0712(.A(KEYINPUT40), .B1(new_n912), .B2(new_n896), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(KEYINPUT40), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  OR2_X1    g0715(.A1(new_n860), .A2(new_n869), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n913), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  AND2_X1   g0717(.A1(new_n911), .A2(new_n454), .ZN(new_n918));
  OR2_X1    g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n917), .A2(new_n918), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n919), .A2(G330), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n902), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n922), .B1(new_n206), .B2(new_n717), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n902), .A2(new_n921), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n838), .B1(new_n923), .B2(new_n924), .ZN(G367));
  NAND2_X1  g0725(.A1(new_n607), .A2(new_n632), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n652), .B1(new_n604), .B2(new_n605), .ZN(new_n927));
  MUX2_X1   g0727(.A(new_n926), .B(new_n632), .S(new_n927), .Z(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(KEYINPUT43), .ZN(new_n930));
  INV_X1    g0730(.A(new_n574), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n578), .B1(new_n931), .B2(new_n652), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n631), .A2(new_n650), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(KEYINPUT42), .B1(new_n665), .B2(new_n935), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n680), .A2(new_n932), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n652), .B1(new_n937), .B2(new_n631), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  NOR3_X1   g0739(.A1(new_n665), .A2(KEYINPUT42), .A3(new_n935), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n930), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n929), .A2(KEYINPUT43), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n941), .B(new_n942), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n662), .A2(new_n935), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n943), .B(new_n944), .ZN(new_n945));
  XNOR2_X1  g0745(.A(KEYINPUT106), .B(KEYINPUT41), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n673), .B(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n667), .A2(new_n934), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT45), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n949), .B(new_n950), .ZN(new_n951));
  OAI211_X1 g0751(.A(new_n666), .B(new_n935), .C1(KEYINPUT107), .C2(KEYINPUT44), .ZN(new_n952));
  NAND2_X1  g0752(.A1(KEYINPUT107), .A2(KEYINPUT44), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n952), .B(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n951), .A2(new_n954), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n662), .A2(KEYINPUT108), .ZN(new_n956));
  OR2_X1    g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n955), .A2(new_n956), .ZN(new_n958));
  XOR2_X1   g0758(.A(new_n658), .B(new_n660), .Z(new_n959));
  XOR2_X1   g0759(.A(new_n959), .B(new_n664), .Z(new_n960));
  NAND4_X1  g0760(.A1(new_n957), .A2(new_n714), .A3(new_n958), .A4(new_n960), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n948), .B1(new_n961), .B2(new_n714), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n945), .B1(new_n962), .B2(new_n719), .ZN(new_n963));
  INV_X1    g0763(.A(new_n786), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n964), .A2(new_n236), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n782), .B1(new_n210), .B2(new_n434), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n720), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  AOI22_X1  g0767(.A1(G58), .A2(new_n755), .B1(new_n750), .B2(G150), .ZN(new_n968));
  INV_X1    g0768(.A(G137), .ZN(new_n969));
  OAI221_X1 g0769(.A(new_n968), .B1(new_n969), .B2(new_n756), .C1(new_n763), .C2(new_n202), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n732), .A2(new_n242), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n812), .A2(G77), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n972), .A2(new_n259), .ZN(new_n973));
  INV_X1    g0773(.A(G143), .ZN(new_n974));
  OAI22_X1  g0774(.A1(new_n773), .A2(new_n768), .B1(new_n775), .B2(new_n974), .ZN(new_n975));
  NOR4_X1   g0775(.A1(new_n970), .A2(new_n971), .A3(new_n973), .A4(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n755), .A2(G116), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT46), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n979), .B(KEYINPUT109), .Z(new_n980));
  AOI22_X1  g0780(.A1(new_n977), .A2(new_n978), .B1(new_n744), .B2(G294), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  XOR2_X1   g0782(.A(new_n982), .B(KEYINPUT110), .Z(new_n983));
  NOR2_X1   g0783(.A1(new_n763), .A2(new_n737), .ZN(new_n984));
  OAI221_X1 g0784(.A(new_n330), .B1(new_n221), .B2(new_n732), .C1(new_n775), .C2(new_n821), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n736), .A2(new_n521), .ZN(new_n986));
  INV_X1    g0786(.A(G317), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n749), .A2(new_n530), .B1(new_n756), .B2(new_n987), .ZN(new_n988));
  NOR4_X1   g0788(.A1(new_n984), .A2(new_n985), .A3(new_n986), .A4(new_n988), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n976), .B1(new_n983), .B2(new_n989), .ZN(new_n990));
  XOR2_X1   g0790(.A(new_n990), .B(KEYINPUT47), .Z(new_n991));
  AOI21_X1  g0791(.A(new_n967), .B1(new_n991), .B2(new_n730), .ZN(new_n992));
  INV_X1    g0792(.A(new_n725), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n992), .B1(new_n993), .B2(new_n929), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n963), .A2(new_n994), .ZN(G387));
  OR2_X1    g0795(.A1(new_n660), .A2(new_n993), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n786), .B1(new_n233), .B2(new_n471), .ZN(new_n997));
  INV_X1    g0797(.A(new_n784), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n997), .B1(new_n675), .B2(new_n998), .ZN(new_n999));
  OR3_X1    g0799(.A1(new_n281), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1000));
  OAI21_X1  g0800(.A(KEYINPUT50), .B1(new_n281), .B2(G50), .ZN(new_n1001));
  AOI21_X1  g0801(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1002));
  NAND4_X1  g0802(.A1(new_n675), .A2(new_n1000), .A3(new_n1001), .A4(new_n1002), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(new_n999), .A2(new_n1003), .B1(new_n221), .B2(new_n670), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n720), .B1(new_n1004), .B2(new_n783), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n775), .A2(new_n768), .B1(new_n732), .B2(new_n434), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n1006), .B1(new_n365), .B2(new_n744), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n751), .A2(new_n242), .B1(new_n756), .B2(new_n283), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1008), .B1(G50), .B2(new_n750), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n986), .B1(G77), .B2(new_n755), .ZN(new_n1010));
  NAND4_X1  g0810(.A1(new_n1007), .A2(new_n1009), .A3(new_n486), .A4(new_n1010), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(G116), .A2(new_n812), .B1(new_n757), .B2(G326), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n754), .A2(new_n459), .B1(new_n732), .B2(new_n737), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n773), .A2(new_n821), .B1(new_n749), .B2(new_n987), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1014), .B1(G322), .B2(new_n740), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1015), .B1(new_n530), .B2(new_n763), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT48), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1013), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1018), .B1(new_n1017), .B2(new_n1016), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT49), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n330), .B(new_n1012), .C1(new_n1019), .C2(new_n1020), .ZN(new_n1021));
  AND2_X1   g0821(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1011), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g0823(.A(KEYINPUT111), .ZN(new_n1024));
  OR2_X1    g0824(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n806), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1005), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n960), .A2(new_n719), .B1(new_n996), .B2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n960), .A2(new_n714), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1029), .A2(KEYINPUT112), .A3(new_n716), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1030), .B1(new_n714), .B2(new_n960), .ZN(new_n1031));
  AOI21_X1  g0831(.A(KEYINPUT112), .B1(new_n1029), .B2(new_n716), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1028), .B1(new_n1031), .B2(new_n1032), .ZN(G393));
  NAND2_X1  g0833(.A1(new_n961), .A2(new_n716), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n955), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1035), .A2(new_n662), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n1036), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n1035), .A2(new_n662), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1029), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  INV_X1    g0839(.A(KEYINPUT114), .ZN(new_n1040));
  OR2_X1    g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1034), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  OR3_X1    g0843(.A1(new_n1037), .A2(new_n718), .A3(new_n1038), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n964), .A2(new_n240), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n782), .B1(new_n521), .B2(new_n210), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n720), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n347), .B1(new_n736), .B2(new_n221), .C1(new_n773), .C2(new_n530), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1048), .B1(G116), .B2(new_n771), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n775), .A2(new_n987), .B1(new_n749), .B2(new_n821), .ZN(new_n1050));
  XOR2_X1   g0850(.A(KEYINPUT113), .B(KEYINPUT52), .Z(new_n1051));
  XNOR2_X1  g0851(.A(new_n1050), .B(new_n1051), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n754), .A2(new_n737), .B1(new_n751), .B2(new_n459), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1053), .B1(G322), .B2(new_n757), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1049), .A2(new_n1052), .A3(new_n1054), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n732), .A2(new_n219), .ZN(new_n1056));
  AOI211_X1 g0856(.A(new_n1056), .B(new_n330), .C1(G50), .C2(new_n744), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n736), .A2(new_n315), .B1(new_n756), .B2(new_n974), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(G68), .B2(new_n755), .ZN(new_n1059));
  OAI211_X1 g0859(.A(new_n1057), .B(new_n1059), .C1(new_n281), .C2(new_n763), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n750), .A2(G159), .B1(G150), .B2(new_n740), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n1061), .B(KEYINPUT51), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1055), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1047), .B1(new_n1063), .B2(new_n730), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1064), .B1(new_n934), .B2(new_n993), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1044), .A2(new_n1065), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n1043), .A2(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n1067), .ZN(G390));
  NAND2_X1  g0868(.A1(new_n894), .A2(new_n886), .ZN(new_n1069));
  NAND4_X1  g0869(.A1(new_n871), .A2(new_n877), .A3(new_n884), .A4(new_n1069), .ZN(new_n1070));
  AND2_X1   g0870(.A1(new_n798), .A2(new_n452), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n889), .B1(new_n711), .B2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n887), .B1(new_n1072), .B2(new_n893), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n916), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1070), .A2(new_n1074), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n800), .A2(new_n657), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n911), .A2(new_n893), .A3(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1075), .A2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(KEYINPUT115), .ZN(new_n1080));
  NOR3_X1   g0880(.A1(new_n515), .A2(new_n616), .A3(new_n650), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n907), .A2(new_n691), .ZN(new_n1082));
  OAI21_X1  g0882(.A(G330), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1083), .A2(KEYINPUT90), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n699), .A2(new_n679), .A3(G330), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n800), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1086), .A2(new_n893), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1070), .A2(new_n1074), .A3(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(KEYINPUT115), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1075), .A2(new_n1089), .A3(new_n1078), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1080), .A2(new_n1088), .A3(new_n1090), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n1091), .A2(new_n718), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n771), .A2(G159), .B1(G137), .B2(new_n744), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(KEYINPUT54), .B(G143), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1093), .B1(new_n763), .B2(new_n1094), .ZN(new_n1095));
  XOR2_X1   g0895(.A(new_n1095), .B(KEYINPUT118), .Z(new_n1096));
  NAND2_X1  g0896(.A1(new_n755), .A2(G150), .ZN(new_n1097));
  OR2_X1    g0897(.A1(new_n1097), .A2(KEYINPUT53), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n1097), .A2(KEYINPUT53), .B1(new_n740), .B2(G128), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n347), .B1(new_n812), .B2(G50), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(G132), .A2(new_n750), .B1(new_n757), .B2(G125), .ZN(new_n1101));
  NAND4_X1  g0901(.A1(new_n1098), .A2(new_n1099), .A3(new_n1100), .A4(new_n1101), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n1096), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1056), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(G107), .A2(new_n744), .B1(new_n740), .B2(G283), .ZN(new_n1105));
  NAND4_X1  g0905(.A1(new_n777), .A2(new_n1104), .A3(new_n1105), .A4(new_n347), .ZN(new_n1106));
  OAI221_X1 g0906(.A(new_n813), .B1(new_n483), .B2(new_n749), .C1(new_n459), .C2(new_n756), .ZN(new_n1107));
  AOI211_X1 g0907(.A(new_n1106), .B(new_n1107), .C1(G97), .C2(new_n764), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n730), .B1(new_n1103), .B2(new_n1108), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n1109), .B(new_n720), .C1(new_n365), .C2(new_n807), .ZN(new_n1110));
  XOR2_X1   g0910(.A(new_n1110), .B(KEYINPUT119), .Z(new_n1111));
  OAI21_X1  g0911(.A(new_n1111), .B1(new_n885), .B2(new_n724), .ZN(new_n1112));
  XOR2_X1   g0912(.A(new_n1112), .B(KEYINPUT120), .Z(new_n1113));
  NOR2_X1   g0913(.A1(new_n1092), .A2(new_n1113), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1077), .B1(new_n1086), .B2(new_n893), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n893), .B1(new_n911), .B2(new_n1076), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n1116), .A2(new_n1072), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n1115), .A2(new_n890), .B1(new_n1087), .B2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n918), .A2(KEYINPUT116), .A3(G330), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n911), .A2(new_n454), .A3(G330), .ZN(new_n1120));
  INV_X1    g0920(.A(KEYINPUT116), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1119), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n900), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  OAI21_X1  g0925(.A(KEYINPUT117), .B1(new_n1118), .B2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT117), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n900), .B1(new_n1122), .B2(new_n1119), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n890), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n799), .B1(new_n700), .B2(new_n701), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1130), .A2(new_n892), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1129), .B1(new_n1131), .B2(new_n1077), .ZN(new_n1132));
  AOI211_X1 g0932(.A(new_n1072), .B(new_n1116), .C1(new_n1086), .C2(new_n893), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n1127), .B(new_n1128), .C1(new_n1132), .C2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1126), .A2(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1091), .A2(new_n1136), .ZN(new_n1137));
  NAND4_X1  g0937(.A1(new_n1135), .A2(new_n1080), .A3(new_n1088), .A4(new_n1090), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1137), .A2(new_n716), .A3(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1114), .A2(new_n1139), .ZN(G378));
  NAND2_X1  g0940(.A1(new_n1138), .A2(new_n1128), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1141), .A2(KEYINPUT122), .ZN(new_n1142));
  INV_X1    g0942(.A(KEYINPUT122), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1138), .A2(new_n1143), .A3(new_n1128), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n917), .A2(G330), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n289), .A2(new_n840), .ZN(new_n1147));
  XOR2_X1   g0947(.A(new_n301), .B(new_n1147), .Z(new_n1148));
  XNOR2_X1  g0948(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(new_n1148), .B(new_n1149), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n1146), .A2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1146), .A2(new_n1150), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n1152), .A2(new_n888), .A3(new_n897), .A4(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1153), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n898), .B1(new_n1155), .B2(new_n1151), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1154), .A2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(KEYINPUT57), .B1(new_n1145), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(KEYINPUT57), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1159), .B1(new_n1154), .B2(new_n1156), .ZN(new_n1160));
  AND3_X1   g0960(.A1(new_n1138), .A2(new_n1143), .A3(new_n1128), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1143), .B1(new_n1138), .B2(new_n1128), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1160), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1163), .A2(new_n716), .ZN(new_n1164));
  OR2_X1    g0964(.A1(new_n1158), .A2(new_n1164), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n720), .B1(G50), .B2(new_n807), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n486), .A2(G41), .ZN(new_n1167));
  AOI211_X1 g0967(.A(G50), .B(new_n1167), .C1(new_n307), .C2(new_n465), .ZN(new_n1168));
  AND2_X1   g0968(.A1(new_n812), .A2(G58), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1169), .B1(G283), .B2(new_n757), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n1170), .B(new_n1167), .C1(new_n434), .C2(new_n751), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n773), .A2(new_n521), .B1(new_n775), .B2(new_n483), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n219), .A2(new_n754), .B1(new_n749), .B2(new_n221), .ZN(new_n1173));
  NOR4_X1   g0973(.A1(new_n1171), .A2(new_n1172), .A3(new_n971), .A4(new_n1173), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1168), .B1(new_n1174), .B2(KEYINPUT58), .ZN(new_n1175));
  OAI22_X1  g0975(.A1(new_n773), .A2(new_n814), .B1(new_n732), .B2(new_n283), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n750), .A2(G128), .ZN(new_n1177));
  OAI221_X1 g0977(.A(new_n1177), .B1(new_n969), .B2(new_n751), .C1(new_n754), .C2(new_n1094), .ZN(new_n1178));
  AOI211_X1 g0978(.A(new_n1176), .B(new_n1178), .C1(G125), .C2(new_n740), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n1180), .A2(KEYINPUT59), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n307), .B(new_n465), .C1(new_n736), .C2(new_n768), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1182), .B1(G124), .B2(new_n757), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT59), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1183), .B1(new_n1179), .B2(new_n1184), .ZN(new_n1185));
  OAI221_X1 g0985(.A(new_n1175), .B1(KEYINPUT58), .B2(new_n1174), .C1(new_n1181), .C2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1166), .B1(new_n1186), .B2(new_n730), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1150), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1187), .B1(new_n1188), .B2(new_n724), .ZN(new_n1189));
  XOR2_X1   g0989(.A(new_n1189), .B(KEYINPUT121), .Z(new_n1190));
  AOI21_X1  g0990(.A(new_n1190), .B1(new_n1157), .B2(new_n719), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1165), .A2(new_n1191), .ZN(G375));
  INV_X1    g0992(.A(new_n1118), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n892), .A2(new_n723), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n720), .B1(G68), .B2(new_n807), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1169), .B1(G128), .B2(new_n757), .ZN(new_n1196));
  OAI22_X1  g0996(.A1(new_n969), .A2(new_n749), .B1(new_n754), .B2(new_n768), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(G150), .B2(new_n752), .ZN(new_n1198));
  OAI22_X1  g0998(.A1(new_n773), .A2(new_n1094), .B1(new_n202), .B2(new_n732), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1199), .B1(G132), .B2(new_n740), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n1196), .A2(new_n486), .A3(new_n1198), .A4(new_n1200), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(G97), .A2(new_n755), .B1(new_n757), .B2(G303), .ZN(new_n1202));
  AND3_X1   g1002(.A1(new_n1202), .A2(new_n347), .A3(new_n972), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(G116), .A2(new_n744), .B1(new_n740), .B2(G294), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n1203), .B(new_n1204), .C1(new_n221), .C2(new_n763), .ZN(new_n1205));
  OAI22_X1  g1005(.A1(new_n749), .A2(new_n737), .B1(new_n732), .B2(new_n434), .ZN(new_n1206));
  XOR2_X1   g1006(.A(new_n1206), .B(KEYINPUT123), .Z(new_n1207));
  OAI21_X1  g1007(.A(new_n1201), .B1(new_n1205), .B2(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1195), .B1(new_n1208), .B2(new_n730), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n1193), .A2(new_n719), .B1(new_n1194), .B2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1118), .A2(new_n1125), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1211), .A2(new_n947), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1210), .B1(new_n1135), .B2(new_n1212), .ZN(G381));
  OR4_X1    g1013(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1214));
  NOR3_X1   g1014(.A1(new_n1214), .A2(G387), .A3(G381), .ZN(new_n1215));
  INV_X1    g1015(.A(G378), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1215), .A2(new_n1216), .A3(new_n1165), .A4(new_n1191), .ZN(G407));
  INV_X1    g1017(.A(G213), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1218), .A2(G343), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(new_n1220));
  NOR3_X1   g1020(.A1(G375), .A2(G378), .A3(new_n1220), .ZN(new_n1221));
  XNOR2_X1  g1021(.A(new_n1221), .B(KEYINPUT124), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(G407), .A2(G213), .A3(new_n1222), .ZN(G409));
  NAND2_X1  g1023(.A1(new_n1067), .A2(G387), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n963), .B(new_n994), .C1(new_n1043), .C2(new_n1066), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  XNOR2_X1  g1026(.A(G393), .B(new_n794), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1226), .A2(new_n1228), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1224), .A2(new_n1227), .A3(new_n1225), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  OAI211_X1 g1031(.A(G378), .B(new_n1191), .C1(new_n1158), .C2(new_n1164), .ZN(new_n1232));
  OAI211_X1 g1032(.A(new_n947), .B(new_n1157), .C1(new_n1161), .C2(new_n1162), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(new_n1191), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(new_n1216), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1232), .A2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1211), .A2(KEYINPUT125), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n673), .B1(new_n1237), .B2(KEYINPUT60), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1238), .B1(KEYINPUT60), .B2(new_n1237), .ZN(new_n1239));
  AND2_X1   g1039(.A1(new_n1135), .A2(new_n1211), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1210), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  OR2_X1    g1041(.A1(new_n1241), .A2(new_n829), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1241), .A2(new_n829), .ZN(new_n1243));
  AND2_X1   g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1236), .A2(new_n1220), .A3(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1231), .B1(new_n1246), .B2(KEYINPUT63), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1236), .A2(new_n1220), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1219), .A2(G2897), .ZN(new_n1249));
  AND3_X1   g1049(.A1(new_n1242), .A2(new_n1243), .A3(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1249), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(KEYINPUT61), .B1(new_n1248), .B2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT63), .ZN(new_n1254));
  AOI21_X1  g1054(.A(KEYINPUT126), .B1(new_n1245), .B2(new_n1254), .ZN(new_n1255));
  AND3_X1   g1055(.A1(new_n1245), .A2(KEYINPUT126), .A3(new_n1254), .ZN(new_n1256));
  OAI211_X1 g1056(.A(new_n1247), .B(new_n1253), .C1(new_n1255), .C2(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1219), .B1(new_n1232), .B2(new_n1235), .ZN(new_n1258));
  AND3_X1   g1058(.A1(new_n1258), .A2(KEYINPUT62), .A3(new_n1244), .ZN(new_n1259));
  AOI21_X1  g1059(.A(KEYINPUT62), .B1(new_n1258), .B2(new_n1244), .ZN(new_n1260));
  OAI211_X1 g1060(.A(new_n1253), .B(KEYINPUT127), .C1(new_n1259), .C2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(new_n1231), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT62), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1245), .A2(new_n1263), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1258), .A2(KEYINPUT62), .A3(new_n1244), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  AOI21_X1  g1066(.A(KEYINPUT127), .B1(new_n1266), .B2(new_n1253), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1257), .B1(new_n1262), .B2(new_n1267), .ZN(G405));
  NAND2_X1  g1068(.A1(G375), .A2(new_n1216), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(new_n1232), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1270), .A2(new_n1244), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1244), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1269), .A2(new_n1272), .A3(new_n1232), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1271), .A2(new_n1273), .ZN(new_n1274));
  XNOR2_X1  g1074(.A(new_n1274), .B(new_n1231), .ZN(G402));
endmodule


