//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 1 1 1 1 1 1 0 0 0 1 1 1 1 0 0 0 0 1 0 0 1 1 1 1 0 0 1 1 1 0 1 1 0 0 0 0 1 0 0 1 0 0 1 0 1 0 1 1 0 0 0 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n709, new_n710, new_n711, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n747, new_n748, new_n749, new_n750, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n800,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n888, new_n889, new_n890,
    new_n892, new_n893, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n945, new_n946, new_n948, new_n949, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n963, new_n964, new_n965, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n974, new_n975, new_n976, new_n977,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n1000, new_n1001;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G197gat), .ZN(new_n203));
  XOR2_X1   g002(.A(KEYINPUT11), .B(G169gat), .Z(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XOR2_X1   g004(.A(new_n205), .B(KEYINPUT12), .Z(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G15gat), .B(G22gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(KEYINPUT92), .ZN(new_n209));
  XNOR2_X1  g008(.A(new_n209), .B(G8gat), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT16), .ZN(new_n211));
  AOI21_X1  g010(.A(G1gat), .B1(new_n208), .B2(new_n211), .ZN(new_n212));
  XOR2_X1   g011(.A(new_n210), .B(new_n212), .Z(new_n213));
  INV_X1    g012(.A(G29gat), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n214), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n215));
  AND2_X1   g014(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n216));
  NOR2_X1   g015(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n215), .B1(new_n218), .B2(G36gat), .ZN(new_n219));
  OR2_X1    g018(.A1(new_n219), .A2(KEYINPUT15), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(KEYINPUT15), .ZN(new_n221));
  XNOR2_X1  g020(.A(G43gat), .B(G50gat), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n220), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  OR2_X1    g022(.A1(new_n221), .A2(new_n222), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT17), .ZN(new_n225));
  AND3_X1   g024(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n225), .B1(new_n223), .B2(new_n224), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n213), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(G229gat), .A2(G233gat), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n210), .B(new_n212), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n223), .A2(new_n224), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n228), .A2(new_n229), .A3(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT18), .ZN(new_n234));
  AND3_X1   g033(.A1(new_n233), .A2(KEYINPUT94), .A3(new_n234), .ZN(new_n235));
  AOI21_X1  g034(.A(KEYINPUT94), .B1(new_n233), .B2(new_n234), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n207), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  AND2_X1   g036(.A1(new_n228), .A2(new_n232), .ZN(new_n238));
  NAND4_X1  g037(.A1(new_n238), .A2(KEYINPUT93), .A3(KEYINPUT18), .A4(new_n229), .ZN(new_n239));
  INV_X1    g038(.A(new_n231), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n213), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(new_n232), .ZN(new_n242));
  XOR2_X1   g041(.A(new_n229), .B(KEYINPUT13), .Z(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT93), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n245), .B1(new_n233), .B2(new_n234), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n239), .A2(new_n244), .A3(new_n246), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n237), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n250));
  NAND4_X1  g049(.A1(new_n239), .A2(new_n246), .A3(new_n250), .A4(new_n244), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(new_n206), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n249), .A2(KEYINPUT95), .A3(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT95), .ZN(new_n254));
  INV_X1    g053(.A(new_n252), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n254), .B1(new_n255), .B2(new_n248), .ZN(new_n256));
  AND2_X1   g055(.A1(new_n253), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(G141gat), .ZN(new_n258));
  INV_X1    g057(.A(G148gat), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(G141gat), .A2(G148gat), .ZN(new_n261));
  AND2_X1   g060(.A1(KEYINPUT76), .A2(KEYINPUT2), .ZN(new_n262));
  NOR2_X1   g061(.A1(KEYINPUT76), .A2(KEYINPUT2), .ZN(new_n263));
  OAI211_X1 g062(.A(new_n260), .B(new_n261), .C1(new_n262), .C2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT75), .ZN(new_n265));
  INV_X1    g064(.A(G155gat), .ZN(new_n266));
  INV_X1    g065(.A(G162gat), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n265), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  OAI21_X1  g067(.A(KEYINPUT75), .B1(G155gat), .B2(G162gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(G155gat), .A2(G162gat), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n264), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n271), .ZN(new_n273));
  NOR2_X1   g072(.A1(G155gat), .A2(G162gat), .ZN(new_n274));
  OAI21_X1  g073(.A(KEYINPUT78), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT77), .ZN(new_n276));
  AND2_X1   g075(.A1(G141gat), .A2(G148gat), .ZN(new_n277));
  NOR2_X1   g076(.A1(G141gat), .A2(G148gat), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n276), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n260), .A2(KEYINPUT77), .A3(new_n261), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n275), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT78), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n282), .B1(G155gat), .B2(G162gat), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT2), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n273), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n272), .B1(new_n281), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(KEYINPUT3), .ZN(new_n287));
  XNOR2_X1  g086(.A(G113gat), .B(G120gat), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT1), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(KEYINPUT68), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  XNOR2_X1  g090(.A(G127gat), .B(G134gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n292), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n294), .B1(new_n288), .B2(new_n290), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  XOR2_X1   g095(.A(KEYINPUT79), .B(KEYINPUT3), .Z(new_n297));
  OAI211_X1 g096(.A(new_n272), .B(new_n297), .C1(new_n281), .C2(new_n285), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n287), .A2(new_n296), .A3(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT4), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n300), .B1(new_n286), .B2(new_n296), .ZN(new_n301));
  INV_X1    g100(.A(new_n286), .ZN(new_n302));
  AND2_X1   g101(.A1(new_n293), .A2(new_n295), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n302), .A2(KEYINPUT4), .A3(new_n303), .ZN(new_n304));
  AND3_X1   g103(.A1(new_n299), .A2(new_n301), .A3(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT81), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT5), .ZN(new_n307));
  NAND2_X1  g106(.A1(G225gat), .A2(G233gat), .ZN(new_n308));
  NAND4_X1  g107(.A1(new_n305), .A2(new_n306), .A3(new_n307), .A4(new_n308), .ZN(new_n309));
  NAND4_X1  g108(.A1(new_n299), .A2(new_n304), .A3(new_n308), .A4(new_n301), .ZN(new_n310));
  OAI21_X1  g109(.A(KEYINPUT81), .B1(new_n310), .B2(KEYINPUT5), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  XNOR2_X1  g111(.A(G1gat), .B(G29gat), .ZN(new_n313));
  XNOR2_X1  g112(.A(new_n313), .B(KEYINPUT0), .ZN(new_n314));
  XNOR2_X1  g113(.A(G57gat), .B(G85gat), .ZN(new_n315));
  XOR2_X1   g114(.A(new_n314), .B(new_n315), .Z(new_n316));
  INV_X1    g115(.A(KEYINPUT80), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n302), .A2(new_n303), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n286), .A2(new_n296), .ZN(new_n319));
  AND2_X1   g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  OAI211_X1 g119(.A(new_n317), .B(KEYINPUT5), .C1(new_n320), .C2(new_n308), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n308), .B1(new_n318), .B2(new_n319), .ZN(new_n322));
  OAI21_X1  g121(.A(KEYINPUT80), .B1(new_n322), .B2(new_n307), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n321), .A2(new_n323), .A3(new_n310), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n312), .A2(new_n316), .A3(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT82), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT6), .ZN(new_n328));
  NAND4_X1  g127(.A1(new_n312), .A2(new_n324), .A3(KEYINPUT82), .A4(new_n316), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n327), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n316), .B1(new_n312), .B2(new_n324), .ZN(new_n331));
  OR2_X1    g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(KEYINPUT6), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(G227gat), .A2(G233gat), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT24), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n337), .A2(G183gat), .A3(G190gat), .ZN(new_n338));
  XNOR2_X1  g137(.A(G183gat), .B(G190gat), .ZN(new_n339));
  OAI211_X1 g138(.A(KEYINPUT66), .B(new_n338), .C1(new_n339), .C2(new_n337), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT25), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n338), .B1(new_n339), .B2(new_n337), .ZN(new_n343));
  NOR2_X1   g142(.A1(G169gat), .A2(G176gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(KEYINPUT23), .ZN(new_n345));
  NAND3_X1  g144(.A1(KEYINPUT65), .A2(G169gat), .A3(G176gat), .ZN(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  AOI21_X1  g146(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n345), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n343), .A2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT64), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n351), .B1(new_n344), .B2(KEYINPUT23), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT23), .ZN(new_n353));
  OAI211_X1 g152(.A(new_n353), .B(KEYINPUT64), .C1(G169gat), .C2(G176gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n342), .A2(new_n350), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(G169gat), .A2(G176gat), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT65), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  AOI22_X1  g158(.A1(new_n359), .A2(new_n346), .B1(KEYINPUT23), .B2(new_n344), .ZN(new_n360));
  INV_X1    g159(.A(G190gat), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n361), .A2(G183gat), .ZN(new_n362));
  INV_X1    g161(.A(G183gat), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n363), .A2(G190gat), .ZN(new_n364));
  OAI21_X1  g163(.A(KEYINPUT24), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  NAND4_X1  g164(.A1(new_n355), .A2(new_n360), .A3(new_n365), .A4(new_n338), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n366), .A2(new_n341), .A3(new_n340), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n356), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n363), .A2(KEYINPUT27), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT27), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(G183gat), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n369), .A2(new_n371), .A3(new_n361), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n372), .A2(KEYINPUT67), .A3(KEYINPUT28), .ZN(new_n373));
  NAND2_X1  g172(.A1(G183gat), .A2(G190gat), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT26), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n344), .A2(new_n375), .ZN(new_n376));
  OAI21_X1  g175(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n377));
  OAI211_X1 g176(.A(new_n376), .B(new_n377), .C1(new_n347), .C2(new_n348), .ZN(new_n378));
  AND3_X1   g177(.A1(new_n373), .A2(new_n374), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n372), .A2(KEYINPUT67), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT28), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n379), .A2(new_n382), .ZN(new_n383));
  AND3_X1   g182(.A1(new_n368), .A2(new_n303), .A3(new_n383), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n303), .B1(new_n368), .B2(new_n383), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n336), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(KEYINPUT32), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT33), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  XOR2_X1   g188(.A(G71gat), .B(G99gat), .Z(new_n390));
  XNOR2_X1  g189(.A(G15gat), .B(G43gat), .ZN(new_n391));
  XNOR2_X1  g190(.A(new_n390), .B(new_n391), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n387), .A2(new_n389), .A3(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT69), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT32), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n342), .B(new_n366), .ZN(new_n396));
  INV_X1    g195(.A(new_n383), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n296), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n368), .A2(new_n303), .A3(new_n383), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n395), .B1(new_n400), .B2(new_n336), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n392), .A2(KEYINPUT33), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n394), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  AND4_X1   g202(.A1(new_n394), .A2(new_n386), .A3(KEYINPUT32), .A4(new_n402), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n393), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT34), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT71), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n406), .B1(new_n335), .B2(new_n407), .ZN(new_n408));
  NOR3_X1   g207(.A1(new_n400), .A2(new_n336), .A3(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n408), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n384), .A2(new_n385), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n410), .B1(new_n411), .B2(new_n335), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n409), .A2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  AND2_X1   g213(.A1(new_n405), .A2(new_n414), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n405), .A2(new_n414), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT35), .ZN(new_n418));
  NAND2_X1  g217(.A1(G197gat), .A2(G204gat), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  NOR2_X1   g219(.A1(G197gat), .A2(G204gat), .ZN(new_n421));
  AND2_X1   g220(.A1(G211gat), .A2(G218gat), .ZN(new_n422));
  OAI22_X1  g221(.A1(new_n420), .A2(new_n421), .B1(new_n422), .B2(KEYINPUT22), .ZN(new_n423));
  NOR2_X1   g222(.A1(G211gat), .A2(G218gat), .ZN(new_n424));
  NOR3_X1   g223(.A1(new_n422), .A2(new_n424), .A3(KEYINPUT73), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT73), .ZN(new_n426));
  INV_X1    g225(.A(G211gat), .ZN(new_n427));
  INV_X1    g226(.A(G218gat), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(G211gat), .A2(G218gat), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n426), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n423), .B1(new_n425), .B2(new_n431), .ZN(new_n432));
  OR2_X1    g231(.A1(G197gat), .A2(G204gat), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT22), .ZN(new_n434));
  AOI22_X1  g233(.A1(new_n433), .A2(new_n419), .B1(new_n434), .B2(new_n430), .ZN(new_n435));
  OAI21_X1  g234(.A(KEYINPUT73), .B1(new_n422), .B2(new_n424), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n429), .A2(new_n426), .A3(new_n430), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n435), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n432), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT29), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n440), .B1(new_n396), .B2(new_n397), .ZN(new_n441));
  INV_X1    g240(.A(G226gat), .ZN(new_n442));
  INV_X1    g241(.A(G233gat), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n441), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  OAI211_X1 g243(.A(G226gat), .B(G233gat), .C1(new_n396), .C2(new_n397), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n439), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n444), .A2(new_n445), .A3(new_n439), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  XOR2_X1   g248(.A(G8gat), .B(G36gat), .Z(new_n450));
  XNOR2_X1  g249(.A(new_n450), .B(KEYINPUT74), .ZN(new_n451));
  XNOR2_X1  g250(.A(G64gat), .B(G92gat), .ZN(new_n452));
  XOR2_X1   g251(.A(new_n451), .B(new_n452), .Z(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n449), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n447), .A2(new_n453), .A3(new_n448), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n455), .A2(new_n456), .A3(KEYINPUT30), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT30), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n449), .A2(new_n458), .A3(new_n454), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n334), .A2(new_n417), .A3(new_n418), .A4(new_n460), .ZN(new_n461));
  XNOR2_X1  g260(.A(G78gat), .B(G106gat), .ZN(new_n462));
  XNOR2_X1  g261(.A(KEYINPUT31), .B(G50gat), .ZN(new_n463));
  XOR2_X1   g262(.A(new_n462), .B(new_n463), .Z(new_n464));
  NAND2_X1  g263(.A1(G228gat), .A2(G233gat), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n432), .A2(new_n440), .A3(new_n438), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(new_n297), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(new_n286), .ZN(new_n468));
  AOI22_X1  g267(.A1(new_n298), .A2(new_n440), .B1(new_n438), .B2(new_n432), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT84), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n298), .A2(new_n440), .ZN(new_n472));
  AND3_X1   g271(.A1(new_n472), .A2(new_n470), .A3(new_n439), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n465), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n472), .A2(new_n439), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n286), .A2(new_n440), .A3(new_n438), .A4(new_n432), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n465), .B1(new_n286), .B2(KEYINPUT3), .ZN(new_n477));
  AND3_X1   g276(.A1(new_n475), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(G22gat), .ZN(new_n480));
  AND3_X1   g279(.A1(new_n474), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n480), .B1(new_n474), .B2(new_n479), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n464), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(KEYINPUT85), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT85), .ZN(new_n485));
  OAI211_X1 g284(.A(new_n485), .B(new_n464), .C1(new_n481), .C2(new_n482), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n482), .A2(new_n464), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n475), .A2(KEYINPUT84), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n469), .A2(new_n470), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n488), .A2(new_n489), .A3(new_n468), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n478), .B1(new_n490), .B2(new_n465), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT86), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n491), .A2(new_n492), .A3(new_n480), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n474), .A2(new_n479), .ZN(new_n494));
  OAI21_X1  g293(.A(KEYINPUT86), .B1(new_n494), .B2(G22gat), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n487), .A2(new_n493), .A3(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n484), .A2(new_n486), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(KEYINPUT87), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT87), .ZN(new_n499));
  NAND4_X1  g298(.A1(new_n484), .A2(new_n499), .A3(new_n496), .A4(new_n486), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(new_n501), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n461), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g302(.A(KEYINPUT70), .B1(new_n412), .B2(new_n409), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n405), .A2(new_n505), .ZN(new_n506));
  OAI211_X1 g305(.A(new_n504), .B(new_n393), .C1(new_n403), .C2(new_n404), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(new_n464), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n510), .B1(new_n491), .B2(new_n480), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n492), .B1(new_n491), .B2(new_n480), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AOI22_X1  g312(.A1(new_n513), .A2(new_n493), .B1(KEYINPUT85), .B2(new_n483), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n499), .B1(new_n514), .B2(new_n486), .ZN(new_n515));
  INV_X1    g314(.A(new_n500), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n509), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(KEYINPUT91), .ZN(new_n518));
  AND2_X1   g317(.A1(new_n457), .A2(new_n459), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT83), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n330), .A2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(new_n331), .ZN(new_n522));
  NAND4_X1  g321(.A1(new_n327), .A2(KEYINPUT83), .A3(new_n328), .A4(new_n329), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n519), .B1(new_n524), .B2(new_n333), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT91), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n501), .A2(new_n526), .A3(new_n509), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n518), .A2(new_n525), .A3(new_n527), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n503), .B1(new_n528), .B2(KEYINPUT35), .ZN(new_n529));
  INV_X1    g328(.A(new_n529), .ZN(new_n530));
  XOR2_X1   g329(.A(KEYINPUT72), .B(KEYINPUT36), .Z(new_n531));
  OAI21_X1  g330(.A(new_n531), .B1(new_n415), .B2(new_n416), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT36), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n532), .B1(new_n533), .B2(new_n508), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n534), .B1(new_n525), .B2(new_n501), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT88), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  OAI211_X1 g336(.A(KEYINPUT88), .B(new_n534), .C1(new_n525), .C2(new_n501), .ZN(new_n538));
  INV_X1    g337(.A(new_n448), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT37), .ZN(new_n540));
  NOR3_X1   g339(.A1(new_n539), .A2(new_n446), .A3(new_n540), .ZN(new_n541));
  OAI21_X1  g340(.A(KEYINPUT90), .B1(new_n541), .B2(new_n454), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n449), .A2(new_n540), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NOR3_X1   g343(.A1(new_n541), .A2(KEYINPUT90), .A3(new_n454), .ZN(new_n545));
  OAI21_X1  g344(.A(KEYINPUT38), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n541), .A2(new_n454), .ZN(new_n547));
  AOI21_X1  g346(.A(KEYINPUT38), .B1(new_n449), .B2(new_n540), .ZN(new_n548));
  AOI22_X1  g347(.A1(new_n547), .A2(new_n548), .B1(new_n454), .B2(new_n449), .ZN(new_n549));
  NAND4_X1  g348(.A1(new_n546), .A2(new_n333), .A3(new_n332), .A4(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(new_n305), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT89), .ZN(new_n552));
  INV_X1    g351(.A(new_n308), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  OAI21_X1  g353(.A(KEYINPUT89), .B1(new_n305), .B2(new_n308), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT39), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n556), .B1(new_n320), .B2(new_n308), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n554), .A2(new_n555), .A3(new_n557), .ZN(new_n558));
  AND2_X1   g357(.A1(new_n554), .A2(new_n555), .ZN(new_n559));
  OAI211_X1 g358(.A(new_n558), .B(new_n316), .C1(new_n559), .C2(KEYINPUT39), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n560), .B(KEYINPUT40), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n519), .A2(new_n561), .A3(new_n522), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n550), .A2(new_n501), .A3(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n537), .A2(new_n538), .A3(new_n563), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n257), .B1(new_n530), .B2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT98), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT97), .ZN(new_n567));
  INV_X1    g366(.A(G57gat), .ZN(new_n568));
  AND2_X1   g367(.A1(new_n568), .A2(G64gat), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n568), .A2(G64gat), .ZN(new_n570));
  AND2_X1   g369(.A1(G71gat), .A2(G78gat), .ZN(new_n571));
  OAI22_X1  g370(.A1(new_n569), .A2(new_n570), .B1(new_n571), .B2(KEYINPUT9), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n567), .B1(new_n572), .B2(KEYINPUT96), .ZN(new_n573));
  XNOR2_X1  g372(.A(G71gat), .B(G78gat), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n572), .A2(new_n567), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n573), .A2(new_n574), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n566), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n578), .ZN(new_n580));
  NAND4_X1  g379(.A1(new_n580), .A2(KEYINPUT98), .A3(new_n576), .A4(new_n575), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n230), .B1(new_n582), .B2(KEYINPUT21), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n577), .A2(new_n578), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n584), .A2(KEYINPUT21), .ZN(new_n585));
  NAND2_X1  g384(.A1(G231gat), .A2(G233gat), .ZN(new_n586));
  XOR2_X1   g385(.A(new_n585), .B(new_n586), .Z(new_n587));
  INV_X1    g386(.A(G127gat), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n587), .A2(new_n588), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n583), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n591), .ZN(new_n593));
  INV_X1    g392(.A(new_n583), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n593), .A2(new_n594), .A3(new_n589), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(G183gat), .B(G211gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n597), .B(KEYINPUT99), .ZN(new_n598));
  XNOR2_X1  g397(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(new_n266), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n598), .B(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n596), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n592), .A2(new_n595), .A3(new_n601), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(G99gat), .A2(G106gat), .ZN(new_n606));
  INV_X1    g405(.A(G85gat), .ZN(new_n607));
  INV_X1    g406(.A(G92gat), .ZN(new_n608));
  AOI22_X1  g407(.A1(KEYINPUT8), .A2(new_n606), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(KEYINPUT100), .ZN(new_n610));
  XOR2_X1   g409(.A(G99gat), .B(G106gat), .Z(new_n611));
  INV_X1    g410(.A(KEYINPUT101), .ZN(new_n612));
  OAI21_X1  g411(.A(KEYINPUT7), .B1(new_n607), .B2(new_n608), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT7), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n614), .A2(G85gat), .A3(G92gat), .ZN(new_n615));
  AOI22_X1  g414(.A1(new_n611), .A2(new_n612), .B1(new_n613), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n610), .A2(new_n616), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n611), .A2(new_n612), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n618), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n610), .A2(new_n620), .A3(new_n616), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT102), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n619), .A2(KEYINPUT102), .A3(new_n621), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n240), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(G232gat), .A2(G233gat), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT41), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  OAI21_X1  g428(.A(KEYINPUT103), .B1(new_n626), .B2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n625), .ZN(new_n631));
  AOI21_X1  g430(.A(KEYINPUT102), .B1(new_n619), .B2(new_n621), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n231), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT103), .ZN(new_n634));
  INV_X1    g433(.A(new_n629), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n633), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n630), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n624), .A2(new_n625), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n226), .A2(new_n227), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n637), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(G190gat), .B(G218gat), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(G134gat), .B(G162gat), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n627), .A2(new_n628), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n645), .B(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n640), .B1(new_n630), .B2(new_n636), .ZN(new_n649));
  INV_X1    g448(.A(new_n643), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n644), .A2(new_n648), .A3(new_n651), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n649), .A2(new_n650), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n651), .B1(new_n653), .B2(KEYINPUT104), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT104), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n649), .A2(new_n655), .A3(new_n650), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  AOI21_X1  g456(.A(KEYINPUT105), .B1(new_n657), .B2(new_n647), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT105), .ZN(new_n659));
  AOI211_X1 g458(.A(new_n659), .B(new_n648), .C1(new_n654), .C2(new_n656), .ZN(new_n660));
  OAI211_X1 g459(.A(new_n605), .B(new_n652), .C1(new_n658), .C2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n661), .A2(KEYINPUT106), .ZN(new_n662));
  AOI211_X1 g461(.A(new_n643), .B(new_n640), .C1(new_n630), .C2(new_n636), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n663), .B1(new_n644), .B2(new_n655), .ZN(new_n664));
  INV_X1    g463(.A(new_n656), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n647), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n666), .A2(new_n659), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n657), .A2(KEYINPUT105), .A3(new_n647), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT106), .ZN(new_n670));
  NAND4_X1  g469(.A1(new_n669), .A2(new_n670), .A3(new_n605), .A4(new_n652), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n584), .A2(new_n619), .A3(new_n621), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n622), .B1(new_n578), .B2(new_n577), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT10), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n638), .A2(KEYINPUT10), .A3(new_n582), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(G230gat), .A2(G233gat), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g479(.A(G120gat), .B(G148gat), .ZN(new_n681));
  XNOR2_X1  g480(.A(G176gat), .B(G204gat), .ZN(new_n682));
  XOR2_X1   g481(.A(new_n681), .B(new_n682), .Z(new_n683));
  OAI211_X1 g482(.A(new_n680), .B(new_n683), .C1(new_n679), .C2(new_n674), .ZN(new_n684));
  INV_X1    g483(.A(new_n683), .ZN(new_n685));
  INV_X1    g484(.A(new_n679), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n686), .B1(new_n676), .B2(new_n677), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n674), .A2(new_n679), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n685), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n684), .A2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  AND3_X1   g490(.A1(new_n662), .A2(new_n671), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n565), .A2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n524), .A2(new_n333), .ZN(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n697), .B(G1gat), .ZN(G1324gat));
  INV_X1    g497(.A(KEYINPUT42), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n565), .A2(new_n519), .A3(new_n692), .ZN(new_n700));
  XOR2_X1   g499(.A(KEYINPUT16), .B(G8gat), .Z(new_n701));
  INV_X1    g500(.A(new_n701), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n699), .B1(new_n700), .B2(new_n702), .ZN(new_n703));
  OR2_X1    g502(.A1(new_n703), .A2(KEYINPUT107), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(KEYINPUT107), .ZN(new_n705));
  NAND4_X1  g504(.A1(new_n694), .A2(KEYINPUT42), .A3(new_n519), .A4(new_n701), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n700), .A2(G8gat), .ZN(new_n707));
  NAND4_X1  g506(.A1(new_n704), .A2(new_n705), .A3(new_n706), .A4(new_n707), .ZN(G1325gat));
  OAI21_X1  g507(.A(G15gat), .B1(new_n693), .B2(new_n534), .ZN(new_n709));
  INV_X1    g508(.A(new_n417), .ZN(new_n710));
  OR2_X1    g509(.A1(new_n710), .A2(G15gat), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n709), .B1(new_n693), .B2(new_n711), .ZN(G1326gat));
  NAND3_X1  g511(.A1(new_n694), .A2(KEYINPUT108), .A3(new_n502), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT108), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n714), .B1(new_n693), .B2(new_n501), .ZN(new_n715));
  XNOR2_X1  g514(.A(KEYINPUT43), .B(G22gat), .ZN(new_n716));
  AND3_X1   g515(.A1(new_n713), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n716), .B1(new_n713), .B2(new_n715), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n717), .A2(new_n718), .ZN(G1327gat));
  OAI21_X1  g518(.A(new_n652), .B1(new_n658), .B2(new_n660), .ZN(new_n720));
  AND2_X1   g519(.A1(new_n562), .A2(new_n501), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n535), .B1(new_n550), .B2(new_n721), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n720), .B1(new_n529), .B2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT44), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(new_n720), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n726), .A2(new_n724), .ZN(new_n727));
  AND3_X1   g526(.A1(new_n537), .A2(new_n538), .A3(new_n563), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n727), .B1(new_n728), .B2(new_n529), .ZN(new_n729));
  AND2_X1   g528(.A1(new_n725), .A2(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(new_n605), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(new_n691), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n249), .A2(new_n252), .ZN(new_n733));
  INV_X1    g532(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(KEYINPUT109), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n730), .A2(new_n736), .ZN(new_n737));
  OAI21_X1  g536(.A(G29gat), .B1(new_n737), .B2(new_n695), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT45), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n726), .A2(new_n732), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n565), .A2(new_n740), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n695), .A2(G29gat), .ZN(new_n742));
  INV_X1    g541(.A(new_n742), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n739), .B1(new_n741), .B2(new_n743), .ZN(new_n744));
  NAND4_X1  g543(.A1(new_n565), .A2(KEYINPUT45), .A3(new_n740), .A4(new_n742), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n738), .A2(new_n744), .A3(new_n745), .ZN(G1328gat));
  OAI21_X1  g545(.A(G36gat), .B1(new_n737), .B2(new_n460), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n460), .A2(G36gat), .ZN(new_n748));
  INV_X1    g547(.A(new_n748), .ZN(new_n749));
  OAI21_X1  g548(.A(KEYINPUT46), .B1(new_n741), .B2(new_n749), .ZN(new_n750));
  OR3_X1    g549(.A1(new_n741), .A2(KEYINPUT46), .A3(new_n749), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n747), .A2(new_n750), .A3(new_n751), .ZN(G1329gat));
  INV_X1    g551(.A(new_n534), .ZN(new_n753));
  NAND4_X1  g552(.A1(new_n730), .A2(G43gat), .A3(new_n753), .A4(new_n736), .ZN(new_n754));
  INV_X1    g553(.A(G43gat), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n755), .B1(new_n741), .B2(new_n710), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(KEYINPUT47), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT47), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n754), .A2(new_n759), .A3(new_n756), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n758), .A2(new_n760), .ZN(G1330gat));
  NAND4_X1  g560(.A1(new_n725), .A2(new_n729), .A3(new_n502), .A4(new_n736), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(G50gat), .ZN(new_n763));
  AOI21_X1  g562(.A(KEYINPUT48), .B1(new_n763), .B2(KEYINPUT111), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n501), .A2(G50gat), .ZN(new_n765));
  XOR2_X1   g564(.A(new_n765), .B(KEYINPUT110), .Z(new_n766));
  NAND3_X1  g565(.A1(new_n565), .A2(new_n740), .A3(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n763), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n764), .A2(new_n768), .ZN(new_n769));
  OAI211_X1 g568(.A(new_n763), .B(new_n767), .C1(KEYINPUT111), .C2(KEYINPUT48), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(G1331gat));
  NAND4_X1  g570(.A1(new_n662), .A2(new_n671), .A3(new_n734), .A4(new_n690), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT112), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n772), .B(new_n773), .ZN(new_n774));
  OAI211_X1 g573(.A(new_n563), .B(new_n534), .C1(new_n525), .C2(new_n501), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n526), .B1(new_n501), .B2(new_n509), .ZN(new_n776));
  AOI211_X1 g575(.A(KEYINPUT91), .B(new_n508), .C1(new_n498), .C2(new_n500), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n418), .B1(new_n778), .B2(new_n525), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n775), .B1(new_n779), .B2(new_n503), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n774), .A2(new_n780), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n781), .A2(new_n695), .ZN(new_n782));
  XNOR2_X1  g581(.A(new_n782), .B(new_n568), .ZN(G1332gat));
  INV_X1    g582(.A(KEYINPUT113), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n772), .B(KEYINPUT112), .ZN(new_n785));
  INV_X1    g584(.A(new_n780), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n784), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n774), .A2(KEYINPUT113), .A3(new_n780), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n787), .A2(new_n519), .A3(new_n788), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n789), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n790));
  XOR2_X1   g589(.A(KEYINPUT49), .B(G64gat), .Z(new_n791));
  OAI21_X1  g590(.A(new_n790), .B1(new_n789), .B2(new_n791), .ZN(G1333gat));
  INV_X1    g591(.A(G71gat), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n534), .A2(new_n793), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n787), .A2(new_n788), .A3(new_n794), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n793), .B1(new_n781), .B2(new_n710), .ZN(new_n796));
  AND3_X1   g595(.A1(new_n795), .A2(KEYINPUT50), .A3(new_n796), .ZN(new_n797));
  AOI21_X1  g596(.A(KEYINPUT50), .B1(new_n795), .B2(new_n796), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n797), .A2(new_n798), .ZN(G1334gat));
  NAND3_X1  g598(.A1(new_n787), .A2(new_n502), .A3(new_n788), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n800), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g600(.A1(new_n605), .A2(new_n733), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(new_n690), .ZN(new_n803));
  XOR2_X1   g602(.A(new_n803), .B(KEYINPUT114), .Z(new_n804));
  AND3_X1   g603(.A1(new_n730), .A2(new_n696), .A3(new_n804), .ZN(new_n805));
  OAI211_X1 g604(.A(new_n720), .B(new_n802), .C1(new_n529), .C2(new_n722), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT51), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND4_X1  g607(.A1(new_n780), .A2(KEYINPUT51), .A3(new_n720), .A4(new_n802), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(new_n810), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n696), .A2(new_n607), .A3(new_n690), .ZN(new_n812));
  OAI22_X1  g611(.A1(new_n805), .A2(new_n607), .B1(new_n811), .B2(new_n812), .ZN(G1336gat));
  NAND4_X1  g612(.A1(new_n725), .A2(new_n729), .A3(new_n519), .A4(new_n804), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(G92gat), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT52), .ZN(new_n816));
  NOR3_X1   g615(.A1(new_n460), .A2(new_n691), .A3(G92gat), .ZN(new_n817));
  INV_X1    g616(.A(new_n817), .ZN(new_n818));
  OAI211_X1 g617(.A(new_n815), .B(new_n816), .C1(new_n811), .C2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT115), .ZN(new_n820));
  AND3_X1   g619(.A1(new_n806), .A2(new_n820), .A3(KEYINPUT51), .ZN(new_n821));
  AOI21_X1  g620(.A(KEYINPUT51), .B1(new_n806), .B2(new_n820), .ZN(new_n822));
  NOR3_X1   g621(.A1(new_n821), .A2(new_n822), .A3(new_n818), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n823), .B1(G92gat), .B2(new_n814), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n819), .B1(new_n824), .B2(new_n816), .ZN(G1337gat));
  INV_X1    g624(.A(G99gat), .ZN(new_n826));
  NAND4_X1  g625(.A1(new_n725), .A2(new_n729), .A3(new_n753), .A4(new_n804), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT116), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n826), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n829), .B1(new_n828), .B2(new_n827), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n417), .A2(new_n826), .A3(new_n690), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n830), .B1(new_n811), .B2(new_n831), .ZN(G1338gat));
  NAND4_X1  g631(.A1(new_n725), .A2(new_n729), .A3(new_n502), .A4(new_n804), .ZN(new_n833));
  AND2_X1   g632(.A1(new_n833), .A2(G106gat), .ZN(new_n834));
  NOR3_X1   g633(.A1(new_n501), .A2(G106gat), .A3(new_n691), .ZN(new_n835));
  XOR2_X1   g634(.A(new_n835), .B(KEYINPUT117), .Z(new_n836));
  NOR3_X1   g635(.A1(new_n821), .A2(new_n822), .A3(new_n836), .ZN(new_n837));
  OAI21_X1  g636(.A(KEYINPUT53), .B1(new_n834), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g637(.A(KEYINPUT53), .B1(new_n810), .B2(new_n835), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n833), .A2(G106gat), .ZN(new_n840));
  AND3_X1   g639(.A1(new_n839), .A2(KEYINPUT118), .A3(new_n840), .ZN(new_n841));
  AOI21_X1  g640(.A(KEYINPUT118), .B1(new_n839), .B2(new_n840), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n838), .B1(new_n841), .B2(new_n842), .ZN(G1339gat));
  NAND3_X1  g642(.A1(new_n676), .A2(new_n677), .A3(new_n686), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n680), .A2(new_n844), .A3(KEYINPUT54), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT54), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n683), .B1(new_n687), .B2(new_n846), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n845), .A2(KEYINPUT55), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(new_n684), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n845), .A2(new_n847), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT55), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT119), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n850), .A2(KEYINPUT119), .A3(new_n851), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n849), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(new_n243), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n241), .A2(new_n232), .A3(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(KEYINPUT120), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT120), .ZN(new_n860));
  NAND4_X1  g659(.A1(new_n241), .A2(new_n232), .A3(new_n860), .A4(new_n857), .ZN(new_n861));
  OAI211_X1 g660(.A(new_n859), .B(new_n861), .C1(new_n238), .C2(new_n229), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n862), .A2(KEYINPUT121), .A3(new_n205), .ZN(new_n863));
  INV_X1    g662(.A(new_n863), .ZN(new_n864));
  AOI21_X1  g663(.A(KEYINPUT121), .B1(new_n862), .B2(new_n205), .ZN(new_n865));
  OAI22_X1  g664(.A1(new_n864), .A2(new_n865), .B1(new_n237), .B2(new_n247), .ZN(new_n866));
  INV_X1    g665(.A(new_n866), .ZN(new_n867));
  AOI22_X1  g666(.A1(new_n856), .A2(new_n733), .B1(new_n690), .B2(new_n867), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n868), .A2(new_n720), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n854), .A2(new_n855), .ZN(new_n870));
  INV_X1    g669(.A(new_n849), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n870), .A2(new_n867), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n872), .B1(new_n669), .B2(new_n652), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n731), .B1(new_n869), .B2(new_n873), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n662), .A2(new_n671), .A3(new_n734), .A4(new_n691), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(new_n778), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n877), .A2(new_n695), .ZN(new_n878));
  AND3_X1   g677(.A1(new_n876), .A2(new_n460), .A3(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(G113gat), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n879), .A2(new_n880), .A3(new_n733), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n502), .B1(new_n874), .B2(new_n875), .ZN(new_n882));
  NOR3_X1   g681(.A1(new_n695), .A2(new_n519), .A3(new_n710), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  OAI21_X1  g683(.A(G113gat), .B1(new_n884), .B2(new_n257), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n881), .A2(new_n885), .ZN(new_n886));
  XNOR2_X1  g685(.A(new_n886), .B(KEYINPUT122), .ZN(G1340gat));
  AOI21_X1  g686(.A(G120gat), .B1(new_n879), .B2(new_n690), .ZN(new_n888));
  INV_X1    g687(.A(G120gat), .ZN(new_n889));
  NOR3_X1   g688(.A1(new_n884), .A2(new_n889), .A3(new_n691), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n888), .A2(new_n890), .ZN(G1341gat));
  NAND3_X1  g690(.A1(new_n879), .A2(new_n588), .A3(new_n605), .ZN(new_n892));
  OAI21_X1  g691(.A(G127gat), .B1(new_n884), .B2(new_n731), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(G1342gat));
  NAND2_X1  g693(.A1(new_n720), .A2(new_n460), .ZN(new_n895));
  XNOR2_X1  g694(.A(new_n895), .B(KEYINPUT123), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n896), .A2(G134gat), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n897), .A2(new_n876), .A3(new_n878), .ZN(new_n898));
  XOR2_X1   g697(.A(new_n898), .B(KEYINPUT56), .Z(new_n899));
  OAI21_X1  g698(.A(G134gat), .B1(new_n884), .B2(new_n726), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(new_n900), .ZN(G1343gat));
  INV_X1    g700(.A(new_n875), .ZN(new_n902));
  OAI21_X1  g701(.A(KEYINPUT124), .B1(new_n866), .B2(new_n691), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n862), .A2(new_n205), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT121), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(new_n863), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT124), .ZN(new_n908));
  NAND4_X1  g707(.A1(new_n907), .A2(new_n249), .A3(new_n908), .A4(new_n690), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n903), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n852), .A2(new_n684), .A3(new_n848), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n911), .B1(new_n253), .B2(new_n256), .ZN(new_n912));
  OAI211_X1 g711(.A(new_n669), .B(new_n652), .C1(new_n910), .C2(new_n912), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n720), .A2(new_n867), .A3(new_n856), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n605), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n502), .B1(new_n902), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(KEYINPUT57), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n501), .B1(new_n874), .B2(new_n875), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT57), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n696), .A2(new_n534), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n921), .A2(new_n519), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n917), .A2(new_n920), .A3(new_n922), .ZN(new_n923));
  OAI21_X1  g722(.A(G141gat), .B1(new_n923), .B2(new_n257), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n918), .A2(new_n922), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n257), .A2(G141gat), .ZN(new_n926));
  AOI21_X1  g725(.A(KEYINPUT58), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n924), .A2(new_n927), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT58), .ZN(new_n929));
  NAND4_X1  g728(.A1(new_n917), .A2(new_n920), .A3(new_n733), .A4(new_n922), .ZN(new_n930));
  AOI22_X1  g729(.A1(new_n930), .A2(G141gat), .B1(new_n925), .B2(new_n926), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n928), .B1(new_n929), .B2(new_n931), .ZN(G1344gat));
  NAND3_X1  g731(.A1(new_n925), .A2(new_n259), .A3(new_n690), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT59), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n934), .A2(G148gat), .ZN(new_n935));
  AND3_X1   g734(.A1(new_n917), .A2(new_n920), .A3(new_n922), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n935), .B1(new_n936), .B2(new_n690), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n876), .A2(new_n502), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n938), .A2(KEYINPUT57), .ZN(new_n939));
  AND4_X1   g738(.A1(new_n257), .A2(new_n662), .A3(new_n671), .A4(new_n691), .ZN(new_n940));
  OAI211_X1 g739(.A(new_n919), .B(new_n502), .C1(new_n940), .C2(new_n915), .ZN(new_n941));
  NAND4_X1  g740(.A1(new_n939), .A2(new_n690), .A3(new_n922), .A4(new_n941), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n934), .B1(new_n942), .B2(G148gat), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n933), .B1(new_n937), .B2(new_n943), .ZN(G1345gat));
  OAI21_X1  g743(.A(G155gat), .B1(new_n923), .B2(new_n731), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n925), .A2(new_n266), .A3(new_n605), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(new_n946), .ZN(G1346gat));
  OAI21_X1  g746(.A(G162gat), .B1(new_n923), .B2(new_n726), .ZN(new_n948));
  OR3_X1    g747(.A1(new_n896), .A2(G162gat), .A3(new_n921), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n948), .B1(new_n938), .B2(new_n949), .ZN(G1347gat));
  NAND2_X1  g749(.A1(new_n695), .A2(new_n519), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n951), .A2(new_n710), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n882), .A2(new_n952), .ZN(new_n953));
  INV_X1    g752(.A(G169gat), .ZN(new_n954));
  NOR3_X1   g753(.A1(new_n953), .A2(new_n954), .A3(new_n257), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT125), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n956), .B1(new_n876), .B2(new_n695), .ZN(new_n957));
  AOI211_X1 g756(.A(KEYINPUT125), .B(new_n696), .C1(new_n874), .C2(new_n875), .ZN(new_n958));
  OR2_X1    g757(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NOR2_X1   g758(.A1(new_n877), .A2(new_n460), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n959), .A2(new_n733), .A3(new_n960), .ZN(new_n961));
  AOI21_X1  g760(.A(new_n955), .B1(new_n961), .B2(new_n954), .ZN(G1348gat));
  OAI21_X1  g761(.A(G176gat), .B1(new_n953), .B2(new_n691), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n959), .A2(new_n960), .ZN(new_n964));
  OR2_X1    g763(.A1(new_n691), .A2(G176gat), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n963), .B1(new_n964), .B2(new_n965), .ZN(G1349gat));
  AND3_X1   g765(.A1(new_n605), .A2(new_n369), .A3(new_n371), .ZN(new_n967));
  OAI211_X1 g766(.A(new_n960), .B(new_n967), .C1(new_n957), .C2(new_n958), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT126), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n882), .A2(new_n605), .A3(new_n952), .ZN(new_n970));
  AOI21_X1  g769(.A(new_n969), .B1(new_n970), .B2(G183gat), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n968), .A2(new_n971), .ZN(new_n972));
  XNOR2_X1  g771(.A(new_n972), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g772(.A(G190gat), .B1(new_n953), .B2(new_n726), .ZN(new_n974));
  AND2_X1   g773(.A1(new_n974), .A2(KEYINPUT61), .ZN(new_n975));
  NOR2_X1   g774(.A1(new_n974), .A2(KEYINPUT61), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n720), .A2(new_n361), .ZN(new_n977));
  OAI22_X1  g776(.A1(new_n975), .A2(new_n976), .B1(new_n964), .B2(new_n977), .ZN(G1351gat));
  NOR2_X1   g777(.A1(new_n951), .A2(new_n753), .ZN(new_n979));
  OAI211_X1 g778(.A(new_n941), .B(new_n979), .C1(new_n919), .C2(new_n918), .ZN(new_n980));
  INV_X1    g779(.A(G197gat), .ZN(new_n981));
  NOR3_X1   g780(.A1(new_n980), .A2(new_n981), .A3(new_n257), .ZN(new_n982));
  NOR3_X1   g781(.A1(new_n753), .A2(new_n460), .A3(new_n501), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n959), .A2(new_n733), .A3(new_n983), .ZN(new_n984));
  AOI21_X1  g783(.A(new_n982), .B1(new_n984), .B2(new_n981), .ZN(G1352gat));
  NOR2_X1   g784(.A1(new_n691), .A2(G204gat), .ZN(new_n986));
  OAI211_X1 g785(.A(new_n983), .B(new_n986), .C1(new_n957), .C2(new_n958), .ZN(new_n987));
  OR2_X1    g786(.A1(new_n987), .A2(KEYINPUT62), .ZN(new_n988));
  OAI21_X1  g787(.A(G204gat), .B1(new_n980), .B2(new_n691), .ZN(new_n989));
  AND3_X1   g788(.A1(new_n987), .A2(KEYINPUT127), .A3(KEYINPUT62), .ZN(new_n990));
  AOI21_X1  g789(.A(KEYINPUT127), .B1(new_n987), .B2(KEYINPUT62), .ZN(new_n991));
  OAI211_X1 g790(.A(new_n988), .B(new_n989), .C1(new_n990), .C2(new_n991), .ZN(G1353gat));
  OAI211_X1 g791(.A(KEYINPUT63), .B(G211gat), .C1(new_n980), .C2(new_n731), .ZN(new_n993));
  INV_X1    g792(.A(new_n993), .ZN(new_n994));
  NAND4_X1  g793(.A1(new_n939), .A2(new_n605), .A3(new_n941), .A4(new_n979), .ZN(new_n995));
  AOI21_X1  g794(.A(KEYINPUT63), .B1(new_n995), .B2(G211gat), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n959), .A2(new_n983), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n605), .A2(new_n427), .ZN(new_n998));
  OAI22_X1  g797(.A1(new_n994), .A2(new_n996), .B1(new_n997), .B2(new_n998), .ZN(G1354gat));
  OAI21_X1  g798(.A(G218gat), .B1(new_n980), .B2(new_n726), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n720), .A2(new_n428), .ZN(new_n1001));
  OAI21_X1  g800(.A(new_n1000), .B1(new_n997), .B2(new_n1001), .ZN(G1355gat));
endmodule


