//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 1 0 1 0 1 0 1 0 1 0 1 0 1 0 0 1 1 1 1 0 0 0 0 1 1 1 0 1 0 0 1 1 1 1 0 0 1 1 1 1 1 1 0 0 1 1 1 1 0 1 1 1 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n710, new_n711, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n790, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n799, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n847, new_n848, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n894, new_n895, new_n897, new_n898,
    new_n900, new_n901, new_n902, new_n903, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n976, new_n977, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1030, new_n1031, new_n1032;
  XNOR2_X1  g000(.A(G8gat), .B(G36gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT77), .ZN(new_n203));
  XNOR2_X1  g002(.A(G64gat), .B(G92gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n205), .B(KEYINPUT78), .ZN(new_n206));
  NAND2_X1  g005(.A1(G226gat), .A2(G233gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT29), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT66), .ZN(new_n210));
  NOR2_X1   g009(.A1(G169gat), .A2(G176gat), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT65), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT23), .ZN(new_n213));
  AOI22_X1  g012(.A1(new_n212), .A2(new_n213), .B1(G169gat), .B2(G176gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(KEYINPUT65), .A2(KEYINPUT23), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n211), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n213), .A2(G176gat), .ZN(new_n217));
  INV_X1    g016(.A(G169gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(KEYINPUT64), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT64), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(G169gat), .ZN(new_n221));
  AND3_X1   g020(.A1(new_n217), .A2(new_n219), .A3(new_n221), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n210), .B1(new_n216), .B2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(G176gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n218), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(G169gat), .A2(G176gat), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n226), .B1(KEYINPUT65), .B2(KEYINPUT23), .ZN(new_n227));
  INV_X1    g026(.A(new_n215), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n225), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(KEYINPUT64), .B(G169gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(new_n217), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n229), .A2(new_n231), .A3(KEYINPUT66), .ZN(new_n232));
  NAND2_X1  g031(.A1(G183gat), .A2(G190gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(KEYINPUT24), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT24), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n235), .A2(G183gat), .A3(G190gat), .ZN(new_n236));
  INV_X1    g035(.A(G183gat), .ZN(new_n237));
  INV_X1    g036(.A(G190gat), .ZN(new_n238));
  AOI22_X1  g037(.A1(new_n234), .A2(new_n236), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(new_n239), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n223), .A2(new_n232), .A3(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT25), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n234), .A2(new_n236), .ZN(new_n244));
  OR2_X1    g043(.A1(KEYINPUT67), .A2(G183gat), .ZN(new_n245));
  NAND2_X1  g044(.A1(KEYINPUT67), .A2(G183gat), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n244), .B1(new_n247), .B2(G190gat), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n242), .B1(new_n217), .B2(new_n218), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n248), .A2(new_n229), .A3(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n243), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT69), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n237), .A2(KEYINPUT27), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT27), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(G183gat), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n253), .A2(new_n255), .A3(new_n238), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(KEYINPUT28), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT26), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n225), .A2(new_n258), .A3(new_n226), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n211), .A2(KEYINPUT26), .ZN(new_n260));
  NAND4_X1  g059(.A1(new_n257), .A2(new_n233), .A3(new_n259), .A4(new_n260), .ZN(new_n261));
  OR2_X1    g060(.A1(KEYINPUT68), .A2(KEYINPUT27), .ZN(new_n262));
  NAND2_X1  g061(.A1(KEYINPUT68), .A2(KEYINPUT27), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n262), .A2(G183gat), .A3(new_n263), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n245), .A2(KEYINPUT27), .A3(new_n246), .ZN(new_n265));
  NOR2_X1   g064(.A1(KEYINPUT28), .A2(G190gat), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n264), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n252), .B1(new_n261), .B2(new_n268), .ZN(new_n269));
  AND3_X1   g068(.A1(new_n259), .A2(new_n233), .A3(new_n260), .ZN(new_n270));
  NAND4_X1  g069(.A1(new_n270), .A2(new_n267), .A3(KEYINPUT69), .A4(new_n257), .ZN(new_n271));
  AND2_X1   g070(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n209), .B1(new_n251), .B2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(new_n250), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n274), .B1(new_n241), .B2(new_n242), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n261), .A2(new_n268), .ZN(new_n276));
  NOR3_X1   g075(.A1(new_n275), .A2(new_n207), .A3(new_n276), .ZN(new_n277));
  AND2_X1   g076(.A1(G211gat), .A2(G218gat), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n278), .A2(KEYINPUT22), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(G197gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(KEYINPUT74), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT74), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(G197gat), .ZN(new_n284));
  AND3_X1   g083(.A1(new_n282), .A2(new_n284), .A3(G204gat), .ZN(new_n285));
  AOI21_X1  g084(.A(G204gat), .B1(new_n282), .B2(new_n284), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n280), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NOR2_X1   g086(.A1(G211gat), .A2(G218gat), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n278), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(G204gat), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n283), .A2(G197gat), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n281), .A2(KEYINPUT74), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n291), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n282), .A2(new_n284), .A3(G204gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n289), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n296), .A2(new_n297), .A3(new_n280), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n290), .A2(new_n298), .ZN(new_n299));
  NOR3_X1   g098(.A1(new_n273), .A2(new_n277), .A3(new_n299), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n208), .B1(new_n275), .B2(new_n276), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT75), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n301), .A2(new_n302), .A3(new_n207), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n251), .A2(new_n272), .ZN(new_n304));
  INV_X1    g103(.A(new_n207), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n303), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(new_n299), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n302), .B1(new_n301), .B2(new_n207), .ZN(new_n309));
  NOR3_X1   g108(.A1(new_n307), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n300), .B1(new_n310), .B2(KEYINPUT76), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n301), .A2(new_n207), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(KEYINPUT75), .ZN(new_n313));
  NAND4_X1  g112(.A1(new_n313), .A2(new_n299), .A3(new_n306), .A4(new_n303), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT76), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n206), .B1(new_n311), .B2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(new_n300), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n207), .B1(new_n251), .B2(new_n272), .ZN(new_n319));
  INV_X1    g118(.A(new_n276), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n229), .A2(new_n231), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n239), .B1(new_n321), .B2(new_n210), .ZN(new_n322));
  AOI21_X1  g121(.A(KEYINPUT25), .B1(new_n322), .B2(new_n232), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n320), .B1(new_n323), .B2(new_n274), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n305), .B1(new_n324), .B2(new_n208), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n319), .B1(new_n325), .B2(new_n302), .ZN(new_n326));
  NAND4_X1  g125(.A1(new_n326), .A2(KEYINPUT76), .A3(new_n299), .A4(new_n313), .ZN(new_n327));
  AND4_X1   g126(.A1(new_n316), .A2(new_n318), .A3(new_n327), .A4(new_n205), .ZN(new_n328));
  OAI21_X1  g127(.A(KEYINPUT30), .B1(new_n317), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT4), .ZN(new_n330));
  NAND2_X1  g129(.A1(G155gat), .A2(G162gat), .ZN(new_n331));
  INV_X1    g130(.A(G155gat), .ZN(new_n332));
  INV_X1    g131(.A(G162gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(G141gat), .ZN(new_n335));
  INV_X1    g134(.A(G148gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(G141gat), .A2(G148gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  OAI211_X1 g138(.A(new_n331), .B(new_n334), .C1(new_n339), .C2(KEYINPUT2), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT79), .ZN(new_n341));
  INV_X1    g140(.A(new_n338), .ZN(new_n342));
  NOR2_X1   g141(.A1(G141gat), .A2(G148gat), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n341), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n337), .A2(KEYINPUT79), .A3(new_n338), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n334), .A2(new_n331), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n344), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT80), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n331), .A2(new_n348), .A3(KEYINPUT2), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n348), .B1(new_n331), .B2(KEYINPUT2), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n340), .B1(new_n347), .B2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT1), .ZN(new_n354));
  INV_X1    g153(.A(G120gat), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(G113gat), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n355), .A2(G113gat), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n354), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(G134gat), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(G127gat), .ZN(new_n361));
  INV_X1    g160(.A(G127gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(G134gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n359), .A2(new_n364), .ZN(new_n365));
  AND3_X1   g164(.A1(new_n361), .A2(new_n363), .A3(new_n354), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT70), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n367), .B1(new_n355), .B2(G113gat), .ZN(new_n368));
  INV_X1    g167(.A(G113gat), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n369), .A2(KEYINPUT70), .A3(G120gat), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n368), .A2(new_n356), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n366), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n365), .A2(new_n372), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n330), .B1(new_n353), .B2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(new_n351), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(new_n349), .ZN(new_n376));
  NAND4_X1  g175(.A1(new_n376), .A2(new_n346), .A3(new_n345), .A4(new_n344), .ZN(new_n377));
  AOI22_X1  g176(.A1(new_n359), .A2(new_n364), .B1(new_n366), .B2(new_n371), .ZN(new_n378));
  NAND4_X1  g177(.A1(new_n377), .A2(new_n378), .A3(KEYINPUT4), .A4(new_n340), .ZN(new_n379));
  XNOR2_X1  g178(.A(KEYINPUT81), .B(KEYINPUT3), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n373), .B1(new_n353), .B2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT3), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n383), .B1(new_n377), .B2(new_n340), .ZN(new_n384));
  OAI211_X1 g183(.A(new_n374), .B(new_n379), .C1(new_n382), .C2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(G225gat), .A2(G233gat), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT5), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n353), .A2(new_n373), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n377), .A2(new_n378), .A3(new_n340), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n386), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  OAI22_X1  g190(.A1(new_n385), .A2(new_n387), .B1(new_n388), .B2(new_n391), .ZN(new_n392));
  XNOR2_X1  g191(.A(G1gat), .B(G29gat), .ZN(new_n393));
  XNOR2_X1  g192(.A(new_n393), .B(KEYINPUT0), .ZN(new_n394));
  XNOR2_X1  g193(.A(G57gat), .B(G85gat), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n394), .B(new_n395), .ZN(new_n396));
  AND2_X1   g195(.A1(new_n374), .A2(new_n379), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n353), .A2(KEYINPUT3), .ZN(new_n398));
  OAI211_X1 g197(.A(new_n398), .B(new_n373), .C1(new_n353), .C2(new_n381), .ZN(new_n399));
  NAND4_X1  g198(.A1(new_n397), .A2(KEYINPUT5), .A3(new_n386), .A4(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n392), .A2(new_n396), .A3(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT6), .ZN(new_n402));
  OAI21_X1  g201(.A(KEYINPUT82), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  AND2_X1   g202(.A1(new_n392), .A2(new_n400), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT82), .ZN(new_n405));
  NAND4_X1  g204(.A1(new_n404), .A2(new_n405), .A3(KEYINPUT6), .A4(new_n396), .ZN(new_n406));
  AND2_X1   g205(.A1(new_n401), .A2(new_n402), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n392), .A2(new_n400), .ZN(new_n408));
  INV_X1    g207(.A(new_n396), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  AOI22_X1  g209(.A1(new_n403), .A2(new_n406), .B1(new_n407), .B2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  NAND4_X1  g211(.A1(new_n316), .A2(new_n318), .A3(new_n327), .A4(new_n205), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT30), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n329), .A2(new_n412), .A3(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(G22gat), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n208), .B1(new_n353), .B2(new_n381), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n308), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(KEYINPUT29), .B1(new_n290), .B2(new_n298), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(new_n353), .ZN(new_n422));
  INV_X1    g221(.A(G228gat), .ZN(new_n423));
  INV_X1    g222(.A(G233gat), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n420), .A2(new_n422), .A3(new_n425), .A4(new_n398), .ZN(new_n426));
  INV_X1    g225(.A(new_n420), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n297), .B1(new_n296), .B2(new_n280), .ZN(new_n428));
  AOI211_X1 g227(.A(new_n289), .B(new_n279), .C1(new_n294), .C2(new_n295), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n208), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(KEYINPUT84), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT84), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n299), .A2(new_n432), .A3(new_n208), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n431), .A2(new_n380), .A3(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n427), .B1(new_n434), .B2(new_n353), .ZN(new_n435));
  OAI211_X1 g234(.A(new_n418), .B(new_n426), .C1(new_n435), .C2(new_n425), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT85), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(new_n353), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n381), .B1(new_n430), .B2(KEYINPUT84), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n439), .B1(new_n440), .B2(new_n433), .ZN(new_n441));
  OAI22_X1  g240(.A1(new_n441), .A2(new_n427), .B1(new_n423), .B2(new_n424), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n442), .A2(KEYINPUT85), .A3(new_n418), .A4(new_n426), .ZN(new_n443));
  XNOR2_X1  g242(.A(G78gat), .B(G106gat), .ZN(new_n444));
  XNOR2_X1  g243(.A(KEYINPUT31), .B(G50gat), .ZN(new_n445));
  XNOR2_X1  g244(.A(new_n444), .B(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(new_n433), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n380), .B1(new_n421), .B2(new_n432), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n353), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n425), .B1(new_n449), .B2(new_n420), .ZN(new_n450));
  INV_X1    g249(.A(new_n426), .ZN(new_n451));
  OAI21_X1  g250(.A(G22gat), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n438), .A2(new_n443), .A3(new_n446), .A4(new_n452), .ZN(new_n453));
  XNOR2_X1  g252(.A(new_n446), .B(KEYINPUT83), .ZN(new_n454));
  INV_X1    g253(.A(new_n436), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n418), .B1(new_n442), .B2(new_n426), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n454), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  AND2_X1   g256(.A1(new_n453), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n251), .A2(new_n272), .A3(new_n373), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n269), .A2(new_n271), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n378), .B1(new_n275), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(G227gat), .A2(G233gat), .ZN(new_n462));
  INV_X1    g261(.A(new_n462), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n459), .A2(new_n461), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(KEYINPUT32), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT33), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  XOR2_X1   g266(.A(G15gat), .B(G43gat), .Z(new_n468));
  XNOR2_X1  g267(.A(G71gat), .B(G99gat), .ZN(new_n469));
  XNOR2_X1  g268(.A(new_n468), .B(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n465), .A2(new_n467), .A3(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(new_n470), .ZN(new_n472));
  OAI211_X1 g271(.A(new_n464), .B(KEYINPUT32), .C1(new_n466), .C2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n373), .B1(new_n251), .B2(new_n272), .ZN(new_n475));
  NOR3_X1   g274(.A1(new_n275), .A2(new_n460), .A3(new_n378), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n462), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(KEYINPUT72), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT34), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n479), .B1(new_n462), .B2(KEYINPUT71), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n463), .B1(new_n459), .B2(new_n461), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT72), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n478), .A2(new_n480), .A3(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(new_n480), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n481), .A2(new_n482), .ZN(new_n486));
  AOI211_X1 g285(.A(KEYINPUT72), .B(new_n463), .C1(new_n459), .C2(new_n461), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n485), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n474), .A2(KEYINPUT73), .A3(new_n484), .A4(new_n488), .ZN(new_n489));
  NOR3_X1   g288(.A1(new_n486), .A2(new_n487), .A3(new_n485), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n480), .B1(new_n478), .B2(new_n483), .ZN(new_n491));
  OAI211_X1 g290(.A(new_n471), .B(new_n473), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT73), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n474), .A2(new_n484), .A3(new_n488), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n492), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  AOI211_X1 g294(.A(KEYINPUT35), .B(new_n458), .C1(new_n489), .C2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n453), .A2(new_n457), .ZN(new_n497));
  AND3_X1   g296(.A1(new_n497), .A2(new_n494), .A3(new_n492), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n498), .A2(new_n412), .A3(new_n329), .A4(new_n415), .ZN(new_n499));
  AOI22_X1  g298(.A1(new_n417), .A2(new_n496), .B1(new_n499), .B2(KEYINPUT35), .ZN(new_n500));
  AND2_X1   g299(.A1(new_n413), .A2(new_n414), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n316), .A2(new_n318), .A3(new_n327), .ZN(new_n502));
  INV_X1    g301(.A(new_n206), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(new_n413), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n501), .B1(new_n505), .B2(KEYINPUT30), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n506), .A2(new_n458), .A3(new_n412), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n329), .A2(new_n415), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n385), .A2(new_n387), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n389), .A2(new_n390), .A3(new_n386), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(KEYINPUT39), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(KEYINPUT86), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(new_n509), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n511), .A2(KEYINPUT86), .ZN(new_n514));
  OAI221_X1 g313(.A(new_n409), .B1(KEYINPUT39), .B2(new_n509), .C1(new_n513), .C2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT40), .ZN(new_n516));
  OR2_X1    g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n515), .A2(new_n516), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n517), .A2(new_n401), .A3(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n502), .A2(KEYINPUT37), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT37), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n311), .A2(new_n522), .A3(new_n316), .ZN(new_n523));
  INV_X1    g322(.A(new_n205), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n521), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(KEYINPUT38), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n411), .A2(new_n413), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n206), .A2(KEYINPUT38), .ZN(new_n528));
  INV_X1    g327(.A(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT87), .ZN(new_n530));
  OAI211_X1 g329(.A(new_n530), .B(new_n308), .C1(new_n307), .C2(new_n309), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(KEYINPUT37), .ZN(new_n532));
  INV_X1    g331(.A(new_n532), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n299), .B1(new_n273), .B2(new_n277), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n534), .A2(KEYINPUT87), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n313), .A2(new_n306), .A3(new_n303), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n535), .B1(new_n536), .B2(new_n308), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n529), .B1(new_n533), .B2(new_n538), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n527), .B1(new_n539), .B2(new_n523), .ZN(new_n540));
  AOI22_X1  g339(.A1(new_n508), .A2(new_n520), .B1(new_n526), .B2(new_n540), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n507), .B1(new_n541), .B2(new_n458), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT36), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n495), .A2(new_n543), .A3(new_n489), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n492), .A2(KEYINPUT36), .A3(new_n494), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n500), .B1(new_n542), .B2(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(G15gat), .B(G22gat), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT16), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n548), .B1(new_n549), .B2(G1gat), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n550), .B1(G1gat), .B2(new_n548), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(G8gat), .ZN(new_n552));
  INV_X1    g351(.A(G8gat), .ZN(new_n553));
  OAI211_X1 g352(.A(new_n550), .B(new_n553), .C1(G1gat), .C2(new_n548), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  XOR2_X1   g355(.A(G43gat), .B(G50gat), .Z(new_n557));
  INV_X1    g356(.A(KEYINPUT15), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(G43gat), .B(G50gat), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n560), .A2(KEYINPUT15), .ZN(new_n561));
  INV_X1    g360(.A(G29gat), .ZN(new_n562));
  INV_X1    g361(.A(G36gat), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NOR2_X1   g363(.A1(G29gat), .A2(G36gat), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n564), .B1(KEYINPUT14), .B2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT14), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n567), .B1(G29gat), .B2(G36gat), .ZN(new_n568));
  NAND4_X1  g367(.A1(new_n559), .A2(new_n561), .A3(new_n566), .A4(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n565), .A2(KEYINPUT14), .ZN(new_n570));
  OAI211_X1 g369(.A(new_n570), .B(new_n568), .C1(new_n562), .C2(new_n563), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n571), .A2(KEYINPUT15), .A3(new_n560), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n569), .A2(KEYINPUT17), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n569), .A2(new_n572), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT17), .ZN(new_n575));
  AOI21_X1  g374(.A(KEYINPUT89), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT89), .ZN(new_n577));
  AOI211_X1 g376(.A(new_n577), .B(KEYINPUT17), .C1(new_n569), .C2(new_n572), .ZN(new_n578));
  OAI211_X1 g377(.A(new_n556), .B(new_n573), .C1(new_n576), .C2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n555), .A2(new_n574), .ZN(new_n580));
  NAND2_X1  g379(.A1(G229gat), .A2(G233gat), .ZN(new_n581));
  NAND4_X1  g380(.A1(new_n579), .A2(KEYINPUT18), .A3(new_n580), .A4(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n555), .B(new_n574), .ZN(new_n583));
  XOR2_X1   g382(.A(new_n581), .B(KEYINPUT13), .Z(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  AND2_X1   g384(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n587));
  XNOR2_X1  g386(.A(KEYINPUT90), .B(KEYINPUT18), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(G113gat), .B(G141gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(KEYINPUT88), .B(KEYINPUT11), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n591), .B(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(G169gat), .B(G197gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n593), .B(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(KEYINPUT12), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n590), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n596), .B1(new_n587), .B2(new_n588), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n586), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT91), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  AOI21_X1  g400(.A(KEYINPUT91), .B1(new_n586), .B2(new_n598), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n597), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n547), .A2(new_n604), .ZN(new_n605));
  XOR2_X1   g404(.A(G57gat), .B(G64gat), .Z(new_n606));
  INV_X1    g405(.A(KEYINPUT9), .ZN(new_n607));
  INV_X1    g406(.A(G71gat), .ZN(new_n608));
  INV_X1    g407(.A(G78gat), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n607), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n606), .A2(new_n610), .ZN(new_n611));
  XOR2_X1   g410(.A(G71gat), .B(G78gat), .Z(new_n612));
  OR2_X1    g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n611), .A2(new_n612), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT21), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(G231gat), .A2(G233gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n617), .B(new_n618), .ZN(new_n619));
  XOR2_X1   g418(.A(G127gat), .B(G155gat), .Z(new_n620));
  XNOR2_X1  g419(.A(new_n620), .B(KEYINPUT20), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n619), .B(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(G183gat), .B(G211gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n622), .B(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n615), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n555), .B1(new_n625), .B2(KEYINPUT21), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(KEYINPUT93), .ZN(new_n627));
  XNOR2_X1  g426(.A(KEYINPUT92), .B(KEYINPUT19), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n627), .B(new_n628), .ZN(new_n629));
  OR2_X1    g428(.A1(new_n624), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n624), .A2(new_n629), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(G85gat), .ZN(new_n634));
  INV_X1    g433(.A(G92gat), .ZN(new_n635));
  OAI21_X1  g434(.A(KEYINPUT94), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT94), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n637), .A2(G85gat), .A3(G92gat), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n636), .A2(new_n638), .A3(KEYINPUT7), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT7), .ZN(new_n640));
  OAI211_X1 g439(.A(KEYINPUT94), .B(new_n640), .C1(new_n634), .C2(new_n635), .ZN(new_n641));
  NAND2_X1  g440(.A1(G99gat), .A2(G106gat), .ZN(new_n642));
  AOI22_X1  g441(.A1(KEYINPUT8), .A2(new_n642), .B1(new_n634), .B2(new_n635), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n639), .A2(new_n641), .A3(new_n643), .ZN(new_n644));
  XOR2_X1   g443(.A(G99gat), .B(G106gat), .Z(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n645), .ZN(new_n647));
  NAND4_X1  g446(.A1(new_n647), .A2(new_n639), .A3(new_n641), .A4(new_n643), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  OAI211_X1 g448(.A(new_n573), .B(new_n649), .C1(new_n576), .C2(new_n578), .ZN(new_n650));
  INV_X1    g449(.A(new_n649), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n651), .A2(new_n574), .ZN(new_n652));
  NAND3_X1  g451(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n653));
  AND3_X1   g452(.A1(new_n652), .A2(KEYINPUT95), .A3(new_n653), .ZN(new_n654));
  AOI21_X1  g453(.A(KEYINPUT95), .B1(new_n652), .B2(new_n653), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n650), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  XOR2_X1   g455(.A(G190gat), .B(G218gat), .Z(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g457(.A(G134gat), .B(G162gat), .ZN(new_n659));
  AOI21_X1  g458(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n659), .B(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n657), .ZN(new_n662));
  OAI211_X1 g461(.A(new_n662), .B(new_n650), .C1(new_n654), .C2(new_n655), .ZN(new_n663));
  AND3_X1   g462(.A1(new_n658), .A2(new_n661), .A3(new_n663), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n661), .B1(new_n658), .B2(new_n663), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n615), .A2(new_n649), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT10), .ZN(new_n668));
  NAND4_X1  g467(.A1(new_n613), .A2(new_n646), .A3(new_n614), .A4(new_n648), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n667), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n625), .A2(new_n651), .A3(KEYINPUT10), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(G230gat), .A2(G233gat), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n673), .B1(new_n667), .B2(new_n669), .ZN(new_n675));
  XNOR2_X1  g474(.A(G120gat), .B(G148gat), .ZN(new_n676));
  XNOR2_X1  g475(.A(G176gat), .B(G204gat), .ZN(new_n677));
  XOR2_X1   g476(.A(new_n676), .B(new_n677), .Z(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n675), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n674), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n673), .B(KEYINPUT96), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n682), .B1(new_n670), .B2(new_n671), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n679), .B1(new_n683), .B2(new_n675), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  NOR3_X1   g484(.A1(new_n633), .A2(new_n666), .A3(new_n685), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n605), .A2(new_n411), .A3(new_n686), .ZN(new_n687));
  XNOR2_X1  g486(.A(KEYINPUT97), .B(G1gat), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n687), .B(new_n688), .ZN(G1324gat));
  NAND3_X1  g488(.A1(new_n605), .A2(new_n508), .A3(new_n686), .ZN(new_n690));
  AND2_X1   g489(.A1(new_n690), .A2(G8gat), .ZN(new_n691));
  XNOR2_X1  g490(.A(KEYINPUT16), .B(G8gat), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  OAI21_X1  g492(.A(KEYINPUT42), .B1(new_n691), .B2(new_n693), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n694), .B1(KEYINPUT42), .B2(new_n693), .ZN(G1325gat));
  NAND2_X1  g494(.A1(new_n605), .A2(new_n686), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n546), .A2(KEYINPUT98), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT98), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n544), .A2(new_n698), .A3(new_n545), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT99), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n697), .A2(new_n699), .A3(KEYINPUT99), .ZN(new_n703));
  AND2_X1   g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  OAI21_X1  g503(.A(G15gat), .B1(new_n696), .B2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(G15gat), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n495), .A2(new_n489), .ZN(new_n707));
  NAND4_X1  g506(.A1(new_n605), .A2(new_n706), .A3(new_n707), .A4(new_n686), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n705), .A2(new_n708), .ZN(G1326gat));
  NOR2_X1   g508(.A1(new_n696), .A2(new_n497), .ZN(new_n710));
  XOR2_X1   g509(.A(KEYINPUT43), .B(G22gat), .Z(new_n711));
  XNOR2_X1  g510(.A(new_n710), .B(new_n711), .ZN(G1327gat));
  INV_X1    g511(.A(new_n685), .ZN(new_n713));
  NAND4_X1  g512(.A1(new_n605), .A2(new_n633), .A3(new_n666), .A4(new_n713), .ZN(new_n714));
  NOR3_X1   g513(.A1(new_n714), .A2(G29gat), .A3(new_n412), .ZN(new_n715));
  XOR2_X1   g514(.A(new_n715), .B(KEYINPUT45), .Z(new_n716));
  INV_X1    g515(.A(new_n666), .ZN(new_n717));
  OAI21_X1  g516(.A(KEYINPUT44), .B1(new_n547), .B2(new_n717), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n717), .A2(KEYINPUT44), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n497), .A2(new_n494), .A3(new_n492), .ZN(new_n720));
  OAI21_X1  g519(.A(KEYINPUT35), .B1(new_n416), .B2(new_n720), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n458), .B1(new_n495), .B2(new_n489), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT35), .ZN(new_n723));
  NAND4_X1  g522(.A1(new_n722), .A2(new_n506), .A3(new_n723), .A4(new_n412), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n721), .A2(new_n724), .A3(KEYINPUT101), .ZN(new_n725));
  AND4_X1   g524(.A1(new_n458), .A2(new_n329), .A3(new_n412), .A4(new_n415), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT38), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n205), .B1(new_n502), .B2(KEYINPUT37), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n727), .B1(new_n728), .B2(new_n523), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n502), .A2(KEYINPUT37), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n528), .B1(new_n532), .B2(new_n537), .ZN(new_n731));
  OAI211_X1 g530(.A(new_n411), .B(new_n413), .C1(new_n730), .C2(new_n731), .ZN(new_n732));
  OAI22_X1  g531(.A1(new_n506), .A2(new_n519), .B1(new_n729), .B2(new_n732), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n726), .B1(new_n733), .B2(new_n497), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n725), .B1(new_n734), .B2(new_n700), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n500), .A2(KEYINPUT101), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n719), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n718), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n685), .B(KEYINPUT100), .ZN(new_n739));
  NOR3_X1   g538(.A1(new_n632), .A2(new_n604), .A3(new_n739), .ZN(new_n740));
  AND2_X1   g539(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  AND2_X1   g540(.A1(new_n741), .A2(new_n411), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n716), .B1(new_n562), .B2(new_n742), .ZN(G1328gat));
  NAND2_X1  g542(.A1(new_n741), .A2(new_n508), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT102), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n563), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n746), .B1(new_n745), .B2(new_n744), .ZN(new_n747));
  NOR3_X1   g546(.A1(new_n714), .A2(G36gat), .A3(new_n506), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(KEYINPUT46), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n747), .A2(new_n749), .ZN(G1329gat));
  INV_X1    g549(.A(G43gat), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n738), .A2(new_n700), .A3(new_n740), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT103), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n751), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n754), .B1(new_n753), .B2(new_n752), .ZN(new_n755));
  INV_X1    g554(.A(new_n707), .ZN(new_n756));
  NOR3_X1   g555(.A1(new_n714), .A2(G43gat), .A3(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT47), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n755), .A2(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(new_n704), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n751), .B1(new_n741), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n758), .B1(new_n762), .B2(new_n757), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n760), .A2(new_n763), .ZN(G1330gat));
  INV_X1    g563(.A(G50gat), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n765), .B1(new_n741), .B2(new_n458), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT48), .ZN(new_n767));
  NOR3_X1   g566(.A1(new_n714), .A2(G50gat), .A3(new_n497), .ZN(new_n768));
  OR3_X1    g567(.A1(new_n766), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n767), .B1(new_n766), .B2(new_n768), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(G1331gat));
  NAND3_X1  g570(.A1(new_n632), .A2(new_n604), .A3(new_n717), .ZN(new_n772));
  INV_X1    g571(.A(new_n739), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n774), .B(KEYINPUT104), .ZN(new_n775));
  INV_X1    g574(.A(new_n699), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n698), .B1(new_n544), .B2(new_n545), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  AOI22_X1  g577(.A1(new_n542), .A2(new_n778), .B1(new_n500), .B2(KEYINPUT101), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n721), .A2(new_n724), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT101), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n775), .B1(new_n779), .B2(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(new_n411), .ZN(new_n784));
  XOR2_X1   g583(.A(KEYINPUT105), .B(G57gat), .Z(new_n785));
  XNOR2_X1  g584(.A(new_n784), .B(new_n785), .ZN(G1332gat));
  AOI21_X1  g585(.A(new_n506), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n787), .B(KEYINPUT106), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n783), .A2(new_n788), .ZN(new_n789));
  NOR2_X1   g588(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n790));
  XOR2_X1   g589(.A(new_n789), .B(new_n790), .Z(G1333gat));
  AOI21_X1  g590(.A(KEYINPUT107), .B1(new_n783), .B2(new_n707), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n792), .A2(G71gat), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n783), .A2(KEYINPUT107), .A3(new_n707), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n704), .A2(new_n608), .ZN(new_n795));
  AOI22_X1  g594(.A1(new_n793), .A2(new_n794), .B1(new_n783), .B2(new_n795), .ZN(new_n796));
  XOR2_X1   g595(.A(KEYINPUT108), .B(KEYINPUT50), .Z(new_n797));
  XNOR2_X1  g596(.A(new_n796), .B(new_n797), .ZN(G1334gat));
  NAND2_X1  g597(.A1(new_n783), .A2(new_n458), .ZN(new_n799));
  XNOR2_X1  g598(.A(new_n799), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g599(.A1(new_n633), .A2(new_n604), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n801), .A2(new_n713), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n738), .A2(new_n802), .ZN(new_n803));
  OAI21_X1  g602(.A(G85gat), .B1(new_n803), .B2(new_n412), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT51), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n801), .A2(new_n805), .ZN(new_n806));
  OAI211_X1 g605(.A(new_n666), .B(new_n806), .C1(new_n735), .C2(new_n736), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(KEYINPUT109), .ZN(new_n808));
  OAI211_X1 g607(.A(new_n782), .B(new_n725), .C1(new_n734), .C2(new_n700), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT109), .ZN(new_n810));
  NAND4_X1  g609(.A1(new_n809), .A2(new_n810), .A3(new_n666), .A4(new_n806), .ZN(new_n811));
  INV_X1    g610(.A(new_n801), .ZN(new_n812));
  OAI211_X1 g611(.A(new_n666), .B(new_n812), .C1(new_n735), .C2(new_n736), .ZN(new_n813));
  AOI22_X1  g612(.A1(new_n808), .A2(new_n811), .B1(new_n805), .B2(new_n813), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n411), .A2(new_n634), .A3(new_n685), .ZN(new_n815));
  XNOR2_X1  g614(.A(new_n815), .B(KEYINPUT110), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n804), .B1(new_n814), .B2(new_n816), .ZN(G1336gat));
  INV_X1    g616(.A(new_n802), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n818), .B1(new_n718), .B2(new_n737), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n635), .B1(new_n819), .B2(new_n508), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n508), .A2(new_n635), .A3(new_n739), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n813), .A2(new_n805), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n821), .B1(new_n822), .B2(new_n807), .ZN(new_n823));
  OAI21_X1  g622(.A(KEYINPUT52), .B1(new_n820), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(KEYINPUT111), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT111), .ZN(new_n826));
  OAI211_X1 g625(.A(new_n826), .B(KEYINPUT52), .C1(new_n820), .C2(new_n823), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT112), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT52), .ZN(new_n830));
  AOI211_X1 g629(.A(new_n506), .B(new_n818), .C1(new_n718), .C2(new_n737), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n830), .B1(new_n831), .B2(new_n635), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n808), .A2(new_n811), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n821), .B1(new_n833), .B2(new_n822), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n829), .B1(new_n832), .B2(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(new_n719), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n836), .B1(new_n779), .B2(new_n782), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT44), .ZN(new_n838));
  INV_X1    g637(.A(new_n546), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n780), .B1(new_n734), .B2(new_n839), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n838), .B1(new_n840), .B2(new_n666), .ZN(new_n841));
  OAI211_X1 g640(.A(new_n508), .B(new_n802), .C1(new_n837), .C2(new_n841), .ZN(new_n842));
  AOI21_X1  g641(.A(KEYINPUT52), .B1(new_n842), .B2(G92gat), .ZN(new_n843));
  OAI211_X1 g642(.A(new_n843), .B(KEYINPUT112), .C1(new_n814), .C2(new_n821), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n835), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n828), .A2(new_n845), .ZN(G1337gat));
  OAI21_X1  g645(.A(G99gat), .B1(new_n803), .B2(new_n704), .ZN(new_n847));
  OR3_X1    g646(.A1(new_n756), .A2(G99gat), .A3(new_n713), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n847), .B1(new_n814), .B2(new_n848), .ZN(G1338gat));
  OAI21_X1  g648(.A(G106gat), .B1(new_n803), .B2(new_n497), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT113), .ZN(new_n851));
  OR3_X1    g650(.A1(new_n773), .A2(new_n497), .A3(G106gat), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n852), .B1(new_n822), .B2(new_n807), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n850), .B1(new_n851), .B2(new_n853), .ZN(new_n854));
  AND2_X1   g653(.A1(new_n853), .A2(new_n851), .ZN(new_n855));
  OAI21_X1  g654(.A(KEYINPUT53), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT53), .ZN(new_n857));
  OAI211_X1 g656(.A(new_n850), .B(new_n857), .C1(new_n814), .C2(new_n852), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n856), .A2(new_n858), .ZN(G1339gat));
  NOR2_X1   g658(.A1(new_n772), .A2(new_n685), .ZN(new_n860));
  INV_X1    g659(.A(new_n682), .ZN(new_n861));
  OAI211_X1 g660(.A(new_n674), .B(KEYINPUT54), .C1(new_n672), .C2(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT55), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT54), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n678), .B1(new_n683), .B2(new_n864), .ZN(new_n865));
  AND3_X1   g664(.A1(new_n862), .A2(new_n863), .A3(new_n865), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n863), .B1(new_n862), .B2(new_n865), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n681), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(new_n666), .ZN(new_n870));
  XNOR2_X1  g669(.A(new_n599), .B(new_n600), .ZN(new_n871));
  INV_X1    g670(.A(new_n595), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n581), .B1(new_n579), .B2(new_n580), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n583), .A2(new_n584), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n872), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  XNOR2_X1  g674(.A(new_n875), .B(KEYINPUT114), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n871), .A2(new_n876), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n870), .A2(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(new_n878), .ZN(new_n879));
  OAI211_X1 g678(.A(new_n876), .B(new_n685), .C1(new_n601), .C2(new_n602), .ZN(new_n880));
  INV_X1    g679(.A(new_n880), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n881), .B1(new_n603), .B2(new_n869), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n879), .B1(new_n882), .B2(new_n666), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n860), .B1(new_n883), .B2(new_n633), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n884), .A2(new_n720), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n508), .A2(new_n412), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(new_n887), .ZN(new_n888));
  AOI21_X1  g687(.A(G113gat), .B1(new_n888), .B2(new_n603), .ZN(new_n889));
  NOR3_X1   g688(.A1(new_n884), .A2(new_n458), .A3(new_n756), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(new_n886), .ZN(new_n891));
  NOR3_X1   g690(.A1(new_n891), .A2(new_n369), .A3(new_n604), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n889), .A2(new_n892), .ZN(G1340gat));
  AOI21_X1  g692(.A(G120gat), .B1(new_n888), .B2(new_n685), .ZN(new_n894));
  NOR3_X1   g693(.A1(new_n891), .A2(new_n355), .A3(new_n773), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n894), .A2(new_n895), .ZN(G1341gat));
  NAND3_X1  g695(.A1(new_n888), .A2(new_n362), .A3(new_n632), .ZN(new_n897));
  OAI21_X1  g696(.A(G127gat), .B1(new_n891), .B2(new_n633), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(G1342gat));
  NOR2_X1   g698(.A1(new_n508), .A2(new_n717), .ZN(new_n900));
  NAND4_X1  g699(.A1(new_n885), .A2(new_n360), .A3(new_n411), .A4(new_n900), .ZN(new_n901));
  XOR2_X1   g700(.A(new_n901), .B(KEYINPUT56), .Z(new_n902));
  OAI21_X1  g701(.A(G134gat), .B1(new_n891), .B2(new_n717), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(new_n903), .ZN(G1343gat));
  OR2_X1    g703(.A1(new_n884), .A2(new_n497), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT57), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n905), .A2(KEYINPUT115), .A3(new_n906), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT115), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n884), .A2(new_n497), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n908), .B1(new_n909), .B2(KEYINPUT57), .ZN(new_n910));
  INV_X1    g709(.A(new_n860), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n868), .A2(KEYINPUT117), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT117), .ZN(new_n913));
  OAI211_X1 g712(.A(new_n913), .B(new_n681), .C1(new_n866), .C2(new_n867), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n912), .A2(new_n603), .A3(new_n914), .ZN(new_n915));
  NAND4_X1  g714(.A1(new_n871), .A2(KEYINPUT116), .A3(new_n685), .A4(new_n876), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT116), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n880), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n915), .A2(new_n916), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n878), .B1(new_n919), .B2(new_n717), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n911), .B1(new_n920), .B2(new_n632), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n497), .A2(new_n906), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n907), .A2(new_n910), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n778), .A2(new_n886), .ZN(new_n925));
  INV_X1    g724(.A(new_n925), .ZN(new_n926));
  AND2_X1   g725(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n335), .B1(new_n927), .B2(new_n603), .ZN(new_n928));
  NOR3_X1   g727(.A1(new_n761), .A2(new_n412), .A3(new_n905), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n929), .A2(new_n506), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n603), .A2(new_n335), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  OAI21_X1  g731(.A(KEYINPUT58), .B1(new_n928), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n924), .A2(new_n926), .ZN(new_n934));
  OAI21_X1  g733(.A(G141gat), .B1(new_n934), .B2(new_n604), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT58), .ZN(new_n936));
  OAI211_X1 g735(.A(new_n935), .B(new_n936), .C1(new_n930), .C2(new_n931), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n933), .A2(new_n937), .ZN(G1344gat));
  INV_X1    g737(.A(new_n930), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n939), .A2(new_n336), .A3(new_n685), .ZN(new_n940));
  AOI211_X1 g739(.A(KEYINPUT59), .B(new_n336), .C1(new_n927), .C2(new_n685), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT59), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT118), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n633), .B1(new_n920), .B2(new_n943), .ZN(new_n944));
  AOI211_X1 g743(.A(KEYINPUT118), .B(new_n878), .C1(new_n919), .C2(new_n717), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n911), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n497), .A2(KEYINPUT57), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g747(.A(KEYINPUT57), .B1(new_n884), .B2(new_n497), .ZN(new_n949));
  AND2_X1   g748(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n950), .A2(new_n685), .A3(new_n926), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n942), .B1(new_n951), .B2(G148gat), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n940), .B1(new_n941), .B2(new_n952), .ZN(G1345gat));
  NAND3_X1  g752(.A1(new_n939), .A2(new_n332), .A3(new_n632), .ZN(new_n954));
  OAI21_X1  g753(.A(G155gat), .B1(new_n934), .B2(new_n633), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(new_n955), .ZN(G1346gat));
  OAI21_X1  g755(.A(G162gat), .B1(new_n934), .B2(new_n717), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n929), .A2(new_n333), .A3(new_n900), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n959), .A2(KEYINPUT119), .ZN(new_n960));
  INV_X1    g759(.A(KEYINPUT119), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n957), .A2(new_n961), .A3(new_n958), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n960), .A2(new_n962), .ZN(G1347gat));
  NOR2_X1   g762(.A1(new_n506), .A2(new_n411), .ZN(new_n964));
  AND2_X1   g763(.A1(new_n885), .A2(new_n964), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n965), .A2(new_n230), .A3(new_n603), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n890), .A2(new_n964), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n967), .A2(KEYINPUT120), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT120), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n890), .A2(new_n969), .A3(new_n964), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n968), .A2(new_n603), .A3(new_n970), .ZN(new_n971));
  INV_X1    g770(.A(KEYINPUT121), .ZN(new_n972));
  AND3_X1   g771(.A1(new_n971), .A2(new_n972), .A3(G169gat), .ZN(new_n973));
  AOI21_X1  g772(.A(new_n972), .B1(new_n971), .B2(G169gat), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n966), .B1(new_n973), .B2(new_n974), .ZN(G1348gat));
  NAND3_X1  g774(.A1(new_n965), .A2(new_n224), .A3(new_n685), .ZN(new_n976));
  AND3_X1   g775(.A1(new_n968), .A2(new_n739), .A3(new_n970), .ZN(new_n977));
  OAI21_X1  g776(.A(new_n976), .B1(new_n977), .B2(new_n224), .ZN(G1349gat));
  INV_X1    g777(.A(KEYINPUT123), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n968), .A2(new_n632), .A3(new_n970), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n980), .A2(new_n247), .ZN(new_n981));
  AND3_X1   g780(.A1(new_n632), .A2(new_n253), .A3(new_n255), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n965), .A2(new_n982), .ZN(new_n983));
  AND2_X1   g782(.A1(KEYINPUT122), .A2(KEYINPUT60), .ZN(new_n984));
  AND4_X1   g783(.A1(new_n979), .A2(new_n981), .A3(new_n983), .A4(new_n984), .ZN(new_n985));
  AOI22_X1  g784(.A1(new_n980), .A2(new_n247), .B1(new_n965), .B2(new_n982), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n986), .A2(new_n979), .ZN(new_n987));
  OAI21_X1  g786(.A(KEYINPUT60), .B1(new_n986), .B2(KEYINPUT122), .ZN(new_n988));
  AOI21_X1  g787(.A(new_n985), .B1(new_n987), .B2(new_n988), .ZN(G1350gat));
  NAND3_X1  g788(.A1(new_n965), .A2(new_n238), .A3(new_n666), .ZN(new_n990));
  NAND3_X1  g789(.A1(new_n968), .A2(new_n666), .A3(new_n970), .ZN(new_n991));
  INV_X1    g790(.A(KEYINPUT61), .ZN(new_n992));
  AND3_X1   g791(.A1(new_n991), .A2(new_n992), .A3(G190gat), .ZN(new_n993));
  AOI21_X1  g792(.A(new_n992), .B1(new_n991), .B2(G190gat), .ZN(new_n994));
  OAI21_X1  g793(.A(new_n990), .B1(new_n993), .B2(new_n994), .ZN(G1351gat));
  AND3_X1   g794(.A1(new_n702), .A2(new_n703), .A3(new_n964), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n996), .A2(new_n909), .ZN(new_n997));
  INV_X1    g796(.A(new_n997), .ZN(new_n998));
  AOI21_X1  g797(.A(G197gat), .B1(new_n998), .B2(new_n603), .ZN(new_n999));
  AND2_X1   g798(.A1(new_n950), .A2(new_n996), .ZN(new_n1000));
  NOR2_X1   g799(.A1(new_n604), .A2(new_n281), .ZN(new_n1001));
  AOI21_X1  g800(.A(new_n999), .B1(new_n1000), .B2(new_n1001), .ZN(G1352gat));
  XNOR2_X1  g801(.A(KEYINPUT124), .B(G204gat), .ZN(new_n1003));
  INV_X1    g802(.A(KEYINPUT125), .ZN(new_n1004));
  INV_X1    g803(.A(KEYINPUT62), .ZN(new_n1005));
  OAI21_X1  g804(.A(new_n1003), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  NOR3_X1   g805(.A1(new_n997), .A2(new_n713), .A3(new_n1006), .ZN(new_n1007));
  NAND2_X1  g806(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1008));
  XNOR2_X1  g807(.A(new_n1007), .B(new_n1008), .ZN(new_n1009));
  AND2_X1   g808(.A1(new_n1000), .A2(new_n739), .ZN(new_n1010));
  OAI21_X1  g809(.A(new_n1009), .B1(new_n1010), .B2(new_n1003), .ZN(G1353gat));
  NAND4_X1  g810(.A1(new_n948), .A2(new_n632), .A3(new_n949), .A4(new_n996), .ZN(new_n1012));
  INV_X1    g811(.A(KEYINPUT126), .ZN(new_n1013));
  INV_X1    g812(.A(KEYINPUT63), .ZN(new_n1014));
  NAND2_X1  g813(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  AND3_X1   g814(.A1(new_n1012), .A2(G211gat), .A3(new_n1015), .ZN(new_n1016));
  AOI21_X1  g815(.A(new_n1015), .B1(new_n1012), .B2(G211gat), .ZN(new_n1017));
  NOR2_X1   g816(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1018));
  NOR3_X1   g817(.A1(new_n1016), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1019));
  NOR3_X1   g818(.A1(new_n997), .A2(G211gat), .A3(new_n633), .ZN(new_n1020));
  OAI21_X1  g819(.A(KEYINPUT127), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g820(.A(new_n1017), .ZN(new_n1022));
  NAND3_X1  g821(.A1(new_n1012), .A2(G211gat), .A3(new_n1015), .ZN(new_n1023));
  INV_X1    g822(.A(new_n1018), .ZN(new_n1024));
  NAND3_X1  g823(.A1(new_n1022), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1025));
  INV_X1    g824(.A(KEYINPUT127), .ZN(new_n1026));
  INV_X1    g825(.A(new_n1020), .ZN(new_n1027));
  NAND3_X1  g826(.A1(new_n1025), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  NAND2_X1  g827(.A1(new_n1021), .A2(new_n1028), .ZN(G1354gat));
  NAND2_X1  g828(.A1(new_n1000), .A2(new_n666), .ZN(new_n1030));
  NAND2_X1  g829(.A1(new_n1030), .A2(G218gat), .ZN(new_n1031));
  OR2_X1    g830(.A1(new_n717), .A2(G218gat), .ZN(new_n1032));
  OAI21_X1  g831(.A(new_n1031), .B1(new_n997), .B2(new_n1032), .ZN(G1355gat));
endmodule


