//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 0 0 0 1 0 1 0 1 1 1 1 0 0 1 0 1 1 0 1 1 1 0 0 0 0 1 1 0 1 1 0 0 1 1 0 1 0 0 0 1 0 0 1 0 0 0 1 0 1 0 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:15 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1326, new_n1327, new_n1328;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  XNOR2_X1  g0003(.A(new_n203), .B(KEYINPUT64), .ZN(new_n204));
  INV_X1    g0004(.A(G77), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n204), .A2(new_n205), .ZN(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  INV_X1    g0008(.A(G226), .ZN(new_n209));
  INV_X1    g0009(.A(G68), .ZN(new_n210));
  INV_X1    g0010(.A(G238), .ZN(new_n211));
  OAI22_X1  g0011(.A1(new_n202), .A2(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT67), .ZN(new_n214));
  AOI211_X1 g0014(.A(new_n212), .B(new_n214), .C1(G77), .C2(G244), .ZN(new_n215));
  INV_X1    g0015(.A(G87), .ZN(new_n216));
  INV_X1    g0016(.A(G250), .ZN(new_n217));
  INV_X1    g0017(.A(G116), .ZN(new_n218));
  INV_X1    g0018(.A(G270), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(G97), .ZN(new_n221));
  INV_X1    g0021(.A(G257), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n208), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT1), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n208), .A2(G13), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n226), .B(G250), .C1(G257), .C2(G264), .ZN(new_n227));
  XOR2_X1   g0027(.A(KEYINPUT65), .B(KEYINPUT0), .Z(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  INV_X1    g0029(.A(new_n201), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n230), .A2(G50), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(new_n232));
  NAND2_X1  g0032(.A1(G1), .A2(G13), .ZN(new_n233));
  INV_X1    g0033(.A(G20), .ZN(new_n234));
  NOR2_X1   g0034(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g0035(.A1(new_n232), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g0036(.A1(new_n229), .A2(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT66), .ZN(new_n238));
  NOR2_X1   g0038(.A1(new_n225), .A2(new_n238), .ZN(G361));
  XNOR2_X1  g0039(.A(KEYINPUT2), .B(G226), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G232), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G238), .B(G244), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n241), .B(new_n242), .Z(new_n243));
  XNOR2_X1  g0043(.A(G250), .B(G257), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(G264), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(new_n219), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n243), .B(new_n246), .Z(G358));
  XNOR2_X1  g0047(.A(G68), .B(G77), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(new_n202), .ZN(new_n249));
  INV_X1    g0049(.A(G58), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G107), .B(G116), .ZN(new_n252));
  XNOR2_X1  g0052(.A(G87), .B(G97), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n251), .B(new_n254), .ZN(G351));
  INV_X1    g0055(.A(KEYINPUT3), .ZN(new_n256));
  INV_X1    g0056(.A(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(KEYINPUT3), .A2(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G1698), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G222), .ZN(new_n262));
  INV_X1    g0062(.A(G223), .ZN(new_n263));
  OAI211_X1 g0063(.A(new_n260), .B(new_n262), .C1(new_n263), .C2(new_n261), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n264), .B1(G77), .B2(new_n260), .ZN(new_n265));
  XNOR2_X1  g0065(.A(new_n265), .B(KEYINPUT69), .ZN(new_n266));
  NAND2_X1  g0066(.A1(G33), .A2(G41), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n267), .A2(G1), .A3(G13), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G1), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n270), .B1(G41), .B2(G45), .ZN(new_n271));
  INV_X1    g0071(.A(G274), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  AND2_X1   g0074(.A1(G33), .A2(G41), .ZN(new_n275));
  NOR2_X1   g0075(.A1(G41), .A2(G45), .ZN(new_n276));
  OAI22_X1  g0076(.A1(new_n275), .A2(new_n233), .B1(new_n276), .B2(G1), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(KEYINPUT68), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT68), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n268), .A2(new_n279), .A3(new_n271), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n274), .B1(new_n282), .B2(new_n209), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n269), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G179), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  XNOR2_X1  g0086(.A(KEYINPUT8), .B(G58), .ZN(new_n287));
  XNOR2_X1  g0087(.A(new_n287), .B(KEYINPUT71), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n257), .A2(G20), .ZN(new_n289));
  NOR2_X1   g0089(.A1(G20), .A2(G33), .ZN(new_n290));
  AOI22_X1  g0090(.A1(new_n288), .A2(new_n289), .B1(G150), .B2(new_n290), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n291), .B1(new_n234), .B2(new_n204), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n233), .B1(new_n208), .B2(new_n257), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(KEYINPUT70), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT70), .ZN(new_n295));
  OAI211_X1 g0095(.A(new_n295), .B(new_n233), .C1(new_n208), .C2(new_n257), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G13), .ZN(new_n298));
  NOR3_X1   g0098(.A1(new_n298), .A2(new_n234), .A3(G1), .ZN(new_n299));
  AOI22_X1  g0099(.A1(new_n292), .A2(new_n297), .B1(new_n202), .B2(new_n299), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n297), .B1(new_n270), .B2(G20), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(G50), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G169), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n304), .B1(new_n269), .B2(new_n283), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n286), .A2(new_n303), .A3(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n284), .A2(G190), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n300), .A2(KEYINPUT9), .A3(new_n302), .ZN(new_n309));
  AND2_X1   g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT10), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT9), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n303), .A2(new_n312), .ZN(new_n313));
  OAI21_X1  g0113(.A(G200), .B1(new_n269), .B2(new_n283), .ZN(new_n314));
  NAND4_X1  g0114(.A1(new_n310), .A2(new_n311), .A3(new_n313), .A4(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n308), .A2(new_n314), .A3(new_n309), .ZN(new_n316));
  INV_X1    g0116(.A(new_n313), .ZN(new_n317));
  OAI21_X1  g0117(.A(KEYINPUT10), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n307), .B1(new_n315), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n261), .A2(G232), .ZN(new_n320));
  OAI211_X1 g0120(.A(new_n260), .B(new_n320), .C1(new_n211), .C2(new_n261), .ZN(new_n321));
  INV_X1    g0121(.A(new_n268), .ZN(new_n322));
  OAI211_X1 g0122(.A(new_n321), .B(new_n322), .C1(G107), .C2(new_n260), .ZN(new_n323));
  INV_X1    g0123(.A(G244), .ZN(new_n324));
  OAI211_X1 g0124(.A(new_n323), .B(new_n274), .C1(new_n282), .C2(new_n324), .ZN(new_n325));
  OR2_X1    g0125(.A1(new_n325), .A2(G179), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n299), .A2(new_n205), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n301), .A2(G77), .ZN(new_n328));
  NAND2_X1  g0128(.A1(G20), .A2(G77), .ZN(new_n329));
  INV_X1    g0129(.A(new_n290), .ZN(new_n330));
  INV_X1    g0130(.A(new_n289), .ZN(new_n331));
  XNOR2_X1  g0131(.A(KEYINPUT15), .B(G87), .ZN(new_n332));
  OAI221_X1 g0132(.A(new_n329), .B1(new_n287), .B2(new_n330), .C1(new_n331), .C2(new_n332), .ZN(new_n333));
  AND3_X1   g0133(.A1(new_n333), .A2(KEYINPUT72), .A3(new_n297), .ZN(new_n334));
  AOI21_X1  g0134(.A(KEYINPUT72), .B1(new_n333), .B2(new_n297), .ZN(new_n335));
  OAI211_X1 g0135(.A(new_n327), .B(new_n328), .C1(new_n334), .C2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n325), .A2(new_n304), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n326), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n336), .ZN(new_n339));
  INV_X1    g0139(.A(G190), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n339), .B1(new_n340), .B2(new_n325), .ZN(new_n341));
  AND2_X1   g0141(.A1(new_n325), .A2(G200), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n319), .A2(new_n338), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(KEYINPUT73), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT73), .ZN(new_n347));
  NAND4_X1  g0147(.A1(new_n319), .A2(new_n347), .A3(new_n338), .A4(new_n344), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT16), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n258), .A2(new_n234), .A3(new_n259), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT7), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND4_X1  g0153(.A1(new_n258), .A2(KEYINPUT7), .A3(new_n234), .A4(new_n259), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n210), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n250), .A2(new_n210), .ZN(new_n356));
  OAI21_X1  g0156(.A(G20), .B1(new_n356), .B2(new_n201), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n290), .A2(G159), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n350), .B1(new_n355), .B2(new_n359), .ZN(new_n360));
  AND2_X1   g0160(.A1(KEYINPUT3), .A2(G33), .ZN(new_n361));
  NOR2_X1   g0161(.A1(KEYINPUT3), .A2(G33), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(KEYINPUT7), .B1(new_n363), .B2(new_n234), .ZN(new_n364));
  INV_X1    g0164(.A(new_n354), .ZN(new_n365));
  OAI21_X1  g0165(.A(G68), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n359), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n366), .A2(KEYINPUT16), .A3(new_n367), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n360), .A2(new_n368), .A3(new_n297), .ZN(new_n369));
  INV_X1    g0169(.A(new_n299), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n288), .A2(new_n370), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n371), .B1(new_n301), .B2(new_n288), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n369), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n263), .A2(new_n261), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n209), .A2(G1698), .ZN(new_n375));
  OAI211_X1 g0175(.A(new_n374), .B(new_n375), .C1(new_n361), .C2(new_n362), .ZN(new_n376));
  NAND2_X1  g0176(.A1(G33), .A2(G87), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n273), .B1(new_n378), .B2(new_n322), .ZN(new_n379));
  AND3_X1   g0179(.A1(new_n268), .A2(G232), .A3(new_n271), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(KEYINPUT75), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n268), .B1(new_n376), .B2(new_n377), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT75), .ZN(new_n384));
  NOR4_X1   g0184(.A1(new_n383), .A2(new_n384), .A3(new_n380), .A4(new_n273), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n304), .B1(new_n382), .B2(new_n385), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n379), .A2(new_n285), .A3(new_n381), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n373), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT18), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n373), .A2(KEYINPUT18), .A3(new_n386), .A4(new_n387), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT17), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n378), .A2(new_n322), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n395), .A2(new_n381), .A3(new_n274), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n396), .A2(G190), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n384), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n379), .A2(KEYINPUT75), .A3(new_n381), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(G200), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n397), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n394), .B1(new_n402), .B2(new_n373), .ZN(new_n403));
  AND2_X1   g0203(.A1(new_n369), .A2(new_n372), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n401), .B1(new_n382), .B2(new_n385), .ZN(new_n405));
  INV_X1    g0205(.A(new_n397), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n404), .A2(new_n407), .A3(KEYINPUT17), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n403), .A2(new_n408), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n393), .A2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  OR2_X1    g0211(.A1(new_n411), .A2(KEYINPUT76), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT13), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n273), .B1(new_n281), .B2(G238), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n209), .A2(new_n261), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n415), .B1(G232), .B2(new_n261), .ZN(new_n416));
  OAI22_X1  g0216(.A1(new_n416), .A2(new_n363), .B1(new_n257), .B2(new_n221), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(new_n322), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n413), .B1(new_n414), .B2(new_n418), .ZN(new_n419));
  AND3_X1   g0219(.A1(new_n268), .A2(new_n279), .A3(new_n271), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n279), .B1(new_n268), .B2(new_n271), .ZN(new_n421));
  OAI21_X1  g0221(.A(G238), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  AND4_X1   g0222(.A1(new_n413), .A2(new_n418), .A3(new_n422), .A4(new_n274), .ZN(new_n423));
  OAI21_X1  g0223(.A(G169), .B1(new_n419), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(KEYINPUT14), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n419), .A2(new_n423), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(G179), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT14), .ZN(new_n428));
  OAI211_X1 g0228(.A(new_n428), .B(G169), .C1(new_n419), .C2(new_n423), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n425), .A2(new_n427), .A3(new_n429), .ZN(new_n430));
  AOI22_X1  g0230(.A1(new_n289), .A2(G77), .B1(G20), .B2(new_n210), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n431), .B1(new_n202), .B2(new_n330), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(new_n297), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(KEYINPUT74), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT74), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n432), .A2(new_n435), .A3(new_n297), .ZN(new_n436));
  AND3_X1   g0236(.A1(new_n434), .A2(KEYINPUT11), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n301), .A2(G68), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT12), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n439), .B1(new_n370), .B2(G68), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n299), .A2(KEYINPUT12), .A3(new_n210), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n438), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  AOI21_X1  g0242(.A(KEYINPUT11), .B1(new_n434), .B2(new_n436), .ZN(new_n443));
  NOR3_X1   g0243(.A1(new_n437), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n430), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n426), .A2(G190), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n444), .B(new_n447), .C1(new_n426), .C2(new_n401), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n449), .B1(new_n411), .B2(KEYINPUT76), .ZN(new_n450));
  AND3_X1   g0250(.A1(new_n349), .A2(new_n412), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n270), .A2(G33), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n294), .A2(new_n370), .A3(new_n296), .A4(new_n452), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n453), .A2(new_n218), .ZN(new_n454));
  OR2_X1    g0254(.A1(KEYINPUT77), .A2(G97), .ZN(new_n455));
  NAND2_X1  g0255(.A1(KEYINPUT77), .A2(G97), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n455), .A2(new_n257), .A3(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT85), .ZN(new_n458));
  NAND2_X1  g0258(.A1(G33), .A2(G283), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n457), .A2(new_n458), .A3(new_n234), .A4(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n218), .A2(G20), .ZN(new_n461));
  AND3_X1   g0261(.A1(new_n460), .A2(new_n293), .A3(new_n461), .ZN(new_n462));
  AND2_X1   g0262(.A1(KEYINPUT77), .A2(G97), .ZN(new_n463));
  NOR2_X1   g0263(.A1(KEYINPUT77), .A2(G97), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g0265(.A(G20), .B1(new_n465), .B2(new_n257), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(new_n459), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(KEYINPUT85), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n462), .A2(new_n468), .A3(KEYINPUT20), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT20), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n460), .A2(new_n293), .A3(new_n461), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n458), .B1(new_n466), .B2(new_n459), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n454), .B1(new_n469), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n299), .A2(new_n218), .ZN(new_n475));
  XOR2_X1   g0275(.A(new_n475), .B(KEYINPUT84), .Z(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n474), .A2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT21), .ZN(new_n479));
  AND2_X1   g0279(.A1(G264), .A2(G1698), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n480), .B1(new_n361), .B2(new_n362), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(KEYINPUT82), .ZN(new_n482));
  OAI211_X1 g0282(.A(G257), .B(new_n261), .C1(new_n361), .C2(new_n362), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n363), .A2(G303), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT82), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n485), .B(new_n480), .C1(new_n361), .C2(new_n362), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n482), .A2(new_n483), .A3(new_n484), .A4(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(KEYINPUT83), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n222), .B1(new_n258), .B2(new_n259), .ZN(new_n489));
  AOI22_X1  g0289(.A1(new_n489), .A2(new_n261), .B1(new_n363), .B2(G303), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT83), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n490), .A2(new_n491), .A3(new_n482), .A4(new_n486), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n488), .A2(new_n492), .A3(new_n322), .ZN(new_n493));
  NOR2_X1   g0293(.A1(KEYINPUT5), .A2(G41), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(KEYINPUT5), .A2(G41), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(G45), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n498), .A2(G1), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n497), .A2(G274), .A3(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(new_n500), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n322), .B1(new_n499), .B2(new_n497), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n501), .B1(G270), .B2(new_n502), .ZN(new_n503));
  AOI211_X1 g0303(.A(new_n479), .B(new_n304), .C1(new_n493), .C2(new_n503), .ZN(new_n504));
  AND3_X1   g0304(.A1(new_n493), .A2(G179), .A3(new_n503), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n478), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT86), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AOI211_X1 g0308(.A(new_n454), .B(new_n476), .C1(new_n469), .C2(new_n473), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n493), .A2(new_n503), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(G169), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n479), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  OAI211_X1 g0312(.A(KEYINPUT86), .B(new_n478), .C1(new_n504), .C2(new_n505), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n510), .A2(G200), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n509), .B(new_n514), .C1(new_n340), .C2(new_n510), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n508), .A2(new_n512), .A3(new_n513), .A4(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT19), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(KEYINPUT80), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT80), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(KEYINPUT19), .ZN(new_n520));
  AND2_X1   g0320(.A1(G33), .A2(G97), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n518), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  AND3_X1   g0322(.A1(new_n522), .A2(KEYINPUT81), .A3(new_n234), .ZN(new_n523));
  AOI21_X1  g0323(.A(KEYINPUT81), .B1(new_n522), .B2(new_n234), .ZN(new_n524));
  NOR3_X1   g0324(.A1(new_n465), .A2(G87), .A3(G107), .ZN(new_n525));
  NOR3_X1   g0325(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n465), .A2(new_n289), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n518), .A2(new_n520), .ZN(new_n528));
  AOI21_X1  g0328(.A(G20), .B1(new_n258), .B2(new_n259), .ZN(new_n529));
  AOI22_X1  g0329(.A1(new_n527), .A2(new_n528), .B1(new_n529), .B2(G68), .ZN(new_n530));
  INV_X1    g0330(.A(new_n530), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n297), .B1(new_n526), .B2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(new_n332), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n533), .A2(new_n370), .ZN(new_n534));
  INV_X1    g0334(.A(new_n534), .ZN(new_n535));
  OR2_X1    g0335(.A1(new_n453), .A2(new_n332), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n532), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n217), .B1(new_n499), .B2(KEYINPUT78), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT79), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT78), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n540), .B1(new_n498), .B2(G1), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n538), .A2(new_n539), .A3(new_n268), .A4(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n270), .A2(KEYINPUT78), .A3(G45), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n268), .A2(new_n541), .A3(G250), .A4(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(KEYINPUT79), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  NOR3_X1   g0346(.A1(new_n498), .A2(new_n272), .A3(G1), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n211), .A2(new_n261), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n324), .A2(G1698), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n548), .B(new_n549), .C1(new_n361), .C2(new_n362), .ZN(new_n550));
  NAND2_X1  g0350(.A1(G33), .A2(G116), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n547), .B1(new_n552), .B2(new_n322), .ZN(new_n553));
  AND2_X1   g0353(.A1(new_n546), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(new_n285), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n546), .A2(new_n553), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(new_n304), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n537), .A2(new_n555), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n522), .A2(new_n234), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT81), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(new_n465), .ZN(new_n562));
  INV_X1    g0362(.A(G107), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n562), .A2(new_n216), .A3(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n522), .A2(KEYINPUT81), .A3(new_n234), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n561), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(new_n530), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n534), .B1(new_n567), .B2(new_n297), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n554), .A2(G190), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n556), .A2(G200), .ZN(new_n570));
  OR2_X1    g0370(.A1(new_n453), .A2(new_n216), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n568), .A2(new_n569), .A3(new_n570), .A4(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n558), .A2(new_n572), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n516), .A2(new_n573), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n234), .A2(G107), .ZN(new_n575));
  XNOR2_X1  g0375(.A(new_n575), .B(KEYINPUT23), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n234), .A2(G33), .A3(G116), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT22), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n578), .B1(new_n529), .B2(G87), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n234), .B(G87), .C1(new_n361), .C2(new_n362), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n580), .A2(KEYINPUT22), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n576), .B(new_n577), .C1(new_n579), .C2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT24), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  XNOR2_X1  g0384(.A(new_n580), .B(KEYINPUT22), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n585), .A2(KEYINPUT24), .A3(new_n576), .A4(new_n577), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n584), .A2(new_n586), .A3(new_n297), .ZN(new_n587));
  OR2_X1    g0387(.A1(new_n453), .A2(new_n563), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n299), .A2(KEYINPUT25), .A3(new_n563), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(KEYINPUT87), .ZN(new_n590));
  AOI21_X1  g0390(.A(KEYINPUT25), .B1(new_n299), .B2(new_n563), .ZN(new_n591));
  XOR2_X1   g0391(.A(new_n590), .B(new_n591), .Z(new_n592));
  AOI21_X1  g0392(.A(new_n217), .B1(new_n258), .B2(new_n259), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(new_n261), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n260), .A2(G257), .A3(G1698), .ZN(new_n595));
  NAND2_X1  g0395(.A1(G33), .A2(G294), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  AOI22_X1  g0397(.A1(new_n597), .A2(new_n322), .B1(G264), .B2(new_n502), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n598), .A2(G190), .A3(new_n500), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n587), .A2(new_n588), .A3(new_n592), .A4(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n597), .A2(new_n322), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n502), .A2(G264), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n601), .A2(new_n500), .A3(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(new_n603), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n604), .A2(new_n401), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n600), .A2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(new_n297), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n330), .A2(new_n205), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n455), .A2(KEYINPUT6), .A3(new_n563), .A4(new_n456), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT6), .ZN(new_n611));
  AND2_X1   g0411(.A1(G97), .A2(G107), .ZN(new_n612));
  NOR2_X1   g0412(.A1(G97), .A2(G107), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n611), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n610), .A2(new_n614), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n609), .B1(new_n615), .B2(G20), .ZN(new_n616));
  OAI21_X1  g0416(.A(G107), .B1(new_n364), .B2(new_n365), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n608), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n453), .A2(new_n221), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n370), .A2(G97), .ZN(new_n620));
  NOR3_X1   g0420(.A1(new_n618), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT4), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n622), .A2(G1698), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n623), .B(G244), .C1(new_n362), .C2(new_n361), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n324), .B1(new_n258), .B2(new_n259), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n624), .B(new_n459), .C1(new_n625), .C2(KEYINPUT4), .ZN(new_n626));
  OAI21_X1  g0426(.A(G250), .B1(new_n361), .B2(new_n362), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n261), .B1(new_n627), .B2(KEYINPUT4), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n322), .B1(new_n626), .B2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(new_n496), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n499), .B1(new_n630), .B2(new_n494), .ZN(new_n631));
  AND3_X1   g0431(.A1(new_n631), .A2(G257), .A3(new_n268), .ZN(new_n632));
  INV_X1    g0432(.A(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n629), .A2(new_n500), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(G200), .ZN(new_n635));
  OAI21_X1  g0435(.A(G1698), .B1(new_n593), .B2(new_n622), .ZN(new_n636));
  OAI21_X1  g0436(.A(G244), .B1(new_n361), .B2(new_n362), .ZN(new_n637));
  AOI22_X1  g0437(.A1(new_n637), .A2(new_n622), .B1(G33), .B2(G283), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n636), .A2(new_n638), .A3(new_n624), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n632), .B1(new_n639), .B2(new_n322), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n640), .A2(G190), .A3(new_n500), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n621), .A2(new_n635), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n634), .A2(new_n304), .ZN(new_n643));
  INV_X1    g0443(.A(new_n619), .ZN(new_n644));
  INV_X1    g0444(.A(new_n620), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n563), .B1(new_n353), .B2(new_n354), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n234), .B1(new_n610), .B2(new_n614), .ZN(new_n647));
  NOR3_X1   g0447(.A1(new_n646), .A2(new_n647), .A3(new_n609), .ZN(new_n648));
  OAI211_X1 g0448(.A(new_n644), .B(new_n645), .C1(new_n648), .C2(new_n608), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n640), .A2(new_n285), .A3(new_n500), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n643), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n642), .A2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n587), .A2(new_n588), .A3(new_n592), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n603), .A2(G169), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT88), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n598), .A2(G179), .A3(new_n500), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n655), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n604), .A2(KEYINPUT88), .A3(G179), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n654), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n607), .A2(new_n653), .A3(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  AND3_X1   g0462(.A1(new_n451), .A2(new_n574), .A3(new_n662), .ZN(G372));
  NAND3_X1  g0463(.A1(new_n506), .A2(new_n512), .A3(new_n660), .ZN(new_n664));
  INV_X1    g0464(.A(new_n569), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n532), .A2(new_n570), .A3(new_n571), .A4(new_n535), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n665), .B1(new_n666), .B2(KEYINPUT89), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT89), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n568), .A2(new_n668), .A3(new_n570), .A4(new_n571), .ZN(new_n669));
  AOI22_X1  g0469(.A1(new_n568), .A2(new_n536), .B1(new_n304), .B2(new_n556), .ZN(new_n670));
  AOI22_X1  g0470(.A1(new_n667), .A2(new_n669), .B1(new_n555), .B2(new_n670), .ZN(new_n671));
  OAI211_X1 g0471(.A(new_n642), .B(new_n651), .C1(new_n600), .C2(new_n605), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  AND3_X1   g0473(.A1(new_n664), .A2(new_n671), .A3(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n558), .ZN(new_n675));
  AOI21_X1  g0475(.A(G169), .B1(new_n640), .B2(new_n500), .ZN(new_n676));
  AND4_X1   g0476(.A1(new_n285), .A2(new_n629), .A3(new_n500), .A4(new_n633), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n558), .A2(new_n678), .A3(new_n572), .A4(new_n649), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n675), .B1(new_n679), .B2(KEYINPUT26), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n666), .A2(KEYINPUT89), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n681), .A2(new_n569), .A3(new_n669), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT26), .ZN(new_n683));
  AND3_X1   g0483(.A1(new_n643), .A2(new_n649), .A3(new_n650), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n682), .A2(new_n683), .A3(new_n558), .A4(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n680), .A2(new_n685), .ZN(new_n686));
  OR2_X1    g0486(.A1(new_n674), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n451), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n338), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n448), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(new_n446), .ZN(new_n691));
  INV_X1    g0491(.A(new_n409), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n393), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  OR2_X1    g0493(.A1(new_n693), .A2(KEYINPUT90), .ZN(new_n694));
  AOI22_X1  g0494(.A1(new_n693), .A2(KEYINPUT90), .B1(new_n318), .B2(new_n315), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n307), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n688), .A2(new_n696), .ZN(G369));
  NAND2_X1  g0497(.A1(new_n506), .A2(new_n512), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n298), .A2(G20), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(new_n270), .ZN(new_n700));
  OR2_X1    g0500(.A1(new_n700), .A2(KEYINPUT27), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(KEYINPUT27), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n701), .A2(G213), .A3(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(G343), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n509), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n698), .A2(new_n707), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n708), .B1(new_n516), .B2(new_n707), .ZN(new_n709));
  XNOR2_X1  g0509(.A(new_n709), .B(KEYINPUT91), .ZN(new_n710));
  AND2_X1   g0510(.A1(new_n654), .A2(new_n705), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n660), .B1(new_n711), .B2(new_n606), .ZN(new_n712));
  INV_X1    g0512(.A(new_n660), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(new_n706), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n710), .A2(G330), .A3(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n508), .A2(new_n512), .A3(new_n513), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n718), .A2(new_n660), .A3(new_n607), .A4(new_n706), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(new_n714), .ZN(new_n720));
  XNOR2_X1  g0520(.A(new_n720), .B(KEYINPUT92), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n717), .A2(new_n721), .ZN(G399));
  INV_X1    g0522(.A(new_n226), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n723), .A2(G41), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(G1), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n525), .A2(new_n218), .ZN(new_n727));
  OAI22_X1  g0527(.A1(new_n726), .A2(new_n727), .B1(new_n231), .B2(new_n725), .ZN(new_n728));
  XNOR2_X1  g0528(.A(new_n728), .B(KEYINPUT28), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n640), .A2(new_n500), .A3(new_n598), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n505), .A2(new_n731), .A3(KEYINPUT30), .A4(new_n554), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT30), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n493), .A2(new_n554), .A3(G179), .A4(new_n503), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n733), .B1(new_n734), .B2(new_n730), .ZN(new_n735));
  AOI21_X1  g0535(.A(G179), .B1(new_n493), .B2(new_n503), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n736), .A2(new_n556), .A3(new_n603), .A4(new_n634), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n732), .A2(new_n735), .A3(new_n737), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n738), .A2(KEYINPUT31), .A3(new_n705), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT93), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n738), .A2(new_n705), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT31), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n741), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n742), .A2(new_n740), .A3(new_n743), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NOR4_X1   g0547(.A1(new_n516), .A2(new_n661), .A3(new_n573), .A4(new_n705), .ZN(new_n748));
  OAI21_X1  g0548(.A(G330), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(KEYINPUT94), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT94), .ZN(new_n751));
  OAI211_X1 g0551(.A(new_n751), .B(G330), .C1(new_n747), .C2(new_n748), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n687), .A2(new_n706), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(KEYINPUT95), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT29), .ZN(new_n756));
  INV_X1    g0556(.A(KEYINPUT95), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n687), .A2(new_n757), .A3(new_n706), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n755), .A2(new_n756), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n682), .A2(new_n558), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(new_n672), .ZN(new_n761));
  NAND4_X1  g0561(.A1(new_n508), .A2(new_n512), .A3(new_n513), .A4(new_n660), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND4_X1  g0563(.A1(new_n684), .A2(new_n558), .A3(new_n683), .A4(new_n572), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(new_n558), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n682), .A2(new_n558), .A3(new_n684), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n765), .B1(KEYINPUT26), .B2(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n763), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(new_n706), .ZN(new_n769));
  INV_X1    g0569(.A(KEYINPUT96), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n768), .A2(KEYINPUT96), .A3(new_n706), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(KEYINPUT29), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n753), .B1(new_n759), .B2(new_n774), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n729), .B1(new_n775), .B2(G1), .ZN(G364));
  AOI21_X1  g0576(.A(new_n726), .B1(G45), .B2(new_n699), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n777), .B1(new_n710), .B2(G330), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n778), .B1(G330), .B2(new_n710), .ZN(new_n779));
  NAND3_X1  g0579(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n780));
  INV_X1    g0580(.A(KEYINPUT98), .ZN(new_n781));
  OR2_X1    g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n780), .A2(new_n781), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n784), .A2(new_n340), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n234), .A2(G190), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n285), .A2(G200), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  OAI22_X1  g0589(.A1(new_n786), .A2(new_n202), .B1(new_n205), .B2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(G179), .A2(G200), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(G190), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(G20), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(G97), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n234), .A2(new_n340), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(new_n788), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n401), .A2(G179), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n797), .A2(new_n787), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n795), .A2(new_n797), .ZN(new_n799));
  OAI221_X1 g0599(.A(new_n260), .B1(new_n798), .B2(new_n563), .C1(new_n216), .C2(new_n799), .ZN(new_n800));
  OAI221_X1 g0600(.A(new_n794), .B1(new_n250), .B2(new_n796), .C1(new_n800), .C2(KEYINPUT100), .ZN(new_n801));
  AOI211_X1 g0601(.A(new_n790), .B(new_n801), .C1(KEYINPUT100), .C2(new_n800), .ZN(new_n802));
  XNOR2_X1  g0602(.A(KEYINPUT99), .B(G159), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n787), .A2(new_n791), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n806), .B(KEYINPUT32), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n782), .A2(new_n340), .A3(new_n783), .ZN(new_n808));
  OAI211_X1 g0608(.A(new_n802), .B(new_n807), .C1(new_n210), .C2(new_n808), .ZN(new_n809));
  XOR2_X1   g0609(.A(new_n809), .B(KEYINPUT101), .Z(new_n810));
  INV_X1    g0610(.A(G303), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n799), .A2(new_n811), .ZN(new_n812));
  XNOR2_X1  g0612(.A(KEYINPUT102), .B(G317), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n813), .B(KEYINPUT33), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n814), .A2(new_n808), .ZN(new_n815));
  INV_X1    g0615(.A(new_n789), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n260), .B1(new_n816), .B2(G311), .ZN(new_n817));
  INV_X1    g0617(.A(G294), .ZN(new_n818));
  INV_X1    g0618(.A(new_n793), .ZN(new_n819));
  INV_X1    g0619(.A(G322), .ZN(new_n820));
  OAI221_X1 g0620(.A(new_n817), .B1(new_n818), .B2(new_n819), .C1(new_n820), .C2(new_n796), .ZN(new_n821));
  INV_X1    g0621(.A(new_n805), .ZN(new_n822));
  AOI211_X1 g0622(.A(new_n815), .B(new_n821), .C1(G329), .C2(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n785), .A2(G326), .ZN(new_n824));
  INV_X1    g0624(.A(G283), .ZN(new_n825));
  OAI211_X1 g0625(.A(new_n823), .B(new_n824), .C1(new_n825), .C2(new_n798), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n810), .B1(new_n812), .B2(new_n826), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n233), .B1(G20), .B2(new_n304), .ZN(new_n828));
  NOR2_X1   g0628(.A1(G13), .A2(G33), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n830), .A2(G20), .ZN(new_n831));
  XOR2_X1   g0631(.A(new_n831), .B(KEYINPUT97), .Z(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n833), .A2(new_n828), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n260), .A2(G355), .A3(new_n226), .ZN(new_n835));
  AND2_X1   g0635(.A1(new_n251), .A2(G45), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n723), .A2(new_n260), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n837), .B1(G45), .B2(new_n231), .ZN(new_n838));
  OAI221_X1 g0638(.A(new_n835), .B1(G116), .B2(new_n226), .C1(new_n836), .C2(new_n838), .ZN(new_n839));
  AOI22_X1  g0639(.A1(new_n827), .A2(new_n828), .B1(new_n834), .B2(new_n839), .ZN(new_n840));
  OAI211_X1 g0640(.A(new_n840), .B(new_n777), .C1(new_n709), .C2(new_n832), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n779), .A2(new_n841), .ZN(G396));
  INV_X1    g0642(.A(new_n777), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n789), .A2(new_n218), .ZN(new_n844));
  AOI22_X1  g0644(.A1(new_n785), .A2(G303), .B1(G97), .B2(new_n793), .ZN(new_n845));
  OAI221_X1 g0645(.A(new_n845), .B1(new_n563), .B2(new_n799), .C1(new_n818), .C2(new_n796), .ZN(new_n846));
  AOI211_X1 g0646(.A(new_n844), .B(new_n846), .C1(G311), .C2(new_n822), .ZN(new_n847));
  INV_X1    g0647(.A(new_n798), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n848), .A2(G87), .ZN(new_n849));
  XOR2_X1   g0649(.A(new_n808), .B(KEYINPUT103), .Z(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(G283), .ZN(new_n851));
  NAND4_X1  g0651(.A1(new_n847), .A2(new_n363), .A3(new_n849), .A4(new_n851), .ZN(new_n852));
  XNOR2_X1  g0652(.A(new_n852), .B(KEYINPUT104), .ZN(new_n853));
  INV_X1    g0653(.A(new_n808), .ZN(new_n854));
  INV_X1    g0654(.A(new_n796), .ZN(new_n855));
  AOI22_X1  g0655(.A1(new_n854), .A2(G150), .B1(G143), .B2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(G137), .ZN(new_n857));
  OAI221_X1 g0657(.A(new_n856), .B1(new_n786), .B2(new_n857), .C1(new_n789), .C2(new_n804), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT34), .ZN(new_n859));
  INV_X1    g0659(.A(new_n799), .ZN(new_n860));
  AOI22_X1  g0660(.A1(new_n858), .A2(new_n859), .B1(G50), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n822), .A2(G132), .ZN(new_n862));
  OAI211_X1 g0662(.A(new_n861), .B(new_n862), .C1(new_n210), .C2(new_n798), .ZN(new_n863));
  OAI221_X1 g0663(.A(new_n260), .B1(new_n250), .B2(new_n819), .C1(new_n858), .C2(new_n859), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n853), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n843), .B1(new_n865), .B2(new_n828), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n828), .A2(new_n829), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n866), .B1(G77), .B2(new_n868), .ZN(new_n869));
  XNOR2_X1  g0669(.A(new_n869), .B(KEYINPUT105), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n338), .A2(new_n705), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n336), .A2(new_n705), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n872), .B1(new_n341), .B2(new_n342), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n871), .B1(new_n873), .B2(new_n338), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n870), .B1(new_n830), .B2(new_n874), .ZN(new_n875));
  XNOR2_X1  g0675(.A(new_n875), .B(KEYINPUT106), .ZN(new_n876));
  INV_X1    g0676(.A(new_n874), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n755), .A2(new_n758), .A3(new_n877), .ZN(new_n878));
  XOR2_X1   g0678(.A(new_n878), .B(KEYINPUT107), .Z(new_n879));
  OAI211_X1 g0679(.A(new_n706), .B(new_n874), .C1(new_n674), .C2(new_n686), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n881), .A2(new_n752), .A3(new_n750), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n879), .A2(new_n753), .A3(new_n880), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n882), .A2(new_n883), .A3(new_n843), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n876), .A2(new_n884), .ZN(G384));
  NAND3_X1  g0685(.A1(new_n451), .A2(new_n759), .A3(new_n774), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(new_n696), .ZN(new_n887));
  OAI21_X1  g0687(.A(KEYINPUT109), .B1(new_n444), .B2(new_n706), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT109), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n445), .A2(new_n889), .A3(new_n705), .ZN(new_n890));
  NAND4_X1  g0690(.A1(new_n446), .A2(new_n448), .A3(new_n888), .A4(new_n890), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n430), .A2(new_n445), .A3(new_n705), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(new_n871), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n880), .A2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT108), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n880), .A2(KEYINPUT108), .A3(new_n895), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n894), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT37), .ZN(new_n901));
  INV_X1    g0701(.A(new_n703), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n373), .A2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT110), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n901), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n404), .A2(new_n407), .ZN(new_n906));
  NAND4_X1  g0706(.A1(new_n905), .A2(new_n906), .A3(new_n388), .A4(new_n903), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n906), .A2(new_n388), .A3(new_n903), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n703), .B1(new_n369), .B2(new_n372), .ZN(new_n909));
  OAI21_X1  g0709(.A(KEYINPUT37), .B1(new_n909), .B2(KEYINPUT110), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  AND2_X1   g0711(.A1(new_n907), .A2(new_n911), .ZN(new_n912));
  OAI211_X1 g0712(.A(new_n912), .B(KEYINPUT38), .C1(new_n410), .C2(new_n903), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT38), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n903), .B1(new_n692), .B2(new_n392), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n907), .A2(new_n911), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n914), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n913), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n900), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n393), .A2(new_n703), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n918), .A2(KEYINPUT39), .ZN(new_n921));
  XNOR2_X1  g0721(.A(KEYINPUT112), .B(KEYINPUT39), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n908), .B(new_n901), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT111), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n409), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n403), .A2(KEYINPUT111), .A3(new_n408), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n925), .A2(new_n392), .A3(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n923), .B1(new_n927), .B2(new_n909), .ZN(new_n928));
  OAI211_X1 g0728(.A(new_n913), .B(new_n922), .C1(new_n928), .C2(KEYINPUT38), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n921), .A2(new_n929), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n446), .A2(new_n705), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  AND3_X1   g0732(.A1(new_n919), .A2(new_n920), .A3(new_n932), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n887), .B(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n893), .A2(new_n874), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n574), .A2(new_n662), .A3(new_n706), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n744), .A2(new_n739), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n935), .B1(new_n936), .B2(new_n938), .ZN(new_n939));
  AOI21_X1  g0739(.A(KEYINPUT40), .B1(new_n939), .B2(new_n918), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n926), .A2(new_n392), .ZN(new_n941));
  AOI21_X1  g0741(.A(KEYINPUT111), .B1(new_n403), .B2(new_n408), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n909), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n908), .B(KEYINPUT37), .ZN(new_n944));
  AOI21_X1  g0744(.A(KEYINPUT38), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NOR3_X1   g0745(.A1(new_n915), .A2(new_n916), .A3(new_n914), .ZN(new_n946));
  OAI21_X1  g0746(.A(KEYINPUT40), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  OAI211_X1 g0747(.A(new_n874), .B(new_n893), .C1(new_n748), .C2(new_n937), .ZN(new_n948));
  OAI21_X1  g0748(.A(KEYINPUT113), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n913), .B1(new_n928), .B2(KEYINPUT38), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT113), .ZN(new_n951));
  NAND4_X1  g0751(.A1(new_n939), .A2(new_n950), .A3(new_n951), .A4(KEYINPUT40), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n940), .B1(new_n949), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n936), .A2(new_n938), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n953), .A2(new_n451), .A3(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(new_n451), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n954), .A2(G330), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n949), .A2(new_n952), .ZN(new_n959));
  INV_X1    g0759(.A(new_n940), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n959), .A2(G330), .A3(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n955), .B1(new_n958), .B2(new_n962), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n934), .B(new_n963), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n964), .B1(new_n270), .B2(new_n699), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n218), .B1(new_n615), .B2(KEYINPUT35), .ZN(new_n966));
  OAI211_X1 g0766(.A(new_n966), .B(new_n235), .C1(KEYINPUT35), .C2(new_n615), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n967), .B(KEYINPUT36), .ZN(new_n968));
  OAI21_X1  g0768(.A(G77), .B1(new_n250), .B2(new_n210), .ZN(new_n969));
  OAI22_X1  g0769(.A1(new_n231), .A2(new_n969), .B1(G50), .B2(new_n210), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n970), .A2(G1), .A3(new_n298), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n965), .A2(new_n968), .A3(new_n971), .ZN(G367));
  NAND2_X1  g0772(.A1(new_n568), .A2(new_n571), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(new_n705), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n671), .A2(new_n974), .ZN(new_n975));
  OR2_X1    g0775(.A1(new_n974), .A2(new_n558), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT43), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n977), .A2(KEYINPUT43), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n653), .B1(new_n621), .B2(new_n706), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n684), .A2(new_n705), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT114), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n984), .B(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(new_n713), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n987), .A2(new_n651), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n988), .B(KEYINPUT115), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n989), .A2(new_n705), .ZN(new_n990));
  OR2_X1    g0790(.A1(new_n719), .A2(new_n982), .ZN(new_n991));
  XOR2_X1   g0791(.A(new_n991), .B(KEYINPUT42), .Z(new_n992));
  INV_X1    g0792(.A(new_n992), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n980), .B(new_n981), .C1(new_n990), .C2(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(new_n717), .ZN(new_n995));
  AND2_X1   g0795(.A1(new_n995), .A2(new_n986), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT115), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n988), .B(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n998), .A2(new_n706), .ZN(new_n999));
  NAND4_X1  g0799(.A1(new_n999), .A2(new_n979), .A3(new_n978), .A4(new_n992), .ZN(new_n1000));
  AND3_X1   g0800(.A1(new_n994), .A2(new_n996), .A3(new_n1000), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n996), .B1(new_n994), .B2(new_n1000), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n724), .B(KEYINPUT41), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n721), .A2(new_n984), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(KEYINPUT45), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n1007), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n721), .A2(new_n984), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(KEYINPUT44), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1008), .A2(new_n717), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT44), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1009), .B(new_n1012), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n995), .B1(new_n1013), .B2(new_n1007), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n710), .A2(G330), .ZN(new_n1015));
  AND2_X1   g0815(.A1(new_n718), .A2(new_n706), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n719), .B1(new_n1016), .B2(new_n716), .ZN(new_n1017));
  XOR2_X1   g0817(.A(new_n1015), .B(new_n1017), .Z(new_n1018));
  NAND4_X1  g0818(.A1(new_n1011), .A2(new_n1014), .A3(new_n775), .A4(new_n1018), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1005), .B1(new_n1019), .B2(new_n775), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n270), .B1(new_n699), .B2(G45), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n1021), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1003), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n799), .A2(new_n218), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n1024), .A2(KEYINPUT46), .B1(G317), .B2(new_n822), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n1025), .B1(KEYINPUT46), .B2(new_n1024), .C1(new_n563), .C2(new_n819), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1026), .B1(G283), .B2(new_n816), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n785), .A2(G311), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n363), .B1(new_n562), .B2(new_n798), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1029), .B1(G303), .B2(new_n855), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1027), .A2(new_n1028), .A3(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1031), .B1(G294), .B2(new_n850), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n850), .A2(new_n803), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n816), .A2(G50), .B1(new_n793), .B2(G68), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n363), .B1(new_n848), .B2(G77), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n785), .A2(G143), .ZN(new_n1036));
  NAND4_X1  g0836(.A1(new_n1033), .A2(new_n1034), .A3(new_n1035), .A4(new_n1036), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1037), .B1(G150), .B2(new_n855), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n799), .A2(new_n250), .B1(new_n805), .B2(new_n857), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1039), .B(KEYINPUT116), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1032), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1041));
  XOR2_X1   g0841(.A(new_n1041), .B(KEYINPUT47), .Z(new_n1042));
  NAND2_X1  g0842(.A1(new_n1042), .A2(new_n828), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n978), .A2(new_n833), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n837), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n834), .B1(new_n226), .B2(new_n332), .C1(new_n246), .C2(new_n1045), .ZN(new_n1046));
  NAND4_X1  g0846(.A1(new_n1043), .A2(new_n777), .A3(new_n1044), .A4(new_n1046), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT117), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1023), .A2(new_n1048), .ZN(G387));
  OR2_X1    g0849(.A1(new_n1018), .A2(new_n775), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1018), .A2(new_n775), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1050), .A2(new_n724), .A3(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1045), .B1(new_n243), .B2(G45), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n210), .A2(new_n205), .ZN(new_n1054));
  NOR3_X1   g0854(.A1(new_n287), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n727), .A2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g0856(.A(KEYINPUT50), .B1(new_n287), .B2(G50), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1056), .A2(new_n498), .A3(new_n1057), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1053), .B1(new_n1054), .B2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n727), .A2(new_n226), .A3(new_n260), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n1059), .B(new_n1060), .C1(G107), .C2(new_n226), .ZN(new_n1061));
  OR2_X1    g0861(.A1(new_n1061), .A2(KEYINPUT118), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1061), .A2(KEYINPUT118), .ZN(new_n1063));
  AND3_X1   g0863(.A1(new_n1062), .A2(new_n834), .A3(new_n1063), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n716), .A2(new_n832), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n850), .A2(G311), .B1(G317), .B2(new_n855), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n1066), .B1(new_n811), .B2(new_n789), .C1(new_n820), .C2(new_n786), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n1067), .B(KEYINPUT48), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n1068), .B1(new_n825), .B2(new_n819), .C1(new_n818), .C2(new_n799), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n1069), .B(KEYINPUT49), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n260), .B1(new_n822), .B2(G326), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n1070), .B(new_n1071), .C1(new_n218), .C2(new_n798), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n799), .A2(new_n205), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(G159), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1074), .B1(new_n786), .B2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n363), .B1(new_n822), .B2(G150), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n819), .A2(new_n332), .B1(new_n796), .B2(new_n202), .ZN(new_n1078));
  OAI221_X1 g0878(.A(new_n1077), .B1(new_n210), .B2(new_n789), .C1(new_n1078), .C2(KEYINPUT119), .ZN(new_n1079));
  AOI211_X1 g0879(.A(new_n1076), .B(new_n1079), .C1(KEYINPUT119), .C2(new_n1078), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n288), .ZN(new_n1081));
  OAI221_X1 g0881(.A(new_n1080), .B1(new_n221), .B2(new_n798), .C1(new_n1081), .C2(new_n808), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1072), .A2(new_n1082), .ZN(new_n1083));
  AOI211_X1 g0883(.A(new_n1064), .B(new_n1065), .C1(new_n1083), .C2(new_n828), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n1084), .A2(new_n777), .B1(new_n1018), .B2(new_n1022), .ZN(new_n1085));
  AOI21_X1  g0885(.A(KEYINPUT120), .B1(new_n1052), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1086), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1052), .A2(new_n1085), .A3(KEYINPUT120), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1087), .A2(new_n1088), .ZN(G393));
  NOR2_X1   g0889(.A1(new_n986), .A2(new_n832), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(new_n1090), .B(KEYINPUT121), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n834), .B1(new_n226), .B2(new_n562), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(new_n254), .B2(new_n837), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n789), .A2(new_n287), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n822), .A2(G143), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n849), .B(new_n1095), .C1(new_n210), .C2(new_n799), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n785), .A2(G150), .B1(G159), .B2(new_n855), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(KEYINPUT122), .B(KEYINPUT51), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1098), .ZN(new_n1099));
  AOI211_X1 g0899(.A(new_n1094), .B(new_n1096), .C1(new_n1097), .C2(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1097), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n363), .B1(new_n1101), .B2(new_n1098), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n793), .A2(G77), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n850), .A2(G50), .ZN(new_n1104));
  NAND4_X1  g0904(.A1(new_n1100), .A2(new_n1102), .A3(new_n1103), .A4(new_n1104), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n785), .A2(G317), .B1(G311), .B2(new_n855), .ZN(new_n1106));
  XOR2_X1   g0906(.A(new_n1106), .B(KEYINPUT52), .Z(new_n1107));
  NAND2_X1  g0907(.A1(new_n816), .A2(G294), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n260), .B1(new_n850), .B2(G303), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n798), .A2(new_n563), .B1(new_n805), .B2(new_n820), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1110), .B1(G116), .B2(new_n793), .ZN(new_n1111));
  NAND4_X1  g0911(.A1(new_n1107), .A2(new_n1108), .A3(new_n1109), .A4(new_n1111), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n799), .A2(new_n825), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1105), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1093), .B1(new_n1114), .B2(new_n828), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1091), .A2(new_n777), .A3(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1011), .A2(new_n1014), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1116), .B1(new_n1117), .B2(new_n1021), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n725), .B1(new_n1117), .B2(new_n1051), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1118), .B1(new_n1019), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(G390));
  OAI211_X1 g0921(.A(new_n886), .B(new_n696), .C1(new_n956), .C2(new_n957), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n894), .B1(new_n957), .B2(new_n877), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n877), .B1(new_n750), .B2(new_n752), .ZN(new_n1124));
  AND2_X1   g0924(.A1(new_n873), .A2(new_n338), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n771), .A2(new_n772), .A3(new_n895), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(new_n1124), .A2(new_n893), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  OR2_X1    g0928(.A1(new_n957), .A2(new_n935), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1129), .B1(new_n1124), .B2(new_n893), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n898), .A2(new_n899), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n1123), .A2(new_n1128), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n1122), .A2(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1127), .A2(new_n1126), .A3(new_n893), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n950), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n1136), .A2(new_n931), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1138));
  AOI211_X1 g0938(.A(new_n877), .B(new_n894), .C1(new_n750), .C2(new_n752), .ZN(new_n1139));
  AND2_X1   g0939(.A1(new_n921), .A2(new_n929), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1140), .B1(new_n900), .B2(new_n931), .ZN(new_n1141));
  AND3_X1   g0941(.A1(new_n1138), .A2(new_n1139), .A3(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1129), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1143), .B1(new_n1138), .B2(new_n1141), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1134), .A2(KEYINPUT123), .A3(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(KEYINPUT123), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1145), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1147), .B1(new_n1133), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1133), .A2(new_n1148), .ZN(new_n1150));
  NAND4_X1  g0950(.A1(new_n1146), .A2(new_n1149), .A3(new_n724), .A4(new_n1150), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(G116), .A2(new_n855), .B1(new_n848), .B2(G68), .ZN(new_n1152));
  OAI221_X1 g0952(.A(new_n1152), .B1(new_n216), .B2(new_n799), .C1(new_n562), .C2(new_n789), .ZN(new_n1153));
  AOI211_X1 g0953(.A(new_n260), .B(new_n1153), .C1(G294), .C2(new_n822), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n850), .A2(G107), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n785), .A2(G283), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n1154), .A2(new_n1103), .A3(new_n1155), .A4(new_n1156), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(G132), .A2(new_n855), .B1(new_n822), .B2(G125), .ZN(new_n1158));
  XOR2_X1   g0958(.A(KEYINPUT54), .B(G143), .Z(new_n1159));
  NAND2_X1  g0959(.A1(new_n816), .A2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1158), .A2(new_n260), .A3(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1161), .B1(G50), .B2(new_n848), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n850), .A2(G137), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n785), .A2(G128), .B1(G159), .B2(new_n793), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1162), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n860), .A2(G150), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(new_n1166), .B(KEYINPUT53), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1157), .B1(new_n1165), .B2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1168), .A2(new_n828), .ZN(new_n1169));
  OAI211_X1 g0969(.A(new_n777), .B(new_n1169), .C1(new_n930), .C2(new_n830), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1170), .B1(new_n1081), .B2(new_n867), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1171), .B1(new_n1148), .B2(new_n1022), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1151), .A2(new_n1172), .ZN(G378));
  NOR2_X1   g0973(.A1(new_n887), .A2(new_n958), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1174), .B1(new_n1145), .B2(new_n1132), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT124), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n919), .A2(new_n920), .A3(new_n932), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n315), .A2(new_n318), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1178), .A2(new_n306), .ZN(new_n1179));
  XOR2_X1   g0979(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1180));
  NAND2_X1  g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n303), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n1182), .A2(new_n703), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1180), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n319), .A2(new_n1184), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1181), .A2(new_n1183), .A3(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1183), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n319), .A2(new_n1184), .ZN(new_n1188));
  AOI211_X1 g0988(.A(new_n307), .B(new_n1180), .C1(new_n315), .C2(new_n318), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1187), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  AND2_X1   g0990(.A1(new_n1186), .A2(new_n1190), .ZN(new_n1191));
  AND4_X1   g0991(.A1(G330), .A2(new_n959), .A3(new_n960), .A4(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1191), .B1(new_n953), .B2(G330), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n1176), .B(new_n1177), .C1(new_n1192), .C2(new_n1193), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1177), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1191), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n961), .A2(new_n1196), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n953), .A2(G330), .A3(new_n1191), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1197), .A2(new_n933), .A3(new_n1198), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1195), .A2(KEYINPUT124), .A3(new_n1199), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n1175), .A2(KEYINPUT57), .A3(new_n1194), .A4(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1201), .A2(new_n724), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1202), .A2(KEYINPUT125), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1195), .A2(new_n1199), .ZN(new_n1204));
  AND2_X1   g1004(.A1(new_n1175), .A2(new_n1204), .ZN(new_n1205));
  OR2_X1    g1005(.A1(new_n1205), .A2(KEYINPUT57), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT125), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1201), .A2(new_n1207), .A3(new_n724), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1203), .A2(new_n1206), .A3(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1204), .A2(new_n1022), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1196), .A2(new_n829), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n854), .A2(G97), .B1(G68), .B2(new_n793), .ZN(new_n1212));
  OAI221_X1 g1012(.A(new_n1212), .B1(new_n563), .B2(new_n796), .C1(new_n332), .C2(new_n789), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n798), .A2(new_n250), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n786), .A2(new_n218), .ZN(new_n1215));
  NOR3_X1   g1015(.A1(new_n1213), .A2(new_n1214), .A3(new_n1215), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n260), .A2(G41), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n822), .A2(G283), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1216), .A2(new_n1074), .A3(new_n1217), .A4(new_n1218), .ZN(new_n1219));
  XOR2_X1   g1019(.A(new_n1219), .B(KEYINPUT58), .Z(new_n1220));
  OAI21_X1  g1020(.A(new_n202), .B1(new_n361), .B2(G41), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n854), .A2(G132), .B1(new_n860), .B2(new_n1159), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n785), .A2(G125), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(G128), .A2(new_n855), .B1(new_n816), .B2(G137), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1222), .A2(new_n1223), .A3(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1225), .B1(G150), .B2(new_n793), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT59), .ZN(new_n1227));
  AOI21_X1  g1027(.A(G33), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(G41), .B1(new_n822), .B2(G124), .ZN(new_n1229));
  OAI211_X1 g1029(.A(new_n1228), .B(new_n1229), .C1(new_n798), .C2(new_n804), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1221), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n828), .B1(new_n1220), .B2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n867), .A2(new_n202), .ZN(new_n1234));
  NAND4_X1  g1034(.A1(new_n1211), .A2(new_n777), .A3(new_n1233), .A4(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1210), .A2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1209), .A2(new_n1237), .ZN(G375));
  AOI22_X1  g1038(.A1(new_n850), .A2(G116), .B1(new_n533), .B2(new_n793), .ZN(new_n1239));
  OAI221_X1 g1039(.A(new_n1239), .B1(new_n205), .B2(new_n798), .C1(new_n818), .C2(new_n786), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n799), .A2(new_n221), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n789), .A2(new_n563), .ZN(new_n1242));
  OAI221_X1 g1042(.A(new_n363), .B1(new_n805), .B2(new_n811), .C1(new_n825), .C2(new_n796), .ZN(new_n1243));
  NOR4_X1   g1043(.A1(new_n1240), .A2(new_n1241), .A3(new_n1242), .A4(new_n1243), .ZN(new_n1244));
  OAI22_X1  g1044(.A1(new_n819), .A2(new_n202), .B1(new_n250), .B2(new_n798), .ZN(new_n1245));
  AOI211_X1 g1045(.A(new_n363), .B(new_n1245), .C1(G128), .C2(new_n822), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n850), .A2(new_n1159), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n785), .A2(G132), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(G137), .A2(new_n855), .B1(new_n860), .B2(G159), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1246), .A2(new_n1247), .A3(new_n1248), .A4(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1250), .B1(G150), .B2(new_n816), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n828), .B1(new_n1244), .B2(new_n1251), .ZN(new_n1252));
  OAI211_X1 g1052(.A(new_n777), .B(new_n1252), .C1(new_n893), .C2(new_n830), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1253), .B1(new_n210), .B2(new_n867), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1132), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1254), .B1(new_n1255), .B2(new_n1022), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1122), .A2(new_n1132), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1257), .A2(new_n1004), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1256), .B1(new_n1258), .B2(new_n1133), .ZN(G381));
  OR2_X1    g1059(.A1(G381), .A2(G384), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(G375), .A2(G378), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1023), .A2(new_n1048), .A3(new_n1120), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n1087), .A2(new_n841), .A3(new_n779), .A4(new_n1088), .ZN(new_n1264));
  OR4_X1    g1064(.A1(new_n1260), .A2(new_n1262), .A3(new_n1263), .A4(new_n1264), .ZN(G407));
  OAI211_X1 g1065(.A(G407), .B(G213), .C1(G343), .C2(new_n1262), .ZN(G409));
  INV_X1    g1066(.A(new_n1088), .ZN(new_n1267));
  OAI21_X1  g1067(.A(G396), .B1(new_n1267), .B2(new_n1086), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1264), .A2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  AND3_X1   g1070(.A1(new_n1023), .A2(new_n1048), .A3(new_n1120), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1120), .B1(new_n1023), .B2(new_n1048), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1270), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(G387), .A2(G390), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1274), .A2(new_n1263), .A3(new_n1269), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1273), .A2(new_n1275), .ZN(new_n1276));
  AND3_X1   g1076(.A1(new_n1201), .A2(new_n1207), .A3(new_n724), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1207), .B1(new_n1201), .B2(new_n724), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1205), .A2(KEYINPUT57), .ZN(new_n1279));
  NOR3_X1   g1079(.A1(new_n1277), .A2(new_n1278), .A3(new_n1279), .ZN(new_n1280));
  OAI21_X1  g1080(.A(G378), .B1(new_n1280), .B2(new_n1236), .ZN(new_n1281));
  INV_X1    g1081(.A(G213), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1282), .A2(G343), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1205), .A2(new_n1004), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1200), .A2(new_n1022), .A3(new_n1194), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1285), .A2(new_n1235), .A3(new_n1286), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(G378), .A2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1288), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1281), .A2(new_n1284), .A3(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1257), .A2(KEYINPUT126), .ZN(new_n1291));
  OAI211_X1 g1091(.A(new_n1134), .B(new_n724), .C1(new_n1291), .C2(KEYINPUT60), .ZN(new_n1292));
  AND2_X1   g1092(.A1(new_n1291), .A2(KEYINPUT60), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1256), .B1(new_n1292), .B2(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(G384), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  OAI211_X1 g1096(.A(G384), .B(new_n1256), .C1(new_n1292), .C2(new_n1293), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1283), .A2(G2897), .ZN(new_n1298));
  AND3_X1   g1098(.A1(new_n1296), .A2(new_n1297), .A3(new_n1298), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1298), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1300));
  NOR2_X1   g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  AOI211_X1 g1101(.A(KEYINPUT61), .B(new_n1276), .C1(new_n1290), .C2(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT127), .ZN(new_n1303));
  AND2_X1   g1103(.A1(new_n1151), .A2(new_n1172), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1304), .B1(new_n1209), .B2(new_n1237), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1306));
  NOR4_X1   g1106(.A1(new_n1305), .A2(new_n1306), .A3(new_n1283), .A4(new_n1288), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1303), .B1(new_n1307), .B2(KEYINPUT63), .ZN(new_n1308));
  AND2_X1   g1108(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1309));
  NAND4_X1  g1109(.A1(new_n1281), .A2(new_n1284), .A3(new_n1289), .A4(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT63), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1310), .A2(KEYINPUT127), .A3(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1307), .A2(KEYINPUT63), .ZN(new_n1313));
  NAND4_X1  g1113(.A1(new_n1302), .A2(new_n1308), .A3(new_n1312), .A4(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1310), .A2(KEYINPUT62), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1283), .B1(G375), .B2(G378), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT62), .ZN(new_n1317));
  NAND4_X1  g1117(.A1(new_n1316), .A2(new_n1317), .A3(new_n1289), .A4(new_n1309), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1315), .A2(new_n1318), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT61), .ZN(new_n1320));
  OR2_X1    g1120(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1321));
  NOR3_X1   g1121(.A1(new_n1305), .A2(new_n1283), .A3(new_n1288), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1320), .B1(new_n1321), .B2(new_n1322), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1276), .B1(new_n1319), .B2(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1314), .A2(new_n1324), .ZN(G405));
  NAND3_X1  g1125(.A1(new_n1262), .A2(new_n1276), .A3(new_n1281), .ZN(new_n1326));
  OAI211_X1 g1126(.A(new_n1273), .B(new_n1275), .C1(new_n1261), .C2(new_n1305), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1326), .A2(new_n1327), .ZN(new_n1328));
  XNOR2_X1  g1128(.A(new_n1328), .B(new_n1309), .ZN(G402));
endmodule


