//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 1 1 0 0 0 1 0 1 1 0 1 0 0 1 1 1 0 0 0 0 0 1 1 0 0 1 0 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1 1 1 0 1 1 0 1 1 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:16 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n556, new_n557,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n607, new_n610, new_n612,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1178, new_n1179,
    new_n1180;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT65), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT66), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AND2_X1   g034(.A1(new_n455), .A2(G2106), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT67), .ZN(new_n461));
  OR2_X1    g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  AOI22_X1  g037(.A1(new_n460), .A2(new_n461), .B1(G567), .B2(new_n457), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(new_n464), .ZN(G319));
  INV_X1    g040(.A(KEYINPUT68), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(KEYINPUT68), .A2(G2104), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n468), .A2(KEYINPUT3), .A3(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n467), .A2(KEYINPUT3), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n473), .A2(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G137), .ZN(new_n475));
  XNOR2_X1  g050(.A(KEYINPUT3), .B(G2104), .ZN(new_n476));
  AOI22_X1  g051(.A1(new_n476), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n477));
  INV_X1    g052(.A(G2105), .ZN(new_n478));
  OR2_X1    g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  AND2_X1   g054(.A1(KEYINPUT68), .A2(G2104), .ZN(new_n480));
  NOR2_X1   g055(.A1(KEYINPUT68), .A2(G2104), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n482), .A2(G2105), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G101), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n475), .A2(new_n479), .A3(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G160));
  NAND2_X1  g061(.A1(new_n474), .A2(G136), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n470), .A2(G2105), .A3(new_n472), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G124), .ZN(new_n490));
  OR2_X1    g065(.A1(G100), .A2(G2105), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n491), .B(G2104), .C1(G112), .C2(new_n478), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n487), .A2(new_n490), .A3(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(G162));
  OR2_X1    g069(.A1(new_n478), .A2(G114), .ZN(new_n495));
  OAI21_X1  g070(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(G126), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n498), .B1(new_n488), .B2(new_n499), .ZN(new_n500));
  AND2_X1   g075(.A1(new_n478), .A2(G138), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n470), .A2(new_n472), .A3(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT69), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n470), .A2(KEYINPUT69), .A3(new_n472), .A4(new_n501), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n504), .A2(KEYINPUT4), .A3(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT4), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n476), .A2(new_n507), .A3(new_n501), .ZN(new_n508));
  AOI211_X1 g083(.A(KEYINPUT70), .B(new_n500), .C1(new_n506), .C2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT70), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n471), .B1(new_n482), .B2(KEYINPUT3), .ZN(new_n511));
  AOI21_X1  g086(.A(KEYINPUT69), .B1(new_n511), .B2(new_n501), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n505), .A2(KEYINPUT4), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n508), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(new_n500), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n510), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n509), .A2(new_n516), .ZN(G164));
  XNOR2_X1  g092(.A(KEYINPUT6), .B(G651), .ZN(new_n518));
  XNOR2_X1  g093(.A(KEYINPUT5), .B(G543), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(G88), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n518), .A2(G543), .ZN(new_n522));
  INV_X1    g097(.A(G50), .ZN(new_n523));
  OAI22_X1  g098(.A1(new_n520), .A2(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n519), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n525));
  INV_X1    g100(.A(G651), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n524), .A2(new_n527), .ZN(G166));
  AOI22_X1  g103(.A1(new_n518), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n529));
  INV_X1    g104(.A(new_n519), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n532), .B(KEYINPUT7), .ZN(new_n533));
  INV_X1    g108(.A(G51), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n533), .B1(new_n522), .B2(new_n534), .ZN(new_n535));
  OR3_X1    g110(.A1(new_n531), .A2(new_n535), .A3(KEYINPUT71), .ZN(new_n536));
  OAI21_X1  g111(.A(KEYINPUT71), .B1(new_n531), .B2(new_n535), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n536), .A2(new_n537), .ZN(G168));
  XNOR2_X1  g113(.A(KEYINPUT72), .B(G90), .ZN(new_n539));
  INV_X1    g114(.A(G52), .ZN(new_n540));
  OAI22_X1  g115(.A1(new_n520), .A2(new_n539), .B1(new_n522), .B2(new_n540), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n519), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n542), .A2(new_n526), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n541), .A2(new_n543), .ZN(G171));
  INV_X1    g119(.A(G81), .ZN(new_n545));
  XNOR2_X1  g120(.A(KEYINPUT73), .B(G43), .ZN(new_n546));
  OAI22_X1  g121(.A1(new_n520), .A2(new_n545), .B1(new_n522), .B2(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(KEYINPUT74), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n547), .B(new_n548), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n519), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n550));
  OR2_X1    g125(.A1(new_n550), .A2(new_n526), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G860), .ZN(G153));
  NAND4_X1  g129(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT8), .ZN(new_n557));
  NAND4_X1  g132(.A1(G319), .A2(G483), .A3(G661), .A4(new_n557), .ZN(G188));
  INV_X1    g133(.A(KEYINPUT75), .ZN(new_n559));
  INV_X1    g134(.A(G53), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n559), .B1(new_n522), .B2(new_n560), .ZN(new_n561));
  OR2_X1    g136(.A1(new_n561), .A2(KEYINPUT9), .ZN(new_n562));
  AND2_X1   g137(.A1(new_n518), .A2(G543), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n563), .A2(KEYINPUT75), .A3(G53), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n564), .A2(KEYINPUT9), .A3(new_n561), .ZN(new_n565));
  AND2_X1   g140(.A1(new_n518), .A2(new_n519), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G91), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n519), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n568));
  OR2_X1    g143(.A1(new_n568), .A2(new_n526), .ZN(new_n569));
  NAND4_X1  g144(.A1(new_n562), .A2(new_n565), .A3(new_n567), .A4(new_n569), .ZN(G299));
  INV_X1    g145(.A(G171), .ZN(G301));
  INV_X1    g146(.A(G168), .ZN(G286));
  INV_X1    g147(.A(G166), .ZN(G303));
  OR2_X1    g148(.A1(new_n519), .A2(G74), .ZN(new_n574));
  AOI22_X1  g149(.A1(G651), .A2(new_n574), .B1(new_n563), .B2(G49), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n566), .A2(G87), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n575), .A2(new_n576), .ZN(G288));
  NAND2_X1  g152(.A1(new_n566), .A2(G86), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n563), .A2(G48), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n519), .A2(G61), .ZN(new_n580));
  NAND2_X1  g155(.A1(G73), .A2(G543), .ZN(new_n581));
  XNOR2_X1  g156(.A(new_n581), .B(KEYINPUT76), .ZN(new_n582));
  AND2_X1   g157(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  OAI211_X1 g158(.A(new_n578), .B(new_n579), .C1(new_n583), .C2(new_n526), .ZN(G305));
  INV_X1    g159(.A(G85), .ZN(new_n585));
  INV_X1    g160(.A(G47), .ZN(new_n586));
  OAI22_X1  g161(.A1(new_n520), .A2(new_n585), .B1(new_n522), .B2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT77), .ZN(new_n588));
  XNOR2_X1  g163(.A(new_n587), .B(new_n588), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n519), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n590));
  OR2_X1    g165(.A1(new_n590), .A2(new_n526), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n589), .A2(new_n591), .ZN(G290));
  INV_X1    g167(.A(G868), .ZN(new_n593));
  NOR2_X1   g168(.A1(G301), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n566), .A2(G92), .ZN(new_n595));
  XOR2_X1   g170(.A(new_n595), .B(KEYINPUT10), .Z(new_n596));
  NAND2_X1  g171(.A1(G79), .A2(G543), .ZN(new_n597));
  XNOR2_X1  g172(.A(KEYINPUT78), .B(G66), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n530), .B2(new_n598), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n599), .A2(G651), .B1(new_n563), .B2(G54), .ZN(new_n600));
  AND3_X1   g175(.A1(new_n596), .A2(KEYINPUT79), .A3(new_n600), .ZN(new_n601));
  AOI21_X1  g176(.A(KEYINPUT79), .B1(new_n596), .B2(new_n600), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(new_n604));
  AOI21_X1  g179(.A(new_n594), .B1(new_n604), .B2(new_n593), .ZN(G284));
  AOI21_X1  g180(.A(new_n594), .B1(new_n604), .B2(new_n593), .ZN(G321));
  NOR2_X1   g181(.A1(G299), .A2(G868), .ZN(new_n607));
  AOI21_X1  g182(.A(new_n607), .B1(G868), .B2(G168), .ZN(G297));
  AOI21_X1  g183(.A(new_n607), .B1(G868), .B2(G168), .ZN(G280));
  NOR2_X1   g184(.A1(new_n603), .A2(G559), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n610), .B1(G860), .B2(new_n604), .ZN(G148));
  NAND2_X1  g186(.A1(new_n552), .A2(new_n593), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n612), .B1(new_n610), .B2(new_n593), .ZN(G323));
  XNOR2_X1  g188(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g189(.A1(new_n483), .A2(new_n476), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT12), .ZN(new_n616));
  XOR2_X1   g191(.A(new_n616), .B(KEYINPUT13), .Z(new_n617));
  INV_X1    g192(.A(KEYINPUT80), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n618), .B2(G2100), .ZN(new_n619));
  INV_X1    g194(.A(G2100), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(KEYINPUT80), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n474), .A2(G135), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n489), .A2(G123), .ZN(new_n623));
  OR2_X1    g198(.A1(G99), .A2(G2105), .ZN(new_n624));
  OAI211_X1 g199(.A(new_n624), .B(G2104), .C1(G111), .C2(new_n478), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n622), .A2(new_n623), .A3(new_n625), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(KEYINPUT81), .Z(new_n627));
  OR2_X1    g202(.A1(new_n627), .A2(G2096), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n627), .A2(G2096), .ZN(new_n629));
  NAND3_X1  g204(.A1(new_n617), .A2(new_n618), .A3(G2100), .ZN(new_n630));
  NAND4_X1  g205(.A1(new_n621), .A2(new_n628), .A3(new_n629), .A4(new_n630), .ZN(G156));
  XNOR2_X1  g206(.A(G2427), .B(G2438), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2430), .ZN(new_n633));
  XNOR2_X1  g208(.A(KEYINPUT15), .B(G2435), .ZN(new_n634));
  OR2_X1    g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n633), .A2(new_n634), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n635), .A2(KEYINPUT14), .A3(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2451), .B(G2454), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT16), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n637), .B(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(G2443), .B(G2446), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(G1341), .B(G1348), .ZN(new_n643));
  INV_X1    g218(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n645), .B(KEYINPUT82), .Z(new_n646));
  OAI21_X1  g221(.A(G14), .B1(new_n642), .B2(new_n644), .ZN(new_n647));
  NOR2_X1   g222(.A1(new_n646), .A2(new_n647), .ZN(G401));
  XOR2_X1   g223(.A(G2084), .B(G2090), .Z(new_n649));
  XNOR2_X1  g224(.A(G2067), .B(G2678), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n650), .B(KEYINPUT83), .Z(new_n651));
  NOR2_X1   g226(.A1(G2072), .A2(G2078), .ZN(new_n652));
  NOR2_X1   g227(.A1(new_n444), .A2(new_n652), .ZN(new_n653));
  AOI21_X1  g228(.A(new_n649), .B1(new_n651), .B2(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(KEYINPUT17), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n654), .B1(new_n651), .B2(new_n655), .ZN(new_n656));
  OAI211_X1 g231(.A(new_n649), .B(new_n650), .C1(new_n444), .C2(new_n652), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n657), .B(KEYINPUT18), .Z(new_n658));
  NAND3_X1  g233(.A1(new_n655), .A2(new_n651), .A3(new_n649), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n656), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(G2096), .B(G2100), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(G227));
  XOR2_X1   g237(.A(G1971), .B(G1976), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT19), .ZN(new_n664));
  XOR2_X1   g239(.A(G1956), .B(G2474), .Z(new_n665));
  XOR2_X1   g240(.A(G1961), .B(G1966), .Z(new_n666));
  AND2_X1   g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT20), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n665), .A2(new_n666), .ZN(new_n670));
  NOR3_X1   g245(.A1(new_n664), .A2(new_n667), .A3(new_n670), .ZN(new_n671));
  AOI21_X1  g246(.A(new_n671), .B1(new_n664), .B2(new_n670), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n674));
  XOR2_X1   g249(.A(new_n673), .B(new_n674), .Z(new_n675));
  XNOR2_X1  g250(.A(G1991), .B(G1996), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1981), .B(G1986), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(G229));
  INV_X1    g255(.A(G16), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n681), .A2(G23), .ZN(new_n682));
  INV_X1    g257(.A(G288), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n682), .B1(new_n683), .B2(new_n681), .ZN(new_n684));
  XNOR2_X1  g259(.A(KEYINPUT33), .B(G1976), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n681), .A2(G22), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n687), .B1(G166), .B2(new_n681), .ZN(new_n688));
  INV_X1    g263(.A(G1971), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  NOR2_X1   g265(.A1(G6), .A2(G16), .ZN(new_n691));
  INV_X1    g266(.A(G305), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n691), .B1(new_n692), .B2(G16), .ZN(new_n693));
  XOR2_X1   g268(.A(KEYINPUT32), .B(G1981), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n686), .A2(new_n690), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n696), .A2(KEYINPUT34), .ZN(new_n697));
  XOR2_X1   g272(.A(new_n697), .B(KEYINPUT85), .Z(new_n698));
  OR2_X1    g273(.A1(new_n696), .A2(KEYINPUT34), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n681), .A2(G24), .ZN(new_n700));
  INV_X1    g275(.A(G290), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n700), .B1(new_n701), .B2(new_n681), .ZN(new_n702));
  XOR2_X1   g277(.A(KEYINPUT84), .B(G1986), .Z(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(G29), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n705), .A2(G25), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n474), .A2(G131), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n489), .A2(G119), .ZN(new_n708));
  OR2_X1    g283(.A1(G95), .A2(G2105), .ZN(new_n709));
  OAI211_X1 g284(.A(new_n709), .B(G2104), .C1(G107), .C2(new_n478), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n707), .A2(new_n708), .A3(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n706), .B1(new_n712), .B2(new_n705), .ZN(new_n713));
  XOR2_X1   g288(.A(KEYINPUT35), .B(G1991), .Z(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  NAND4_X1  g290(.A1(new_n698), .A2(new_n699), .A3(new_n704), .A4(new_n715), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(KEYINPUT36), .Z(new_n717));
  NAND2_X1  g292(.A1(new_n705), .A2(G35), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(G162), .B2(new_n705), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT29), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n720), .A2(G2090), .ZN(new_n721));
  NOR2_X1   g296(.A1(G4), .A2(G16), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(new_n604), .B2(G16), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(G1348), .ZN(new_n724));
  AND2_X1   g299(.A1(new_n705), .A2(G33), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n474), .A2(G139), .ZN(new_n726));
  NAND3_X1  g301(.A1(new_n478), .A2(G103), .A3(G2104), .ZN(new_n727));
  XOR2_X1   g302(.A(new_n727), .B(KEYINPUT25), .Z(new_n728));
  NAND2_X1  g303(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT87), .ZN(new_n730));
  AOI22_X1  g305(.A1(new_n476), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n730), .B1(new_n478), .B2(new_n731), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n725), .B1(new_n732), .B2(G29), .ZN(new_n733));
  AOI211_X1 g308(.A(new_n721), .B(new_n724), .C1(new_n442), .C2(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n681), .A2(G20), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT23), .ZN(new_n736));
  INV_X1    g311(.A(G299), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n736), .B1(new_n737), .B2(new_n681), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(G1956), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(G2090), .B2(new_n720), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT92), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n705), .A2(G27), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G164), .B2(new_n705), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(G2078), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n741), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n681), .A2(G21), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(G168), .B2(new_n681), .ZN(new_n747));
  XOR2_X1   g322(.A(KEYINPUT86), .B(KEYINPUT28), .Z(new_n748));
  NAND2_X1  g323(.A1(new_n705), .A2(G26), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n474), .A2(G140), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n489), .A2(G128), .ZN(new_n752));
  OR2_X1    g327(.A1(G104), .A2(G2105), .ZN(new_n753));
  OAI211_X1 g328(.A(new_n753), .B(G2104), .C1(G116), .C2(new_n478), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n751), .A2(new_n752), .A3(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(new_n755), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n750), .B1(new_n756), .B2(new_n705), .ZN(new_n757));
  AOI22_X1  g332(.A1(new_n747), .A2(G1966), .B1(new_n757), .B2(G2067), .ZN(new_n758));
  OAI221_X1 g333(.A(new_n758), .B1(G2067), .B2(new_n757), .C1(new_n733), .C2(new_n442), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n681), .A2(G19), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(new_n553), .B2(new_n681), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(G1341), .ZN(new_n762));
  INV_X1    g337(.A(KEYINPUT24), .ZN(new_n763));
  OR2_X1    g338(.A1(new_n763), .A2(G34), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n763), .A2(G34), .ZN(new_n765));
  AOI21_X1  g340(.A(G29), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(new_n485), .B2(G29), .ZN(new_n767));
  XOR2_X1   g342(.A(KEYINPUT88), .B(G2084), .Z(new_n768));
  XNOR2_X1  g343(.A(new_n767), .B(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(KEYINPUT30), .ZN(new_n770));
  INV_X1    g345(.A(KEYINPUT91), .ZN(new_n771));
  AND3_X1   g346(.A1(new_n771), .A2(new_n770), .A3(G28), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n771), .B1(new_n770), .B2(G28), .ZN(new_n773));
  OAI221_X1 g348(.A(new_n705), .B1(new_n770), .B2(G28), .C1(new_n772), .C2(new_n773), .ZN(new_n774));
  XNOR2_X1  g349(.A(KEYINPUT31), .B(G11), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n681), .A2(G5), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G171), .B2(new_n681), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n776), .B1(new_n778), .B2(G1961), .ZN(new_n779));
  OAI211_X1 g354(.A(new_n769), .B(new_n779), .C1(G1961), .C2(new_n778), .ZN(new_n780));
  OAI22_X1  g355(.A1(new_n627), .A2(new_n705), .B1(new_n747), .B2(G1966), .ZN(new_n781));
  NOR4_X1   g356(.A1(new_n759), .A2(new_n762), .A3(new_n780), .A4(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n705), .A2(G32), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n474), .A2(G141), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n784), .B(KEYINPUT89), .Z(new_n785));
  NAND2_X1  g360(.A1(new_n489), .A2(G129), .ZN(new_n786));
  NAND3_X1  g361(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(KEYINPUT26), .Z(new_n788));
  NAND2_X1  g363(.A1(new_n483), .A2(G105), .ZN(new_n789));
  AND4_X1   g364(.A1(new_n785), .A2(new_n786), .A3(new_n788), .A4(new_n789), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n783), .B1(new_n790), .B2(new_n705), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT90), .ZN(new_n792));
  XNOR2_X1  g367(.A(KEYINPUT27), .B(G1996), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NAND4_X1  g369(.A1(new_n734), .A2(new_n745), .A3(new_n782), .A4(new_n794), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n717), .A2(new_n795), .ZN(G311));
  INV_X1    g371(.A(G311), .ZN(G150));
  NAND2_X1  g372(.A1(new_n604), .A2(G559), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT38), .ZN(new_n799));
  INV_X1    g374(.A(G93), .ZN(new_n800));
  INV_X1    g375(.A(G55), .ZN(new_n801));
  OAI22_X1  g376(.A1(new_n520), .A2(new_n800), .B1(new_n522), .B2(new_n801), .ZN(new_n802));
  AOI22_X1  g377(.A1(new_n519), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n803), .A2(new_n526), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  INV_X1    g380(.A(new_n805), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n552), .B(new_n806), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n799), .B(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(KEYINPUT39), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  XOR2_X1   g385(.A(new_n810), .B(KEYINPUT94), .Z(new_n811));
  XOR2_X1   g386(.A(KEYINPUT93), .B(G860), .Z(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(new_n808), .B2(new_n809), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n806), .A2(new_n812), .ZN(new_n815));
  XOR2_X1   g390(.A(new_n815), .B(KEYINPUT37), .Z(new_n816));
  NAND2_X1  g391(.A1(new_n814), .A2(new_n816), .ZN(G145));
  XNOR2_X1  g392(.A(new_n790), .B(new_n732), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n489), .A2(G130), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n478), .A2(G118), .ZN(new_n820));
  OAI21_X1  g395(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n819), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n822), .B1(G142), .B2(new_n474), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(new_n616), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n818), .B(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n514), .A2(new_n515), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(new_n755), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(new_n712), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n825), .B(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n627), .B(new_n493), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(new_n485), .ZN(new_n831));
  XNOR2_X1  g406(.A(KEYINPUT95), .B(KEYINPUT96), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n831), .B(new_n832), .ZN(new_n833));
  AND2_X1   g408(.A1(new_n829), .A2(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(G37), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n835), .B1(new_n829), .B2(new_n833), .ZN(new_n836));
  OR2_X1    g411(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g413(.A(new_n610), .B(new_n807), .Z(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT41), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n596), .A2(new_n600), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n842), .A2(new_n737), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT98), .ZN(new_n844));
  INV_X1    g419(.A(new_n844), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n842), .A2(new_n737), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT97), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n841), .B1(new_n845), .B2(new_n847), .ZN(new_n848));
  XOR2_X1   g423(.A(new_n846), .B(KEYINPUT97), .Z(new_n849));
  NAND3_X1  g424(.A1(new_n849), .A2(KEYINPUT41), .A3(new_n844), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT99), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n848), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  OAI211_X1 g427(.A(KEYINPUT99), .B(new_n841), .C1(new_n845), .C2(new_n847), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n840), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n839), .B1(new_n847), .B2(new_n845), .ZN(new_n855));
  XNOR2_X1  g430(.A(G303), .B(G288), .ZN(new_n856));
  NAND2_X1  g431(.A1(G290), .A2(new_n692), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n589), .A2(G305), .A3(new_n591), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n856), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n856), .A2(new_n857), .A3(new_n858), .ZN(new_n861));
  AOI21_X1  g436(.A(KEYINPUT42), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  AOI21_X1  g437(.A(KEYINPUT100), .B1(new_n860), .B2(new_n861), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n860), .A2(KEYINPUT100), .A3(new_n861), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n862), .B1(new_n866), .B2(KEYINPUT42), .ZN(new_n867));
  AND3_X1   g442(.A1(new_n854), .A2(new_n855), .A3(new_n867), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n867), .B1(new_n854), .B2(new_n855), .ZN(new_n869));
  OAI21_X1  g444(.A(G868), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n870), .B1(G868), .B2(new_n805), .ZN(G295));
  OAI21_X1  g446(.A(new_n870), .B1(G868), .B2(new_n805), .ZN(G331));
  INV_X1    g447(.A(KEYINPUT44), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n848), .A2(new_n850), .ZN(new_n874));
  XNOR2_X1  g449(.A(G168), .B(G171), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n807), .B(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n845), .A2(new_n847), .ZN(new_n878));
  OR2_X1    g453(.A1(new_n878), .A2(new_n876), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT102), .ZN(new_n881));
  INV_X1    g456(.A(new_n865), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n881), .B1(new_n882), .B2(new_n863), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n864), .A2(new_n865), .A3(KEYINPUT102), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(G37), .B1(new_n880), .B2(new_n886), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n852), .A2(new_n853), .A3(new_n876), .ZN(new_n888));
  NAND4_X1  g463(.A1(new_n888), .A2(new_n865), .A3(new_n879), .A4(new_n864), .ZN(new_n889));
  XNOR2_X1  g464(.A(KEYINPUT101), .B(KEYINPUT43), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n887), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n889), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT103), .ZN(new_n893));
  AND2_X1   g468(.A1(new_n888), .A2(new_n879), .ZN(new_n894));
  OAI211_X1 g469(.A(new_n893), .B(new_n835), .C1(new_n894), .C2(new_n885), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n885), .B1(new_n888), .B2(new_n879), .ZN(new_n896));
  OAI21_X1  g471(.A(KEYINPUT103), .B1(new_n896), .B2(G37), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n892), .B1(new_n895), .B2(new_n897), .ZN(new_n898));
  OAI211_X1 g473(.A(new_n873), .B(new_n891), .C1(new_n898), .C2(new_n890), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n889), .A2(new_n890), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n900), .B1(new_n895), .B2(new_n897), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT43), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n902), .B1(new_n887), .B2(new_n889), .ZN(new_n903));
  OAI21_X1  g478(.A(KEYINPUT44), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  AND2_X1   g479(.A1(new_n899), .A2(new_n904), .ZN(G397));
  AOI21_X1  g480(.A(G1384), .B1(new_n514), .B2(new_n515), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n906), .A2(KEYINPUT45), .ZN(new_n907));
  NAND4_X1  g482(.A1(new_n475), .A2(new_n479), .A3(G40), .A4(new_n484), .ZN(new_n908));
  INV_X1    g483(.A(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  XOR2_X1   g485(.A(new_n755), .B(G2067), .Z(new_n911));
  XNOR2_X1  g486(.A(new_n911), .B(KEYINPUT104), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n910), .B1(new_n912), .B2(new_n790), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n910), .A2(G1996), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n913), .B1(KEYINPUT46), .B2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n914), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT46), .ZN(new_n917));
  AOI21_X1  g492(.A(KEYINPUT124), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n916), .A2(KEYINPUT124), .A3(new_n917), .ZN(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n915), .B1(new_n918), .B2(new_n920), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n921), .B(KEYINPUT47), .ZN(new_n922));
  INV_X1    g497(.A(G1996), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n912), .A2(new_n923), .ZN(new_n924));
  AOI22_X1  g499(.A1(new_n913), .A2(new_n924), .B1(new_n790), .B2(new_n914), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n712), .A2(new_n714), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n926), .B(KEYINPUT123), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n928), .B1(G2067), .B2(new_n755), .ZN(new_n929));
  INV_X1    g504(.A(new_n910), .ZN(new_n930));
  XOR2_X1   g505(.A(new_n711), .B(new_n714), .Z(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n925), .A2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  NOR3_X1   g509(.A1(new_n910), .A2(G1986), .A3(G290), .ZN(new_n935));
  XOR2_X1   g510(.A(new_n935), .B(KEYINPUT48), .Z(new_n936));
  AOI22_X1  g511(.A1(new_n929), .A2(new_n930), .B1(new_n934), .B2(new_n936), .ZN(new_n937));
  AND2_X1   g512(.A1(new_n922), .A2(new_n937), .ZN(new_n938));
  XNOR2_X1  g513(.A(G290), .B(G1986), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n933), .B1(new_n930), .B2(new_n939), .ZN(new_n940));
  NOR2_X1   g515(.A1(G305), .A2(G1981), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT109), .ZN(new_n942));
  OAI21_X1  g517(.A(KEYINPUT49), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT49), .ZN(new_n944));
  OAI211_X1 g519(.A(KEYINPUT109), .B(new_n944), .C1(G305), .C2(G1981), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(G1981), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n692), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  OAI211_X1 g524(.A(new_n943), .B(new_n945), .C1(new_n947), .C2(new_n692), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n906), .A2(new_n909), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(G8), .ZN(new_n953));
  INV_X1    g528(.A(G1976), .ZN(new_n954));
  OAI211_X1 g529(.A(new_n952), .B(G8), .C1(new_n954), .C2(G288), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT52), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n956), .B1(new_n683), .B2(G1976), .ZN(new_n957));
  OAI22_X1  g532(.A1(new_n951), .A2(new_n953), .B1(new_n955), .B2(new_n957), .ZN(new_n958));
  AND2_X1   g533(.A1(new_n955), .A2(KEYINPUT52), .ZN(new_n959));
  OR2_X1    g534(.A1(new_n959), .A2(KEYINPUT108), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(KEYINPUT108), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n958), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  OAI211_X1 g537(.A(G303), .B(G8), .C1(KEYINPUT106), .C2(KEYINPUT55), .ZN(new_n963));
  XNOR2_X1  g538(.A(KEYINPUT106), .B(KEYINPUT55), .ZN(new_n964));
  INV_X1    g539(.A(G8), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n964), .B1(G166), .B2(new_n965), .ZN(new_n966));
  AND2_X1   g541(.A1(new_n963), .A2(new_n966), .ZN(new_n967));
  XNOR2_X1  g542(.A(new_n967), .B(KEYINPUT107), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT50), .ZN(new_n969));
  INV_X1    g544(.A(G1384), .ZN(new_n970));
  INV_X1    g545(.A(new_n508), .ZN(new_n971));
  AND2_X1   g546(.A1(new_n505), .A2(KEYINPUT4), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n971), .B1(new_n972), .B2(new_n504), .ZN(new_n973));
  OAI211_X1 g548(.A(new_n969), .B(new_n970), .C1(new_n973), .C2(new_n500), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(new_n909), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n970), .B1(new_n509), .B2(new_n516), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n975), .B1(new_n976), .B2(KEYINPUT50), .ZN(new_n977));
  INV_X1    g552(.A(G2090), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n977), .A2(KEYINPUT105), .A3(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n908), .B1(new_n906), .B2(KEYINPUT45), .ZN(new_n980));
  OAI21_X1  g555(.A(KEYINPUT70), .B1(new_n973), .B2(new_n500), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n514), .A2(new_n510), .A3(new_n515), .ZN(new_n982));
  AOI21_X1  g557(.A(G1384), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n980), .B1(new_n983), .B2(KEYINPUT45), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(new_n689), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n979), .A2(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(KEYINPUT105), .B1(new_n977), .B2(new_n978), .ZN(new_n987));
  OAI211_X1 g562(.A(G8), .B(new_n968), .C1(new_n986), .C2(new_n987), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n970), .B1(new_n973), .B2(new_n500), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n908), .B1(new_n989), .B2(KEYINPUT50), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n990), .B1(new_n976), .B2(KEYINPUT50), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n991), .A2(G2090), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT45), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n976), .A2(new_n993), .ZN(new_n994));
  AOI21_X1  g569(.A(G1971), .B1(new_n994), .B2(new_n980), .ZN(new_n995));
  OAI21_X1  g570(.A(G8), .B1(new_n992), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(new_n967), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n962), .A2(new_n988), .A3(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT119), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n976), .A2(KEYINPUT50), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n908), .B1(new_n906), .B2(new_n969), .ZN(new_n1001));
  AOI21_X1  g576(.A(G1961), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  OAI211_X1 g577(.A(KEYINPUT45), .B(new_n970), .C1(new_n509), .C2(new_n516), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n908), .B1(new_n989), .B2(new_n993), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT53), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n1005), .A2(G2078), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1003), .A2(new_n1004), .A3(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n999), .B1(new_n1002), .B2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1001), .B1(new_n983), .B2(new_n969), .ZN(new_n1010));
  INV_X1    g585(.A(G1961), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1012), .A2(KEYINPUT119), .A3(new_n1007), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1009), .A2(new_n1013), .ZN(new_n1014));
  OAI211_X1 g589(.A(new_n443), .B(new_n980), .C1(new_n983), .C2(KEYINPUT45), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(new_n1005), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT120), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1015), .A2(KEYINPUT120), .A3(new_n1005), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1014), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(G171), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n998), .A2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n536), .A2(G8), .A3(new_n537), .ZN(new_n1024));
  XOR2_X1   g599(.A(new_n1024), .B(KEYINPUT117), .Z(new_n1025));
  INV_X1    g600(.A(KEYINPUT118), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT51), .ZN(new_n1027));
  INV_X1    g602(.A(G2084), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1029));
  INV_X1    g604(.A(G1966), .ZN(new_n1030));
  AOI22_X1  g605(.A1(new_n977), .A2(new_n1028), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  OAI221_X1 g606(.A(new_n1025), .B1(new_n1026), .B2(new_n1027), .C1(new_n1031), .C2(new_n965), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1033));
  OAI211_X1 g608(.A(new_n1028), .B(new_n1001), .C1(new_n983), .C2(new_n969), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1025), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n965), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1037), .B1(new_n1038), .B2(new_n1036), .ZN(new_n1039));
  OAI21_X1  g614(.A(KEYINPUT51), .B1(new_n1038), .B2(KEYINPUT118), .ZN(new_n1040));
  OAI211_X1 g615(.A(new_n1032), .B(KEYINPUT62), .C1(new_n1039), .C2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1032), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT62), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1023), .A2(new_n1041), .A3(new_n1044), .ZN(new_n1045));
  OR2_X1    g620(.A1(new_n986), .A2(new_n987), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n962), .A2(new_n1046), .A3(G8), .A4(new_n968), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n683), .A2(new_n954), .ZN(new_n1048));
  XNOR2_X1  g623(.A(new_n1048), .B(KEYINPUT110), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1049), .B1(new_n949), .B2(new_n950), .ZN(new_n1050));
  OAI211_X1 g625(.A(G8), .B(new_n952), .C1(new_n1050), .C2(new_n941), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1047), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT112), .ZN(new_n1054));
  AOI21_X1  g629(.A(G1348), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n952), .A2(G2067), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1054), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  OAI221_X1 g632(.A(KEYINPUT112), .B1(G2067), .B2(new_n952), .C1(new_n977), .C2(G1348), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1057), .A2(new_n1058), .A3(new_n604), .ZN(new_n1059));
  NAND3_X1  g634(.A1(G299), .A2(KEYINPUT111), .A3(KEYINPUT57), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1060), .ZN(new_n1061));
  AOI21_X1  g636(.A(KEYINPUT57), .B1(G299), .B2(KEYINPUT111), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(G1956), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n991), .A2(new_n1064), .ZN(new_n1065));
  XNOR2_X1  g640(.A(KEYINPUT56), .B(G2072), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n994), .A2(new_n980), .A3(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1063), .B1(new_n1065), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1059), .A2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1065), .A2(new_n1063), .A3(new_n1067), .ZN(new_n1071));
  AND2_X1   g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  OAI211_X1 g647(.A(new_n923), .B(new_n980), .C1(new_n983), .C2(KEYINPUT45), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT113), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n994), .A2(KEYINPUT113), .A3(new_n923), .A4(new_n980), .ZN(new_n1076));
  XOR2_X1   g651(.A(KEYINPUT58), .B(G1341), .Z(new_n1077));
  NAND2_X1  g652(.A1(new_n952), .A2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1075), .A2(new_n1076), .A3(new_n1078), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n552), .A2(KEYINPUT114), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1079), .A2(KEYINPUT59), .A3(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT59), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1065), .A2(new_n1067), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1063), .ZN(new_n1086));
  AOI21_X1  g661(.A(KEYINPUT61), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  OR2_X1    g662(.A1(KEYINPUT115), .A2(KEYINPUT61), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1071), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1090));
  OAI211_X1 g665(.A(new_n1071), .B(new_n1088), .C1(new_n1068), .C2(KEYINPUT61), .ZN(new_n1091));
  AND4_X1   g666(.A1(new_n1081), .A2(new_n1084), .A3(new_n1090), .A4(new_n1091), .ZN(new_n1092));
  OAI21_X1  g667(.A(KEYINPUT60), .B1(new_n603), .B2(KEYINPUT116), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(G1348), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1056), .B1(new_n1010), .B2(new_n1095), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1096), .A2(KEYINPUT112), .ZN(new_n1097));
  AOI211_X1 g672(.A(new_n1054), .B(new_n1056), .C1(new_n1010), .C2(new_n1095), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1094), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT116), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n604), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1093), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1101), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT60), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1057), .A2(new_n1058), .A3(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1102), .A2(new_n1105), .A3(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1072), .B1(new_n1092), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT54), .ZN(new_n1110));
  AOI21_X1  g685(.A(G301), .B1(new_n1014), .B2(new_n1020), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n906), .A2(KEYINPUT45), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1004), .A2(KEYINPUT121), .A3(new_n1112), .A4(new_n1006), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT121), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1006), .B1(new_n989), .B2(new_n993), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n909), .B1(new_n906), .B2(KEYINPUT45), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1114), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  OAI211_X1 g692(.A(new_n1113), .B(new_n1117), .C1(new_n977), .C2(G1961), .ZN(new_n1118));
  AOI211_X1 g693(.A(G171), .B(new_n1118), .C1(new_n1018), .C2(new_n1019), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1110), .B1(new_n1111), .B2(new_n1119), .ZN(new_n1120));
  AND3_X1   g695(.A1(new_n962), .A2(new_n988), .A3(new_n997), .ZN(new_n1121));
  AND3_X1   g696(.A1(new_n1015), .A2(KEYINPUT120), .A3(new_n1005), .ZN(new_n1122));
  AOI21_X1  g697(.A(KEYINPUT120), .B1(new_n1015), .B2(new_n1005), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  OAI21_X1  g699(.A(G171), .B1(new_n1124), .B2(new_n1118), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1014), .A2(new_n1020), .A3(G301), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1125), .A2(new_n1126), .A3(KEYINPUT54), .ZN(new_n1127));
  AOI221_X4 g702(.A(new_n1036), .B1(KEYINPUT118), .B2(KEYINPUT51), .C1(new_n1035), .C2(G8), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1040), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1025), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1038), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1130), .B1(new_n1131), .B2(new_n1025), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1128), .B1(new_n1129), .B2(new_n1132), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1120), .A2(new_n1121), .A3(new_n1127), .A4(new_n1133), .ZN(new_n1134));
  OAI211_X1 g709(.A(new_n1045), .B(new_n1053), .C1(new_n1109), .C2(new_n1134), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1131), .A2(G286), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1121), .A2(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT63), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  OAI21_X1  g714(.A(G8), .B1(new_n986), .B2(new_n987), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1140), .A2(new_n967), .ZN(new_n1141));
  NOR3_X1   g716(.A1(new_n1131), .A2(new_n1138), .A3(G286), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1141), .A2(new_n988), .A3(new_n962), .A4(new_n1142), .ZN(new_n1143));
  AND2_X1   g718(.A1(new_n1139), .A2(new_n1143), .ZN(new_n1144));
  OAI211_X1 g719(.A(KEYINPUT122), .B(new_n940), .C1(new_n1135), .C2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1107), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1148));
  AOI211_X1 g723(.A(new_n1101), .B(new_n1093), .C1(new_n1057), .C2(new_n1058), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1084), .A2(new_n1090), .A3(new_n1081), .A4(new_n1091), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1147), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  AND2_X1   g727(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1153));
  AND2_X1   g728(.A1(new_n1127), .A2(new_n1133), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1152), .A2(new_n1153), .A3(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1041), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1026), .B1(new_n1031), .B2(new_n965), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1025), .B1(new_n1031), .B2(new_n965), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1157), .A2(new_n1158), .A3(KEYINPUT51), .A4(new_n1037), .ZN(new_n1159));
  AOI21_X1  g734(.A(KEYINPUT62), .B1(new_n1159), .B2(new_n1032), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n1156), .A2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1052), .B1(new_n1161), .B2(new_n1023), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1139), .A2(new_n1143), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1155), .A2(new_n1162), .A3(new_n1163), .ZN(new_n1164));
  AOI21_X1  g739(.A(KEYINPUT122), .B1(new_n1164), .B2(new_n940), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n938), .B1(new_n1146), .B2(new_n1165), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g741(.A1(G227), .A2(new_n464), .ZN(new_n1168));
  XOR2_X1   g742(.A(new_n1168), .B(KEYINPUT125), .Z(new_n1169));
  NAND2_X1  g743(.A1(new_n679), .A2(new_n1169), .ZN(new_n1170));
  NOR2_X1   g744(.A1(new_n1170), .A2(G401), .ZN(new_n1171));
  INV_X1    g745(.A(KEYINPUT126), .ZN(new_n1172));
  NOR2_X1   g746(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  NOR3_X1   g747(.A1(new_n1170), .A2(KEYINPUT126), .A3(G401), .ZN(new_n1174));
  OAI21_X1  g748(.A(new_n837), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  OR2_X1    g749(.A1(new_n898), .A2(new_n890), .ZN(new_n1176));
  AOI21_X1  g750(.A(new_n1175), .B1(new_n1176), .B2(new_n891), .ZN(G308));
  OR2_X1    g751(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1178));
  NOR2_X1   g752(.A1(new_n898), .A2(new_n890), .ZN(new_n1179));
  INV_X1    g753(.A(new_n891), .ZN(new_n1180));
  OAI211_X1 g754(.A(new_n1178), .B(new_n837), .C1(new_n1179), .C2(new_n1180), .ZN(G225));
endmodule


