

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588;

  INV_X1 U323 ( .A(n536), .ZN(n527) );
  AND2_X1 U324 ( .A1(n571), .A2(n477), .ZN(n478) );
  XOR2_X2 U325 ( .A(n326), .B(n325), .Z(n579) );
  XNOR2_X1 U326 ( .A(n308), .B(KEYINPUT70), .ZN(n335) );
  XNOR2_X1 U327 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n308) );
  XNOR2_X1 U328 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U329 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U330 ( .A(n348), .B(n347), .ZN(n352) );
  XNOR2_X1 U331 ( .A(n408), .B(n388), .ZN(n389) );
  XNOR2_X1 U332 ( .A(n472), .B(KEYINPUT123), .ZN(n473) );
  XNOR2_X1 U333 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U334 ( .A(KEYINPUT81), .B(KEYINPUT17), .ZN(n382) );
  XNOR2_X1 U335 ( .A(n474), .B(n473), .ZN(n571) );
  XNOR2_X1 U336 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U337 ( .A(n383), .B(n382), .ZN(n385) );
  XOR2_X1 U338 ( .A(n393), .B(n392), .Z(n536) );
  XOR2_X1 U339 ( .A(n458), .B(KEYINPUT76), .Z(n566) );
  XNOR2_X1 U340 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U341 ( .A(n451), .B(G36GAT), .ZN(n452) );
  XNOR2_X1 U342 ( .A(n484), .B(n483), .ZN(G1349GAT) );
  XNOR2_X1 U343 ( .A(n453), .B(n452), .ZN(G1329GAT) );
  XOR2_X1 U344 ( .A(KEYINPUT68), .B(G22GAT), .Z(n292) );
  XNOR2_X1 U345 ( .A(G169GAT), .B(G141GAT), .ZN(n291) );
  XNOR2_X1 U346 ( .A(n292), .B(n291), .ZN(n296) );
  XOR2_X1 U347 ( .A(KEYINPUT29), .B(KEYINPUT69), .Z(n294) );
  XNOR2_X1 U348 ( .A(KEYINPUT30), .B(KEYINPUT66), .ZN(n293) );
  XNOR2_X1 U349 ( .A(n294), .B(n293), .ZN(n295) );
  XNOR2_X1 U350 ( .A(n296), .B(n295), .ZN(n307) );
  XOR2_X1 U351 ( .A(G197GAT), .B(G50GAT), .Z(n298) );
  XOR2_X1 U352 ( .A(G113GAT), .B(G15GAT), .Z(n386) );
  XOR2_X1 U353 ( .A(G8GAT), .B(G1GAT), .Z(n340) );
  XNOR2_X1 U354 ( .A(n386), .B(n340), .ZN(n297) );
  XNOR2_X1 U355 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U356 ( .A(n299), .B(G43GAT), .Z(n305) );
  XNOR2_X1 U357 ( .A(G29GAT), .B(KEYINPUT7), .ZN(n300) );
  XNOR2_X1 U358 ( .A(n300), .B(KEYINPUT8), .ZN(n354) );
  XOR2_X1 U359 ( .A(n354), .B(KEYINPUT67), .Z(n302) );
  NAND2_X1 U360 ( .A1(G229GAT), .A2(G233GAT), .ZN(n301) );
  XNOR2_X1 U361 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U362 ( .A(n303), .B(G36GAT), .ZN(n304) );
  XNOR2_X1 U363 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U364 ( .A(n307), .B(n306), .Z(n510) );
  INV_X1 U365 ( .A(n510), .ZN(n574) );
  XOR2_X1 U366 ( .A(G148GAT), .B(G78GAT), .Z(n361) );
  XNOR2_X1 U367 ( .A(n335), .B(n361), .ZN(n310) );
  AND2_X1 U368 ( .A1(G230GAT), .A2(G233GAT), .ZN(n309) );
  XNOR2_X1 U369 ( .A(n310), .B(n309), .ZN(n311) );
  XNOR2_X1 U370 ( .A(n311), .B(KEYINPUT31), .ZN(n313) );
  XOR2_X1 U371 ( .A(G204GAT), .B(G64GAT), .Z(n396) );
  XOR2_X1 U372 ( .A(n396), .B(KEYINPUT32), .Z(n312) );
  XNOR2_X1 U373 ( .A(n313), .B(n312), .ZN(n317) );
  XOR2_X1 U374 ( .A(KEYINPUT73), .B(KEYINPUT72), .Z(n315) );
  XNOR2_X1 U375 ( .A(KEYINPUT33), .B(KEYINPUT71), .ZN(n314) );
  XOR2_X1 U376 ( .A(n315), .B(n314), .Z(n316) );
  XNOR2_X1 U377 ( .A(n317), .B(n316), .ZN(n326) );
  XNOR2_X1 U378 ( .A(G71GAT), .B(G176GAT), .ZN(n318) );
  XNOR2_X1 U379 ( .A(n318), .B(G120GAT), .ZN(n380) );
  INV_X1 U380 ( .A(G92GAT), .ZN(n319) );
  NAND2_X1 U381 ( .A1(G85GAT), .A2(n319), .ZN(n322) );
  INV_X1 U382 ( .A(G85GAT), .ZN(n320) );
  NAND2_X1 U383 ( .A1(n320), .A2(G92GAT), .ZN(n321) );
  NAND2_X1 U384 ( .A1(n322), .A2(n321), .ZN(n324) );
  XNOR2_X1 U385 ( .A(G99GAT), .B(G106GAT), .ZN(n323) );
  XNOR2_X1 U386 ( .A(n324), .B(n323), .ZN(n348) );
  XNOR2_X1 U387 ( .A(n380), .B(n348), .ZN(n325) );
  INV_X1 U388 ( .A(n579), .ZN(n464) );
  NAND2_X1 U389 ( .A1(n574), .A2(n464), .ZN(n490) );
  XOR2_X1 U390 ( .A(KEYINPUT12), .B(G64GAT), .Z(n328) );
  XNOR2_X1 U391 ( .A(G15GAT), .B(G71GAT), .ZN(n327) );
  XNOR2_X1 U392 ( .A(n328), .B(n327), .ZN(n332) );
  XOR2_X1 U393 ( .A(KEYINPUT77), .B(KEYINPUT14), .Z(n330) );
  XNOR2_X1 U394 ( .A(KEYINPUT79), .B(KEYINPUT15), .ZN(n329) );
  XNOR2_X1 U395 ( .A(n330), .B(n329), .ZN(n331) );
  XNOR2_X1 U396 ( .A(n332), .B(n331), .ZN(n344) );
  XOR2_X1 U397 ( .A(G78GAT), .B(G211GAT), .Z(n334) );
  XNOR2_X1 U398 ( .A(G183GAT), .B(G127GAT), .ZN(n333) );
  XNOR2_X1 U399 ( .A(n334), .B(n333), .ZN(n339) );
  XOR2_X1 U400 ( .A(n335), .B(KEYINPUT78), .Z(n337) );
  NAND2_X1 U401 ( .A1(G231GAT), .A2(G233GAT), .ZN(n336) );
  XNOR2_X1 U402 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U403 ( .A(n339), .B(n338), .Z(n342) );
  XOR2_X1 U404 ( .A(G22GAT), .B(G155GAT), .Z(n360) );
  XNOR2_X1 U405 ( .A(n340), .B(n360), .ZN(n341) );
  XNOR2_X1 U406 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U407 ( .A(n344), .B(n343), .Z(n485) );
  INV_X1 U408 ( .A(n485), .ZN(n582) );
  NAND2_X1 U409 ( .A1(G232GAT), .A2(G233GAT), .ZN(n346) );
  INV_X1 U410 ( .A(KEYINPUT11), .ZN(n345) );
  XOR2_X1 U411 ( .A(KEYINPUT10), .B(KEYINPUT74), .Z(n350) );
  XNOR2_X1 U412 ( .A(KEYINPUT75), .B(KEYINPUT9), .ZN(n349) );
  XOR2_X1 U413 ( .A(n350), .B(n349), .Z(n351) );
  XNOR2_X1 U414 ( .A(n352), .B(n351), .ZN(n358) );
  XNOR2_X1 U415 ( .A(G43GAT), .B(G190GAT), .ZN(n353) );
  XNOR2_X1 U416 ( .A(n353), .B(G134GAT), .ZN(n381) );
  XNOR2_X1 U417 ( .A(n354), .B(n381), .ZN(n356) );
  XOR2_X1 U418 ( .A(G50GAT), .B(G162GAT), .Z(n364) );
  XOR2_X1 U419 ( .A(G36GAT), .B(G218GAT), .Z(n394) );
  XOR2_X1 U420 ( .A(n364), .B(n394), .Z(n355) );
  INV_X1 U421 ( .A(n359), .ZN(n458) );
  XNOR2_X1 U422 ( .A(KEYINPUT36), .B(n566), .ZN(n584) );
  XOR2_X1 U423 ( .A(n361), .B(n360), .Z(n363) );
  NAND2_X1 U424 ( .A1(G228GAT), .A2(G233GAT), .ZN(n362) );
  XNOR2_X1 U425 ( .A(n363), .B(n362), .ZN(n365) );
  XOR2_X1 U426 ( .A(n365), .B(n364), .Z(n373) );
  XOR2_X1 U427 ( .A(KEYINPUT23), .B(KEYINPUT83), .Z(n367) );
  XNOR2_X1 U428 ( .A(G218GAT), .B(G106GAT), .ZN(n366) );
  XNOR2_X1 U429 ( .A(n367), .B(n366), .ZN(n371) );
  XOR2_X1 U430 ( .A(KEYINPUT22), .B(KEYINPUT84), .Z(n369) );
  XNOR2_X1 U431 ( .A(G204GAT), .B(KEYINPUT24), .ZN(n368) );
  XNOR2_X1 U432 ( .A(n369), .B(n368), .ZN(n370) );
  XNOR2_X1 U433 ( .A(n371), .B(n370), .ZN(n372) );
  XNOR2_X1 U434 ( .A(n373), .B(n372), .ZN(n379) );
  XOR2_X1 U435 ( .A(G211GAT), .B(KEYINPUT21), .Z(n375) );
  XNOR2_X1 U436 ( .A(G197GAT), .B(KEYINPUT85), .ZN(n374) );
  XNOR2_X1 U437 ( .A(n375), .B(n374), .ZN(n395) );
  XOR2_X1 U438 ( .A(KEYINPUT2), .B(KEYINPUT86), .Z(n377) );
  XNOR2_X1 U439 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n376) );
  XNOR2_X1 U440 ( .A(n377), .B(n376), .ZN(n424) );
  XOR2_X1 U441 ( .A(n395), .B(n424), .Z(n378) );
  XNOR2_X1 U442 ( .A(n379), .B(n378), .ZN(n475) );
  XNOR2_X1 U443 ( .A(n381), .B(n380), .ZN(n393) );
  XOR2_X1 U444 ( .A(KEYINPUT0), .B(G127GAT), .Z(n420) );
  XNOR2_X1 U445 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n383) );
  XOR2_X1 U446 ( .A(G169GAT), .B(G183GAT), .Z(n384) );
  XNOR2_X1 U447 ( .A(n385), .B(n384), .ZN(n408) );
  XOR2_X1 U448 ( .A(KEYINPUT20), .B(G99GAT), .Z(n387) );
  XOR2_X1 U449 ( .A(n420), .B(n389), .Z(n391) );
  NAND2_X1 U450 ( .A1(G227GAT), .A2(G233GAT), .ZN(n390) );
  XNOR2_X1 U451 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U452 ( .A(n395), .B(n394), .ZN(n397) );
  XNOR2_X1 U453 ( .A(n397), .B(n396), .ZN(n401) );
  XOR2_X1 U454 ( .A(KEYINPUT92), .B(KEYINPUT93), .Z(n399) );
  NAND2_X1 U455 ( .A1(G226GAT), .A2(G233GAT), .ZN(n398) );
  XNOR2_X1 U456 ( .A(n399), .B(n398), .ZN(n400) );
  XOR2_X1 U457 ( .A(n401), .B(n400), .Z(n406) );
  XOR2_X1 U458 ( .A(G92GAT), .B(G176GAT), .Z(n403) );
  XNOR2_X1 U459 ( .A(G8GAT), .B(G190GAT), .ZN(n402) );
  XNOR2_X1 U460 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U461 ( .A(n404), .B(KEYINPUT91), .ZN(n405) );
  XNOR2_X1 U462 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U463 ( .A(n408), .B(n407), .ZN(n524) );
  NOR2_X1 U464 ( .A1(n527), .A2(n524), .ZN(n409) );
  XNOR2_X1 U465 ( .A(n409), .B(KEYINPUT96), .ZN(n410) );
  NOR2_X1 U466 ( .A1(n475), .A2(n410), .ZN(n411) );
  XNOR2_X1 U467 ( .A(KEYINPUT25), .B(n411), .ZN(n415) );
  XOR2_X1 U468 ( .A(KEYINPUT26), .B(KEYINPUT95), .Z(n413) );
  NAND2_X1 U469 ( .A1(n527), .A2(n475), .ZN(n412) );
  XNOR2_X1 U470 ( .A(n413), .B(n412), .ZN(n573) );
  XNOR2_X1 U471 ( .A(KEYINPUT27), .B(n524), .ZN(n441) );
  OR2_X1 U472 ( .A1(n573), .A2(n441), .ZN(n414) );
  AND2_X1 U473 ( .A1(n415), .A2(n414), .ZN(n416) );
  XNOR2_X1 U474 ( .A(n416), .B(KEYINPUT97), .ZN(n439) );
  XOR2_X1 U475 ( .A(G85GAT), .B(G162GAT), .Z(n418) );
  XNOR2_X1 U476 ( .A(G29GAT), .B(G134GAT), .ZN(n417) );
  XNOR2_X1 U477 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U478 ( .A(n420), .B(n419), .Z(n422) );
  NAND2_X1 U479 ( .A1(G225GAT), .A2(G233GAT), .ZN(n421) );
  XNOR2_X1 U480 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U481 ( .A(n423), .B(KEYINPUT88), .Z(n426) );
  XNOR2_X1 U482 ( .A(n424), .B(KEYINPUT89), .ZN(n425) );
  XNOR2_X1 U483 ( .A(n426), .B(n425), .ZN(n430) );
  XOR2_X1 U484 ( .A(G155GAT), .B(G148GAT), .Z(n428) );
  XNOR2_X1 U485 ( .A(G113GAT), .B(G120GAT), .ZN(n427) );
  XNOR2_X1 U486 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U487 ( .A(n430), .B(n429), .Z(n438) );
  XOR2_X1 U488 ( .A(KEYINPUT90), .B(KEYINPUT1), .Z(n432) );
  XNOR2_X1 U489 ( .A(KEYINPUT4), .B(KEYINPUT6), .ZN(n431) );
  XNOR2_X1 U490 ( .A(n432), .B(n431), .ZN(n436) );
  XOR2_X1 U491 ( .A(KEYINPUT5), .B(KEYINPUT87), .Z(n434) );
  XNOR2_X1 U492 ( .A(G1GAT), .B(G57GAT), .ZN(n433) );
  XNOR2_X1 U493 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U494 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U495 ( .A(n438), .B(n437), .ZN(n570) );
  NAND2_X1 U496 ( .A1(n439), .A2(n570), .ZN(n446) );
  XOR2_X1 U497 ( .A(KEYINPUT82), .B(n536), .Z(n444) );
  XOR2_X1 U498 ( .A(KEYINPUT28), .B(KEYINPUT65), .Z(n440) );
  XOR2_X1 U499 ( .A(n475), .B(n440), .Z(n531) );
  INV_X1 U500 ( .A(n531), .ZN(n539) );
  NOR2_X1 U501 ( .A1(n570), .A2(n441), .ZN(n442) );
  XOR2_X1 U502 ( .A(KEYINPUT94), .B(n442), .Z(n534) );
  NOR2_X1 U503 ( .A1(n539), .A2(n534), .ZN(n443) );
  NAND2_X1 U504 ( .A1(n444), .A2(n443), .ZN(n445) );
  NAND2_X1 U505 ( .A1(n446), .A2(n445), .ZN(n488) );
  NAND2_X1 U506 ( .A1(n584), .A2(n488), .ZN(n447) );
  NOR2_X1 U507 ( .A1(n582), .A2(n447), .ZN(n449) );
  XNOR2_X1 U508 ( .A(KEYINPUT37), .B(KEYINPUT102), .ZN(n448) );
  XNOR2_X1 U509 ( .A(n449), .B(n448), .ZN(n522) );
  NOR2_X1 U510 ( .A1(n490), .A2(n522), .ZN(n450) );
  XOR2_X1 U511 ( .A(KEYINPUT38), .B(n450), .Z(n508) );
  NOR2_X1 U512 ( .A1(n508), .A2(n524), .ZN(n453) );
  XNOR2_X1 U513 ( .A(KEYINPUT103), .B(KEYINPUT104), .ZN(n451) );
  XOR2_X1 U514 ( .A(KEYINPUT41), .B(n579), .Z(n454) );
  XOR2_X1 U515 ( .A(KEYINPUT107), .B(n454), .Z(n543) );
  XNOR2_X1 U516 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n471) );
  XOR2_X1 U517 ( .A(KEYINPUT113), .B(KEYINPUT47), .Z(n461) );
  XNOR2_X1 U518 ( .A(KEYINPUT46), .B(KEYINPUT112), .ZN(n456) );
  NAND2_X1 U519 ( .A1(n574), .A2(n454), .ZN(n455) );
  XNOR2_X1 U520 ( .A(n456), .B(n455), .ZN(n457) );
  AND2_X1 U521 ( .A1(n457), .A2(n485), .ZN(n459) );
  NAND2_X1 U522 ( .A1(n459), .A2(n458), .ZN(n460) );
  XNOR2_X1 U523 ( .A(n461), .B(n460), .ZN(n469) );
  NAND2_X1 U524 ( .A1(n582), .A2(n584), .ZN(n463) );
  XOR2_X1 U525 ( .A(KEYINPUT45), .B(KEYINPUT114), .Z(n462) );
  XNOR2_X1 U526 ( .A(n463), .B(n462), .ZN(n465) );
  NAND2_X1 U527 ( .A1(n465), .A2(n464), .ZN(n466) );
  XNOR2_X1 U528 ( .A(n466), .B(KEYINPUT115), .ZN(n467) );
  AND2_X1 U529 ( .A1(n510), .A2(n467), .ZN(n468) );
  NOR2_X1 U530 ( .A1(n469), .A2(n468), .ZN(n470) );
  XNOR2_X1 U531 ( .A(n471), .B(n470), .ZN(n535) );
  NOR2_X1 U532 ( .A1(n535), .A2(n524), .ZN(n474) );
  INV_X1 U533 ( .A(KEYINPUT54), .ZN(n472) );
  INV_X1 U534 ( .A(n475), .ZN(n476) );
  AND2_X1 U535 ( .A1(n570), .A2(n476), .ZN(n477) );
  XNOR2_X1 U536 ( .A(n478), .B(KEYINPUT55), .ZN(n479) );
  NOR2_X1 U537 ( .A1(n527), .A2(n479), .ZN(n480) );
  XNOR2_X1 U538 ( .A(KEYINPUT124), .B(n480), .ZN(n567) );
  NAND2_X1 U539 ( .A1(n543), .A2(n567), .ZN(n484) );
  XOR2_X1 U540 ( .A(G176GAT), .B(KEYINPUT125), .Z(n482) );
  XOR2_X1 U541 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n481) );
  NOR2_X1 U542 ( .A1(n566), .A2(n485), .ZN(n487) );
  XNOR2_X1 U543 ( .A(KEYINPUT80), .B(KEYINPUT16), .ZN(n486) );
  XNOR2_X1 U544 ( .A(n487), .B(n486), .ZN(n489) );
  NAND2_X1 U545 ( .A1(n489), .A2(n488), .ZN(n512) );
  OR2_X1 U546 ( .A1(n490), .A2(n512), .ZN(n499) );
  NOR2_X1 U547 ( .A1(n570), .A2(n499), .ZN(n492) );
  XNOR2_X1 U548 ( .A(KEYINPUT98), .B(KEYINPUT34), .ZN(n491) );
  XNOR2_X1 U549 ( .A(n492), .B(n491), .ZN(n493) );
  XOR2_X1 U550 ( .A(G1GAT), .B(n493), .Z(G1324GAT) );
  NOR2_X1 U551 ( .A1(n524), .A2(n499), .ZN(n495) );
  XNOR2_X1 U552 ( .A(KEYINPUT99), .B(KEYINPUT100), .ZN(n494) );
  XNOR2_X1 U553 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U554 ( .A(G8GAT), .B(n496), .ZN(G1325GAT) );
  NOR2_X1 U555 ( .A1(n527), .A2(n499), .ZN(n498) );
  XNOR2_X1 U556 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n497) );
  XNOR2_X1 U557 ( .A(n498), .B(n497), .ZN(G1326GAT) );
  NOR2_X1 U558 ( .A1(n531), .A2(n499), .ZN(n500) );
  XOR2_X1 U559 ( .A(G22GAT), .B(n500), .Z(G1327GAT) );
  NOR2_X1 U560 ( .A1(n570), .A2(n508), .ZN(n503) );
  XOR2_X1 U561 ( .A(G29GAT), .B(KEYINPUT101), .Z(n501) );
  XNOR2_X1 U562 ( .A(KEYINPUT39), .B(n501), .ZN(n502) );
  XNOR2_X1 U563 ( .A(n503), .B(n502), .ZN(G1328GAT) );
  XOR2_X1 U564 ( .A(KEYINPUT40), .B(KEYINPUT106), .Z(n505) );
  XNOR2_X1 U565 ( .A(G43GAT), .B(KEYINPUT105), .ZN(n504) );
  XNOR2_X1 U566 ( .A(n505), .B(n504), .ZN(n507) );
  NOR2_X1 U567 ( .A1(n527), .A2(n508), .ZN(n506) );
  XOR2_X1 U568 ( .A(n507), .B(n506), .Z(G1330GAT) );
  NOR2_X1 U569 ( .A1(n508), .A2(n531), .ZN(n509) );
  XOR2_X1 U570 ( .A(G50GAT), .B(n509), .Z(G1331GAT) );
  NAND2_X1 U571 ( .A1(n543), .A2(n510), .ZN(n511) );
  XNOR2_X1 U572 ( .A(n511), .B(KEYINPUT108), .ZN(n521) );
  NOR2_X1 U573 ( .A1(n521), .A2(n512), .ZN(n513) );
  XNOR2_X1 U574 ( .A(KEYINPUT109), .B(n513), .ZN(n518) );
  NOR2_X1 U575 ( .A1(n570), .A2(n518), .ZN(n514) );
  XOR2_X1 U576 ( .A(KEYINPUT42), .B(n514), .Z(n515) );
  XNOR2_X1 U577 ( .A(G57GAT), .B(n515), .ZN(G1332GAT) );
  NOR2_X1 U578 ( .A1(n524), .A2(n518), .ZN(n516) );
  XOR2_X1 U579 ( .A(G64GAT), .B(n516), .Z(G1333GAT) );
  NOR2_X1 U580 ( .A1(n527), .A2(n518), .ZN(n517) );
  XOR2_X1 U581 ( .A(G71GAT), .B(n517), .Z(G1334GAT) );
  NOR2_X1 U582 ( .A1(n531), .A2(n518), .ZN(n520) );
  XNOR2_X1 U583 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n519) );
  XNOR2_X1 U584 ( .A(n520), .B(n519), .ZN(G1335GAT) );
  OR2_X1 U585 ( .A1(n522), .A2(n521), .ZN(n530) );
  NOR2_X1 U586 ( .A1(n570), .A2(n530), .ZN(n523) );
  XOR2_X1 U587 ( .A(G85GAT), .B(n523), .Z(G1336GAT) );
  NOR2_X1 U588 ( .A1(n524), .A2(n530), .ZN(n525) );
  XOR2_X1 U589 ( .A(KEYINPUT110), .B(n525), .Z(n526) );
  XNOR2_X1 U590 ( .A(G92GAT), .B(n526), .ZN(G1337GAT) );
  NOR2_X1 U591 ( .A1(n527), .A2(n530), .ZN(n529) );
  XNOR2_X1 U592 ( .A(G99GAT), .B(KEYINPUT111), .ZN(n528) );
  XNOR2_X1 U593 ( .A(n529), .B(n528), .ZN(G1338GAT) );
  NOR2_X1 U594 ( .A1(n531), .A2(n530), .ZN(n532) );
  XOR2_X1 U595 ( .A(KEYINPUT44), .B(n532), .Z(n533) );
  XNOR2_X1 U596 ( .A(G106GAT), .B(n533), .ZN(G1339GAT) );
  XOR2_X1 U597 ( .A(KEYINPUT117), .B(KEYINPUT118), .Z(n541) );
  NOR2_X1 U598 ( .A1(n535), .A2(n534), .ZN(n551) );
  NAND2_X1 U599 ( .A1(n551), .A2(n536), .ZN(n537) );
  XNOR2_X1 U600 ( .A(KEYINPUT116), .B(n537), .ZN(n538) );
  NOR2_X1 U601 ( .A1(n539), .A2(n538), .ZN(n548) );
  NAND2_X1 U602 ( .A1(n548), .A2(n574), .ZN(n540) );
  XNOR2_X1 U603 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U604 ( .A(G113GAT), .B(n542), .ZN(G1340GAT) );
  XOR2_X1 U605 ( .A(G120GAT), .B(KEYINPUT49), .Z(n545) );
  NAND2_X1 U606 ( .A1(n548), .A2(n543), .ZN(n544) );
  XNOR2_X1 U607 ( .A(n545), .B(n544), .ZN(G1341GAT) );
  NAND2_X1 U608 ( .A1(n548), .A2(n582), .ZN(n546) );
  XNOR2_X1 U609 ( .A(n546), .B(KEYINPUT50), .ZN(n547) );
  XNOR2_X1 U610 ( .A(G127GAT), .B(n547), .ZN(G1342GAT) );
  XOR2_X1 U611 ( .A(G134GAT), .B(KEYINPUT51), .Z(n550) );
  NAND2_X1 U612 ( .A1(n548), .A2(n566), .ZN(n549) );
  XNOR2_X1 U613 ( .A(n550), .B(n549), .ZN(G1343GAT) );
  INV_X1 U614 ( .A(n551), .ZN(n552) );
  NOR2_X1 U615 ( .A1(n552), .A2(n573), .ZN(n561) );
  AND2_X1 U616 ( .A1(n574), .A2(n561), .ZN(n553) );
  XOR2_X1 U617 ( .A(G141GAT), .B(n553), .Z(G1344GAT) );
  XOR2_X1 U618 ( .A(KEYINPUT120), .B(KEYINPUT53), .Z(n555) );
  NAND2_X1 U619 ( .A1(n561), .A2(n454), .ZN(n554) );
  XNOR2_X1 U620 ( .A(n555), .B(n554), .ZN(n556) );
  XOR2_X1 U621 ( .A(n556), .B(KEYINPUT52), .Z(n558) );
  XNOR2_X1 U622 ( .A(G148GAT), .B(KEYINPUT119), .ZN(n557) );
  XNOR2_X1 U623 ( .A(n558), .B(n557), .ZN(G1345GAT) );
  XOR2_X1 U624 ( .A(G155GAT), .B(KEYINPUT121), .Z(n560) );
  NAND2_X1 U625 ( .A1(n561), .A2(n582), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n560), .B(n559), .ZN(G1346GAT) );
  NAND2_X1 U627 ( .A1(n359), .A2(n561), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n562), .B(KEYINPUT122), .ZN(n563) );
  XNOR2_X1 U629 ( .A(G162GAT), .B(n563), .ZN(G1347GAT) );
  NAND2_X1 U630 ( .A1(n574), .A2(n567), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n564), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U632 ( .A1(n567), .A2(n582), .ZN(n565) );
  XNOR2_X1 U633 ( .A(n565), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U634 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n568), .B(KEYINPUT58), .ZN(n569) );
  XNOR2_X1 U636 ( .A(G190GAT), .B(n569), .ZN(G1351GAT) );
  XNOR2_X1 U637 ( .A(KEYINPUT59), .B(KEYINPUT126), .ZN(n578) );
  XOR2_X1 U638 ( .A(G197GAT), .B(KEYINPUT60), .Z(n576) );
  NAND2_X1 U639 ( .A1(n571), .A2(n570), .ZN(n572) );
  NOR2_X1 U640 ( .A1(n573), .A2(n572), .ZN(n585) );
  NAND2_X1 U641 ( .A1(n585), .A2(n574), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(G1352GAT) );
  XOR2_X1 U644 ( .A(G204GAT), .B(KEYINPUT61), .Z(n581) );
  NAND2_X1 U645 ( .A1(n585), .A2(n579), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(G1353GAT) );
  NAND2_X1 U647 ( .A1(n585), .A2(n582), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n583), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U649 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n587) );
  NAND2_X1 U650 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U651 ( .A(n587), .B(n586), .ZN(n588) );
  XNOR2_X1 U652 ( .A(G218GAT), .B(n588), .ZN(G1355GAT) );
endmodule

