//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 0 1 1 1 1 0 1 0 1 0 1 0 0 1 1 1 1 1 1 0 0 1 0 0 1 1 1 0 0 1 0 0 1 0 1 0 0 1 1 1 0 0 0 1 0 1 1 1 0 0 0 1 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:44 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n449, new_n452, new_n453, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n546, new_n547, new_n548, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n567, new_n568, new_n569,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n617, new_n620, new_n622, new_n623, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n830, new_n831, new_n832, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1180, new_n1181, new_n1182;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT65), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT66), .B(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  INV_X1    g026(.A(G2106), .ZN(new_n452));
  NOR2_X1   g027(.A1(new_n449), .A2(new_n452), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT67), .ZN(G217));
  NOR4_X1   g029(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT2), .ZN(new_n456));
  NOR4_X1   g031(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(new_n457), .ZN(G261));
  INV_X1    g033(.A(G261), .ZN(G325));
  INV_X1    g034(.A(G567), .ZN(new_n460));
  OAI22_X1  g035(.A1(new_n456), .A2(new_n452), .B1(new_n460), .B2(new_n457), .ZN(new_n461));
  XNOR2_X1  g036(.A(new_n461), .B(KEYINPUT68), .ZN(G319));
  INV_X1    g037(.A(G125), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n463), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(KEYINPUT69), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT69), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n471), .A2(G113), .A3(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  OAI21_X1  g048(.A(G2105), .B1(new_n468), .B2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G2104), .ZN(new_n476));
  INV_X1    g051(.A(G101), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g053(.A(G2105), .B1(new_n466), .B2(new_n467), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n478), .B1(new_n479), .B2(G137), .ZN(new_n480));
  AND2_X1   g055(.A1(new_n474), .A2(new_n480), .ZN(G160));
  XNOR2_X1  g056(.A(KEYINPUT3), .B(G2104), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G2105), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(KEYINPUT70), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT70), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n482), .A2(new_n485), .A3(G2105), .ZN(new_n486));
  AND2_X1   g061(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G124), .ZN(new_n488));
  XNOR2_X1  g063(.A(new_n488), .B(KEYINPUT71), .ZN(new_n489));
  OAI21_X1  g064(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(G112), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n490), .B1(new_n491), .B2(G2105), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n492), .B1(G136), .B2(new_n479), .ZN(new_n493));
  AND2_X1   g068(.A1(new_n489), .A2(new_n493), .ZN(G162));
  AND2_X1   g069(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n495));
  NOR2_X1   g070(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n496));
  OAI211_X1 g071(.A(G126), .B(G2105), .C1(new_n495), .C2(new_n496), .ZN(new_n497));
  OR2_X1    g072(.A1(G102), .A2(G2105), .ZN(new_n498));
  INV_X1    g073(.A(G114), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(G2105), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n498), .A2(new_n500), .A3(G2104), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n497), .A2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(G138), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n503), .A2(G2105), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n504), .B1(new_n495), .B2(new_n496), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(KEYINPUT4), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT4), .ZN(new_n507));
  OAI211_X1 g082(.A(new_n504), .B(new_n507), .C1(new_n496), .C2(new_n495), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n502), .B1(new_n506), .B2(new_n508), .ZN(G164));
  INV_X1    g084(.A(G543), .ZN(new_n510));
  OR2_X1    g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G50), .ZN(new_n514));
  XNOR2_X1  g089(.A(KEYINPUT5), .B(G543), .ZN(new_n515));
  XNOR2_X1  g090(.A(KEYINPUT6), .B(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(G88), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n515), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n519));
  INV_X1    g094(.A(G651), .ZN(new_n520));
  OAI221_X1 g095(.A(new_n514), .B1(new_n517), .B2(new_n518), .C1(new_n519), .C2(new_n520), .ZN(G303));
  INV_X1    g096(.A(G303), .ZN(G166));
  NAND3_X1  g097(.A1(new_n515), .A2(G63), .A3(G651), .ZN(new_n523));
  XOR2_X1   g098(.A(new_n523), .B(KEYINPUT72), .Z(new_n524));
  NAND2_X1  g099(.A1(new_n513), .A2(G51), .ZN(new_n525));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  XNOR2_X1  g101(.A(new_n526), .B(KEYINPUT7), .ZN(new_n527));
  INV_X1    g102(.A(G89), .ZN(new_n528));
  OAI211_X1 g103(.A(new_n525), .B(new_n527), .C1(new_n528), .C2(new_n517), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n524), .A2(new_n529), .ZN(G168));
  INV_X1    g105(.A(G90), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n516), .A2(G543), .ZN(new_n532));
  INV_X1    g107(.A(G52), .ZN(new_n533));
  OAI22_X1  g108(.A1(new_n517), .A2(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n515), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n535), .A2(new_n520), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n534), .A2(new_n536), .ZN(G171));
  INV_X1    g112(.A(G81), .ZN(new_n538));
  XOR2_X1   g113(.A(KEYINPUT73), .B(G43), .Z(new_n539));
  OAI22_X1  g114(.A1(new_n517), .A2(new_n538), .B1(new_n532), .B2(new_n539), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n515), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n541), .A2(new_n520), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G860), .ZN(G153));
  NAND4_X1  g119(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g120(.A1(G1), .A2(G3), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT8), .ZN(new_n547));
  NAND4_X1  g122(.A1(G319), .A2(G483), .A3(G661), .A4(new_n547), .ZN(new_n548));
  XOR2_X1   g123(.A(new_n548), .B(KEYINPUT74), .Z(G188));
  NAND3_X1  g124(.A1(new_n516), .A2(G53), .A3(G543), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT9), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n550), .B(new_n551), .ZN(new_n552));
  AND2_X1   g127(.A1(new_n515), .A2(new_n516), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G91), .ZN(new_n554));
  NAND2_X1  g129(.A1(G78), .A2(G543), .ZN(new_n555));
  AND2_X1   g130(.A1(KEYINPUT5), .A2(G543), .ZN(new_n556));
  NOR2_X1   g131(.A1(KEYINPUT5), .A2(G543), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(G65), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n555), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G651), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n554), .A2(new_n561), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n552), .A2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(new_n563), .ZN(G299));
  INV_X1    g139(.A(G171), .ZN(G301));
  INV_X1    g140(.A(G168), .ZN(G286));
  NAND2_X1  g141(.A1(new_n513), .A2(G49), .ZN(new_n567));
  OAI21_X1  g142(.A(G651), .B1(new_n515), .B2(G74), .ZN(new_n568));
  INV_X1    g143(.A(G87), .ZN(new_n569));
  OAI211_X1 g144(.A(new_n567), .B(new_n568), .C1(new_n569), .C2(new_n517), .ZN(G288));
  NAND3_X1  g145(.A1(new_n553), .A2(KEYINPUT77), .A3(G86), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT77), .ZN(new_n572));
  INV_X1    g147(.A(G86), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n572), .B1(new_n517), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  OAI21_X1  g150(.A(G61), .B1(new_n556), .B2(new_n557), .ZN(new_n576));
  NAND2_X1  g151(.A1(G73), .A2(G543), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  AOI21_X1  g153(.A(KEYINPUT75), .B1(new_n578), .B2(G651), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT75), .ZN(new_n580));
  AOI211_X1 g155(.A(new_n580), .B(new_n520), .C1(new_n576), .C2(new_n577), .ZN(new_n581));
  OAI21_X1  g156(.A(KEYINPUT76), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n515), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n580), .B1(new_n583), .B2(new_n520), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT76), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n578), .A2(KEYINPUT75), .A3(G651), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n575), .B1(new_n582), .B2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT78), .ZN(new_n589));
  INV_X1    g164(.A(G48), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n532), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n513), .A2(KEYINPUT78), .A3(G48), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n588), .A2(new_n593), .ZN(G305));
  AOI22_X1  g169(.A1(new_n553), .A2(G85), .B1(G47), .B2(new_n513), .ZN(new_n595));
  XNOR2_X1  g170(.A(new_n595), .B(KEYINPUT79), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n515), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n597));
  OR2_X1    g172(.A1(new_n597), .A2(new_n520), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n596), .A2(new_n598), .ZN(G290));
  INV_X1    g174(.A(G868), .ZN(new_n600));
  NOR2_X1   g175(.A1(G171), .A2(new_n600), .ZN(new_n601));
  XNOR2_X1  g176(.A(new_n601), .B(KEYINPUT80), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT81), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n553), .A2(new_n603), .A3(G92), .ZN(new_n604));
  INV_X1    g179(.A(G92), .ZN(new_n605));
  OAI21_X1  g180(.A(KEYINPUT81), .B1(new_n517), .B2(new_n605), .ZN(new_n606));
  AOI21_X1  g181(.A(KEYINPUT10), .B1(new_n604), .B2(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(new_n607), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n604), .A2(KEYINPUT10), .A3(new_n606), .ZN(new_n609));
  NAND2_X1  g184(.A1(G79), .A2(G543), .ZN(new_n610));
  INV_X1    g185(.A(G66), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n558), .B2(new_n611), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n612), .A2(G651), .B1(G54), .B2(new_n513), .ZN(new_n613));
  AND3_X1   g188(.A1(new_n608), .A2(new_n609), .A3(new_n613), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n602), .B1(G868), .B2(new_n614), .ZN(G321));
  XNOR2_X1  g190(.A(G321), .B(KEYINPUT82), .ZN(G284));
  NAND2_X1  g191(.A1(G299), .A2(new_n600), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n617), .B1(G168), .B2(new_n600), .ZN(G280));
  XNOR2_X1  g193(.A(G280), .B(KEYINPUT83), .ZN(G297));
  INV_X1    g194(.A(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n614), .B1(new_n620), .B2(G860), .ZN(G148));
  NAND2_X1  g196(.A1(new_n614), .A2(new_n620), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n622), .A2(G868), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n623), .B1(G868), .B2(new_n543), .ZN(G323));
  XNOR2_X1  g199(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g200(.A1(new_n475), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(KEYINPUT12), .Z(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(KEYINPUT13), .Z(new_n628));
  INV_X1    g203(.A(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n487), .A2(G123), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n479), .A2(G135), .ZN(new_n631));
  NOR2_X1   g206(.A1(new_n475), .A2(G111), .ZN(new_n632));
  OAI21_X1  g207(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n633));
  OAI211_X1 g208(.A(new_n630), .B(new_n631), .C1(new_n632), .C2(new_n633), .ZN(new_n634));
  AOI22_X1  g209(.A1(G2100), .A2(new_n629), .B1(new_n634), .B2(G2096), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n634), .A2(G2096), .ZN(new_n636));
  OAI211_X1 g211(.A(new_n635), .B(new_n636), .C1(G2100), .C2(new_n629), .ZN(G156));
  XNOR2_X1  g212(.A(G2427), .B(G2438), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2430), .ZN(new_n639));
  XNOR2_X1  g214(.A(KEYINPUT15), .B(G2435), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n639), .A2(new_n640), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n641), .A2(new_n642), .A3(KEYINPUT14), .ZN(new_n643));
  XOR2_X1   g218(.A(G1341), .B(G1348), .Z(new_n644));
  XNOR2_X1  g219(.A(G2443), .B(G2446), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n643), .B(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(G2451), .B(G2454), .Z(new_n648));
  XNOR2_X1  g223(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  OR2_X1    g225(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n647), .A2(new_n650), .ZN(new_n652));
  AND3_X1   g227(.A1(new_n651), .A2(G14), .A3(new_n652), .ZN(G401));
  XOR2_X1   g228(.A(G2067), .B(G2678), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT85), .ZN(new_n655));
  XOR2_X1   g230(.A(G2072), .B(G2078), .Z(new_n656));
  XOR2_X1   g231(.A(G2084), .B(G2090), .Z(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  NOR3_X1   g233(.A1(new_n655), .A2(new_n656), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT18), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n655), .A2(new_n656), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n656), .B(KEYINPUT17), .ZN(new_n662));
  OAI211_X1 g237(.A(new_n661), .B(new_n658), .C1(new_n655), .C2(new_n662), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n662), .A2(new_n655), .A3(new_n657), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n660), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(G2096), .B(G2100), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(G227));
  XOR2_X1   g242(.A(G1971), .B(G1976), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT19), .ZN(new_n669));
  XOR2_X1   g244(.A(G1956), .B(G2474), .Z(new_n670));
  XOR2_X1   g245(.A(G1961), .B(G1966), .Z(new_n671));
  AND2_X1   g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  INV_X1    g248(.A(KEYINPUT20), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n670), .A2(new_n671), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n672), .A2(new_n676), .ZN(new_n677));
  MUX2_X1   g252(.A(new_n677), .B(new_n676), .S(new_n669), .Z(new_n678));
  NOR2_X1   g253(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT86), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n679), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1981), .B(G1986), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT87), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n682), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1991), .B(G1996), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(G229));
  INV_X1    g262(.A(G16), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n688), .A2(G5), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n689), .B1(G171), .B2(new_n688), .ZN(new_n690));
  XOR2_X1   g265(.A(new_n690), .B(KEYINPUT98), .Z(new_n691));
  INV_X1    g266(.A(G1961), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(G29), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n694), .A2(G32), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n479), .A2(G141), .ZN(new_n696));
  NAND3_X1  g271(.A1(new_n475), .A2(G105), .A3(G2104), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(KEYINPUT26), .ZN(new_n699));
  NAND3_X1  g274(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT96), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n698), .B1(new_n699), .B2(new_n701), .ZN(new_n702));
  OR2_X1    g277(.A1(new_n701), .A2(new_n699), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n487), .A2(G129), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n695), .B1(new_n707), .B2(new_n694), .ZN(new_n708));
  XNOR2_X1  g283(.A(KEYINPUT27), .B(G1996), .ZN(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n693), .B1(new_n708), .B2(new_n710), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n694), .A2(KEYINPUT88), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n694), .A2(KEYINPUT88), .ZN(new_n713));
  AND2_X1   g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT24), .B(G34), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT95), .ZN(new_n717));
  NAND2_X1  g292(.A1(G160), .A2(G29), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(G2084), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n721), .B(KEYINPUT99), .Z(new_n722));
  OR2_X1    g297(.A1(new_n708), .A2(new_n710), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n711), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n614), .A2(G16), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(G4), .B2(G16), .ZN(new_n726));
  INV_X1    g301(.A(G1348), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g303(.A(KEYINPUT31), .B(G11), .ZN(new_n729));
  INV_X1    g304(.A(KEYINPUT30), .ZN(new_n730));
  AND2_X1   g305(.A1(new_n730), .A2(G28), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n694), .B1(new_n730), .B2(G28), .ZN(new_n732));
  OAI221_X1 g307(.A(new_n729), .B1(new_n731), .B2(new_n732), .C1(new_n634), .C2(new_n714), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n714), .A2(G27), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT100), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n506), .A2(new_n508), .ZN(new_n736));
  INV_X1    g311(.A(new_n502), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(new_n714), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n735), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n733), .B1(new_n443), .B2(new_n740), .ZN(new_n741));
  OAI221_X1 g316(.A(new_n741), .B1(new_n443), .B2(new_n740), .C1(new_n720), .C2(new_n719), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n694), .A2(G33), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n475), .A2(G103), .A3(G2104), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT25), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n482), .A2(G127), .ZN(new_n746));
  NAND2_X1  g321(.A1(G115), .A2(G2104), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n475), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  AOI211_X1 g323(.A(new_n745), .B(new_n748), .C1(G139), .C2(new_n479), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n743), .B1(new_n749), .B2(new_n694), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(new_n442), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n688), .A2(G19), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT94), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(new_n543), .B2(new_n688), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(G1341), .ZN(new_n755));
  INV_X1    g330(.A(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n751), .A2(new_n756), .ZN(new_n757));
  NOR4_X1   g332(.A1(new_n724), .A2(new_n728), .A3(new_n742), .A4(new_n757), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n739), .A2(G35), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(G162), .B2(new_n739), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT29), .ZN(new_n761));
  INV_X1    g336(.A(G2090), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n761), .B(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n688), .A2(G21), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(G168), .B2(new_n688), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(KEYINPUT97), .Z(new_n766));
  NOR2_X1   g341(.A1(new_n766), .A2(G1966), .ZN(new_n767));
  AND2_X1   g342(.A1(new_n766), .A2(G1966), .ZN(new_n768));
  AOI211_X1 g343(.A(new_n767), .B(new_n768), .C1(new_n727), .C2(new_n726), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n688), .A2(G20), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT23), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(new_n563), .B2(new_n688), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(G1956), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n714), .A2(G26), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(KEYINPUT28), .Z(new_n775));
  NAND2_X1  g350(.A1(new_n487), .A2(G128), .ZN(new_n776));
  OAI21_X1  g351(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n777));
  INV_X1    g352(.A(G116), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n777), .B1(new_n778), .B2(G2105), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(G140), .B2(new_n479), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n776), .A2(new_n780), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n775), .B1(new_n781), .B2(G29), .ZN(new_n782));
  INV_X1    g357(.A(G2067), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  AOI211_X1 g359(.A(new_n773), .B(new_n784), .C1(new_n692), .C2(new_n691), .ZN(new_n785));
  NAND4_X1  g360(.A1(new_n758), .A2(new_n763), .A3(new_n769), .A4(new_n785), .ZN(new_n786));
  AND2_X1   g361(.A1(new_n688), .A2(G6), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(G305), .B2(G16), .ZN(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT32), .B(G1981), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(KEYINPUT90), .ZN(new_n791));
  OR2_X1    g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n790), .A2(new_n791), .ZN(new_n793));
  NOR2_X1   g368(.A1(G16), .A2(G22), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(G166), .B2(G16), .ZN(new_n795));
  XOR2_X1   g370(.A(KEYINPUT92), .B(G1971), .Z(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  MUX2_X1   g372(.A(G23), .B(G288), .S(G16), .Z(new_n798));
  XNOR2_X1  g373(.A(KEYINPUT33), .B(G1976), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT91), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n798), .B(new_n800), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n797), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n792), .A2(new_n793), .A3(new_n802), .ZN(new_n803));
  XNOR2_X1  g378(.A(KEYINPUT93), .B(KEYINPUT34), .ZN(new_n804));
  INV_X1    g379(.A(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  NAND4_X1  g381(.A1(new_n792), .A2(new_n793), .A3(new_n802), .A4(new_n804), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n688), .A2(G24), .ZN(new_n809));
  XOR2_X1   g384(.A(new_n809), .B(KEYINPUT89), .Z(new_n810));
  INV_X1    g385(.A(G290), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n810), .B1(new_n811), .B2(new_n688), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(G1986), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n739), .A2(G25), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n487), .A2(G119), .ZN(new_n815));
  OAI21_X1  g390(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n816));
  INV_X1    g391(.A(G107), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n816), .B1(new_n817), .B2(G2105), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n818), .B1(G131), .B2(new_n479), .ZN(new_n819));
  AND2_X1   g394(.A1(new_n815), .A2(new_n819), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n814), .B1(new_n820), .B2(new_n739), .ZN(new_n821));
  XOR2_X1   g396(.A(KEYINPUT35), .B(G1991), .Z(new_n822));
  XOR2_X1   g397(.A(new_n821), .B(new_n822), .Z(new_n823));
  NOR2_X1   g398(.A1(new_n813), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n808), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n825), .A2(KEYINPUT36), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT36), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n808), .A2(new_n827), .A3(new_n824), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n786), .B1(new_n826), .B2(new_n828), .ZN(G311));
  INV_X1    g404(.A(new_n786), .ZN(new_n830));
  INV_X1    g405(.A(new_n828), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n827), .B1(new_n808), .B2(new_n824), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n830), .B1(new_n831), .B2(new_n832), .ZN(G150));
  NAND2_X1  g408(.A1(new_n614), .A2(G559), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT38), .ZN(new_n835));
  INV_X1    g410(.A(G93), .ZN(new_n836));
  INV_X1    g411(.A(G55), .ZN(new_n837));
  OAI22_X1  g412(.A1(new_n517), .A2(new_n836), .B1(new_n532), .B2(new_n837), .ZN(new_n838));
  AOI22_X1  g413(.A1(new_n515), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n839), .A2(new_n520), .ZN(new_n840));
  OR2_X1    g415(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n841), .B1(new_n542), .B2(new_n540), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n838), .A2(new_n840), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n543), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n835), .B(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT39), .ZN(new_n847));
  AOI21_X1  g422(.A(G860), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n848), .B1(new_n847), .B2(new_n846), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n841), .A2(G860), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n850), .B(KEYINPUT37), .Z(new_n851));
  NAND2_X1  g426(.A1(new_n849), .A2(new_n851), .ZN(G145));
  AND2_X1   g427(.A1(new_n776), .A2(new_n780), .ZN(new_n853));
  AND2_X1   g428(.A1(new_n702), .A2(new_n703), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n853), .A2(new_n854), .A3(new_n705), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n781), .B1(new_n704), .B2(new_n706), .ZN(new_n856));
  AND3_X1   g431(.A1(new_n855), .A2(G164), .A3(new_n856), .ZN(new_n857));
  AOI21_X1  g432(.A(G164), .B1(new_n855), .B2(new_n856), .ZN(new_n858));
  OAI211_X1 g433(.A(KEYINPUT101), .B(new_n749), .C1(new_n857), .C2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n855), .A2(new_n856), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n860), .A2(new_n738), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n749), .A2(KEYINPUT101), .ZN(new_n862));
  OR2_X1    g437(.A1(new_n749), .A2(KEYINPUT101), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n855), .A2(G164), .A3(new_n856), .ZN(new_n864));
  NAND4_X1  g439(.A1(new_n861), .A2(new_n862), .A3(new_n863), .A4(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n859), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n487), .A2(G130), .ZN(new_n867));
  OAI21_X1  g442(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n868));
  INV_X1    g443(.A(G118), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n868), .B1(new_n869), .B2(G2105), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n870), .B1(G142), .B2(new_n479), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n867), .A2(new_n871), .ZN(new_n872));
  AND3_X1   g447(.A1(new_n815), .A2(KEYINPUT102), .A3(new_n819), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n627), .ZN(new_n875));
  AOI21_X1  g450(.A(KEYINPUT102), .B1(new_n815), .B2(new_n819), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n874), .A2(new_n875), .A3(new_n877), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n627), .B1(new_n873), .B2(new_n876), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n872), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n878), .A2(new_n879), .A3(new_n872), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n866), .A2(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n634), .B(G160), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(G162), .ZN(new_n886));
  NAND4_X1  g461(.A1(new_n859), .A2(new_n865), .A3(new_n881), .A4(new_n882), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n884), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(G37), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n886), .B1(new_n884), .B2(new_n887), .ZN(new_n891));
  OAI21_X1  g466(.A(KEYINPUT103), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n884), .A2(new_n887), .ZN(new_n893));
  INV_X1    g468(.A(new_n886), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT103), .ZN(new_n896));
  NAND4_X1  g471(.A1(new_n895), .A2(new_n896), .A3(new_n889), .A4(new_n888), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n892), .A2(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n892), .A2(new_n897), .A3(new_n899), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(G395));
  XNOR2_X1  g478(.A(G305), .B(G290), .ZN(new_n904));
  XNOR2_X1  g479(.A(G303), .B(G288), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n905), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n811), .A2(G305), .ZN(new_n908));
  AOI21_X1  g483(.A(G290), .B1(new_n593), .B2(new_n588), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n907), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n906), .A2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT107), .ZN(new_n912));
  OAI21_X1  g487(.A(KEYINPUT106), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  OR2_X1    g488(.A1(new_n913), .A2(KEYINPUT42), .ZN(new_n914));
  OAI211_X1 g489(.A(new_n913), .B(KEYINPUT42), .C1(KEYINPUT106), .C2(new_n911), .ZN(new_n915));
  INV_X1    g490(.A(new_n613), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n607), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(new_n609), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n918), .A2(G299), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n563), .B1(new_n917), .B2(new_n609), .ZN(new_n920));
  OAI21_X1  g495(.A(KEYINPUT41), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n614), .A2(new_n563), .ZN(new_n922));
  INV_X1    g497(.A(new_n920), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT41), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n922), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT105), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n921), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  OAI211_X1 g502(.A(KEYINPUT105), .B(KEYINPUT41), .C1(new_n919), .C2(new_n920), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n622), .B(new_n845), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n919), .A2(new_n920), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n931), .B1(new_n930), .B2(new_n932), .ZN(new_n933));
  AND3_X1   g508(.A1(new_n914), .A2(new_n915), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n933), .B1(new_n914), .B2(new_n915), .ZN(new_n935));
  OAI21_X1  g510(.A(G868), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n936), .B1(G868), .B2(new_n843), .ZN(G295));
  OAI21_X1  g512(.A(new_n936), .B1(G868), .B2(new_n843), .ZN(G331));
  NAND3_X1  g513(.A1(new_n842), .A2(G301), .A3(new_n844), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(G301), .B1(new_n842), .B2(new_n844), .ZN(new_n941));
  NOR3_X1   g516(.A1(new_n940), .A2(new_n941), .A3(G286), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n845), .A2(G171), .ZN(new_n943));
  AOI21_X1  g518(.A(G168), .B1(new_n943), .B2(new_n939), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n945), .A2(new_n927), .A3(new_n928), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n932), .B1(new_n942), .B2(new_n944), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n946), .A2(new_n911), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(new_n889), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n911), .B1(new_n946), .B2(new_n947), .ZN(new_n950));
  OAI21_X1  g525(.A(KEYINPUT43), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT44), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n921), .A2(new_n925), .A3(KEYINPUT108), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT108), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n932), .A2(new_n954), .A3(new_n924), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n945), .A2(new_n953), .A3(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(new_n947), .ZN(new_n957));
  INV_X1    g532(.A(new_n911), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT43), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n959), .A2(new_n960), .A3(new_n889), .A4(new_n948), .ZN(new_n961));
  AND3_X1   g536(.A1(new_n951), .A2(new_n952), .A3(new_n961), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n911), .B1(new_n956), .B2(new_n947), .ZN(new_n963));
  OAI21_X1  g538(.A(KEYINPUT43), .B1(new_n949), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(KEYINPUT109), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT109), .ZN(new_n966));
  OAI211_X1 g541(.A(new_n966), .B(KEYINPUT43), .C1(new_n949), .C2(new_n963), .ZN(new_n967));
  OR3_X1    g542(.A1(new_n949), .A2(KEYINPUT43), .A3(new_n950), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n965), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n962), .B1(new_n969), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g545(.A(KEYINPUT45), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n971), .B1(G164), .B2(G1384), .ZN(new_n972));
  INV_X1    g547(.A(G1384), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n738), .A2(KEYINPUT45), .A3(new_n973), .ZN(new_n974));
  AND3_X1   g549(.A1(new_n474), .A2(new_n480), .A3(G40), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n972), .A2(new_n974), .A3(new_n443), .A4(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT125), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(KEYINPUT53), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT53), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n976), .A2(new_n977), .A3(new_n980), .ZN(new_n981));
  OAI21_X1  g556(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT50), .ZN(new_n983));
  INV_X1    g558(.A(new_n508), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n507), .B1(new_n482), .B2(new_n504), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  OAI211_X1 g561(.A(new_n983), .B(new_n973), .C1(new_n986), .C2(new_n502), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n982), .A2(new_n975), .A3(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n988), .A2(new_n692), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n979), .A2(new_n981), .A3(new_n989), .ZN(new_n990));
  AOI21_X1  g565(.A(KEYINPUT126), .B1(new_n990), .B2(G171), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT54), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n990), .A2(G171), .ZN(new_n993));
  AOI22_X1  g568(.A1(new_n978), .A2(KEYINPUT53), .B1(new_n692), .B2(new_n988), .ZN(new_n994));
  AOI21_X1  g569(.A(G301), .B1(new_n994), .B2(new_n981), .ZN(new_n995));
  OAI22_X1  g570(.A1(new_n991), .A2(new_n992), .B1(new_n993), .B2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(new_n995), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n994), .A2(G301), .A3(new_n981), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n997), .A2(KEYINPUT126), .A3(KEYINPUT54), .A4(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n996), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(G1976), .ZN(new_n1001));
  NOR2_X1   g576(.A1(G288), .A2(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g577(.A(new_n1002), .B(KEYINPUT113), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n474), .A2(new_n480), .A3(G40), .ZN(new_n1004));
  NOR3_X1   g579(.A1(new_n1004), .A2(G164), .A3(G1384), .ZN(new_n1005));
  INV_X1    g580(.A(G8), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1003), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(KEYINPUT52), .ZN(new_n1009));
  AOI21_X1  g584(.A(KEYINPUT52), .B1(G288), .B2(new_n1001), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1003), .A2(new_n1007), .A3(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(G1981), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n579), .A2(new_n581), .ZN(new_n1014));
  XNOR2_X1  g589(.A(KEYINPUT114), .B(G86), .ZN(new_n1015));
  AOI22_X1  g590(.A1(new_n591), .A2(new_n592), .B1(new_n553), .B2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1013), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(G1981), .B1(new_n591), .B2(new_n592), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1017), .B1(new_n588), .B2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1007), .B1(new_n1019), .B2(KEYINPUT49), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n582), .A2(new_n587), .ZN(new_n1021));
  INV_X1    g596(.A(new_n575), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1021), .A2(new_n1022), .A3(new_n1018), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1017), .ZN(new_n1024));
  AND3_X1   g599(.A1(new_n1023), .A2(KEYINPUT49), .A3(new_n1024), .ZN(new_n1025));
  OAI21_X1  g600(.A(KEYINPUT115), .B1(new_n1020), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT49), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1019), .A2(KEYINPUT49), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT115), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1029), .A2(new_n1030), .A3(new_n1031), .A4(new_n1007), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1012), .B1(new_n1026), .B2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n972), .A2(new_n974), .A3(new_n975), .ZN(new_n1034));
  INV_X1    g609(.A(G1966), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n982), .A2(new_n987), .A3(new_n720), .A4(new_n975), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1036), .A2(G168), .A3(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(G8), .ZN(new_n1039));
  AOI21_X1  g614(.A(G168), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1040));
  OAI21_X1  g615(.A(KEYINPUT51), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT51), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1038), .A2(new_n1042), .A3(G8), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1041), .A2(new_n1043), .ZN(new_n1044));
  XNOR2_X1  g619(.A(KEYINPUT112), .B(KEYINPUT55), .ZN(new_n1045));
  NAND3_X1  g620(.A1(G303), .A2(G8), .A3(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1046), .ZN(new_n1047));
  AOI22_X1  g622(.A1(G303), .A2(G8), .B1(KEYINPUT112), .B2(KEYINPUT55), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n982), .A2(new_n987), .A3(new_n762), .A4(new_n975), .ZN(new_n1050));
  XNOR2_X1  g625(.A(KEYINPUT111), .B(G1971), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1034), .A2(new_n1051), .ZN(new_n1052));
  AOI211_X1 g627(.A(new_n1006), .B(new_n1049), .C1(new_n1050), .C2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n988), .A2(KEYINPUT116), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT116), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n982), .A2(new_n987), .A3(new_n1055), .A4(new_n975), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1054), .A2(new_n762), .A3(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(new_n1052), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(G8), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1053), .B1(new_n1059), .B2(new_n1049), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1033), .A2(new_n1044), .A3(new_n1060), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1000), .A2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g637(.A(G1384), .B1(new_n736), .B2(new_n737), .ZN(new_n1063));
  AND3_X1   g638(.A1(new_n1063), .A2(new_n975), .A3(new_n783), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1064), .B1(new_n988), .B2(new_n727), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1065), .A2(KEYINPUT123), .A3(KEYINPUT60), .ZN(new_n1066));
  AOI211_X1 g641(.A(KEYINPUT123), .B(new_n614), .C1(new_n1065), .C2(KEYINPUT60), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n975), .B1(new_n1063), .B2(new_n983), .ZN(new_n1068));
  NOR3_X1   g643(.A1(G164), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n727), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1064), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1070), .A2(KEYINPUT60), .A3(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT123), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n918), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1066), .B1(new_n1067), .B2(new_n1074), .ZN(new_n1075));
  OR2_X1    g650(.A1(new_n1065), .A2(KEYINPUT60), .ZN(new_n1076));
  AND3_X1   g651(.A1(new_n1075), .A2(KEYINPUT124), .A3(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(KEYINPUT124), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT61), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT118), .ZN(new_n1080));
  OAI211_X1 g655(.A(new_n1080), .B(KEYINPUT57), .C1(new_n552), .C2(new_n562), .ZN(new_n1081));
  XNOR2_X1  g656(.A(new_n550), .B(KEYINPUT9), .ZN(new_n1082));
  AOI22_X1  g657(.A1(G91), .A2(new_n553), .B1(new_n560), .B2(G651), .ZN(new_n1083));
  OR2_X1    g658(.A1(new_n1080), .A2(KEYINPUT57), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1080), .A2(KEYINPUT57), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1082), .A2(new_n1083), .A3(new_n1084), .A4(new_n1085), .ZN(new_n1086));
  AND2_X1   g661(.A1(new_n1081), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(G1956), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n988), .A2(new_n1088), .ZN(new_n1089));
  XNOR2_X1  g664(.A(KEYINPUT56), .B(G2072), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n972), .A2(new_n974), .A3(new_n975), .A4(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1087), .A2(new_n1089), .A3(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1087), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1079), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(G1996), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n972), .A2(new_n974), .A3(new_n1096), .A4(new_n975), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1063), .A2(new_n975), .ZN(new_n1098));
  XOR2_X1   g673(.A(KEYINPUT58), .B(G1341), .Z(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1097), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(new_n543), .ZN(new_n1102));
  XOR2_X1   g677(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n1103));
  XNOR2_X1  g678(.A(new_n1102), .B(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1094), .A2(KEYINPUT120), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT120), .ZN(new_n1106));
  AND3_X1   g681(.A1(new_n972), .A2(new_n974), .A3(new_n975), .ZN(new_n1107));
  AOI22_X1  g682(.A1(new_n1107), .A2(new_n1090), .B1(new_n988), .B2(new_n1088), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1106), .B1(new_n1108), .B2(new_n1087), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1105), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT122), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1092), .A2(new_n1111), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1087), .A2(new_n1089), .A3(KEYINPUT122), .A4(new_n1091), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1112), .A2(KEYINPUT61), .A3(new_n1113), .ZN(new_n1114));
  OAI211_X1 g689(.A(new_n1095), .B(new_n1104), .C1(new_n1110), .C2(new_n1114), .ZN(new_n1115));
  NOR3_X1   g690(.A1(new_n1077), .A2(new_n1078), .A3(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1110), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1065), .A2(new_n918), .ZN(new_n1118));
  XNOR2_X1  g693(.A(new_n1118), .B(KEYINPUT119), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1093), .B1(new_n1117), .B2(new_n1119), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1062), .B1(new_n1116), .B2(new_n1120), .ZN(new_n1121));
  AOI211_X1 g696(.A(new_n1006), .B(G286), .C1(new_n1036), .C2(new_n1037), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(KEYINPUT63), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1123), .A2(new_n1053), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1006), .B1(new_n1052), .B2(new_n1050), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1049), .ZN(new_n1126));
  OAI211_X1 g701(.A(new_n1033), .B(new_n1124), .C1(new_n1125), .C2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1033), .A2(new_n1060), .A3(new_n1122), .ZN(new_n1128));
  AND2_X1   g703(.A1(new_n1128), .A2(KEYINPUT117), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT117), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1033), .A2(new_n1060), .A3(new_n1130), .A4(new_n1122), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT63), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1127), .B1(new_n1129), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1033), .A2(new_n1053), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1023), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1026), .A2(new_n1032), .ZN(new_n1137));
  NOR2_X1   g712(.A1(G288), .A2(G1976), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1136), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1007), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1135), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  AND2_X1   g716(.A1(new_n1033), .A2(new_n1060), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT62), .ZN(new_n1143));
  AND3_X1   g718(.A1(new_n1041), .A2(new_n1143), .A3(new_n1043), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1143), .B1(new_n1041), .B2(new_n1043), .ZN(new_n1145));
  NOR3_X1   g720(.A1(new_n1144), .A2(new_n1145), .A3(new_n997), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1141), .B1(new_n1142), .B2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1121), .A2(new_n1134), .A3(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(G1986), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n972), .A2(new_n1004), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n811), .A2(new_n1149), .A3(new_n1150), .ZN(new_n1151));
  NAND3_X1  g726(.A1(G290), .A2(new_n1150), .A3(G1986), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  XNOR2_X1  g728(.A(new_n1153), .B(KEYINPUT110), .ZN(new_n1154));
  XNOR2_X1  g729(.A(new_n707), .B(G1996), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n781), .A2(G2067), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n853), .A2(new_n783), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1155), .A2(new_n1156), .A3(new_n1157), .ZN(new_n1158));
  XNOR2_X1  g733(.A(new_n820), .B(new_n822), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1150), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  AND2_X1   g735(.A1(new_n1154), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1148), .A2(new_n1161), .ZN(new_n1162));
  XNOR2_X1  g737(.A(new_n1151), .B(KEYINPUT48), .ZN(new_n1163));
  AND2_X1   g738(.A1(new_n1160), .A2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1157), .A2(new_n1156), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT46), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n707), .B1(new_n1166), .B2(G1996), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1150), .B1(new_n1165), .B2(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT127), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1150), .A2(new_n1096), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1169), .B1(new_n1170), .B2(new_n1166), .ZN(new_n1171));
  AOI211_X1 g746(.A(KEYINPUT127), .B(KEYINPUT46), .C1(new_n1150), .C2(new_n1096), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1168), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  XOR2_X1   g748(.A(new_n1173), .B(KEYINPUT47), .Z(new_n1174));
  NAND2_X1  g749(.A1(new_n820), .A2(new_n822), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1157), .B1(new_n1158), .B2(new_n1175), .ZN(new_n1176));
  AOI211_X1 g751(.A(new_n1164), .B(new_n1174), .C1(new_n1150), .C2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1162), .A2(new_n1177), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g753(.A(G319), .ZN(new_n1180));
  NOR4_X1   g754(.A1(G229), .A2(new_n1180), .A3(G401), .A4(G227), .ZN(new_n1181));
  NAND2_X1  g755(.A1(new_n951), .A2(new_n961), .ZN(new_n1182));
  AND3_X1   g756(.A1(new_n1181), .A2(new_n898), .A3(new_n1182), .ZN(G308));
  NAND3_X1  g757(.A1(new_n1181), .A2(new_n898), .A3(new_n1182), .ZN(G225));
endmodule


