

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584;

  XNOR2_X1 U322 ( .A(n444), .B(KEYINPUT115), .ZN(n523) );
  XNOR2_X1 U323 ( .A(n465), .B(n464), .ZN(n482) );
  INV_X1 U324 ( .A(KEYINPUT98), .ZN(n464) );
  INV_X1 U325 ( .A(n523), .ZN(n526) );
  XOR2_X1 U326 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n290) );
  XOR2_X1 U327 ( .A(n312), .B(n365), .Z(n291) );
  XOR2_X1 U328 ( .A(KEYINPUT40), .B(n495), .Z(n292) );
  AND2_X1 U329 ( .A1(n456), .A2(n455), .ZN(n457) );
  INV_X1 U330 ( .A(KEYINPUT112), .ZN(n416) );
  NOR2_X1 U331 ( .A1(n550), .A2(n531), .ZN(n427) );
  XNOR2_X1 U332 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U333 ( .A(n306), .B(n305), .ZN(n307) );
  AND2_X1 U334 ( .A1(n510), .A2(n487), .ZN(n488) );
  XNOR2_X1 U335 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U336 ( .A(n448), .B(n447), .ZN(G1341GAT) );
  XOR2_X1 U337 ( .A(KEYINPUT0), .B(G127GAT), .Z(n294) );
  XNOR2_X1 U338 ( .A(KEYINPUT81), .B(G120GAT), .ZN(n293) );
  XNOR2_X1 U339 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U340 ( .A(G113GAT), .B(n295), .Z(n344) );
  XNOR2_X1 U341 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n296) );
  XNOR2_X1 U342 ( .A(n290), .B(n296), .ZN(n312) );
  XOR2_X1 U343 ( .A(G190GAT), .B(G134GAT), .Z(n365) );
  XNOR2_X1 U344 ( .A(G43GAT), .B(G99GAT), .ZN(n297) );
  XNOR2_X1 U345 ( .A(n291), .B(n297), .ZN(n306) );
  XOR2_X1 U346 ( .A(KEYINPUT82), .B(KEYINPUT20), .Z(n299) );
  XNOR2_X1 U347 ( .A(G15GAT), .B(G71GAT), .ZN(n298) );
  XNOR2_X1 U348 ( .A(n299), .B(n298), .ZN(n300) );
  XNOR2_X1 U349 ( .A(n300), .B(KEYINPUT65), .ZN(n304) );
  XOR2_X1 U350 ( .A(G183GAT), .B(G176GAT), .Z(n302) );
  NAND2_X1 U351 ( .A1(G227GAT), .A2(G233GAT), .ZN(n301) );
  XOR2_X1 U352 ( .A(n302), .B(n301), .Z(n303) );
  XOR2_X1 U353 ( .A(n344), .B(n307), .Z(n455) );
  INV_X1 U354 ( .A(n455), .ZN(n550) );
  XOR2_X1 U355 ( .A(KEYINPUT76), .B(G211GAT), .Z(n309) );
  XNOR2_X1 U356 ( .A(G8GAT), .B(G183GAT), .ZN(n308) );
  XNOR2_X1 U357 ( .A(n309), .B(n308), .ZN(n352) );
  XOR2_X1 U358 ( .A(G176GAT), .B(G64GAT), .Z(n392) );
  XOR2_X1 U359 ( .A(n352), .B(n392), .Z(n311) );
  XNOR2_X1 U360 ( .A(G36GAT), .B(G92GAT), .ZN(n310) );
  XNOR2_X1 U361 ( .A(n311), .B(n310), .ZN(n316) );
  XOR2_X1 U362 ( .A(n312), .B(KEYINPUT94), .Z(n314) );
  NAND2_X1 U363 ( .A1(G226GAT), .A2(G233GAT), .ZN(n313) );
  XNOR2_X1 U364 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U365 ( .A(n316), .B(n315), .Z(n324) );
  XOR2_X1 U366 ( .A(KEYINPUT84), .B(G218GAT), .Z(n318) );
  XNOR2_X1 U367 ( .A(KEYINPUT85), .B(KEYINPUT21), .ZN(n317) );
  XNOR2_X1 U368 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U369 ( .A(G197GAT), .B(n319), .Z(n429) );
  XOR2_X1 U370 ( .A(KEYINPUT93), .B(KEYINPUT92), .Z(n321) );
  XNOR2_X1 U371 ( .A(G190GAT), .B(G204GAT), .ZN(n320) );
  XNOR2_X1 U372 ( .A(n321), .B(n320), .ZN(n322) );
  XNOR2_X1 U373 ( .A(n429), .B(n322), .ZN(n323) );
  XNOR2_X1 U374 ( .A(n324), .B(n323), .ZN(n543) );
  XNOR2_X1 U375 ( .A(n543), .B(KEYINPUT95), .ZN(n325) );
  XNOR2_X1 U376 ( .A(n325), .B(KEYINPUT27), .ZN(n453) );
  XOR2_X1 U377 ( .A(KEYINPUT88), .B(KEYINPUT1), .Z(n327) );
  XNOR2_X1 U378 ( .A(KEYINPUT89), .B(KEYINPUT6), .ZN(n326) );
  XNOR2_X1 U379 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U380 ( .A(KEYINPUT4), .B(n328), .Z(n330) );
  NAND2_X1 U381 ( .A1(G225GAT), .A2(G233GAT), .ZN(n329) );
  XNOR2_X1 U382 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U383 ( .A(n331), .B(KEYINPUT90), .Z(n336) );
  XOR2_X1 U384 ( .A(KEYINPUT2), .B(G162GAT), .Z(n333) );
  XNOR2_X1 U385 ( .A(KEYINPUT86), .B(G155GAT), .ZN(n332) );
  XNOR2_X1 U386 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U387 ( .A(KEYINPUT3), .B(n334), .Z(n428) );
  XNOR2_X1 U388 ( .A(n428), .B(KEYINPUT91), .ZN(n335) );
  XNOR2_X1 U389 ( .A(n336), .B(n335), .ZN(n340) );
  XOR2_X1 U390 ( .A(G85GAT), .B(G148GAT), .Z(n338) );
  XNOR2_X1 U391 ( .A(G29GAT), .B(G134GAT), .ZN(n337) );
  XNOR2_X1 U392 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U393 ( .A(n340), .B(n339), .Z(n346) );
  XOR2_X1 U394 ( .A(KEYINPUT5), .B(G57GAT), .Z(n342) );
  XNOR2_X1 U395 ( .A(G141GAT), .B(G1GAT), .ZN(n341) );
  XNOR2_X1 U396 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U397 ( .A(n344), .B(n343), .ZN(n345) );
  XNOR2_X1 U398 ( .A(n346), .B(n345), .ZN(n545) );
  XNOR2_X1 U399 ( .A(KEYINPUT113), .B(KEYINPUT48), .ZN(n425) );
  XOR2_X1 U400 ( .A(KEYINPUT71), .B(KEYINPUT13), .Z(n348) );
  XNOR2_X1 U401 ( .A(G71GAT), .B(G57GAT), .ZN(n347) );
  XNOR2_X1 U402 ( .A(n348), .B(n347), .ZN(n387) );
  XOR2_X1 U403 ( .A(G15GAT), .B(G1GAT), .Z(n402) );
  XOR2_X1 U404 ( .A(n387), .B(n402), .Z(n350) );
  NAND2_X1 U405 ( .A1(G231GAT), .A2(G233GAT), .ZN(n349) );
  XNOR2_X1 U406 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U407 ( .A(n351), .B(KEYINPUT78), .Z(n354) );
  XNOR2_X1 U408 ( .A(n352), .B(KEYINPUT12), .ZN(n353) );
  XNOR2_X1 U409 ( .A(n354), .B(n353), .ZN(n362) );
  XOR2_X1 U410 ( .A(G78GAT), .B(G155GAT), .Z(n356) );
  XNOR2_X1 U411 ( .A(G22GAT), .B(G127GAT), .ZN(n355) );
  XNOR2_X1 U412 ( .A(n356), .B(n355), .ZN(n360) );
  XOR2_X1 U413 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n358) );
  XNOR2_X1 U414 ( .A(G64GAT), .B(KEYINPUT77), .ZN(n357) );
  XNOR2_X1 U415 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U416 ( .A(n360), .B(n359), .Z(n361) );
  XOR2_X1 U417 ( .A(n362), .B(n361), .Z(n466) );
  INV_X1 U418 ( .A(n466), .ZN(n578) );
  XOR2_X1 U419 ( .A(KEYINPUT73), .B(G92GAT), .Z(n364) );
  XNOR2_X1 U420 ( .A(G99GAT), .B(G85GAT), .ZN(n363) );
  XNOR2_X1 U421 ( .A(n364), .B(n363), .ZN(n388) );
  XOR2_X1 U422 ( .A(n388), .B(G162GAT), .Z(n367) );
  XNOR2_X1 U423 ( .A(n365), .B(G218GAT), .ZN(n366) );
  XNOR2_X1 U424 ( .A(n367), .B(n366), .ZN(n371) );
  XOR2_X1 U425 ( .A(KEYINPUT75), .B(KEYINPUT9), .Z(n369) );
  NAND2_X1 U426 ( .A1(G232GAT), .A2(G233GAT), .ZN(n368) );
  XNOR2_X1 U427 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U428 ( .A(n371), .B(n370), .Z(n376) );
  XOR2_X1 U429 ( .A(KEYINPUT10), .B(KEYINPUT11), .Z(n373) );
  XNOR2_X1 U430 ( .A(G50GAT), .B(G106GAT), .ZN(n372) );
  XNOR2_X1 U431 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U432 ( .A(n374), .B(KEYINPUT64), .ZN(n375) );
  XNOR2_X1 U433 ( .A(n376), .B(n375), .ZN(n381) );
  XOR2_X1 U434 ( .A(KEYINPUT7), .B(G43GAT), .Z(n378) );
  XNOR2_X1 U435 ( .A(G36GAT), .B(G29GAT), .ZN(n377) );
  XNOR2_X1 U436 ( .A(n378), .B(n377), .ZN(n379) );
  XNOR2_X1 U437 ( .A(KEYINPUT8), .B(n379), .ZN(n412) );
  INV_X1 U438 ( .A(n412), .ZN(n380) );
  XOR2_X2 U439 ( .A(n381), .B(n380), .Z(n564) );
  XNOR2_X1 U440 ( .A(n564), .B(KEYINPUT36), .ZN(n581) );
  NOR2_X1 U441 ( .A1(n578), .A2(n581), .ZN(n383) );
  XNOR2_X1 U442 ( .A(KEYINPUT66), .B(KEYINPUT45), .ZN(n382) );
  XNOR2_X1 U443 ( .A(n383), .B(n382), .ZN(n400) );
  XOR2_X1 U444 ( .A(KEYINPUT33), .B(KEYINPUT32), .Z(n385) );
  NAND2_X1 U445 ( .A1(G230GAT), .A2(G233GAT), .ZN(n384) );
  XNOR2_X1 U446 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U447 ( .A(n386), .B(KEYINPUT74), .Z(n390) );
  XNOR2_X1 U448 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U449 ( .A(n390), .B(n389), .ZN(n391) );
  XOR2_X1 U450 ( .A(n391), .B(KEYINPUT31), .Z(n394) );
  XNOR2_X1 U451 ( .A(G120GAT), .B(n392), .ZN(n393) );
  XNOR2_X1 U452 ( .A(n394), .B(n393), .ZN(n399) );
  XOR2_X1 U453 ( .A(G148GAT), .B(G106GAT), .Z(n396) );
  XNOR2_X1 U454 ( .A(G204GAT), .B(G78GAT), .ZN(n395) );
  XNOR2_X1 U455 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U456 ( .A(KEYINPUT72), .B(n397), .ZN(n432) );
  INV_X1 U457 ( .A(n432), .ZN(n398) );
  XOR2_X1 U458 ( .A(n399), .B(n398), .Z(n575) );
  NAND2_X1 U459 ( .A1(n400), .A2(n575), .ZN(n415) );
  XNOR2_X1 U460 ( .A(G50GAT), .B(G22GAT), .ZN(n401) );
  XNOR2_X1 U461 ( .A(n401), .B(G141GAT), .ZN(n437) );
  XOR2_X1 U462 ( .A(n437), .B(n402), .Z(n404) );
  NAND2_X1 U463 ( .A1(G229GAT), .A2(G233GAT), .ZN(n403) );
  XNOR2_X1 U464 ( .A(n404), .B(n403), .ZN(n408) );
  XOR2_X1 U465 ( .A(KEYINPUT68), .B(KEYINPUT30), .Z(n406) );
  XNOR2_X1 U466 ( .A(KEYINPUT69), .B(KEYINPUT29), .ZN(n405) );
  XNOR2_X1 U467 ( .A(n406), .B(n405), .ZN(n407) );
  XOR2_X1 U468 ( .A(n408), .B(n407), .Z(n414) );
  XOR2_X1 U469 ( .A(G8GAT), .B(G197GAT), .Z(n410) );
  XNOR2_X1 U470 ( .A(G169GAT), .B(G113GAT), .ZN(n409) );
  XNOR2_X1 U471 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U472 ( .A(n412), .B(n411), .Z(n413) );
  XNOR2_X1 U473 ( .A(n414), .B(n413), .ZN(n572) );
  XOR2_X1 U474 ( .A(n572), .B(KEYINPUT70), .Z(n551) );
  NOR2_X1 U475 ( .A1(n415), .A2(n551), .ZN(n417) );
  XNOR2_X1 U476 ( .A(n417), .B(n416), .ZN(n423) );
  XOR2_X1 U477 ( .A(KEYINPUT111), .B(n578), .Z(n559) );
  NAND2_X1 U478 ( .A1(n564), .A2(n559), .ZN(n420) );
  XOR2_X1 U479 ( .A(KEYINPUT41), .B(n575), .Z(n536) );
  NOR2_X1 U480 ( .A1(n572), .A2(n536), .ZN(n418) );
  XNOR2_X1 U481 ( .A(n418), .B(KEYINPUT46), .ZN(n419) );
  NOR2_X1 U482 ( .A1(n420), .A2(n419), .ZN(n421) );
  XNOR2_X1 U483 ( .A(KEYINPUT47), .B(n421), .ZN(n422) );
  NAND2_X1 U484 ( .A1(n423), .A2(n422), .ZN(n424) );
  XNOR2_X1 U485 ( .A(n425), .B(n424), .ZN(n542) );
  NOR2_X1 U486 ( .A1(n545), .A2(n542), .ZN(n426) );
  NAND2_X1 U487 ( .A1(n453), .A2(n426), .ZN(n531) );
  XNOR2_X1 U488 ( .A(KEYINPUT114), .B(n427), .ZN(n443) );
  XNOR2_X1 U489 ( .A(n429), .B(n428), .ZN(n441) );
  XOR2_X1 U490 ( .A(KEYINPUT87), .B(KEYINPUT24), .Z(n431) );
  XNOR2_X1 U491 ( .A(KEYINPUT83), .B(G211GAT), .ZN(n430) );
  XNOR2_X1 U492 ( .A(n431), .B(n430), .ZN(n433) );
  XNOR2_X1 U493 ( .A(n433), .B(n432), .ZN(n439) );
  XOR2_X1 U494 ( .A(KEYINPUT22), .B(KEYINPUT23), .Z(n435) );
  NAND2_X1 U495 ( .A1(G228GAT), .A2(G233GAT), .ZN(n434) );
  XNOR2_X1 U496 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U497 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U498 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U499 ( .A(n441), .B(n440), .ZN(n547) );
  XNOR2_X1 U500 ( .A(n547), .B(KEYINPUT67), .ZN(n442) );
  XNOR2_X1 U501 ( .A(n442), .B(KEYINPUT28), .ZN(n517) );
  NAND2_X1 U502 ( .A1(n443), .A2(n517), .ZN(n444) );
  XNOR2_X1 U503 ( .A(n536), .B(KEYINPUT105), .ZN(n554) );
  NAND2_X1 U504 ( .A1(n523), .A2(n554), .ZN(n448) );
  XOR2_X1 U505 ( .A(KEYINPUT116), .B(KEYINPUT49), .Z(n446) );
  XOR2_X1 U506 ( .A(G120GAT), .B(KEYINPUT117), .Z(n445) );
  AND2_X1 U507 ( .A1(n551), .A2(n575), .ZN(n487) );
  NAND2_X1 U508 ( .A1(n517), .A2(n453), .ZN(n449) );
  NOR2_X1 U509 ( .A1(n455), .A2(n449), .ZN(n450) );
  NOR2_X1 U510 ( .A1(n545), .A2(n450), .ZN(n463) );
  XOR2_X1 U511 ( .A(KEYINPUT96), .B(KEYINPUT26), .Z(n452) );
  NAND2_X1 U512 ( .A1(n547), .A2(n550), .ZN(n451) );
  XNOR2_X1 U513 ( .A(n452), .B(n451), .ZN(n570) );
  NAND2_X1 U514 ( .A1(n453), .A2(n570), .ZN(n454) );
  NAND2_X1 U515 ( .A1(n545), .A2(n454), .ZN(n461) );
  INV_X1 U516 ( .A(n543), .ZN(n456) );
  XOR2_X1 U517 ( .A(KEYINPUT97), .B(n457), .Z(n458) );
  NOR2_X1 U518 ( .A1(n547), .A2(n458), .ZN(n459) );
  XOR2_X1 U519 ( .A(KEYINPUT25), .B(n459), .Z(n460) );
  NOR2_X1 U520 ( .A1(n461), .A2(n460), .ZN(n462) );
  NOR2_X1 U521 ( .A1(n463), .A2(n462), .ZN(n465) );
  XOR2_X1 U522 ( .A(KEYINPUT80), .B(KEYINPUT79), .Z(n468) );
  NAND2_X1 U523 ( .A1(n466), .A2(n564), .ZN(n467) );
  XNOR2_X1 U524 ( .A(n468), .B(n467), .ZN(n469) );
  XNOR2_X1 U525 ( .A(n469), .B(KEYINPUT16), .ZN(n470) );
  NOR2_X1 U526 ( .A1(n482), .A2(n470), .ZN(n499) );
  NAND2_X1 U527 ( .A1(n487), .A2(n499), .ZN(n479) );
  NOR2_X1 U528 ( .A1(n545), .A2(n479), .ZN(n472) );
  XNOR2_X1 U529 ( .A(KEYINPUT34), .B(KEYINPUT99), .ZN(n471) );
  XNOR2_X1 U530 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U531 ( .A(G1GAT), .B(n473), .ZN(G1324GAT) );
  NOR2_X1 U532 ( .A1(n543), .A2(n479), .ZN(n474) );
  XOR2_X1 U533 ( .A(G8GAT), .B(n474), .Z(G1325GAT) );
  NOR2_X1 U534 ( .A1(n479), .A2(n550), .ZN(n478) );
  XOR2_X1 U535 ( .A(KEYINPUT100), .B(KEYINPUT101), .Z(n476) );
  XNOR2_X1 U536 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n475) );
  XNOR2_X1 U537 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U538 ( .A(n478), .B(n477), .ZN(G1326GAT) );
  NOR2_X1 U539 ( .A1(n517), .A2(n479), .ZN(n480) );
  XOR2_X1 U540 ( .A(KEYINPUT102), .B(n480), .Z(n481) );
  XNOR2_X1 U541 ( .A(G22GAT), .B(n481), .ZN(G1327GAT) );
  XNOR2_X1 U542 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n491) );
  INV_X1 U543 ( .A(KEYINPUT38), .ZN(n489) );
  INV_X1 U544 ( .A(KEYINPUT37), .ZN(n486) );
  NOR2_X1 U545 ( .A1(n482), .A2(n581), .ZN(n483) );
  NAND2_X1 U546 ( .A1(n578), .A2(n483), .ZN(n484) );
  XNOR2_X1 U547 ( .A(n484), .B(KEYINPUT103), .ZN(n485) );
  XNOR2_X1 U548 ( .A(n486), .B(n485), .ZN(n510) );
  XNOR2_X1 U549 ( .A(n489), .B(n488), .ZN(n496) );
  NOR2_X1 U550 ( .A1(n545), .A2(n496), .ZN(n490) );
  XNOR2_X1 U551 ( .A(n491), .B(n490), .ZN(G1328GAT) );
  INV_X1 U552 ( .A(KEYINPUT104), .ZN(n493) );
  NOR2_X1 U553 ( .A1(n543), .A2(n496), .ZN(n492) );
  XNOR2_X1 U554 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U555 ( .A(G36GAT), .B(n494), .ZN(G1329GAT) );
  NOR2_X1 U556 ( .A1(n496), .A2(n550), .ZN(n495) );
  XNOR2_X1 U557 ( .A(G43GAT), .B(n292), .ZN(G1330GAT) );
  NOR2_X1 U558 ( .A1(n517), .A2(n496), .ZN(n497) );
  XOR2_X1 U559 ( .A(G50GAT), .B(n497), .Z(G1331GAT) );
  NAND2_X1 U560 ( .A1(n554), .A2(n572), .ZN(n498) );
  XOR2_X1 U561 ( .A(n498), .B(KEYINPUT106), .Z(n511) );
  NAND2_X1 U562 ( .A1(n499), .A2(n511), .ZN(n507) );
  NOR2_X1 U563 ( .A1(n545), .A2(n507), .ZN(n501) );
  XNOR2_X1 U564 ( .A(KEYINPUT107), .B(KEYINPUT42), .ZN(n500) );
  XNOR2_X1 U565 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U566 ( .A(G57GAT), .B(n502), .ZN(G1332GAT) );
  NOR2_X1 U567 ( .A1(n543), .A2(n507), .ZN(n504) );
  XNOR2_X1 U568 ( .A(KEYINPUT108), .B(KEYINPUT109), .ZN(n503) );
  XNOR2_X1 U569 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U570 ( .A(G64GAT), .B(n505), .ZN(G1333GAT) );
  NOR2_X1 U571 ( .A1(n550), .A2(n507), .ZN(n506) );
  XOR2_X1 U572 ( .A(G71GAT), .B(n506), .Z(G1334GAT) );
  NOR2_X1 U573 ( .A1(n517), .A2(n507), .ZN(n509) );
  XNOR2_X1 U574 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n508) );
  XNOR2_X1 U575 ( .A(n509), .B(n508), .ZN(G1335GAT) );
  NAND2_X1 U576 ( .A1(n511), .A2(n510), .ZN(n516) );
  NOR2_X1 U577 ( .A1(n545), .A2(n516), .ZN(n512) );
  XOR2_X1 U578 ( .A(KEYINPUT110), .B(n512), .Z(n513) );
  XNOR2_X1 U579 ( .A(G85GAT), .B(n513), .ZN(G1336GAT) );
  NOR2_X1 U580 ( .A1(n543), .A2(n516), .ZN(n514) );
  XOR2_X1 U581 ( .A(G92GAT), .B(n514), .Z(G1337GAT) );
  NOR2_X1 U582 ( .A1(n550), .A2(n516), .ZN(n515) );
  XOR2_X1 U583 ( .A(G99GAT), .B(n515), .Z(G1338GAT) );
  NOR2_X1 U584 ( .A1(n517), .A2(n516), .ZN(n518) );
  XOR2_X1 U585 ( .A(KEYINPUT44), .B(n518), .Z(n519) );
  XNOR2_X1 U586 ( .A(G106GAT), .B(n519), .ZN(G1339GAT) );
  NAND2_X1 U587 ( .A1(n551), .A2(n523), .ZN(n520) );
  XNOR2_X1 U588 ( .A(G113GAT), .B(n520), .ZN(G1340GAT) );
  XOR2_X1 U589 ( .A(KEYINPUT50), .B(KEYINPUT118), .Z(n522) );
  XNOR2_X1 U590 ( .A(G127GAT), .B(KEYINPUT119), .ZN(n521) );
  XNOR2_X1 U591 ( .A(n522), .B(n521), .ZN(n525) );
  NOR2_X1 U592 ( .A1(n559), .A2(n526), .ZN(n524) );
  XOR2_X1 U593 ( .A(n525), .B(n524), .Z(G1342GAT) );
  NOR2_X1 U594 ( .A1(n526), .A2(n564), .ZN(n530) );
  XOR2_X1 U595 ( .A(KEYINPUT120), .B(KEYINPUT51), .Z(n528) );
  XNOR2_X1 U596 ( .A(G134GAT), .B(KEYINPUT121), .ZN(n527) );
  XNOR2_X1 U597 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U598 ( .A(n530), .B(n529), .ZN(G1343GAT) );
  INV_X1 U599 ( .A(n531), .ZN(n532) );
  NAND2_X1 U600 ( .A1(n532), .A2(n570), .ZN(n540) );
  NOR2_X1 U601 ( .A1(n572), .A2(n540), .ZN(n533) );
  XOR2_X1 U602 ( .A(G141GAT), .B(n533), .Z(G1344GAT) );
  XOR2_X1 U603 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n535) );
  XNOR2_X1 U604 ( .A(G148GAT), .B(KEYINPUT122), .ZN(n534) );
  XNOR2_X1 U605 ( .A(n535), .B(n534), .ZN(n538) );
  NOR2_X1 U606 ( .A1(n536), .A2(n540), .ZN(n537) );
  XOR2_X1 U607 ( .A(n538), .B(n537), .Z(G1345GAT) );
  NOR2_X1 U608 ( .A1(n578), .A2(n540), .ZN(n539) );
  XOR2_X1 U609 ( .A(G155GAT), .B(n539), .Z(G1346GAT) );
  NOR2_X1 U610 ( .A1(n564), .A2(n540), .ZN(n541) );
  XOR2_X1 U611 ( .A(G162GAT), .B(n541), .Z(G1347GAT) );
  XOR2_X1 U612 ( .A(G169GAT), .B(KEYINPUT123), .Z(n553) );
  NOR2_X1 U613 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U614 ( .A(KEYINPUT54), .B(n544), .ZN(n546) );
  NAND2_X1 U615 ( .A1(n546), .A2(n545), .ZN(n569) );
  NOR2_X1 U616 ( .A1(n547), .A2(n569), .ZN(n548) );
  XNOR2_X1 U617 ( .A(n548), .B(KEYINPUT55), .ZN(n549) );
  NOR2_X1 U618 ( .A1(n550), .A2(n549), .ZN(n558) );
  NAND2_X1 U619 ( .A1(n558), .A2(n551), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n553), .B(n552), .ZN(G1348GAT) );
  XOR2_X1 U621 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n556) );
  NAND2_X1 U622 ( .A1(n558), .A2(n554), .ZN(n555) );
  XNOR2_X1 U623 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U624 ( .A(G176GAT), .B(n557), .ZN(G1349GAT) );
  INV_X1 U625 ( .A(n558), .ZN(n563) );
  NOR2_X1 U626 ( .A1(n559), .A2(n563), .ZN(n560) );
  XOR2_X1 U627 ( .A(G183GAT), .B(n560), .Z(G1350GAT) );
  XOR2_X1 U628 ( .A(KEYINPUT124), .B(KEYINPUT58), .Z(n562) );
  XNOR2_X1 U629 ( .A(G190GAT), .B(KEYINPUT125), .ZN(n561) );
  XNOR2_X1 U630 ( .A(n562), .B(n561), .ZN(n566) );
  NOR2_X1 U631 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U632 ( .A(n566), .B(n565), .Z(G1351GAT) );
  XOR2_X1 U633 ( .A(KEYINPUT59), .B(KEYINPUT126), .Z(n568) );
  XNOR2_X1 U634 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n567) );
  XNOR2_X1 U635 ( .A(n568), .B(n567), .ZN(n574) );
  INV_X1 U636 ( .A(n569), .ZN(n571) );
  NAND2_X1 U637 ( .A1(n571), .A2(n570), .ZN(n580) );
  NOR2_X1 U638 ( .A1(n572), .A2(n580), .ZN(n573) );
  XOR2_X1 U639 ( .A(n574), .B(n573), .Z(G1352GAT) );
  NOR2_X1 U640 ( .A1(n575), .A2(n580), .ZN(n577) );
  XNOR2_X1 U641 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1353GAT) );
  NOR2_X1 U643 ( .A1(n578), .A2(n580), .ZN(n579) );
  XOR2_X1 U644 ( .A(G211GAT), .B(n579), .Z(G1354GAT) );
  NOR2_X1 U645 ( .A1(n581), .A2(n580), .ZN(n583) );
  XNOR2_X1 U646 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U648 ( .A(G218GAT), .B(n584), .ZN(G1355GAT) );
endmodule

