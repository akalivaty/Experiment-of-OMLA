//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 1 0 0 1 1 1 1 1 0 1 1 1 0 0 0 0 1 0 1 0 1 1 0 1 1 0 1 1 1 0 1 1 0 0 0 0 1 1 1 1 0 0 0 0 1 0 0 1 1 0 0 0 0 0 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:58 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n714, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n738, new_n739, new_n741,
    new_n742, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n783, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n813, new_n814, new_n815, new_n816, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G134), .ZN(new_n190));
  OAI21_X1  g004(.A(KEYINPUT11), .B1(new_n190), .B2(G137), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT11), .ZN(new_n192));
  INV_X1    g006(.A(G137), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n192), .A2(new_n193), .A3(G134), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n191), .A2(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n190), .A2(G137), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  OAI21_X1  g011(.A(KEYINPUT68), .B1(new_n197), .B2(G131), .ZN(new_n198));
  AOI22_X1  g012(.A1(new_n191), .A2(new_n194), .B1(new_n190), .B2(G137), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT68), .ZN(new_n200));
  INV_X1    g014(.A(G131), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n199), .A2(new_n200), .A3(new_n201), .ZN(new_n202));
  AOI22_X1  g016(.A1(new_n198), .A2(new_n202), .B1(G131), .B2(new_n197), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n203), .A2(KEYINPUT85), .ZN(new_n204));
  XNOR2_X1  g018(.A(KEYINPUT65), .B(G146), .ZN(new_n205));
  OAI21_X1  g019(.A(KEYINPUT66), .B1(new_n205), .B2(G143), .ZN(new_n206));
  INV_X1    g020(.A(G146), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(KEYINPUT65), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT65), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G146), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT66), .ZN(new_n212));
  INV_X1    g026(.A(G143), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n211), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n207), .A2(G143), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n206), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n208), .A2(new_n210), .A3(G143), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(KEYINPUT1), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G128), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n216), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n213), .A2(G146), .ZN(new_n221));
  INV_X1    g035(.A(G128), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n222), .A2(KEYINPUT1), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n217), .A2(new_n221), .A3(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT70), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND4_X1  g040(.A1(new_n217), .A2(KEYINPUT70), .A3(new_n221), .A4(new_n223), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(G104), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(G107), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n229), .A2(G107), .ZN(new_n232));
  OAI21_X1  g046(.A(G101), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  OAI21_X1  g047(.A(KEYINPUT3), .B1(new_n229), .B2(G107), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT3), .ZN(new_n235));
  INV_X1    g049(.A(G107), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n235), .A2(new_n236), .A3(G104), .ZN(new_n237));
  INV_X1    g051(.A(G101), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n234), .A2(new_n237), .A3(new_n238), .A4(new_n230), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n233), .A2(new_n239), .ZN(new_n240));
  AND3_X1   g054(.A1(new_n220), .A2(new_n228), .A3(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n217), .A2(new_n221), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n215), .A2(KEYINPUT1), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G128), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n240), .B1(new_n228), .B2(new_n245), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n204), .B1(new_n241), .B2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT12), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  OAI211_X1 g063(.A(new_n204), .B(KEYINPUT12), .C1(new_n241), .C2(new_n246), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  AOI22_X1  g065(.A1(new_n216), .A2(new_n219), .B1(new_n226), .B2(new_n227), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n239), .A2(new_n233), .A3(KEYINPUT10), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT67), .ZN(new_n255));
  NAND2_X1  g069(.A1(KEYINPUT0), .A2(G128), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n256), .A2(KEYINPUT64), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT64), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n258), .B1(KEYINPUT0), .B2(G128), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n257), .B1(new_n256), .B2(new_n259), .ZN(new_n260));
  AOI21_X1  g074(.A(G143), .B1(new_n208), .B2(new_n210), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n215), .B1(new_n261), .B2(new_n212), .ZN(new_n262));
  NOR3_X1   g076(.A1(new_n205), .A2(KEYINPUT66), .A3(G143), .ZN(new_n263));
  OAI211_X1 g077(.A(new_n255), .B(new_n260), .C1(new_n262), .C2(new_n263), .ZN(new_n264));
  OR2_X1    g078(.A1(new_n242), .A2(new_n256), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n255), .B1(new_n216), .B2(new_n260), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n234), .A2(new_n237), .A3(new_n230), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(G101), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n270), .A2(KEYINPUT83), .A3(KEYINPUT4), .A4(new_n239), .ZN(new_n271));
  AND3_X1   g085(.A1(new_n270), .A2(KEYINPUT4), .A3(new_n239), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT4), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n269), .A2(new_n273), .A3(G101), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT83), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n271), .B1(new_n272), .B2(new_n276), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n254), .B1(new_n268), .B2(new_n277), .ZN(new_n278));
  OAI21_X1  g092(.A(KEYINPUT84), .B1(new_n246), .B2(KEYINPUT10), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT84), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT10), .ZN(new_n281));
  AOI22_X1  g095(.A1(new_n226), .A2(new_n227), .B1(new_n242), .B2(new_n244), .ZN(new_n282));
  OAI211_X1 g096(.A(new_n280), .B(new_n281), .C1(new_n282), .C2(new_n240), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n279), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n278), .A2(new_n284), .A3(new_n203), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n251), .A2(new_n285), .ZN(new_n286));
  AND2_X1   g100(.A1(KEYINPUT72), .A2(G953), .ZN(new_n287));
  NOR2_X1   g101(.A1(KEYINPUT72), .A2(G953), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(G227), .ZN(new_n290));
  XOR2_X1   g104(.A(G110), .B(G140), .Z(new_n291));
  XNOR2_X1  g105(.A(new_n290), .B(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n286), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n197), .A2(G131), .ZN(new_n294));
  AND3_X1   g108(.A1(new_n199), .A2(new_n200), .A3(new_n201), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n200), .B1(new_n199), .B2(new_n201), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n294), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  AND2_X1   g111(.A1(new_n279), .A2(new_n283), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n260), .B1(new_n262), .B2(new_n263), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(KEYINPUT67), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n300), .A2(new_n265), .A3(new_n264), .ZN(new_n301));
  INV_X1    g115(.A(new_n277), .ZN(new_n302));
  OAI22_X1  g116(.A1(new_n301), .A2(new_n302), .B1(new_n252), .B2(new_n253), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n297), .B1(new_n298), .B2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(new_n292), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n304), .A2(new_n305), .A3(new_n285), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n293), .A2(G469), .A3(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT86), .ZN(new_n308));
  INV_X1    g122(.A(G469), .ZN(new_n309));
  INV_X1    g123(.A(G902), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n307), .A2(new_n308), .A3(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n308), .B1(new_n307), .B2(new_n312), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n251), .A2(new_n285), .A3(new_n305), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n305), .B1(new_n304), .B2(new_n285), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT87), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n317), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  AND3_X1   g134(.A1(new_n278), .A2(new_n284), .A3(new_n203), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n203), .B1(new_n278), .B2(new_n284), .ZN(new_n322));
  OAI211_X1 g136(.A(new_n319), .B(new_n292), .C1(new_n321), .C2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  OAI211_X1 g138(.A(new_n309), .B(new_n310), .C1(new_n320), .C2(new_n324), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n189), .B1(new_n316), .B2(new_n325), .ZN(new_n326));
  OAI21_X1  g140(.A(G214), .B1(G237), .B2(G902), .ZN(new_n327));
  XOR2_X1   g141(.A(new_n327), .B(KEYINPUT88), .Z(new_n328));
  OAI21_X1  g142(.A(G125), .B1(new_n266), .B2(new_n267), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT89), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n301), .A2(KEYINPUT89), .A3(G125), .ZN(new_n332));
  INV_X1    g146(.A(G125), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n252), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n331), .A2(new_n332), .A3(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(G224), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n336), .A2(G953), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(new_n337), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n331), .A2(new_n332), .A3(new_n339), .A4(new_n334), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(G119), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(G116), .ZN(new_n343));
  OAI21_X1  g157(.A(G113), .B1(new_n343), .B2(KEYINPUT5), .ZN(new_n344));
  XNOR2_X1  g158(.A(G116), .B(G119), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n344), .B1(KEYINPUT5), .B2(new_n345), .ZN(new_n346));
  XOR2_X1   g160(.A(G116), .B(G119), .Z(new_n347));
  XNOR2_X1  g161(.A(KEYINPUT2), .B(G113), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NOR3_X1   g163(.A1(new_n346), .A2(new_n240), .A3(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT71), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n345), .A2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(new_n348), .ZN(new_n353));
  XNOR2_X1  g167(.A(new_n352), .B(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n350), .B1(new_n277), .B2(new_n355), .ZN(new_n356));
  XNOR2_X1  g170(.A(G110), .B(G122), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n357), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n270), .A2(KEYINPUT4), .A3(new_n239), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n360), .A2(new_n275), .A3(new_n274), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n354), .B1(new_n361), .B2(new_n271), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n359), .B1(new_n362), .B2(new_n350), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n358), .A2(new_n363), .A3(KEYINPUT6), .ZN(new_n364));
  OR3_X1    g178(.A1(new_n356), .A2(KEYINPUT6), .A3(new_n357), .ZN(new_n365));
  AND2_X1   g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n341), .A2(new_n366), .ZN(new_n367));
  AND2_X1   g181(.A1(new_n331), .A2(new_n332), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n368), .A2(KEYINPUT7), .A3(new_n339), .A4(new_n334), .ZN(new_n369));
  XOR2_X1   g183(.A(new_n357), .B(KEYINPUT8), .Z(new_n370));
  NOR2_X1   g184(.A1(new_n346), .A2(new_n349), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n370), .B1(new_n371), .B2(new_n240), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n345), .A2(KEYINPUT5), .ZN(new_n373));
  OR2_X1    g187(.A1(new_n373), .A2(KEYINPUT90), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n344), .B1(new_n373), .B2(KEYINPUT90), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n349), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n372), .B1(new_n240), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n358), .A2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT91), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n334), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n252), .A2(KEYINPUT91), .A3(new_n333), .ZN(new_n381));
  NAND4_X1  g195(.A1(new_n331), .A2(new_n332), .A3(new_n380), .A4(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT7), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n337), .B1(KEYINPUT92), .B2(new_n383), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n384), .B1(KEYINPUT92), .B2(new_n383), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n378), .B1(new_n382), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n369), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n367), .A2(new_n387), .A3(new_n310), .ZN(new_n388));
  OAI21_X1  g202(.A(G210), .B1(G237), .B2(G902), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  NAND4_X1  g205(.A1(new_n367), .A2(new_n387), .A3(new_n310), .A4(new_n389), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n328), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  OR2_X1    g207(.A1(KEYINPUT72), .A2(G953), .ZN(new_n394));
  INV_X1    g208(.A(G237), .ZN(new_n395));
  NAND2_X1  g209(.A1(KEYINPUT72), .A2(G953), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n394), .A2(G214), .A3(new_n395), .A4(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(new_n213), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n289), .A2(G143), .A3(G214), .A4(new_n395), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(G131), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT17), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n398), .A2(new_n399), .A3(new_n201), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n401), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT16), .ZN(new_n405));
  INV_X1    g219(.A(G140), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n405), .A2(new_n406), .A3(G125), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(G125), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n333), .A2(G140), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n407), .B1(new_n410), .B2(new_n405), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(new_n207), .ZN(new_n412));
  OAI211_X1 g226(.A(G146), .B(new_n407), .C1(new_n410), .C2(new_n405), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n412), .A2(KEYINPUT78), .A3(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT78), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n411), .A2(new_n415), .A3(new_n207), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n400), .A2(KEYINPUT17), .A3(G131), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n404), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT94), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n205), .A2(new_n408), .A3(new_n409), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n410), .A2(G146), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n420), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n421), .A2(new_n422), .A3(new_n420), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(KEYINPUT18), .A2(G131), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n398), .A2(new_n399), .A3(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n427), .ZN(new_n429));
  AOI21_X1  g243(.A(KEYINPUT93), .B1(new_n400), .B2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT93), .ZN(new_n431));
  AOI211_X1 g245(.A(new_n431), .B(new_n427), .C1(new_n398), .C2(new_n399), .ZN(new_n432));
  OAI211_X1 g246(.A(new_n426), .B(new_n428), .C1(new_n430), .C2(new_n432), .ZN(new_n433));
  XNOR2_X1  g247(.A(G113), .B(G122), .ZN(new_n434));
  XNOR2_X1  g248(.A(new_n434), .B(new_n229), .ZN(new_n435));
  XNOR2_X1  g249(.A(new_n435), .B(KEYINPUT95), .ZN(new_n436));
  AND3_X1   g250(.A1(new_n419), .A2(new_n433), .A3(new_n436), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n435), .B1(new_n419), .B2(new_n433), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n310), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(G475), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT20), .ZN(new_n441));
  INV_X1    g255(.A(new_n435), .ZN(new_n442));
  AND3_X1   g256(.A1(new_n421), .A2(new_n422), .A3(new_n420), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n428), .B1(new_n443), .B2(new_n423), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n400), .A2(new_n429), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(new_n431), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n400), .A2(KEYINPUT93), .A3(new_n429), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n444), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  XNOR2_X1  g262(.A(new_n410), .B(KEYINPUT19), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n413), .B1(new_n449), .B2(new_n211), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n450), .B1(new_n401), .B2(new_n403), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n442), .B1(new_n448), .B2(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n419), .A2(new_n433), .A3(new_n436), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NOR2_X1   g268(.A1(G475), .A2(G902), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n441), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(new_n455), .ZN(new_n457));
  AOI211_X1 g271(.A(KEYINPUT20), .B(new_n457), .C1(new_n452), .C2(new_n453), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n440), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT98), .ZN(new_n460));
  XNOR2_X1  g274(.A(G116), .B(G122), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(new_n236), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT14), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(G122), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n465), .A2(G116), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n236), .B1(new_n466), .B2(KEYINPUT14), .ZN(new_n467));
  AOI22_X1  g281(.A1(new_n460), .A2(new_n462), .B1(new_n464), .B2(new_n467), .ZN(new_n468));
  OAI21_X1  g282(.A(KEYINPUT96), .B1(new_n213), .B2(G128), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT96), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n470), .A2(new_n222), .A3(G143), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n213), .A2(G128), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n472), .A2(new_n190), .A3(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n190), .B1(new_n472), .B2(new_n473), .ZN(new_n476));
  OAI221_X1 g290(.A(new_n468), .B1(new_n460), .B2(new_n462), .C1(new_n475), .C2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT13), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n473), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n213), .A2(KEYINPUT13), .A3(G128), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n472), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  OR2_X1    g295(.A1(new_n461), .A2(new_n236), .ZN(new_n482));
  AOI22_X1  g296(.A1(new_n481), .A2(G134), .B1(new_n482), .B2(new_n462), .ZN(new_n483));
  AOI21_X1  g297(.A(KEYINPUT97), .B1(new_n483), .B2(new_n474), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n481), .A2(G134), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n482), .A2(new_n462), .ZN(new_n486));
  AND4_X1   g300(.A1(KEYINPUT97), .A2(new_n485), .A3(new_n486), .A4(new_n474), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n477), .B1(new_n484), .B2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(G217), .ZN(new_n489));
  NOR3_X1   g303(.A1(new_n187), .A2(new_n489), .A3(G953), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(new_n490), .ZN(new_n492));
  OAI211_X1 g306(.A(new_n477), .B(new_n492), .C1(new_n484), .C2(new_n487), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n491), .A2(new_n310), .A3(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(G478), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n495), .A2(KEYINPUT15), .ZN(new_n496));
  XNOR2_X1  g310(.A(new_n494), .B(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(G952), .ZN(new_n498));
  AOI211_X1 g312(.A(G953), .B(new_n498), .C1(G234), .C2(G237), .ZN(new_n499));
  AOI211_X1 g313(.A(new_n310), .B(new_n289), .C1(G234), .C2(G237), .ZN(new_n500));
  XNOR2_X1  g314(.A(KEYINPUT21), .B(G898), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n499), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NOR3_X1   g316(.A1(new_n459), .A2(new_n497), .A3(new_n502), .ZN(new_n503));
  AND2_X1   g317(.A1(new_n393), .A2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT32), .ZN(new_n505));
  XNOR2_X1  g319(.A(KEYINPUT26), .B(G101), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n289), .A2(G210), .A3(new_n395), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(KEYINPUT27), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n508), .A2(KEYINPUT27), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n507), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(new_n511), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n513), .A2(new_n509), .A3(new_n506), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n220), .A2(new_n228), .ZN(new_n517));
  OR2_X1    g331(.A1(new_n196), .A2(KEYINPUT69), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n193), .A2(G134), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n196), .A2(KEYINPUT69), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n518), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  AOI22_X1  g335(.A1(new_n198), .A2(new_n202), .B1(G131), .B2(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n355), .B1(new_n517), .B2(new_n522), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n300), .A2(new_n297), .A3(new_n265), .A4(new_n264), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n517), .A2(new_n522), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n354), .B1(new_n524), .B2(new_n527), .ZN(new_n528));
  OAI21_X1  g342(.A(KEYINPUT28), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT28), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n525), .A2(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n516), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT31), .ZN(new_n533));
  AOI21_X1  g347(.A(KEYINPUT73), .B1(new_n525), .B2(new_n516), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT73), .ZN(new_n535));
  AOI211_X1 g349(.A(new_n535), .B(new_n515), .C1(new_n523), .C2(new_n524), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n524), .A2(new_n527), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(KEYINPUT30), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT30), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n524), .A2(new_n527), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n354), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n533), .B1(new_n537), .B2(new_n542), .ZN(new_n543));
  NOR3_X1   g357(.A1(new_n266), .A2(new_n203), .A3(new_n267), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n521), .A2(G131), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n545), .B1(new_n295), .B2(new_n296), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n354), .B1(new_n252), .B2(new_n546), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n516), .B1(new_n544), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(new_n535), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n525), .A2(KEYINPUT73), .A3(new_n516), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(new_n541), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n540), .B1(new_n524), .B2(new_n527), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n355), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n551), .A2(KEYINPUT31), .A3(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n532), .B1(new_n543), .B2(new_n555), .ZN(new_n556));
  NOR2_X1   g370(.A1(G472), .A2(G902), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n505), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT75), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n558), .A2(new_n505), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n560), .B1(new_n556), .B2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(new_n532), .ZN(new_n564));
  NOR3_X1   g378(.A1(new_n537), .A2(new_n533), .A3(new_n542), .ZN(new_n565));
  AOI21_X1  g379(.A(KEYINPUT31), .B1(new_n551), .B2(new_n554), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n564), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n567), .A2(KEYINPUT75), .A3(new_n561), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT74), .ZN(new_n569));
  AOI22_X1  g383(.A1(new_n538), .A2(new_n355), .B1(new_n524), .B2(new_n523), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n569), .B1(new_n570), .B2(new_n530), .ZN(new_n571));
  OAI211_X1 g385(.A(KEYINPUT74), .B(KEYINPUT28), .C1(new_n526), .C2(new_n528), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT29), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n515), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n571), .A2(new_n531), .A3(new_n572), .A4(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n529), .A2(new_n531), .A3(new_n516), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(new_n573), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n516), .B1(new_n554), .B2(new_n525), .ZN(new_n578));
  OAI211_X1 g392(.A(new_n575), .B(new_n310), .C1(new_n577), .C2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(G472), .ZN(new_n580));
  NAND4_X1  g394(.A1(new_n559), .A2(new_n563), .A3(new_n568), .A4(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n489), .B1(G234), .B2(new_n310), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n222), .A2(G119), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n342), .A2(G128), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(G110), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(KEYINPUT24), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT24), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(G110), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT76), .ZN(new_n591));
  AND3_X1   g405(.A1(new_n588), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n591), .B1(new_n588), .B2(new_n590), .ZN(new_n593));
  OAI211_X1 g407(.A(KEYINPUT79), .B(new_n586), .C1(new_n592), .C2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT23), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n595), .B1(new_n342), .B2(G128), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n222), .A2(KEYINPUT23), .A3(G119), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n596), .A2(new_n597), .A3(new_n585), .ZN(new_n598));
  OR2_X1    g412(.A1(new_n598), .A2(G110), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n594), .A2(new_n599), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n589), .A2(G110), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n587), .A2(KEYINPUT24), .ZN(new_n602));
  OAI21_X1  g416(.A(KEYINPUT76), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n588), .A2(new_n590), .A3(new_n591), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  AOI21_X1  g419(.A(KEYINPUT79), .B1(new_n605), .B2(new_n586), .ZN(new_n606));
  OAI21_X1  g420(.A(KEYINPUT80), .B1(new_n600), .B2(new_n606), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n586), .B1(new_n592), .B2(new_n593), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT79), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT80), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n610), .A2(new_n611), .A3(new_n599), .A4(new_n594), .ZN(new_n612));
  AND2_X1   g426(.A1(new_n413), .A2(new_n421), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n607), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT82), .ZN(new_n615));
  OR2_X1    g429(.A1(new_n605), .A2(new_n586), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT77), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n587), .B1(new_n598), .B2(new_n617), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n618), .B1(new_n617), .B2(new_n598), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n414), .A2(new_n616), .A3(new_n619), .A4(new_n416), .ZN(new_n620));
  AND3_X1   g434(.A1(new_n614), .A2(new_n615), .A3(new_n620), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n615), .B1(new_n614), .B2(new_n620), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n289), .A2(G221), .A3(G234), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n623), .B(KEYINPUT81), .ZN(new_n624));
  XNOR2_X1  g438(.A(KEYINPUT22), .B(G137), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n624), .B(new_n625), .ZN(new_n626));
  NOR3_X1   g440(.A1(new_n621), .A2(new_n622), .A3(new_n626), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n626), .A2(new_n614), .A3(new_n615), .A4(new_n620), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n310), .B1(new_n627), .B2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT25), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n614), .A2(new_n620), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(KEYINPUT82), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n614), .A2(new_n615), .A3(new_n620), .ZN(new_n635));
  INV_X1    g449(.A(new_n626), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n634), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(new_n628), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n638), .A2(KEYINPUT25), .A3(new_n310), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n583), .B1(new_n632), .B2(new_n639), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n582), .A2(G902), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n638), .A2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n326), .A2(new_n504), .A3(new_n581), .A4(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(G101), .ZN(G3));
  OAI21_X1  g460(.A(G472), .B1(new_n556), .B2(G902), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n567), .A2(new_n557), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  AOI21_X1  g463(.A(KEYINPUT25), .B1(new_n638), .B2(new_n310), .ZN(new_n650));
  AOI211_X1 g464(.A(new_n631), .B(G902), .C1(new_n637), .C2(new_n628), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n582), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(new_n642), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n649), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n326), .A2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(new_n327), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n656), .B1(new_n391), .B2(new_n392), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n494), .A2(new_n495), .ZN(new_n658));
  INV_X1    g472(.A(KEYINPUT33), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n491), .A2(new_n659), .A3(new_n493), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT99), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n491), .A2(KEYINPUT99), .A3(new_n659), .A4(new_n493), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n490), .A2(KEYINPUT100), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n659), .B1(new_n488), .B2(new_n664), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n665), .B1(new_n488), .B2(new_n664), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n662), .A2(new_n663), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n310), .A2(G478), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n658), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(new_n459), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n670), .A2(new_n502), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n657), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n655), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(KEYINPUT34), .B(G104), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(G6));
  NAND2_X1  g489(.A1(new_n391), .A2(new_n392), .ZN(new_n676));
  OAI211_X1 g490(.A(new_n497), .B(new_n440), .C1(new_n456), .C2(new_n458), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n677), .A2(new_n502), .ZN(new_n678));
  AND3_X1   g492(.A1(new_n676), .A2(new_n327), .A3(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n326), .A2(new_n654), .A3(new_n679), .ZN(new_n680));
  XOR2_X1   g494(.A(KEYINPUT35), .B(G107), .Z(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(G9));
  NOR2_X1   g496(.A1(new_n626), .A2(KEYINPUT36), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(new_n633), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(new_n641), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n652), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n686), .A2(new_n647), .A3(new_n648), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n326), .A2(new_n504), .A3(new_n688), .ZN(new_n689));
  XOR2_X1   g503(.A(KEYINPUT37), .B(G110), .Z(new_n690));
  XNOR2_X1  g504(.A(new_n689), .B(new_n690), .ZN(G12));
  INV_X1    g505(.A(G900), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n499), .B1(new_n500), .B2(new_n692), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n677), .A2(new_n693), .ZN(new_n694));
  AND3_X1   g508(.A1(new_n657), .A2(new_n686), .A3(new_n694), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n695), .A2(new_n326), .A3(new_n581), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G128), .ZN(G30));
  XOR2_X1   g511(.A(new_n693), .B(KEYINPUT39), .Z(new_n698));
  NAND2_X1  g512(.A1(new_n326), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(KEYINPUT40), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT40), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n326), .A2(new_n701), .A3(new_n698), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n537), .A2(new_n542), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n570), .A2(new_n516), .ZN(new_n704));
  OAI21_X1  g518(.A(new_n310), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(G472), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n559), .A2(new_n563), .A3(new_n568), .A4(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(new_n686), .ZN(new_n708));
  AND2_X1   g522(.A1(new_n459), .A2(new_n497), .ZN(new_n709));
  AND4_X1   g523(.A1(new_n327), .A2(new_n707), .A3(new_n708), .A4(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n676), .B(KEYINPUT38), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n700), .A2(new_n702), .A3(new_n710), .A4(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G143), .ZN(G45));
  INV_X1    g527(.A(new_n693), .ZN(new_n714));
  AND3_X1   g528(.A1(new_n669), .A2(new_n459), .A3(new_n714), .ZN(new_n715));
  AND4_X1   g529(.A1(new_n676), .A2(new_n686), .A3(new_n715), .A4(new_n327), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n326), .A2(new_n716), .A3(new_n581), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G146), .ZN(G48));
  INV_X1    g532(.A(KEYINPUT101), .ZN(new_n719));
  INV_X1    g533(.A(new_n325), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n292), .B1(new_n321), .B2(new_n322), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(KEYINPUT87), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n722), .A2(new_n323), .A3(new_n317), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n309), .B1(new_n723), .B2(new_n310), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n720), .A2(new_n724), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n725), .A2(new_n188), .A3(new_n657), .A4(new_n671), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n581), .A2(new_n644), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n719), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  AND2_X1   g542(.A1(new_n581), .A2(new_n644), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n310), .B1(new_n320), .B2(new_n324), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(G469), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n731), .A2(new_n188), .A3(new_n325), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n732), .A2(new_n672), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n729), .A2(new_n733), .A3(KEYINPUT101), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n728), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(KEYINPUT41), .B(G113), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n735), .B(new_n736), .ZN(G15));
  NOR3_X1   g551(.A1(new_n720), .A2(new_n724), .A3(new_n189), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n738), .A2(new_n679), .A3(new_n581), .A4(new_n644), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G116), .ZN(G18));
  AND2_X1   g554(.A1(new_n686), .A2(new_n503), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n738), .A2(new_n581), .A3(new_n657), .A4(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G119), .ZN(G21));
  NAND2_X1  g557(.A1(new_n543), .A2(new_n555), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n571), .A2(new_n531), .A3(new_n572), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n745), .A2(new_n515), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(new_n557), .ZN(new_n748));
  AND3_X1   g562(.A1(new_n644), .A2(new_n647), .A3(new_n748), .ZN(new_n749));
  AND3_X1   g563(.A1(new_n676), .A2(new_n327), .A3(new_n709), .ZN(new_n750));
  INV_X1    g564(.A(new_n502), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n749), .A2(new_n738), .A3(new_n750), .A4(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G122), .ZN(G24));
  AND4_X1   g567(.A1(new_n647), .A2(new_n686), .A3(new_n748), .A4(new_n715), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n754), .A2(new_n738), .A3(KEYINPUT102), .A4(new_n657), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT102), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n657), .A2(new_n731), .A3(new_n188), .A4(new_n325), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n686), .A2(new_n748), .A3(new_n647), .A4(new_n715), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n756), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n755), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G125), .ZN(G27));
  NAND2_X1  g575(.A1(new_n567), .A2(new_n561), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n559), .A2(new_n580), .A3(new_n762), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n763), .A2(new_n644), .A3(new_n715), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n391), .A2(new_n392), .A3(new_n327), .ZN(new_n765));
  INV_X1    g579(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n321), .A2(new_n322), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT103), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n767), .A2(new_n768), .A3(new_n305), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n306), .A2(KEYINPUT103), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n769), .A2(new_n770), .A3(G469), .A4(new_n293), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n325), .A2(new_n312), .A3(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n766), .A2(new_n772), .A3(new_n188), .ZN(new_n773));
  OAI21_X1  g587(.A(KEYINPUT42), .B1(new_n764), .B2(new_n773), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n391), .A2(new_n188), .A3(new_n392), .A4(new_n327), .ZN(new_n775));
  AND2_X1   g589(.A1(new_n771), .A2(new_n312), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n775), .B1(new_n325), .B2(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(new_n715), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n778), .A2(KEYINPUT42), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n777), .A2(new_n581), .A3(new_n644), .A4(new_n779), .ZN(new_n780));
  AND2_X1   g594(.A1(new_n774), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G131), .ZN(G33));
  NAND3_X1  g596(.A1(new_n729), .A2(new_n694), .A3(new_n777), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G134), .ZN(G36));
  NAND2_X1  g598(.A1(new_n293), .A2(new_n306), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT45), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n309), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n769), .A2(new_n770), .A3(new_n293), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n787), .B1(new_n788), .B2(new_n786), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n789), .A2(new_n312), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT46), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n720), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n789), .A2(KEYINPUT104), .A3(KEYINPUT46), .A4(new_n312), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n789), .A2(KEYINPUT46), .A3(new_n312), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT104), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n792), .A2(new_n793), .A3(new_n796), .ZN(new_n797));
  AND3_X1   g611(.A1(new_n797), .A2(new_n188), .A3(new_n698), .ZN(new_n798));
  OR2_X1    g612(.A1(new_n459), .A2(KEYINPUT105), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n459), .A2(KEYINPUT105), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n799), .A2(new_n669), .A3(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(KEYINPUT43), .ZN(new_n802));
  INV_X1    g616(.A(new_n459), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT43), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n669), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n802), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n806), .A2(new_n649), .A3(new_n686), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT44), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n765), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n798), .B(new_n809), .C1(new_n808), .C2(new_n807), .ZN(new_n810));
  XNOR2_X1  g624(.A(KEYINPUT106), .B(G137), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n810), .B(new_n811), .ZN(G39));
  NOR4_X1   g626(.A1(new_n581), .A2(new_n644), .A3(new_n778), .A4(new_n765), .ZN(new_n813));
  AND3_X1   g627(.A1(new_n797), .A2(KEYINPUT47), .A3(new_n188), .ZN(new_n814));
  AOI21_X1  g628(.A(KEYINPUT47), .B1(new_n797), .B2(new_n188), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n813), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(G140), .ZN(G42));
  INV_X1    g631(.A(KEYINPUT54), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT53), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT52), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n755), .A2(new_n759), .ZN(new_n821));
  AND2_X1   g635(.A1(new_n693), .A2(KEYINPUT107), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n188), .B1(new_n693), .B2(KEYINPUT107), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n686), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n750), .A2(new_n824), .A3(new_n707), .A4(new_n772), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n696), .A2(new_n717), .A3(new_n825), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n820), .B1(new_n821), .B2(new_n826), .ZN(new_n827));
  OAI211_X1 g641(.A(new_n581), .B(new_n326), .C1(new_n695), .C2(new_n716), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n760), .A2(KEYINPUT52), .A3(new_n828), .A4(new_n825), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n777), .A2(new_n754), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n459), .A2(new_n497), .A3(new_n693), .ZN(new_n832));
  INV_X1    g646(.A(new_n685), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n832), .B1(new_n640), .B2(new_n833), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n834), .A2(new_n765), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n305), .B1(new_n251), .B2(new_n285), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n836), .B1(new_n305), .B2(new_n767), .ZN(new_n837));
  OAI211_X1 g651(.A(KEYINPUT86), .B(G469), .C1(new_n837), .C2(G902), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n325), .A2(new_n838), .A3(new_n313), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n835), .A2(new_n581), .A3(new_n188), .A4(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n777), .A2(new_n581), .A3(new_n644), .ZN(new_n841));
  INV_X1    g655(.A(new_n694), .ZN(new_n842));
  OAI211_X1 g656(.A(new_n831), .B(new_n840), .C1(new_n841), .C2(new_n842), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n502), .B1(new_n670), .B2(new_n677), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n326), .A2(new_n654), .A3(new_n393), .A4(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n645), .A2(new_n845), .A3(new_n689), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n843), .A2(new_n846), .ZN(new_n847));
  AND3_X1   g661(.A1(new_n752), .A2(new_n739), .A3(new_n742), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n847), .A2(new_n735), .A3(new_n781), .A4(new_n848), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n819), .B1(new_n830), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n827), .A2(new_n829), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n781), .A2(new_n735), .A3(new_n848), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n839), .A2(new_n188), .A3(new_n393), .A4(new_n503), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n853), .B1(new_n727), .B2(new_n687), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n839), .A2(new_n188), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n393), .A2(new_n844), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n644), .A2(new_n648), .A3(new_n647), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n854), .A2(new_n858), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n840), .A2(new_n831), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n859), .A2(KEYINPUT53), .A3(new_n783), .A4(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(new_n861), .ZN(new_n862));
  AND4_X1   g676(.A1(KEYINPUT108), .A2(new_n851), .A3(new_n852), .A4(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n781), .A2(new_n735), .A3(new_n848), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n864), .A2(new_n861), .ZN(new_n865));
  AOI21_X1  g679(.A(KEYINPUT108), .B1(new_n865), .B2(new_n851), .ZN(new_n866));
  OAI211_X1 g680(.A(new_n818), .B(new_n850), .C1(new_n863), .C2(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n862), .A2(new_n852), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n868), .A2(new_n830), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n859), .A2(new_n783), .A3(new_n860), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n864), .A2(new_n870), .ZN(new_n871));
  AOI21_X1  g685(.A(KEYINPUT53), .B1(new_n871), .B2(new_n851), .ZN(new_n872));
  OAI21_X1  g686(.A(KEYINPUT54), .B1(new_n869), .B2(new_n872), .ZN(new_n873));
  AND3_X1   g687(.A1(new_n806), .A2(new_n499), .A3(new_n749), .ZN(new_n874));
  INV_X1    g688(.A(new_n757), .ZN(new_n875));
  AOI211_X1 g689(.A(new_n498), .B(G953), .C1(new_n874), .C2(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(new_n499), .ZN(new_n877));
  NOR4_X1   g691(.A1(new_n775), .A2(new_n720), .A3(new_n724), .A4(new_n877), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n707), .A2(new_n653), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n763), .A2(new_n644), .ZN(new_n881));
  AND3_X1   g695(.A1(new_n878), .A2(new_n881), .A3(new_n806), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT48), .ZN(new_n883));
  AND2_X1   g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n882), .A2(new_n883), .ZN(new_n885));
  OAI221_X1 g699(.A(new_n876), .B1(new_n670), .B2(new_n880), .C1(new_n884), .C2(new_n885), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n669), .A2(new_n459), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n878), .A2(new_n879), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n878), .A2(new_n806), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n686), .A2(new_n748), .A3(new_n647), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n888), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NOR3_X1   g705(.A1(new_n711), .A2(new_n327), .A3(new_n732), .ZN(new_n892));
  OAI211_X1 g706(.A(new_n874), .B(new_n892), .C1(KEYINPUT110), .C2(KEYINPUT50), .ZN(new_n893));
  NOR2_X1   g707(.A1(KEYINPUT110), .A2(KEYINPUT50), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n806), .A2(new_n499), .A3(new_n749), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT38), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n676), .B(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n897), .A2(new_n656), .A3(new_n738), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n894), .B1(new_n895), .B2(new_n898), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n891), .B1(new_n893), .B2(new_n899), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n189), .B1(new_n725), .B2(KEYINPUT109), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n901), .B1(KEYINPUT109), .B2(new_n725), .ZN(new_n902));
  NOR3_X1   g716(.A1(new_n814), .A2(new_n815), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n874), .A2(new_n766), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n900), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n905), .A2(KEYINPUT51), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT51), .ZN(new_n907));
  OAI211_X1 g721(.A(new_n900), .B(new_n907), .C1(new_n903), .C2(new_n904), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n886), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n867), .A2(new_n873), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(KEYINPUT111), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT111), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n867), .A2(new_n909), .A3(new_n873), .A4(new_n912), .ZN(new_n913));
  NOR2_X1   g727(.A1(G952), .A2(G953), .ZN(new_n914));
  XOR2_X1   g728(.A(new_n914), .B(KEYINPUT112), .Z(new_n915));
  NAND3_X1  g729(.A1(new_n911), .A2(new_n913), .A3(new_n915), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n725), .B(KEYINPUT49), .ZN(new_n917));
  NOR3_X1   g731(.A1(new_n801), .A2(new_n189), .A3(new_n328), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n917), .A2(new_n897), .A3(new_n879), .A4(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n916), .A2(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT113), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n916), .A2(KEYINPUT113), .A3(new_n919), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n922), .A2(new_n923), .ZN(G75));
  INV_X1    g738(.A(KEYINPUT56), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n850), .B1(new_n863), .B2(new_n866), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(G902), .ZN(new_n927));
  INV_X1    g741(.A(G210), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n925), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n341), .B(new_n366), .ZN(new_n930));
  XNOR2_X1  g744(.A(KEYINPUT114), .B(KEYINPUT55), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n930), .B(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n929), .A2(new_n933), .ZN(new_n934));
  OAI211_X1 g748(.A(new_n925), .B(new_n932), .C1(new_n927), .C2(new_n928), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n289), .A2(G952), .ZN(new_n936));
  INV_X1    g750(.A(new_n936), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n934), .A2(new_n935), .A3(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT115), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n934), .A2(KEYINPUT115), .A3(new_n935), .A4(new_n937), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n940), .A2(new_n941), .ZN(G51));
  INV_X1    g756(.A(new_n723), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n926), .A2(KEYINPUT54), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(new_n867), .ZN(new_n945));
  XNOR2_X1  g759(.A(KEYINPUT116), .B(KEYINPUT57), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n946), .B(new_n311), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n943), .B1(new_n945), .B2(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT117), .ZN(new_n949));
  OR2_X1    g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n927), .A2(new_n789), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n951), .B1(new_n948), .B2(new_n949), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n936), .B1(new_n950), .B2(new_n952), .ZN(G54));
  NAND4_X1  g767(.A1(new_n926), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n954));
  INV_X1    g768(.A(new_n454), .ZN(new_n955));
  AND2_X1   g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n954), .A2(new_n955), .ZN(new_n957));
  NOR3_X1   g771(.A1(new_n956), .A2(new_n957), .A3(new_n936), .ZN(G60));
  XNOR2_X1  g772(.A(new_n667), .B(KEYINPUT118), .ZN(new_n959));
  NAND2_X1  g773(.A1(G478), .A2(G902), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n960), .B(KEYINPUT59), .ZN(new_n961));
  AND3_X1   g775(.A1(new_n945), .A2(new_n959), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n867), .A2(new_n873), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n959), .B1(new_n963), .B2(new_n961), .ZN(new_n964));
  NOR3_X1   g778(.A1(new_n962), .A2(new_n936), .A3(new_n964), .ZN(G63));
  INV_X1    g779(.A(KEYINPUT108), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n966), .B1(new_n868), .B2(new_n830), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n865), .A2(KEYINPUT108), .A3(new_n851), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n872), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(G217), .A2(G902), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n970), .B(KEYINPUT60), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n936), .B1(new_n972), .B2(new_n684), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n973), .A2(KEYINPUT120), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n972), .A2(new_n684), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n638), .B(KEYINPUT119), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n976), .B1(new_n969), .B2(new_n971), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n975), .A2(new_n937), .A3(new_n977), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n974), .A2(new_n978), .A3(KEYINPUT61), .ZN(new_n979));
  INV_X1    g793(.A(KEYINPUT61), .ZN(new_n980));
  OAI211_X1 g794(.A(new_n973), .B(new_n977), .C1(KEYINPUT120), .C2(new_n980), .ZN(new_n981));
  AND2_X1   g795(.A1(new_n979), .A2(new_n981), .ZN(G66));
  NAND3_X1  g796(.A1(new_n735), .A2(new_n848), .A3(new_n859), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n983), .A2(new_n289), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n984), .B(KEYINPUT121), .Z(new_n985));
  OAI21_X1  g799(.A(G953), .B1(new_n501), .B2(new_n336), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g801(.A(G898), .ZN(new_n988));
  INV_X1    g802(.A(new_n289), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n366), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n990), .B(KEYINPUT122), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n987), .B(new_n991), .ZN(G69));
  AOI21_X1  g806(.A(new_n289), .B1(G227), .B2(G900), .ZN(new_n993));
  INV_X1    g807(.A(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT126), .ZN(new_n995));
  AND2_X1   g809(.A1(new_n670), .A2(new_n677), .ZN(new_n996));
  NOR4_X1   g810(.A1(new_n699), .A2(new_n727), .A3(new_n765), .A4(new_n996), .ZN(new_n997));
  AND2_X1   g811(.A1(new_n760), .A2(new_n828), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n998), .A2(new_n712), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n997), .B1(new_n999), .B2(KEYINPUT62), .ZN(new_n1000));
  INV_X1    g814(.A(KEYINPUT62), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n998), .A2(new_n712), .A3(new_n1001), .ZN(new_n1002));
  NAND4_X1  g816(.A1(new_n1000), .A2(new_n810), .A3(new_n816), .A4(new_n1002), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1003), .A2(new_n289), .ZN(new_n1004));
  NOR2_X1   g818(.A1(new_n552), .A2(new_n553), .ZN(new_n1005));
  XOR2_X1   g819(.A(new_n449), .B(KEYINPUT123), .Z(new_n1006));
  XNOR2_X1  g820(.A(new_n1005), .B(new_n1006), .ZN(new_n1007));
  XOR2_X1   g821(.A(new_n1007), .B(KEYINPUT124), .Z(new_n1008));
  INV_X1    g822(.A(new_n1008), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1004), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1010), .A2(KEYINPUT125), .ZN(new_n1011));
  INV_X1    g825(.A(KEYINPUT125), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n1004), .A2(new_n1012), .A3(new_n1009), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n989), .A2(G900), .ZN(new_n1015));
  AND3_X1   g829(.A1(new_n998), .A2(new_n781), .A3(new_n783), .ZN(new_n1016));
  NAND3_X1  g830(.A1(new_n798), .A2(new_n750), .A3(new_n881), .ZN(new_n1017));
  NAND4_X1  g831(.A1(new_n1016), .A2(new_n810), .A3(new_n816), .A4(new_n1017), .ZN(new_n1018));
  OAI211_X1 g832(.A(new_n1007), .B(new_n1015), .C1(new_n1018), .C2(new_n989), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n995), .B1(new_n1014), .B2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g834(.A(new_n1012), .B1(new_n1004), .B2(new_n1009), .ZN(new_n1021));
  AOI211_X1 g835(.A(KEYINPUT125), .B(new_n1008), .C1(new_n1003), .C2(new_n289), .ZN(new_n1022));
  OAI211_X1 g836(.A(new_n995), .B(new_n1019), .C1(new_n1021), .C2(new_n1022), .ZN(new_n1023));
  INV_X1    g837(.A(new_n1023), .ZN(new_n1024));
  OAI21_X1  g838(.A(new_n994), .B1(new_n1020), .B2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g839(.A(new_n1019), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1026), .A2(KEYINPUT126), .ZN(new_n1027));
  NAND3_X1  g841(.A1(new_n1027), .A2(new_n993), .A3(new_n1023), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n1025), .A2(new_n1028), .ZN(G72));
  NAND2_X1  g843(.A1(G472), .A2(G902), .ZN(new_n1030));
  XOR2_X1   g844(.A(new_n1030), .B(KEYINPUT63), .Z(new_n1031));
  OAI21_X1  g845(.A(new_n1031), .B1(new_n1018), .B2(new_n983), .ZN(new_n1032));
  NOR2_X1   g846(.A1(new_n542), .A2(new_n526), .ZN(new_n1033));
  NAND3_X1  g847(.A1(new_n1032), .A2(new_n515), .A3(new_n1033), .ZN(new_n1034));
  OAI221_X1 g848(.A(new_n1031), .B1(new_n703), .B2(new_n578), .C1(new_n869), .C2(new_n872), .ZN(new_n1035));
  NAND3_X1  g849(.A1(new_n1034), .A2(new_n1035), .A3(new_n937), .ZN(new_n1036));
  OAI21_X1  g850(.A(new_n1031), .B1(new_n1003), .B2(new_n983), .ZN(new_n1037));
  XNOR2_X1  g851(.A(new_n1037), .B(KEYINPUT127), .ZN(new_n1038));
  NOR2_X1   g852(.A1(new_n1033), .A2(new_n515), .ZN(new_n1039));
  AOI21_X1  g853(.A(new_n1036), .B1(new_n1038), .B2(new_n1039), .ZN(G57));
endmodule


