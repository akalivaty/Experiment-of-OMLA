//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 0 0 1 0 1 1 1 1 1 0 0 1 0 1 0 0 1 0 0 0 1 0 0 0 1 0 1 1 0 1 0 1 1 1 1 1 0 1 0 1 1 0 0 1 0 1 1 1 1 0 0 0 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:49 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n689, new_n690, new_n691, new_n692,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n750, new_n751, new_n752, new_n753, new_n755, new_n756, new_n757,
    new_n759, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n792, new_n793, new_n794, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n844, new_n846, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n910,
    new_n911, new_n912, new_n913, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n928, new_n929, new_n930, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n945, new_n946, new_n947, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n955, new_n956, new_n957;
  INV_X1    g000(.A(KEYINPUT76), .ZN(new_n202));
  INV_X1    g001(.A(G141gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n203), .A2(G148gat), .ZN(new_n204));
  INV_X1    g003(.A(G148gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n205), .A2(G141gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(KEYINPUT70), .A2(KEYINPUT2), .ZN(new_n207));
  AND2_X1   g006(.A1(KEYINPUT70), .A2(KEYINPUT2), .ZN(new_n208));
  OAI22_X1  g007(.A1(new_n204), .A2(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  XOR2_X1   g008(.A(G155gat), .B(G162gat), .Z(new_n210));
  INV_X1    g009(.A(KEYINPUT71), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n211), .B1(new_n203), .B2(G148gat), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n205), .A2(KEYINPUT71), .A3(G141gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n203), .A2(G148gat), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n212), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT2), .ZN(new_n216));
  INV_X1    g015(.A(G155gat), .ZN(new_n217));
  INV_X1    g016(.A(G162gat), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n216), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(G155gat), .A2(G162gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  AOI22_X1  g020(.A1(new_n209), .A2(new_n210), .B1(new_n215), .B2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT3), .ZN(new_n223));
  AOI21_X1  g022(.A(KEYINPUT29), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(G211gat), .A2(G218gat), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT22), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NOR2_X1   g026(.A1(G197gat), .A2(G204gat), .ZN(new_n228));
  AND2_X1   g027(.A1(G197gat), .A2(G204gat), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n227), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  XOR2_X1   g029(.A(G211gat), .B(G218gat), .Z(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(G211gat), .B(G218gat), .ZN(new_n233));
  XNOR2_X1  g032(.A(G197gat), .B(G204gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n233), .A2(new_n234), .A3(new_n227), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n232), .A2(new_n235), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n202), .B1(new_n224), .B2(new_n236), .ZN(new_n237));
  XNOR2_X1  g036(.A(G141gat), .B(G148gat), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n208), .A2(new_n207), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n210), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n215), .A2(new_n221), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n240), .A2(new_n241), .A3(new_n223), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT29), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n236), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n244), .A2(KEYINPUT76), .A3(new_n245), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n240), .A2(new_n241), .A3(KEYINPUT72), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  AOI21_X1  g047(.A(KEYINPUT72), .B1(new_n240), .B2(new_n241), .ZN(new_n249));
  AOI21_X1  g048(.A(KEYINPUT29), .B1(new_n232), .B2(new_n235), .ZN(new_n250));
  OAI22_X1  g049(.A1(new_n248), .A2(new_n249), .B1(new_n250), .B2(KEYINPUT3), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n237), .A2(new_n246), .A3(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(G228gat), .A2(G233gat), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(G22gat), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n230), .A2(new_n231), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n233), .B1(new_n227), .B2(new_n234), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n243), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n222), .B1(new_n258), .B2(new_n223), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n236), .B1(new_n242), .B2(new_n243), .ZN(new_n260));
  NOR3_X1   g059(.A1(new_n259), .A2(new_n260), .A3(new_n253), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n254), .A2(new_n255), .A3(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n261), .B1(new_n252), .B2(new_n253), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n265), .A2(new_n255), .ZN(new_n266));
  XNOR2_X1  g065(.A(G78gat), .B(G106gat), .ZN(new_n267));
  INV_X1    g066(.A(G50gat), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n267), .B(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(KEYINPUT75), .B(KEYINPUT31), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n269), .B(new_n270), .ZN(new_n271));
  NOR3_X1   g070(.A1(new_n264), .A2(new_n266), .A3(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT77), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n263), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT78), .ZN(new_n276));
  INV_X1    g075(.A(new_n253), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n244), .A2(new_n245), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT72), .ZN(new_n279));
  AND2_X1   g078(.A1(new_n215), .A2(new_n221), .ZN(new_n280));
  XNOR2_X1  g079(.A(G155gat), .B(G162gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n205), .A2(G141gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(new_n214), .ZN(new_n283));
  XNOR2_X1  g082(.A(KEYINPUT70), .B(KEYINPUT2), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n281), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n279), .B1(new_n280), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(new_n247), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n258), .A2(new_n223), .ZN(new_n288));
  AOI22_X1  g087(.A1(new_n278), .A2(new_n202), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n277), .B1(new_n289), .B2(new_n246), .ZN(new_n290));
  OAI211_X1 g089(.A(new_n276), .B(G22gat), .C1(new_n290), .C2(new_n261), .ZN(new_n291));
  OAI21_X1  g090(.A(KEYINPUT78), .B1(new_n265), .B2(new_n255), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n265), .A2(KEYINPUT77), .A3(new_n255), .ZN(new_n293));
  NAND4_X1  g092(.A1(new_n275), .A2(new_n291), .A3(new_n292), .A4(new_n293), .ZN(new_n294));
  AND3_X1   g093(.A1(new_n294), .A2(KEYINPUT79), .A3(new_n271), .ZN(new_n295));
  AOI21_X1  g094(.A(KEYINPUT79), .B1(new_n294), .B2(new_n271), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n273), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT69), .ZN(new_n298));
  NAND2_X1  g097(.A1(G183gat), .A2(G190gat), .ZN(new_n299));
  INV_X1    g098(.A(G169gat), .ZN(new_n300));
  INV_X1    g099(.A(G176gat), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n300), .A2(new_n301), .A3(KEYINPUT26), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT26), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n303), .B1(G169gat), .B2(G176gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(G169gat), .A2(G176gat), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  OAI211_X1 g105(.A(new_n299), .B(new_n302), .C1(new_n304), .C2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(G183gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(KEYINPUT27), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT27), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(G183gat), .ZN(new_n311));
  INV_X1    g110(.A(G190gat), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n309), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT28), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  XNOR2_X1  g114(.A(KEYINPUT27), .B(G183gat), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n316), .A2(KEYINPUT28), .A3(new_n312), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n307), .B1(new_n315), .B2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n299), .A2(KEYINPUT24), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT24), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n321), .A2(G183gat), .A3(G190gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT66), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n324), .B1(G183gat), .B2(G190gat), .ZN(new_n325));
  NOR2_X1   g124(.A1(G183gat), .A2(G190gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(KEYINPUT66), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n323), .A2(new_n325), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n305), .A2(KEYINPUT23), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n300), .A2(new_n301), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n300), .A2(new_n301), .A3(KEYINPUT23), .ZN(new_n332));
  AND2_X1   g131(.A1(new_n332), .A2(KEYINPUT25), .ZN(new_n333));
  AND3_X1   g132(.A1(new_n328), .A2(new_n331), .A3(new_n333), .ZN(new_n334));
  AND2_X1   g133(.A1(KEYINPUT65), .A2(G176gat), .ZN(new_n335));
  NOR2_X1   g134(.A1(KEYINPUT65), .A2(G176gat), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n300), .A2(KEYINPUT23), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  AOI22_X1  g138(.A1(new_n337), .A2(new_n339), .B1(new_n330), .B2(new_n329), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n326), .B1(new_n320), .B2(new_n322), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  AOI21_X1  g141(.A(KEYINPUT25), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n319), .B1(new_n334), .B2(new_n343), .ZN(new_n344));
  AOI22_X1  g143(.A1(new_n344), .A2(new_n243), .B1(G226gat), .B2(G233gat), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT25), .ZN(new_n346));
  XNOR2_X1  g145(.A(KEYINPUT65), .B(G176gat), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n331), .B1(new_n347), .B2(new_n338), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n346), .B1(new_n348), .B2(new_n341), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n328), .A2(new_n331), .A3(new_n333), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n318), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(G226gat), .ZN(new_n352));
  INV_X1    g151(.A(G233gat), .ZN(new_n353));
  NOR3_X1   g152(.A1(new_n351), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  NOR3_X1   g153(.A1(new_n345), .A2(new_n354), .A3(new_n245), .ZN(new_n355));
  OAI22_X1  g154(.A1(new_n351), .A2(KEYINPUT29), .B1(new_n352), .B2(new_n353), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n344), .A2(G226gat), .A3(G233gat), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n236), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n355), .A2(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(G8gat), .B(G36gat), .ZN(new_n360));
  XNOR2_X1  g159(.A(G64gat), .B(G92gat), .ZN(new_n361));
  XOR2_X1   g160(.A(new_n360), .B(new_n361), .Z(new_n362));
  OAI21_X1  g161(.A(new_n298), .B1(new_n359), .B2(new_n362), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n245), .B1(new_n345), .B2(new_n354), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n356), .A2(new_n357), .A3(new_n236), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(new_n362), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n366), .A2(KEYINPUT69), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n363), .A2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT30), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n359), .A2(new_n370), .A3(new_n362), .ZN(new_n371));
  OAI21_X1  g170(.A(KEYINPUT30), .B1(new_n366), .B2(new_n367), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n369), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n240), .A2(new_n241), .ZN(new_n375));
  INV_X1    g174(.A(G113gat), .ZN(new_n376));
  INV_X1    g175(.A(G120gat), .ZN(new_n377));
  AOI21_X1  g176(.A(KEYINPUT1), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(G134gat), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(G127gat), .ZN(new_n380));
  INV_X1    g179(.A(G127gat), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(G134gat), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n378), .A2(new_n380), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n376), .A2(KEYINPUT67), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT67), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(G113gat), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n377), .B1(new_n384), .B2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT1), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n388), .B1(G113gat), .B2(G120gat), .ZN(new_n389));
  AND2_X1   g188(.A1(G113gat), .A2(G120gat), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  XNOR2_X1  g190(.A(G127gat), .B(G134gat), .ZN(new_n392));
  OAI22_X1  g191(.A1(new_n383), .A2(new_n387), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n375), .A2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT74), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n394), .B(new_n395), .ZN(new_n396));
  OAI21_X1  g195(.A(KEYINPUT73), .B1(new_n375), .B2(new_n393), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT73), .ZN(new_n398));
  INV_X1    g197(.A(new_n392), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n399), .B1(new_n389), .B2(new_n390), .ZN(new_n400));
  AND2_X1   g199(.A1(new_n384), .A2(new_n386), .ZN(new_n401));
  OAI211_X1 g200(.A(new_n378), .B(new_n392), .C1(new_n401), .C2(new_n377), .ZN(new_n402));
  NAND4_X1  g201(.A1(new_n222), .A2(new_n398), .A3(new_n400), .A4(new_n402), .ZN(new_n403));
  AND2_X1   g202(.A1(new_n397), .A2(new_n403), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n396), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(G225gat), .A2(G233gat), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n405), .A2(KEYINPUT5), .A3(new_n407), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n397), .A2(new_n403), .A3(KEYINPUT4), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n375), .A2(KEYINPUT3), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n410), .A2(new_n393), .A3(new_n242), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT68), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n393), .A2(new_n414), .ZN(new_n415));
  OAI221_X1 g214(.A(KEYINPUT68), .B1(new_n391), .B2(new_n392), .C1(new_n383), .C2(new_n387), .ZN(new_n416));
  NAND4_X1  g215(.A1(new_n286), .A2(new_n247), .A3(new_n415), .A4(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT4), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(KEYINPUT5), .B1(new_n413), .B2(new_n419), .ZN(new_n420));
  OAI211_X1 g219(.A(KEYINPUT5), .B(new_n411), .C1(new_n417), .C2(new_n418), .ZN(new_n421));
  AOI21_X1  g220(.A(KEYINPUT4), .B1(new_n397), .B2(new_n403), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n406), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n408), .B1(new_n420), .B2(new_n423), .ZN(new_n424));
  XNOR2_X1  g223(.A(G1gat), .B(G29gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(new_n425), .B(KEYINPUT0), .ZN(new_n426));
  XNOR2_X1  g225(.A(G57gat), .B(G85gat), .ZN(new_n427));
  XOR2_X1   g226(.A(new_n426), .B(new_n427), .Z(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n424), .A2(KEYINPUT6), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n424), .A2(new_n429), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT6), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n419), .A2(new_n409), .A3(new_n411), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT5), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  AND2_X1   g234(.A1(new_n411), .A2(KEYINPUT5), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n415), .A2(new_n416), .ZN(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n248), .A2(new_n249), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n438), .A2(new_n439), .A3(KEYINPUT4), .ZN(new_n440));
  OAI211_X1 g239(.A(new_n436), .B(new_n440), .C1(KEYINPUT4), .C2(new_n404), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n435), .A2(new_n441), .A3(new_n406), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n442), .A2(new_n428), .A3(new_n408), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n431), .A2(new_n432), .A3(new_n443), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n374), .B1(new_n430), .B2(new_n444), .ZN(new_n445));
  XOR2_X1   g244(.A(G15gat), .B(G43gat), .Z(new_n446));
  XNOR2_X1  g245(.A(G71gat), .B(G99gat), .ZN(new_n447));
  XNOR2_X1  g246(.A(new_n446), .B(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(G227gat), .A2(G233gat), .ZN(new_n450));
  XOR2_X1   g249(.A(new_n450), .B(KEYINPUT64), .Z(new_n451));
  NOR2_X1   g250(.A1(new_n344), .A2(new_n437), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n349), .A2(new_n350), .ZN(new_n453));
  AOI22_X1  g252(.A1(new_n453), .A2(new_n319), .B1(new_n415), .B2(new_n416), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n451), .B1(new_n452), .B2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT33), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n449), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n340), .A2(new_n342), .ZN(new_n458));
  AND3_X1   g257(.A1(new_n331), .A2(KEYINPUT25), .A3(new_n332), .ZN(new_n459));
  AOI22_X1  g258(.A1(new_n458), .A2(new_n346), .B1(new_n459), .B2(new_n328), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n437), .B1(new_n460), .B2(new_n318), .ZN(new_n461));
  NAND4_X1  g260(.A1(new_n453), .A2(new_n415), .A3(new_n416), .A4(new_n319), .ZN(new_n462));
  INV_X1    g261(.A(new_n451), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n461), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(KEYINPUT34), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT34), .ZN(new_n466));
  NAND4_X1  g265(.A1(new_n461), .A2(new_n462), .A3(new_n466), .A4(new_n463), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n457), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n461), .A2(new_n462), .ZN(new_n470));
  AOI21_X1  g269(.A(KEYINPUT33), .B1(new_n470), .B2(new_n451), .ZN(new_n471));
  OAI211_X1 g270(.A(new_n465), .B(new_n467), .C1(new_n471), .C2(new_n449), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n455), .A2(KEYINPUT32), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  AND3_X1   g273(.A1(new_n469), .A2(new_n472), .A3(new_n474), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n474), .B1(new_n469), .B2(new_n472), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n297), .A2(new_n445), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(KEYINPUT35), .ZN(new_n479));
  AOI22_X1  g278(.A1(new_n363), .A2(new_n368), .B1(new_n371), .B2(new_n372), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT35), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n469), .A2(new_n472), .A3(new_n474), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n469), .A2(new_n472), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(new_n473), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n480), .A2(new_n481), .A3(new_n482), .A4(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT83), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n430), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n428), .B1(new_n442), .B2(new_n408), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n488), .A2(KEYINPUT83), .A3(KEYINPUT6), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n485), .B1(new_n444), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(new_n297), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT36), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n493), .B1(new_n475), .B2(new_n476), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n484), .A2(KEYINPUT36), .A3(new_n482), .ZN(new_n495));
  AND2_X1   g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n294), .A2(new_n271), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT79), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n294), .A2(KEYINPUT79), .A3(new_n271), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n272), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n444), .A2(new_n430), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(new_n480), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n496), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n366), .A2(new_n367), .ZN(new_n505));
  OAI21_X1  g304(.A(KEYINPUT37), .B1(new_n355), .B2(new_n358), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT37), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n364), .A2(new_n507), .A3(new_n365), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT38), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n506), .A2(new_n508), .A3(new_n509), .A4(new_n367), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(KEYINPUT82), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n507), .B1(new_n364), .B2(new_n365), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n512), .A2(new_n362), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT82), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n513), .A2(new_n514), .A3(new_n509), .A4(new_n508), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n505), .B1(new_n511), .B2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT84), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n517), .B1(new_n512), .B2(new_n362), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n506), .A2(KEYINPUT84), .A3(new_n367), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n518), .A2(new_n519), .A3(new_n508), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(KEYINPUT38), .ZN(new_n521));
  NAND4_X1  g320(.A1(new_n516), .A2(new_n490), .A3(new_n444), .A4(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT39), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n433), .A2(KEYINPUT80), .A3(new_n407), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  AOI21_X1  g324(.A(KEYINPUT80), .B1(new_n433), .B2(new_n407), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n523), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n433), .A2(new_n407), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT80), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n523), .B1(new_n405), .B2(new_n406), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n530), .A2(new_n531), .A3(new_n524), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n527), .A2(new_n532), .A3(new_n428), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT40), .ZN(new_n534));
  OAI21_X1  g333(.A(KEYINPUT81), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n488), .B1(new_n369), .B2(new_n373), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n530), .A2(new_n524), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n429), .B1(new_n537), .B2(new_n523), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT81), .ZN(new_n539));
  NAND4_X1  g338(.A1(new_n538), .A2(new_n539), .A3(KEYINPUT40), .A4(new_n532), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n533), .A2(new_n534), .ZN(new_n541));
  NAND4_X1  g340(.A1(new_n535), .A2(new_n536), .A3(new_n540), .A4(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n522), .A2(new_n542), .A3(new_n297), .ZN(new_n543));
  AOI22_X1  g342(.A1(new_n479), .A2(new_n492), .B1(new_n504), .B2(new_n543), .ZN(new_n544));
  OR2_X1    g343(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n545));
  NAND2_X1  g344(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n546));
  AOI21_X1  g345(.A(G36gat), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(G29gat), .ZN(new_n548));
  AND3_X1   g347(.A1(new_n548), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n549));
  OR2_X1    g348(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT86), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  XNOR2_X1  g351(.A(G43gat), .B(G50gat), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n553), .A2(KEYINPUT15), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  NAND4_X1  g354(.A1(new_n550), .A2(new_n551), .A3(KEYINPUT15), .A4(new_n553), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT15), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT87), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n553), .A2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(G43gat), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n560), .A2(KEYINPUT87), .A3(G50gat), .ZN(new_n561));
  NAND4_X1  g360(.A1(new_n550), .A2(new_n557), .A3(new_n559), .A4(new_n561), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n555), .A2(new_n556), .A3(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT88), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND4_X1  g364(.A1(new_n555), .A2(new_n556), .A3(KEYINPUT88), .A4(new_n562), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(G15gat), .B(G22gat), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT16), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n568), .B1(new_n569), .B2(G1gat), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n570), .B1(G1gat), .B2(new_n568), .ZN(new_n571));
  INV_X1    g370(.A(G8gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  OR2_X1    g372(.A1(new_n567), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT17), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n565), .A2(new_n575), .A3(new_n566), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n563), .A2(KEYINPUT17), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n576), .A2(new_n573), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(G229gat), .A2(G233gat), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n574), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT18), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND4_X1  g381(.A1(new_n574), .A2(new_n578), .A3(KEYINPUT18), .A4(new_n579), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n567), .B(new_n573), .ZN(new_n584));
  XOR2_X1   g383(.A(new_n579), .B(KEYINPUT13), .Z(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n582), .A2(new_n583), .A3(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(G113gat), .B(G141gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(KEYINPUT85), .B(KEYINPUT11), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n588), .B(new_n589), .ZN(new_n590));
  XOR2_X1   g389(.A(G169gat), .B(G197gat), .Z(new_n591));
  XNOR2_X1  g390(.A(new_n590), .B(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n592), .B(KEYINPUT12), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n587), .A2(new_n594), .ZN(new_n595));
  NAND4_X1  g394(.A1(new_n582), .A2(new_n583), .A3(new_n586), .A4(new_n593), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n544), .A2(new_n598), .ZN(new_n599));
  AND2_X1   g398(.A1(G232gat), .A2(G233gat), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n600), .A2(KEYINPUT41), .ZN(new_n601));
  XNOR2_X1  g400(.A(G134gat), .B(G162gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(G85gat), .A2(G92gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(KEYINPUT7), .ZN(new_n606));
  XNOR2_X1  g405(.A(G99gat), .B(G106gat), .ZN(new_n607));
  NAND2_X1  g406(.A1(G99gat), .A2(G106gat), .ZN(new_n608));
  INV_X1    g407(.A(G85gat), .ZN(new_n609));
  INV_X1    g408(.A(G92gat), .ZN(new_n610));
  AOI22_X1  g409(.A1(KEYINPUT8), .A2(new_n608), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  AND3_X1   g410(.A1(new_n606), .A2(new_n607), .A3(new_n611), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n607), .B1(new_n606), .B2(new_n611), .ZN(new_n613));
  OAI211_X1 g412(.A(new_n576), .B(new_n577), .C1(new_n612), .C2(new_n613), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n612), .A2(new_n613), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n565), .A2(new_n566), .A3(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(G190gat), .B(G218gat), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT93), .ZN(new_n618));
  AOI22_X1  g417(.A1(new_n617), .A2(new_n618), .B1(KEYINPUT41), .B2(new_n600), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n614), .A2(new_n616), .A3(new_n619), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n617), .A2(new_n618), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n621), .B(KEYINPUT94), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n620), .A2(new_n622), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n604), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n625), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n627), .A2(new_n603), .A3(new_n623), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT90), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n630), .A2(KEYINPUT89), .A3(G57gat), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n631), .B1(KEYINPUT89), .B2(G57gat), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n632), .A2(G64gat), .ZN(new_n633));
  AOI21_X1  g432(.A(G64gat), .B1(new_n630), .B2(G57gat), .ZN(new_n634));
  NAND2_X1  g433(.A1(G71gat), .A2(G78gat), .ZN(new_n635));
  INV_X1    g434(.A(G71gat), .ZN(new_n636));
  INV_X1    g435(.A(G78gat), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n636), .A2(new_n637), .A3(KEYINPUT9), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n634), .B1(new_n635), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n633), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n636), .A2(new_n637), .ZN(new_n641));
  OAI21_X1  g440(.A(KEYINPUT9), .B1(G57gat), .B2(G64gat), .ZN(new_n642));
  AND2_X1   g441(.A1(G57gat), .A2(G64gat), .ZN(new_n643));
  OAI211_X1 g442(.A(new_n635), .B(new_n641), .C1(new_n642), .C2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n640), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT21), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  XOR2_X1   g446(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n648));
  XNOR2_X1  g447(.A(new_n647), .B(new_n648), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n573), .B1(new_n646), .B2(new_n645), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(G127gat), .B(G155gat), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n652), .B(KEYINPUT92), .ZN(new_n653));
  NAND2_X1  g452(.A1(G231gat), .A2(G233gat), .ZN(new_n654));
  XOR2_X1   g453(.A(new_n654), .B(KEYINPUT91), .Z(new_n655));
  XNOR2_X1  g454(.A(new_n653), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(G183gat), .B(G211gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n651), .B(new_n658), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n629), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(G230gat), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n662), .A2(new_n353), .ZN(new_n663));
  INV_X1    g462(.A(new_n645), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(new_n615), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT10), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n645), .B1(new_n613), .B2(new_n612), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n665), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n664), .A2(new_n615), .A3(KEYINPUT10), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n663), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  XNOR2_X1  g470(.A(G120gat), .B(G148gat), .ZN(new_n672));
  XNOR2_X1  g471(.A(G176gat), .B(G204gat), .ZN(new_n673));
  XOR2_X1   g472(.A(new_n672), .B(new_n673), .Z(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n663), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n676), .B1(new_n665), .B2(new_n667), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n675), .B1(new_n677), .B2(KEYINPUT95), .ZN(new_n678));
  OAI211_X1 g477(.A(new_n671), .B(new_n678), .C1(KEYINPUT95), .C2(new_n677), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n675), .B1(new_n670), .B2(new_n677), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n661), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n599), .A2(new_n682), .ZN(new_n683));
  OR2_X1    g482(.A1(new_n502), .A2(KEYINPUT96), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n502), .A2(KEYINPUT96), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  XOR2_X1   g486(.A(new_n687), .B(G1gat), .Z(G1324gat));
  NOR2_X1   g487(.A1(new_n683), .A2(new_n480), .ZN(new_n689));
  XOR2_X1   g488(.A(KEYINPUT16), .B(G8gat), .Z(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n691), .B1(new_n572), .B2(new_n689), .ZN(new_n692));
  MUX2_X1   g491(.A(new_n691), .B(new_n692), .S(KEYINPUT42), .Z(G1325gat));
  NAND2_X1  g492(.A1(new_n494), .A2(new_n495), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(KEYINPUT97), .ZN(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  OAI21_X1  g495(.A(G15gat), .B1(new_n683), .B2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n477), .ZN(new_n698));
  OR2_X1    g497(.A1(new_n698), .A2(G15gat), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n697), .B1(new_n683), .B2(new_n699), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n700), .B(KEYINPUT98), .ZN(G1326gat));
  NOR2_X1   g500(.A1(new_n683), .A2(new_n297), .ZN(new_n702));
  XOR2_X1   g501(.A(KEYINPUT43), .B(G22gat), .Z(new_n703));
  XNOR2_X1  g502(.A(new_n702), .B(new_n703), .ZN(G1327gat));
  INV_X1    g503(.A(new_n544), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(new_n629), .ZN(new_n706));
  INV_X1    g505(.A(new_n681), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n597), .A2(new_n659), .A3(new_n707), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(new_n686), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n709), .A2(new_n548), .A3(new_n710), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n711), .B(KEYINPUT45), .ZN(new_n712));
  INV_X1    g511(.A(new_n629), .ZN(new_n713));
  OAI21_X1  g512(.A(KEYINPUT44), .B1(new_n544), .B2(new_n713), .ZN(new_n714));
  XNOR2_X1  g513(.A(KEYINPUT99), .B(KEYINPUT44), .ZN(new_n715));
  AND2_X1   g514(.A1(new_n504), .A2(new_n543), .ZN(new_n716));
  AOI22_X1  g515(.A1(new_n478), .A2(KEYINPUT35), .B1(new_n491), .B2(new_n297), .ZN(new_n717));
  OAI211_X1 g516(.A(new_n629), .B(new_n715), .C1(new_n716), .C2(new_n717), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n708), .B1(new_n714), .B2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(new_n719), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n720), .A2(new_n686), .ZN(new_n721));
  AND2_X1   g520(.A1(new_n721), .A2(KEYINPUT100), .ZN(new_n722));
  OAI21_X1  g521(.A(G29gat), .B1(new_n721), .B2(KEYINPUT100), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n712), .B1(new_n722), .B2(new_n723), .ZN(G1328gat));
  INV_X1    g523(.A(new_n659), .ZN(new_n725));
  NOR4_X1   g524(.A1(new_n725), .A2(new_n480), .A3(G36gat), .A4(new_n681), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n599), .A2(new_n629), .A3(new_n726), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n727), .A2(KEYINPUT46), .ZN(new_n728));
  XOR2_X1   g527(.A(new_n728), .B(KEYINPUT102), .Z(new_n729));
  OAI21_X1  g528(.A(G36gat), .B1(new_n720), .B2(new_n480), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n727), .A2(KEYINPUT46), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(KEYINPUT101), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n729), .A2(new_n730), .A3(new_n732), .ZN(G1329gat));
  OAI21_X1  g532(.A(G43gat), .B1(new_n720), .B2(new_n694), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n709), .A2(new_n560), .A3(new_n477), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n734), .A2(KEYINPUT47), .A3(new_n735), .ZN(new_n736));
  OAI21_X1  g535(.A(G43gat), .B1(new_n720), .B2(new_n696), .ZN(new_n737));
  AND2_X1   g536(.A1(new_n737), .A2(new_n735), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n736), .B1(new_n738), .B2(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g538(.A1(new_n709), .A2(new_n268), .A3(new_n501), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n720), .A2(new_n297), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n740), .B1(new_n741), .B2(new_n268), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT103), .ZN(new_n743));
  AOI21_X1  g542(.A(KEYINPUT48), .B1(new_n740), .B2(new_n743), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n742), .B(new_n744), .ZN(G1331gat));
  NOR4_X1   g544(.A1(new_n544), .A2(new_n597), .A3(new_n661), .A4(new_n707), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(new_n710), .ZN(new_n747));
  XNOR2_X1  g546(.A(KEYINPUT89), .B(G57gat), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n747), .B(new_n748), .ZN(G1332gat));
  AOI21_X1  g548(.A(new_n480), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n746), .A2(new_n750), .ZN(new_n751));
  XOR2_X1   g550(.A(new_n751), .B(KEYINPUT104), .Z(new_n752));
  NOR2_X1   g551(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n752), .B(new_n753), .ZN(G1333gat));
  AOI21_X1  g553(.A(new_n636), .B1(new_n746), .B2(new_n695), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n698), .A2(G71gat), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n755), .B1(new_n746), .B2(new_n756), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g557(.A1(new_n746), .A2(new_n501), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n759), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g559(.A1(new_n714), .A2(new_n718), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n597), .A2(new_n725), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(new_n681), .ZN(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  AOI21_X1  g563(.A(KEYINPUT105), .B1(new_n761), .B2(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT105), .ZN(new_n766));
  AOI211_X1 g565(.A(new_n766), .B(new_n763), .C1(new_n714), .C2(new_n718), .ZN(new_n767));
  NOR3_X1   g566(.A1(new_n765), .A2(new_n767), .A3(new_n686), .ZN(new_n768));
  AND2_X1   g567(.A1(new_n768), .A2(KEYINPUT106), .ZN(new_n769));
  OAI21_X1  g568(.A(G85gat), .B1(new_n768), .B2(KEYINPUT106), .ZN(new_n770));
  NOR4_X1   g569(.A1(new_n544), .A2(new_n597), .A3(new_n725), .A4(new_n713), .ZN(new_n771));
  XOR2_X1   g570(.A(new_n771), .B(KEYINPUT51), .Z(new_n772));
  NOR3_X1   g571(.A1(new_n686), .A2(G85gat), .A3(new_n707), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n773), .B(KEYINPUT107), .ZN(new_n774));
  OAI22_X1  g573(.A1(new_n769), .A2(new_n770), .B1(new_n772), .B2(new_n774), .ZN(G1336gat));
  NAND2_X1  g574(.A1(new_n761), .A2(new_n764), .ZN(new_n776));
  OAI21_X1  g575(.A(G92gat), .B1(new_n776), .B2(new_n480), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT52), .ZN(new_n778));
  NOR3_X1   g577(.A1(new_n480), .A2(G92gat), .A3(new_n707), .ZN(new_n779));
  INV_X1    g578(.A(new_n779), .ZN(new_n780));
  OAI211_X1 g579(.A(new_n777), .B(new_n778), .C1(new_n772), .C2(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n776), .A2(new_n766), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n761), .A2(KEYINPUT105), .A3(new_n764), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n782), .A2(new_n374), .A3(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(new_n771), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT109), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n786), .A2(KEYINPUT51), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n785), .B(new_n787), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n779), .B(KEYINPUT108), .ZN(new_n789));
  AOI22_X1  g588(.A1(new_n784), .A2(G92gat), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n781), .B1(new_n790), .B2(new_n778), .ZN(G1337gat));
  NOR3_X1   g590(.A1(new_n765), .A2(new_n767), .A3(new_n696), .ZN(new_n792));
  INV_X1    g591(.A(G99gat), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n477), .A2(new_n793), .A3(new_n681), .ZN(new_n794));
  OAI22_X1  g593(.A1(new_n792), .A2(new_n793), .B1(new_n772), .B2(new_n794), .ZN(G1338gat));
  NOR3_X1   g594(.A1(new_n765), .A2(new_n767), .A3(new_n297), .ZN(new_n796));
  INV_X1    g595(.A(G106gat), .ZN(new_n797));
  OAI21_X1  g596(.A(KEYINPUT110), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n782), .A2(new_n501), .A3(new_n783), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT110), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n799), .A2(new_n800), .A3(G106gat), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n501), .A2(new_n797), .A3(new_n681), .ZN(new_n802));
  INV_X1    g601(.A(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n788), .A2(new_n803), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n798), .A2(new_n801), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(KEYINPUT53), .ZN(new_n806));
  OAI21_X1  g605(.A(G106gat), .B1(new_n776), .B2(new_n297), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT53), .ZN(new_n808));
  OAI211_X1 g607(.A(new_n807), .B(new_n808), .C1(new_n772), .C2(new_n802), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n806), .A2(new_n809), .ZN(G1339gat));
  NAND3_X1  g609(.A1(new_n668), .A2(new_n663), .A3(new_n669), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(KEYINPUT111), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT111), .ZN(new_n813));
  NAND4_X1  g612(.A1(new_n668), .A2(new_n813), .A3(new_n663), .A4(new_n669), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n812), .A2(new_n671), .A3(KEYINPUT54), .A4(new_n814), .ZN(new_n815));
  XOR2_X1   g614(.A(KEYINPUT112), .B(KEYINPUT54), .Z(new_n816));
  AOI21_X1  g615(.A(new_n674), .B1(new_n670), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT55), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n815), .A2(KEYINPUT55), .A3(new_n817), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n820), .A2(new_n679), .A3(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT113), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n820), .A2(KEYINPUT113), .A3(new_n679), .A4(new_n821), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n597), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n584), .A2(new_n585), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n579), .B1(new_n574), .B2(new_n578), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n592), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  AND3_X1   g628(.A1(new_n596), .A2(new_n829), .A3(new_n681), .ZN(new_n830));
  INV_X1    g629(.A(new_n830), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n629), .B1(new_n826), .B2(new_n831), .ZN(new_n832));
  AND2_X1   g631(.A1(new_n596), .A2(new_n829), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n629), .A2(new_n824), .A3(new_n825), .A4(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(new_n834), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n659), .B1(new_n832), .B2(new_n835), .ZN(new_n836));
  NOR4_X1   g635(.A1(new_n629), .A2(new_n597), .A3(new_n659), .A4(new_n681), .ZN(new_n837));
  INV_X1    g636(.A(new_n837), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n501), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  NOR3_X1   g638(.A1(new_n686), .A2(new_n374), .A3(new_n698), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n841), .A2(new_n598), .ZN(new_n842));
  MUX2_X1   g641(.A(G113gat), .B(new_n401), .S(new_n842), .Z(G1340gat));
  NOR2_X1   g642(.A1(new_n841), .A2(new_n707), .ZN(new_n844));
  XNOR2_X1  g643(.A(new_n844), .B(new_n377), .ZN(G1341gat));
  NOR2_X1   g644(.A1(new_n841), .A2(new_n659), .ZN(new_n846));
  XNOR2_X1  g645(.A(new_n846), .B(new_n381), .ZN(G1342gat));
  NAND3_X1  g646(.A1(new_n839), .A2(new_n629), .A3(new_n840), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n848), .A2(G134gat), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n848), .A2(G134gat), .ZN(new_n850));
  XOR2_X1   g649(.A(KEYINPUT114), .B(KEYINPUT56), .Z(new_n851));
  AOI21_X1  g650(.A(new_n849), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n852), .B1(new_n850), .B2(new_n851), .ZN(G1343gat));
  INV_X1    g652(.A(KEYINPUT119), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT58), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n836), .A2(new_n838), .ZN(new_n856));
  NOR4_X1   g655(.A1(new_n695), .A2(new_n686), .A3(new_n374), .A4(new_n297), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n598), .A2(G141gat), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n856), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT117), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND4_X1  g660(.A1(new_n856), .A2(KEYINPUT117), .A3(new_n857), .A4(new_n858), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n297), .B1(new_n836), .B2(new_n838), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT57), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NOR3_X1   g665(.A1(new_n686), .A2(new_n374), .A3(new_n496), .ZN(new_n867));
  XNOR2_X1  g666(.A(new_n867), .B(KEYINPUT115), .ZN(new_n868));
  INV_X1    g667(.A(new_n822), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n830), .B1(new_n869), .B2(new_n597), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n834), .B1(new_n870), .B2(new_n629), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n837), .B1(new_n871), .B2(new_n659), .ZN(new_n872));
  OAI21_X1  g671(.A(KEYINPUT57), .B1(new_n872), .B2(new_n297), .ZN(new_n873));
  NAND4_X1  g672(.A1(new_n866), .A2(new_n597), .A3(new_n868), .A4(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(G141gat), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT116), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n863), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n874), .A2(KEYINPUT116), .A3(G141gat), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n855), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  XNOR2_X1  g678(.A(KEYINPUT118), .B(KEYINPUT58), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n875), .A2(new_n859), .A3(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(new_n881), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n854), .B1(new_n879), .B2(new_n882), .ZN(new_n883));
  AND3_X1   g682(.A1(new_n874), .A2(KEYINPUT116), .A3(G141gat), .ZN(new_n884));
  AOI21_X1  g683(.A(KEYINPUT116), .B1(new_n874), .B2(G141gat), .ZN(new_n885));
  NOR3_X1   g684(.A1(new_n884), .A2(new_n885), .A3(new_n863), .ZN(new_n886));
  OAI211_X1 g685(.A(KEYINPUT119), .B(new_n881), .C1(new_n886), .C2(new_n855), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n883), .A2(new_n887), .ZN(G1344gat));
  XOR2_X1   g687(.A(new_n837), .B(KEYINPUT120), .Z(new_n889));
  OR2_X1    g688(.A1(new_n870), .A2(new_n629), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n629), .A2(new_n869), .A3(new_n833), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n725), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  OAI211_X1 g691(.A(new_n865), .B(new_n501), .C1(new_n889), .C2(new_n892), .ZN(new_n893));
  AND2_X1   g692(.A1(new_n868), .A2(new_n681), .ZN(new_n894));
  OAI211_X1 g693(.A(new_n893), .B(new_n894), .C1(new_n864), .C2(new_n865), .ZN(new_n895));
  AND2_X1   g694(.A1(new_n895), .A2(KEYINPUT121), .ZN(new_n896));
  OAI21_X1  g695(.A(G148gat), .B1(new_n895), .B2(KEYINPUT121), .ZN(new_n897));
  OAI21_X1  g696(.A(KEYINPUT59), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n205), .A2(KEYINPUT59), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n866), .A2(new_n868), .A3(new_n873), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n899), .B1(new_n900), .B2(new_n707), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n898), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n856), .A2(new_n857), .ZN(new_n903));
  INV_X1    g702(.A(new_n903), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n904), .A2(new_n205), .A3(new_n681), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n902), .A2(new_n905), .ZN(G1345gat));
  OAI21_X1  g705(.A(G155gat), .B1(new_n900), .B2(new_n659), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n904), .A2(new_n217), .A3(new_n725), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(G1346gat));
  OR2_X1    g708(.A1(new_n900), .A2(new_n713), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n218), .B1(new_n910), .B2(KEYINPUT122), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n911), .B1(KEYINPUT122), .B2(new_n910), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n904), .A2(new_n218), .A3(new_n629), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(new_n913), .ZN(G1347gat));
  AOI21_X1  g713(.A(new_n710), .B1(new_n836), .B2(new_n838), .ZN(new_n915));
  AND4_X1   g714(.A1(new_n374), .A2(new_n915), .A3(new_n297), .A4(new_n477), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n916), .A2(new_n300), .A3(new_n597), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n686), .A2(new_n374), .ZN(new_n918));
  XNOR2_X1  g717(.A(new_n918), .B(KEYINPUT123), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n919), .A2(new_n698), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(new_n839), .ZN(new_n921));
  OAI21_X1  g720(.A(G169gat), .B1(new_n921), .B2(new_n598), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n917), .A2(new_n922), .ZN(new_n923));
  XNOR2_X1  g722(.A(new_n923), .B(KEYINPUT124), .ZN(G1348gat));
  AOI21_X1  g723(.A(G176gat), .B1(new_n916), .B2(new_n681), .ZN(new_n925));
  NOR3_X1   g724(.A1(new_n921), .A2(new_n337), .A3(new_n707), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n925), .A2(new_n926), .ZN(G1349gat));
  NAND3_X1  g726(.A1(new_n916), .A2(new_n316), .A3(new_n725), .ZN(new_n928));
  OAI21_X1  g727(.A(G183gat), .B1(new_n921), .B2(new_n659), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  XNOR2_X1  g729(.A(new_n930), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g730(.A1(new_n916), .A2(new_n312), .A3(new_n629), .ZN(new_n932));
  XNOR2_X1  g731(.A(new_n932), .B(KEYINPUT125), .ZN(new_n933));
  OAI21_X1  g732(.A(G190gat), .B1(new_n921), .B2(new_n713), .ZN(new_n934));
  XOR2_X1   g733(.A(KEYINPUT126), .B(KEYINPUT61), .Z(new_n935));
  XNOR2_X1  g734(.A(new_n934), .B(new_n935), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n933), .A2(new_n936), .ZN(G1351gat));
  NOR2_X1   g736(.A1(new_n919), .A2(new_n695), .ZN(new_n938));
  OAI211_X1 g737(.A(new_n893), .B(new_n938), .C1(new_n864), .C2(new_n865), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n597), .A2(G197gat), .ZN(new_n940));
  NAND4_X1  g739(.A1(new_n915), .A2(new_n374), .A3(new_n501), .A4(new_n696), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n941), .A2(new_n598), .ZN(new_n942));
  OAI22_X1  g741(.A1(new_n939), .A2(new_n940), .B1(G197gat), .B2(new_n942), .ZN(new_n943));
  INV_X1    g742(.A(new_n943), .ZN(G1352gat));
  NOR3_X1   g743(.A1(new_n941), .A2(G204gat), .A3(new_n707), .ZN(new_n945));
  XNOR2_X1  g744(.A(new_n945), .B(KEYINPUT62), .ZN(new_n946));
  OAI21_X1  g745(.A(G204gat), .B1(new_n939), .B2(new_n707), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n947), .ZN(G1353gat));
  OR3_X1    g747(.A1(new_n941), .A2(G211gat), .A3(new_n659), .ZN(new_n949));
  OR2_X1    g748(.A1(new_n939), .A2(new_n659), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n950), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n951));
  INV_X1    g750(.A(new_n951), .ZN(new_n952));
  AOI21_X1  g751(.A(KEYINPUT63), .B1(new_n950), .B2(G211gat), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n949), .B1(new_n952), .B2(new_n953), .ZN(G1354gat));
  OAI21_X1  g753(.A(G218gat), .B1(new_n939), .B2(new_n713), .ZN(new_n955));
  OR2_X1    g754(.A1(new_n713), .A2(G218gat), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n955), .B1(new_n941), .B2(new_n956), .ZN(new_n957));
  XNOR2_X1  g756(.A(new_n957), .B(KEYINPUT127), .ZN(G1355gat));
endmodule


