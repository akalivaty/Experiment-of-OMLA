

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579;

  INV_X1 U321 ( .A(KEYINPUT66), .ZN(n291) );
  XNOR2_X1 U322 ( .A(KEYINPUT113), .B(KEYINPUT48), .ZN(n413) );
  XNOR2_X1 U323 ( .A(n292), .B(n291), .ZN(n293) );
  XNOR2_X1 U324 ( .A(n414), .B(n413), .ZN(n519) );
  XNOR2_X1 U325 ( .A(n294), .B(n293), .ZN(n298) );
  NOR2_X1 U326 ( .A1(n512), .A2(n447), .ZN(n555) );
  XNOR2_X1 U327 ( .A(G169GAT), .B(KEYINPUT120), .ZN(n448) );
  XNOR2_X1 U328 ( .A(n449), .B(n448), .ZN(G1348GAT) );
  XOR2_X1 U329 ( .A(G141GAT), .B(G22GAT), .Z(n348) );
  XOR2_X1 U330 ( .A(G1GAT), .B(KEYINPUT71), .Z(n290) );
  XNOR2_X1 U331 ( .A(G15GAT), .B(G8GAT), .ZN(n289) );
  XNOR2_X1 U332 ( .A(n290), .B(n289), .ZN(n396) );
  XOR2_X1 U333 ( .A(n348), .B(n396), .Z(n294) );
  NAND2_X1 U334 ( .A1(G229GAT), .A2(G233GAT), .ZN(n292) );
  XOR2_X1 U335 ( .A(G29GAT), .B(G43GAT), .Z(n296) );
  XNOR2_X1 U336 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n295) );
  XNOR2_X1 U337 ( .A(n296), .B(n295), .ZN(n355) );
  XNOR2_X1 U338 ( .A(n355), .B(KEYINPUT30), .ZN(n297) );
  XNOR2_X1 U339 ( .A(n298), .B(n297), .ZN(n302) );
  XOR2_X1 U340 ( .A(G113GAT), .B(G50GAT), .Z(n300) );
  XNOR2_X1 U341 ( .A(G169GAT), .B(G36GAT), .ZN(n299) );
  XNOR2_X1 U342 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U343 ( .A(n302), .B(n301), .Z(n310) );
  XOR2_X1 U344 ( .A(KEYINPUT70), .B(KEYINPUT72), .Z(n304) );
  XNOR2_X1 U345 ( .A(KEYINPUT68), .B(KEYINPUT69), .ZN(n303) );
  XNOR2_X1 U346 ( .A(n304), .B(n303), .ZN(n308) );
  XOR2_X1 U347 ( .A(KEYINPUT29), .B(KEYINPUT67), .Z(n306) );
  XNOR2_X1 U348 ( .A(G197GAT), .B(KEYINPUT65), .ZN(n305) );
  XNOR2_X1 U349 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U350 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U351 ( .A(n310), .B(n309), .ZN(n564) );
  XNOR2_X1 U352 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n311) );
  XNOR2_X1 U353 ( .A(n311), .B(KEYINPUT88), .ZN(n312) );
  XOR2_X1 U354 ( .A(n312), .B(KEYINPUT17), .Z(n314) );
  XNOR2_X1 U355 ( .A(G169GAT), .B(G183GAT), .ZN(n313) );
  XNOR2_X1 U356 ( .A(n314), .B(n313), .ZN(n416) );
  XOR2_X1 U357 ( .A(G190GAT), .B(G99GAT), .Z(n316) );
  XOR2_X1 U358 ( .A(G120GAT), .B(G71GAT), .Z(n368) );
  XNOR2_X1 U359 ( .A(n368), .B(KEYINPUT86), .ZN(n315) );
  XNOR2_X1 U360 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U361 ( .A(n416), .B(n317), .Z(n319) );
  NAND2_X1 U362 ( .A1(G227GAT), .A2(G233GAT), .ZN(n318) );
  XNOR2_X1 U363 ( .A(n319), .B(n318), .ZN(n323) );
  XOR2_X1 U364 ( .A(G176GAT), .B(KEYINPUT85), .Z(n321) );
  XNOR2_X1 U365 ( .A(G43GAT), .B(G15GAT), .ZN(n320) );
  XNOR2_X1 U366 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U367 ( .A(n323), .B(n322), .Z(n331) );
  XOR2_X1 U368 ( .A(KEYINPUT84), .B(G134GAT), .Z(n325) );
  XNOR2_X1 U369 ( .A(KEYINPUT0), .B(G127GAT), .ZN(n324) );
  XNOR2_X1 U370 ( .A(n325), .B(n324), .ZN(n326) );
  XOR2_X1 U371 ( .A(G113GAT), .B(n326), .Z(n444) );
  XOR2_X1 U372 ( .A(KEYINPUT87), .B(KEYINPUT20), .Z(n328) );
  XNOR2_X1 U373 ( .A(KEYINPUT90), .B(KEYINPUT89), .ZN(n327) );
  XNOR2_X1 U374 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U375 ( .A(n444), .B(n329), .ZN(n330) );
  XNOR2_X1 U376 ( .A(n331), .B(n330), .ZN(n512) );
  XNOR2_X1 U377 ( .A(KEYINPUT94), .B(KEYINPUT92), .ZN(n332) );
  XNOR2_X1 U378 ( .A(n332), .B(G155GAT), .ZN(n333) );
  XOR2_X1 U379 ( .A(n333), .B(KEYINPUT93), .Z(n335) );
  XNOR2_X1 U380 ( .A(KEYINPUT2), .B(KEYINPUT3), .ZN(n334) );
  XNOR2_X1 U381 ( .A(n335), .B(n334), .ZN(n440) );
  XOR2_X1 U382 ( .A(G148GAT), .B(G106GAT), .Z(n337) );
  XNOR2_X1 U383 ( .A(KEYINPUT75), .B(G78GAT), .ZN(n336) );
  XNOR2_X1 U384 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U385 ( .A(KEYINPUT76), .B(n338), .Z(n381) );
  XNOR2_X1 U386 ( .A(n440), .B(n381), .ZN(n352) );
  XOR2_X1 U387 ( .A(KEYINPUT24), .B(G204GAT), .Z(n340) );
  XNOR2_X1 U388 ( .A(KEYINPUT23), .B(KEYINPUT22), .ZN(n339) );
  XNOR2_X1 U389 ( .A(n340), .B(n339), .ZN(n344) );
  XOR2_X1 U390 ( .A(KEYINPUT21), .B(G218GAT), .Z(n342) );
  XNOR2_X1 U391 ( .A(KEYINPUT91), .B(G211GAT), .ZN(n341) );
  XNOR2_X1 U392 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U393 ( .A(G197GAT), .B(n343), .Z(n415) );
  XOR2_X1 U394 ( .A(n344), .B(n415), .Z(n350) );
  XOR2_X1 U395 ( .A(G50GAT), .B(G162GAT), .Z(n362) );
  XOR2_X1 U396 ( .A(n362), .B(KEYINPUT95), .Z(n346) );
  NAND2_X1 U397 ( .A1(G228GAT), .A2(G233GAT), .ZN(n345) );
  XNOR2_X1 U398 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U399 ( .A(n348), .B(n347), .ZN(n349) );
  XNOR2_X1 U400 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U401 ( .A(n352), .B(n351), .ZN(n455) );
  XOR2_X1 U402 ( .A(KEYINPUT9), .B(KEYINPUT64), .Z(n354) );
  XNOR2_X1 U403 ( .A(G218GAT), .B(KEYINPUT10), .ZN(n353) );
  XNOR2_X1 U404 ( .A(n354), .B(n353), .ZN(n366) );
  XOR2_X1 U405 ( .A(G99GAT), .B(G85GAT), .Z(n367) );
  XOR2_X1 U406 ( .A(n367), .B(n355), .Z(n357) );
  NAND2_X1 U407 ( .A1(G232GAT), .A2(G233GAT), .ZN(n356) );
  XNOR2_X1 U408 ( .A(n357), .B(n356), .ZN(n361) );
  XOR2_X1 U409 ( .A(KEYINPUT11), .B(G92GAT), .Z(n359) );
  XNOR2_X1 U410 ( .A(G134GAT), .B(G106GAT), .ZN(n358) );
  XNOR2_X1 U411 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U412 ( .A(n361), .B(n360), .Z(n364) );
  XOR2_X1 U413 ( .A(G36GAT), .B(G190GAT), .Z(n421) );
  XNOR2_X1 U414 ( .A(n362), .B(n421), .ZN(n363) );
  XNOR2_X1 U415 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U416 ( .A(n366), .B(n365), .ZN(n556) );
  XNOR2_X1 U417 ( .A(n368), .B(n367), .ZN(n371) );
  XOR2_X1 U418 ( .A(KEYINPUT73), .B(KEYINPUT74), .Z(n370) );
  XNOR2_X1 U419 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n369) );
  XNOR2_X1 U420 ( .A(n370), .B(n369), .ZN(n400) );
  XNOR2_X1 U421 ( .A(n371), .B(n400), .ZN(n377) );
  XOR2_X1 U422 ( .A(G64GAT), .B(G92GAT), .Z(n373) );
  XNOR2_X1 U423 ( .A(G176GAT), .B(G204GAT), .ZN(n372) );
  XNOR2_X1 U424 ( .A(n373), .B(n372), .ZN(n417) );
  XOR2_X1 U425 ( .A(KEYINPUT33), .B(n417), .Z(n375) );
  NAND2_X1 U426 ( .A1(G230GAT), .A2(G233GAT), .ZN(n374) );
  XNOR2_X1 U427 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U428 ( .A(n377), .B(n376), .Z(n383) );
  XOR2_X1 U429 ( .A(KEYINPUT77), .B(KEYINPUT31), .Z(n379) );
  XNOR2_X1 U430 ( .A(KEYINPUT32), .B(KEYINPUT78), .ZN(n378) );
  XNOR2_X1 U431 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U432 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U433 ( .A(n383), .B(n382), .ZN(n567) );
  XOR2_X1 U434 ( .A(n567), .B(KEYINPUT41), .Z(n551) );
  NAND2_X1 U435 ( .A1(n564), .A2(n551), .ZN(n384) );
  XNOR2_X1 U436 ( .A(n384), .B(KEYINPUT46), .ZN(n405) );
  XOR2_X1 U437 ( .A(KEYINPUT83), .B(KEYINPUT14), .Z(n386) );
  XNOR2_X1 U438 ( .A(KEYINPUT12), .B(KEYINPUT80), .ZN(n385) );
  XNOR2_X1 U439 ( .A(n386), .B(n385), .ZN(n404) );
  XOR2_X1 U440 ( .A(G211GAT), .B(G155GAT), .Z(n388) );
  XNOR2_X1 U441 ( .A(G22GAT), .B(G71GAT), .ZN(n387) );
  XNOR2_X1 U442 ( .A(n388), .B(n387), .ZN(n392) );
  XOR2_X1 U443 ( .A(KEYINPUT15), .B(KEYINPUT79), .Z(n390) );
  XNOR2_X1 U444 ( .A(G78GAT), .B(G64GAT), .ZN(n389) );
  XNOR2_X1 U445 ( .A(n390), .B(n389), .ZN(n391) );
  XOR2_X1 U446 ( .A(n392), .B(n391), .Z(n398) );
  XOR2_X1 U447 ( .A(G183GAT), .B(G127GAT), .Z(n394) );
  NAND2_X1 U448 ( .A1(G231GAT), .A2(G233GAT), .ZN(n393) );
  XNOR2_X1 U449 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U450 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U451 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U452 ( .A(n399), .B(KEYINPUT81), .Z(n402) );
  XNOR2_X1 U453 ( .A(n400), .B(KEYINPUT82), .ZN(n401) );
  XNOR2_X1 U454 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U455 ( .A(n404), .B(n403), .Z(n544) );
  NAND2_X1 U456 ( .A1(n405), .A2(n544), .ZN(n406) );
  NOR2_X1 U457 ( .A1(n556), .A2(n406), .ZN(n407) );
  XNOR2_X1 U458 ( .A(KEYINPUT47), .B(n407), .ZN(n412) );
  INV_X1 U459 ( .A(n556), .ZN(n535) );
  XNOR2_X1 U460 ( .A(KEYINPUT36), .B(n535), .ZN(n577) );
  NOR2_X1 U461 ( .A1(n544), .A2(n577), .ZN(n408) );
  XNOR2_X1 U462 ( .A(KEYINPUT45), .B(n408), .ZN(n410) );
  NOR2_X1 U463 ( .A1(n564), .A2(n567), .ZN(n409) );
  NAND2_X1 U464 ( .A1(n410), .A2(n409), .ZN(n411) );
  NAND2_X1 U465 ( .A1(n412), .A2(n411), .ZN(n414) );
  XNOR2_X1 U466 ( .A(n416), .B(n415), .ZN(n425) );
  XOR2_X1 U467 ( .A(n417), .B(KEYINPUT97), .Z(n419) );
  NAND2_X1 U468 ( .A1(G226GAT), .A2(G233GAT), .ZN(n418) );
  XNOR2_X1 U469 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U470 ( .A(n420), .B(KEYINPUT98), .Z(n423) );
  XNOR2_X1 U471 ( .A(G8GAT), .B(n421), .ZN(n422) );
  XNOR2_X1 U472 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U473 ( .A(n425), .B(n424), .ZN(n509) );
  XOR2_X1 U474 ( .A(KEYINPUT119), .B(n509), .Z(n426) );
  NOR2_X1 U475 ( .A1(n519), .A2(n426), .ZN(n427) );
  XNOR2_X1 U476 ( .A(n427), .B(KEYINPUT54), .ZN(n445) );
  XOR2_X1 U477 ( .A(G57GAT), .B(G148GAT), .Z(n429) );
  XNOR2_X1 U478 ( .A(G141GAT), .B(G1GAT), .ZN(n428) );
  XNOR2_X1 U479 ( .A(n429), .B(n428), .ZN(n433) );
  XOR2_X1 U480 ( .A(KEYINPUT1), .B(KEYINPUT4), .Z(n431) );
  XNOR2_X1 U481 ( .A(KEYINPUT96), .B(KEYINPUT6), .ZN(n430) );
  XNOR2_X1 U482 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U483 ( .A(n433), .B(n432), .Z(n442) );
  XOR2_X1 U484 ( .A(G85GAT), .B(G162GAT), .Z(n435) );
  XNOR2_X1 U485 ( .A(G29GAT), .B(G120GAT), .ZN(n434) );
  XNOR2_X1 U486 ( .A(n435), .B(n434), .ZN(n436) );
  XOR2_X1 U487 ( .A(KEYINPUT5), .B(n436), .Z(n438) );
  NAND2_X1 U488 ( .A1(G225GAT), .A2(G233GAT), .ZN(n437) );
  XNOR2_X1 U489 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U490 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U491 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U492 ( .A(n444), .B(n443), .ZN(n506) );
  NAND2_X1 U493 ( .A1(n445), .A2(n506), .ZN(n562) );
  NOR2_X1 U494 ( .A1(n455), .A2(n562), .ZN(n446) );
  XNOR2_X1 U495 ( .A(n446), .B(KEYINPUT55), .ZN(n447) );
  NAND2_X1 U496 ( .A1(n564), .A2(n555), .ZN(n449) );
  INV_X1 U497 ( .A(n564), .ZN(n524) );
  NOR2_X1 U498 ( .A1(n567), .A2(n524), .ZN(n479) );
  INV_X1 U499 ( .A(n512), .ZN(n522) );
  XNOR2_X1 U500 ( .A(n509), .B(KEYINPUT27), .ZN(n457) );
  NOR2_X1 U501 ( .A1(n457), .A2(n506), .ZN(n450) );
  XNOR2_X1 U502 ( .A(n450), .B(KEYINPUT99), .ZN(n518) );
  XNOR2_X1 U503 ( .A(n455), .B(KEYINPUT28), .ZN(n521) );
  NOR2_X1 U504 ( .A1(n518), .A2(n521), .ZN(n451) );
  XOR2_X1 U505 ( .A(n451), .B(KEYINPUT100), .Z(n452) );
  NOR2_X1 U506 ( .A1(n522), .A2(n452), .ZN(n462) );
  INV_X1 U507 ( .A(n506), .ZN(n494) );
  NOR2_X1 U508 ( .A1(n512), .A2(n509), .ZN(n453) );
  NOR2_X1 U509 ( .A1(n455), .A2(n453), .ZN(n454) );
  XOR2_X1 U510 ( .A(KEYINPUT25), .B(n454), .Z(n459) );
  NAND2_X1 U511 ( .A1(n455), .A2(n512), .ZN(n456) );
  XNOR2_X1 U512 ( .A(n456), .B(KEYINPUT26), .ZN(n563) );
  NOR2_X1 U513 ( .A1(n457), .A2(n563), .ZN(n458) );
  NOR2_X1 U514 ( .A1(n459), .A2(n458), .ZN(n460) );
  NOR2_X1 U515 ( .A1(n494), .A2(n460), .ZN(n461) );
  NOR2_X1 U516 ( .A1(n462), .A2(n461), .ZN(n475) );
  NOR2_X1 U517 ( .A1(n544), .A2(n556), .ZN(n463) );
  XOR2_X1 U518 ( .A(KEYINPUT16), .B(n463), .Z(n464) );
  NOR2_X1 U519 ( .A1(n475), .A2(n464), .ZN(n492) );
  NAND2_X1 U520 ( .A1(n479), .A2(n492), .ZN(n465) );
  XNOR2_X1 U521 ( .A(KEYINPUT101), .B(n465), .ZN(n473) );
  NAND2_X1 U522 ( .A1(n473), .A2(n494), .ZN(n466) );
  XNOR2_X1 U523 ( .A(n466), .B(KEYINPUT34), .ZN(n467) );
  XNOR2_X1 U524 ( .A(G1GAT), .B(n467), .ZN(G1324GAT) );
  INV_X1 U525 ( .A(n509), .ZN(n497) );
  NAND2_X1 U526 ( .A1(n497), .A2(n473), .ZN(n468) );
  XNOR2_X1 U527 ( .A(n468), .B(KEYINPUT102), .ZN(n469) );
  XNOR2_X1 U528 ( .A(G8GAT), .B(n469), .ZN(G1325GAT) );
  XOR2_X1 U529 ( .A(KEYINPUT103), .B(KEYINPUT35), .Z(n471) );
  NAND2_X1 U530 ( .A1(n473), .A2(n522), .ZN(n470) );
  XNOR2_X1 U531 ( .A(n471), .B(n470), .ZN(n472) );
  XOR2_X1 U532 ( .A(G15GAT), .B(n472), .Z(G1326GAT) );
  NAND2_X1 U533 ( .A1(n521), .A2(n473), .ZN(n474) );
  XNOR2_X1 U534 ( .A(n474), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U535 ( .A(KEYINPUT38), .B(KEYINPUT105), .Z(n481) );
  NOR2_X1 U536 ( .A1(n577), .A2(n475), .ZN(n476) );
  NAND2_X1 U537 ( .A1(n544), .A2(n476), .ZN(n477) );
  XNOR2_X1 U538 ( .A(KEYINPUT37), .B(n477), .ZN(n478) );
  XNOR2_X1 U539 ( .A(KEYINPUT104), .B(n478), .ZN(n504) );
  NAND2_X1 U540 ( .A1(n479), .A2(n504), .ZN(n480) );
  XNOR2_X1 U541 ( .A(n481), .B(n480), .ZN(n489) );
  NOR2_X1 U542 ( .A1(n489), .A2(n506), .ZN(n482) );
  XNOR2_X1 U543 ( .A(n482), .B(KEYINPUT39), .ZN(n483) );
  XNOR2_X1 U544 ( .A(G29GAT), .B(n483), .ZN(G1328GAT) );
  NOR2_X1 U545 ( .A1(n509), .A2(n489), .ZN(n484) );
  XOR2_X1 U546 ( .A(KEYINPUT106), .B(n484), .Z(n485) );
  XNOR2_X1 U547 ( .A(G36GAT), .B(n485), .ZN(G1329GAT) );
  XNOR2_X1 U548 ( .A(KEYINPUT107), .B(KEYINPUT40), .ZN(n487) );
  NOR2_X1 U549 ( .A1(n512), .A2(n489), .ZN(n486) );
  XNOR2_X1 U550 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U551 ( .A(G43GAT), .B(n488), .ZN(G1330GAT) );
  INV_X1 U552 ( .A(n521), .ZN(n515) );
  NOR2_X1 U553 ( .A1(n515), .A2(n489), .ZN(n490) );
  XOR2_X1 U554 ( .A(G50GAT), .B(n490), .Z(n491) );
  XNOR2_X1 U555 ( .A(KEYINPUT108), .B(n491), .ZN(G1331GAT) );
  XNOR2_X1 U556 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n496) );
  INV_X1 U557 ( .A(n551), .ZN(n527) );
  NOR2_X1 U558 ( .A1(n564), .A2(n527), .ZN(n505) );
  NAND2_X1 U559 ( .A1(n505), .A2(n492), .ZN(n493) );
  XNOR2_X1 U560 ( .A(n493), .B(KEYINPUT109), .ZN(n501) );
  NAND2_X1 U561 ( .A1(n494), .A2(n501), .ZN(n495) );
  XNOR2_X1 U562 ( .A(n496), .B(n495), .ZN(G1332GAT) );
  NAND2_X1 U563 ( .A1(n497), .A2(n501), .ZN(n498) );
  XNOR2_X1 U564 ( .A(n498), .B(KEYINPUT110), .ZN(n499) );
  XNOR2_X1 U565 ( .A(G64GAT), .B(n499), .ZN(G1333GAT) );
  NAND2_X1 U566 ( .A1(n522), .A2(n501), .ZN(n500) );
  XNOR2_X1 U567 ( .A(n500), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U568 ( .A(G78GAT), .B(KEYINPUT43), .Z(n503) );
  NAND2_X1 U569 ( .A1(n501), .A2(n521), .ZN(n502) );
  XNOR2_X1 U570 ( .A(n503), .B(n502), .ZN(G1335GAT) );
  NAND2_X1 U571 ( .A1(n505), .A2(n504), .ZN(n514) );
  NOR2_X1 U572 ( .A1(n506), .A2(n514), .ZN(n508) );
  XNOR2_X1 U573 ( .A(G85GAT), .B(KEYINPUT111), .ZN(n507) );
  XNOR2_X1 U574 ( .A(n508), .B(n507), .ZN(G1336GAT) );
  NOR2_X1 U575 ( .A1(n509), .A2(n514), .ZN(n510) );
  XOR2_X1 U576 ( .A(KEYINPUT112), .B(n510), .Z(n511) );
  XNOR2_X1 U577 ( .A(G92GAT), .B(n511), .ZN(G1337GAT) );
  NOR2_X1 U578 ( .A1(n512), .A2(n514), .ZN(n513) );
  XOR2_X1 U579 ( .A(G99GAT), .B(n513), .Z(G1338GAT) );
  NOR2_X1 U580 ( .A1(n515), .A2(n514), .ZN(n516) );
  XOR2_X1 U581 ( .A(KEYINPUT44), .B(n516), .Z(n517) );
  XNOR2_X1 U582 ( .A(G106GAT), .B(n517), .ZN(G1339GAT) );
  NOR2_X1 U583 ( .A1(n519), .A2(n518), .ZN(n520) );
  XOR2_X1 U584 ( .A(KEYINPUT114), .B(n520), .Z(n539) );
  NOR2_X1 U585 ( .A1(n539), .A2(n521), .ZN(n523) );
  NAND2_X1 U586 ( .A1(n523), .A2(n522), .ZN(n534) );
  NOR2_X1 U587 ( .A1(n524), .A2(n534), .ZN(n526) );
  XNOR2_X1 U588 ( .A(G113GAT), .B(KEYINPUT115), .ZN(n525) );
  XNOR2_X1 U589 ( .A(n526), .B(n525), .ZN(G1340GAT) );
  NOR2_X1 U590 ( .A1(n527), .A2(n534), .ZN(n529) );
  XNOR2_X1 U591 ( .A(KEYINPUT49), .B(KEYINPUT116), .ZN(n528) );
  XNOR2_X1 U592 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U593 ( .A(G120GAT), .B(n530), .ZN(G1341GAT) );
  NOR2_X1 U594 ( .A1(n544), .A2(n534), .ZN(n532) );
  XNOR2_X1 U595 ( .A(KEYINPUT117), .B(KEYINPUT50), .ZN(n531) );
  XNOR2_X1 U596 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U597 ( .A(G127GAT), .B(n533), .ZN(G1342GAT) );
  NOR2_X1 U598 ( .A1(n535), .A2(n534), .ZN(n537) );
  XNOR2_X1 U599 ( .A(KEYINPUT118), .B(KEYINPUT51), .ZN(n536) );
  XNOR2_X1 U600 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U601 ( .A(G134GAT), .B(n538), .ZN(G1343GAT) );
  NOR2_X1 U602 ( .A1(n563), .A2(n539), .ZN(n546) );
  NAND2_X1 U603 ( .A1(n564), .A2(n546), .ZN(n540) );
  XNOR2_X1 U604 ( .A(G141GAT), .B(n540), .ZN(G1344GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n542) );
  NAND2_X1 U606 ( .A1(n546), .A2(n551), .ZN(n541) );
  XNOR2_X1 U607 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U608 ( .A(G148GAT), .B(n543), .ZN(G1345GAT) );
  INV_X1 U609 ( .A(n544), .ZN(n570) );
  NAND2_X1 U610 ( .A1(n570), .A2(n546), .ZN(n545) );
  XNOR2_X1 U611 ( .A(n545), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U612 ( .A1(n556), .A2(n546), .ZN(n547) );
  XNOR2_X1 U613 ( .A(n547), .B(G162GAT), .ZN(G1347GAT) );
  XOR2_X1 U614 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n549) );
  XNOR2_X1 U615 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n548) );
  XNOR2_X1 U616 ( .A(n549), .B(n548), .ZN(n550) );
  XOR2_X1 U617 ( .A(KEYINPUT56), .B(n550), .Z(n553) );
  NAND2_X1 U618 ( .A1(n555), .A2(n551), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n553), .B(n552), .ZN(G1349GAT) );
  NAND2_X1 U620 ( .A1(n570), .A2(n555), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n554), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U622 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U623 ( .A(n557), .B(KEYINPUT58), .ZN(n558) );
  XNOR2_X1 U624 ( .A(G190GAT), .B(n558), .ZN(G1351GAT) );
  XOR2_X1 U625 ( .A(KEYINPUT124), .B(KEYINPUT60), .Z(n560) );
  XNOR2_X1 U626 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(n561) );
  XOR2_X1 U628 ( .A(KEYINPUT123), .B(n561), .Z(n566) );
  NOR2_X1 U629 ( .A1(n563), .A2(n562), .ZN(n575) );
  NAND2_X1 U630 ( .A1(n575), .A2(n564), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n566), .B(n565), .ZN(G1352GAT) );
  XOR2_X1 U632 ( .A(G204GAT), .B(KEYINPUT61), .Z(n569) );
  NAND2_X1 U633 ( .A1(n575), .A2(n567), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n569), .B(n568), .ZN(G1353GAT) );
  XOR2_X1 U635 ( .A(G211GAT), .B(KEYINPUT125), .Z(n572) );
  NAND2_X1 U636 ( .A1(n575), .A2(n570), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(G1354GAT) );
  XOR2_X1 U638 ( .A(KEYINPUT126), .B(KEYINPUT127), .Z(n574) );
  XNOR2_X1 U639 ( .A(G218GAT), .B(KEYINPUT62), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(n579) );
  INV_X1 U641 ( .A(n575), .ZN(n576) );
  NOR2_X1 U642 ( .A1(n577), .A2(n576), .ZN(n578) );
  XOR2_X1 U643 ( .A(n579), .B(n578), .Z(G1355GAT) );
endmodule

