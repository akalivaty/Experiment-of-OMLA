

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585;

  XNOR2_X1 U326 ( .A(n384), .B(n383), .ZN(n551) );
  NOR2_X1 U327 ( .A1(n435), .A2(n524), .ZN(n568) );
  XNOR2_X1 U328 ( .A(n382), .B(n381), .ZN(n383) );
  INV_X1 U329 ( .A(G169GAT), .ZN(n455) );
  XOR2_X1 U330 ( .A(n467), .B(KEYINPUT28), .Z(n522) );
  XNOR2_X1 U331 ( .A(n455), .B(KEYINPUT120), .ZN(n456) );
  XNOR2_X1 U332 ( .A(n457), .B(n456), .ZN(G1348GAT) );
  XOR2_X1 U333 ( .A(KEYINPUT65), .B(KEYINPUT64), .Z(n295) );
  XNOR2_X1 U334 ( .A(G197GAT), .B(KEYINPUT29), .ZN(n294) );
  XNOR2_X1 U335 ( .A(n295), .B(n294), .ZN(n299) );
  XOR2_X1 U336 ( .A(G50GAT), .B(G36GAT), .Z(n297) );
  XOR2_X1 U337 ( .A(G113GAT), .B(G1GAT), .Z(n426) );
  XNOR2_X1 U338 ( .A(n426), .B(KEYINPUT66), .ZN(n296) );
  XNOR2_X1 U339 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U340 ( .A(n299), .B(n298), .Z(n301) );
  NAND2_X1 U341 ( .A1(G229GAT), .A2(G233GAT), .ZN(n300) );
  XNOR2_X1 U342 ( .A(n301), .B(n300), .ZN(n305) );
  XOR2_X1 U343 ( .A(G15GAT), .B(KEYINPUT67), .Z(n303) );
  XNOR2_X1 U344 ( .A(G169GAT), .B(G22GAT), .ZN(n302) );
  XNOR2_X1 U345 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U346 ( .A(n305), .B(n304), .Z(n313) );
  XOR2_X1 U347 ( .A(KEYINPUT8), .B(KEYINPUT7), .Z(n307) );
  XNOR2_X1 U348 ( .A(G43GAT), .B(G29GAT), .ZN(n306) );
  XNOR2_X1 U349 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U350 ( .A(KEYINPUT68), .B(n308), .ZN(n381) );
  XOR2_X1 U351 ( .A(KEYINPUT30), .B(G141GAT), .Z(n310) );
  XNOR2_X1 U352 ( .A(G8GAT), .B(KEYINPUT69), .ZN(n309) );
  XNOR2_X1 U353 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U354 ( .A(n381), .B(n311), .Z(n312) );
  XNOR2_X1 U355 ( .A(n313), .B(n312), .ZN(n569) );
  XOR2_X1 U356 ( .A(KEYINPUT21), .B(KEYINPUT89), .Z(n315) );
  XNOR2_X1 U357 ( .A(G197GAT), .B(G204GAT), .ZN(n314) );
  XNOR2_X1 U358 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U359 ( .A(G211GAT), .B(n316), .Z(n400) );
  XOR2_X1 U360 ( .A(G50GAT), .B(G162GAT), .Z(n368) );
  XOR2_X1 U361 ( .A(KEYINPUT2), .B(KEYINPUT3), .Z(n318) );
  XNOR2_X1 U362 ( .A(G141GAT), .B(KEYINPUT90), .ZN(n317) );
  XNOR2_X1 U363 ( .A(n318), .B(n317), .ZN(n413) );
  XOR2_X1 U364 ( .A(n368), .B(n413), .Z(n320) );
  NAND2_X1 U365 ( .A1(G228GAT), .A2(G233GAT), .ZN(n319) );
  XNOR2_X1 U366 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U367 ( .A(n400), .B(n321), .ZN(n332) );
  XOR2_X1 U368 ( .A(KEYINPUT91), .B(KEYINPUT22), .Z(n323) );
  XNOR2_X1 U369 ( .A(KEYINPUT92), .B(KEYINPUT23), .ZN(n322) );
  XNOR2_X1 U370 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U371 ( .A(G22GAT), .B(G155GAT), .Z(n344) );
  XOR2_X1 U372 ( .A(n324), .B(n344), .Z(n326) );
  XNOR2_X1 U373 ( .A(G218GAT), .B(G106GAT), .ZN(n325) );
  XNOR2_X1 U374 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U375 ( .A(n327), .B(KEYINPUT24), .Z(n330) );
  XNOR2_X1 U376 ( .A(G78GAT), .B(KEYINPUT72), .ZN(n328) );
  XNOR2_X1 U377 ( .A(n328), .B(G148GAT), .ZN(n351) );
  XNOR2_X1 U378 ( .A(n351), .B(KEYINPUT88), .ZN(n329) );
  XNOR2_X1 U379 ( .A(n330), .B(n329), .ZN(n331) );
  XNOR2_X1 U380 ( .A(n332), .B(n331), .ZN(n467) );
  XOR2_X1 U381 ( .A(KEYINPUT111), .B(KEYINPUT47), .Z(n387) );
  XOR2_X1 U382 ( .A(KEYINPUT12), .B(G211GAT), .Z(n334) );
  NAND2_X1 U383 ( .A1(G231GAT), .A2(G233GAT), .ZN(n333) );
  XNOR2_X1 U384 ( .A(n334), .B(n333), .ZN(n338) );
  XOR2_X1 U385 ( .A(KEYINPUT81), .B(KEYINPUT14), .Z(n336) );
  XNOR2_X1 U386 ( .A(KEYINPUT15), .B(KEYINPUT80), .ZN(n335) );
  XNOR2_X1 U387 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U388 ( .A(n338), .B(n337), .Z(n343) );
  XOR2_X1 U389 ( .A(G64GAT), .B(G78GAT), .Z(n340) );
  XNOR2_X1 U390 ( .A(G1GAT), .B(G8GAT), .ZN(n339) );
  XNOR2_X1 U391 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U392 ( .A(G183GAT), .B(n341), .ZN(n342) );
  XNOR2_X1 U393 ( .A(n343), .B(n342), .ZN(n345) );
  XOR2_X1 U394 ( .A(n345), .B(n344), .Z(n349) );
  XOR2_X1 U395 ( .A(G15GAT), .B(G127GAT), .Z(n440) );
  XOR2_X1 U396 ( .A(G57GAT), .B(KEYINPUT70), .Z(n347) );
  XNOR2_X1 U397 ( .A(G71GAT), .B(KEYINPUT13), .ZN(n346) );
  XNOR2_X1 U398 ( .A(n347), .B(n346), .ZN(n352) );
  XNOR2_X1 U399 ( .A(n440), .B(n352), .ZN(n348) );
  XOR2_X1 U400 ( .A(n349), .B(n348), .Z(n557) );
  INV_X1 U401 ( .A(n557), .ZN(n577) );
  XNOR2_X1 U402 ( .A(G99GAT), .B(G85GAT), .ZN(n350) );
  XNOR2_X1 U403 ( .A(n350), .B(G106GAT), .ZN(n380) );
  XNOR2_X1 U404 ( .A(n380), .B(n351), .ZN(n365) );
  XOR2_X1 U405 ( .A(G176GAT), .B(G64GAT), .Z(n397) );
  XOR2_X1 U406 ( .A(n397), .B(KEYINPUT73), .Z(n354) );
  XNOR2_X1 U407 ( .A(G92GAT), .B(n352), .ZN(n353) );
  XNOR2_X1 U408 ( .A(n354), .B(n353), .ZN(n358) );
  XOR2_X1 U409 ( .A(KEYINPUT32), .B(KEYINPUT71), .Z(n356) );
  NAND2_X1 U410 ( .A1(G230GAT), .A2(G233GAT), .ZN(n355) );
  XNOR2_X1 U411 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U412 ( .A(n358), .B(n357), .Z(n363) );
  XOR2_X1 U413 ( .A(KEYINPUT33), .B(G204GAT), .Z(n360) );
  XNOR2_X1 U414 ( .A(G120GAT), .B(KEYINPUT31), .ZN(n359) );
  XNOR2_X1 U415 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U416 ( .A(n361), .B(KEYINPUT74), .ZN(n362) );
  XNOR2_X1 U417 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U418 ( .A(n365), .B(n364), .ZN(n573) );
  XOR2_X1 U419 ( .A(KEYINPUT41), .B(n573), .Z(n497) );
  INV_X1 U420 ( .A(n497), .ZN(n553) );
  NOR2_X1 U421 ( .A1(n569), .A2(n553), .ZN(n366) );
  XNOR2_X1 U422 ( .A(n366), .B(KEYINPUT46), .ZN(n367) );
  NOR2_X1 U423 ( .A1(n577), .A2(n367), .ZN(n385) );
  XOR2_X1 U424 ( .A(KEYINPUT76), .B(KEYINPUT11), .Z(n370) );
  XOR2_X1 U425 ( .A(G134GAT), .B(KEYINPUT77), .Z(n425) );
  XNOR2_X1 U426 ( .A(n425), .B(n368), .ZN(n369) );
  XOR2_X1 U427 ( .A(n370), .B(n369), .Z(n374) );
  XOR2_X1 U428 ( .A(G218GAT), .B(G92GAT), .Z(n372) );
  XNOR2_X1 U429 ( .A(G190GAT), .B(KEYINPUT78), .ZN(n371) );
  XNOR2_X1 U430 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U431 ( .A(G36GAT), .B(n373), .Z(n407) );
  XNOR2_X1 U432 ( .A(n374), .B(n407), .ZN(n376) );
  NAND2_X1 U433 ( .A1(G232GAT), .A2(G233GAT), .ZN(n375) );
  XNOR2_X1 U434 ( .A(n376), .B(n375), .ZN(n377) );
  NAND2_X1 U435 ( .A1(n377), .A2(KEYINPUT9), .ZN(n379) );
  OR2_X1 U436 ( .A1(n377), .A2(KEYINPUT9), .ZN(n378) );
  NAND2_X1 U437 ( .A1(n379), .A2(n378), .ZN(n384) );
  XOR2_X1 U438 ( .A(n380), .B(KEYINPUT10), .Z(n382) );
  NAND2_X1 U439 ( .A1(n385), .A2(n551), .ZN(n386) );
  XNOR2_X1 U440 ( .A(n387), .B(n386), .ZN(n392) );
  XNOR2_X1 U441 ( .A(n551), .B(KEYINPUT79), .ZN(n560) );
  XNOR2_X1 U442 ( .A(KEYINPUT36), .B(n560), .ZN(n580) );
  NAND2_X1 U443 ( .A1(n577), .A2(n580), .ZN(n388) );
  XNOR2_X1 U444 ( .A(KEYINPUT45), .B(n388), .ZN(n389) );
  NOR2_X1 U445 ( .A1(n389), .A2(n573), .ZN(n390) );
  AND2_X1 U446 ( .A1(n569), .A2(n390), .ZN(n391) );
  NOR2_X1 U447 ( .A1(n392), .A2(n391), .ZN(n393) );
  XNOR2_X1 U448 ( .A(n393), .B(KEYINPUT48), .ZN(n526) );
  XOR2_X1 U449 ( .A(KEYINPUT97), .B(KEYINPUT98), .Z(n395) );
  XNOR2_X1 U450 ( .A(G8GAT), .B(KEYINPUT99), .ZN(n394) );
  XNOR2_X1 U451 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X1 U452 ( .A(n397), .B(n396), .Z(n399) );
  NAND2_X1 U453 ( .A1(G226GAT), .A2(G233GAT), .ZN(n398) );
  XNOR2_X1 U454 ( .A(n399), .B(n398), .ZN(n401) );
  XOR2_X1 U455 ( .A(n401), .B(n400), .Z(n409) );
  XOR2_X1 U456 ( .A(KEYINPUT85), .B(KEYINPUT19), .Z(n403) );
  XNOR2_X1 U457 ( .A(KEYINPUT17), .B(KEYINPUT86), .ZN(n402) );
  XNOR2_X1 U458 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U459 ( .A(n404), .B(G183GAT), .Z(n406) );
  XNOR2_X1 U460 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n405) );
  XNOR2_X1 U461 ( .A(n406), .B(n405), .ZN(n451) );
  XNOR2_X1 U462 ( .A(n451), .B(n407), .ZN(n408) );
  XNOR2_X1 U463 ( .A(n409), .B(n408), .ZN(n511) );
  XNOR2_X1 U464 ( .A(n511), .B(KEYINPUT119), .ZN(n410) );
  NOR2_X1 U465 ( .A1(n526), .A2(n410), .ZN(n411) );
  XOR2_X1 U466 ( .A(KEYINPUT54), .B(n411), .Z(n435) );
  XNOR2_X1 U467 ( .A(G120GAT), .B(KEYINPUT0), .ZN(n412) );
  XNOR2_X1 U468 ( .A(n412), .B(KEYINPUT82), .ZN(n443) );
  XNOR2_X1 U469 ( .A(n443), .B(n413), .ZN(n434) );
  XOR2_X1 U470 ( .A(KEYINPUT93), .B(G155GAT), .Z(n415) );
  XNOR2_X1 U471 ( .A(G127GAT), .B(G57GAT), .ZN(n414) );
  XNOR2_X1 U472 ( .A(n415), .B(n414), .ZN(n419) );
  XOR2_X1 U473 ( .A(KEYINPUT5), .B(KEYINPUT4), .Z(n417) );
  XNOR2_X1 U474 ( .A(KEYINPUT6), .B(KEYINPUT1), .ZN(n416) );
  XNOR2_X1 U475 ( .A(n417), .B(n416), .ZN(n418) );
  XOR2_X1 U476 ( .A(n419), .B(n418), .Z(n424) );
  XOR2_X1 U477 ( .A(KEYINPUT94), .B(KEYINPUT96), .Z(n421) );
  NAND2_X1 U478 ( .A1(G225GAT), .A2(G233GAT), .ZN(n420) );
  XNOR2_X1 U479 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U480 ( .A(KEYINPUT95), .B(n422), .ZN(n423) );
  XNOR2_X1 U481 ( .A(n424), .B(n423), .ZN(n430) );
  XOR2_X1 U482 ( .A(G162GAT), .B(n425), .Z(n428) );
  XNOR2_X1 U483 ( .A(n426), .B(G85GAT), .ZN(n427) );
  XNOR2_X1 U484 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U485 ( .A(n430), .B(n429), .Z(n432) );
  XNOR2_X1 U486 ( .A(G29GAT), .B(G148GAT), .ZN(n431) );
  XNOR2_X1 U487 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U488 ( .A(n434), .B(n433), .ZN(n524) );
  NAND2_X1 U489 ( .A1(n467), .A2(n568), .ZN(n436) );
  XNOR2_X1 U490 ( .A(KEYINPUT55), .B(n436), .ZN(n454) );
  XOR2_X1 U491 ( .A(G176GAT), .B(G134GAT), .Z(n438) );
  XNOR2_X1 U492 ( .A(G113GAT), .B(G190GAT), .ZN(n437) );
  XNOR2_X1 U493 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U494 ( .A(n439), .B(G99GAT), .Z(n442) );
  XNOR2_X1 U495 ( .A(G43GAT), .B(n440), .ZN(n441) );
  XNOR2_X1 U496 ( .A(n442), .B(n441), .ZN(n447) );
  XOR2_X1 U497 ( .A(KEYINPUT84), .B(n443), .Z(n445) );
  NAND2_X1 U498 ( .A1(G227GAT), .A2(G233GAT), .ZN(n444) );
  XNOR2_X1 U499 ( .A(n445), .B(n444), .ZN(n446) );
  XOR2_X1 U500 ( .A(n447), .B(n446), .Z(n453) );
  XOR2_X1 U501 ( .A(KEYINPUT87), .B(KEYINPUT83), .Z(n449) );
  XNOR2_X1 U502 ( .A(G71GAT), .B(KEYINPUT20), .ZN(n448) );
  XNOR2_X1 U503 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U504 ( .A(n451), .B(n450), .ZN(n452) );
  XOR2_X1 U505 ( .A(n453), .B(n452), .Z(n521) );
  INV_X1 U506 ( .A(n521), .ZN(n514) );
  NAND2_X1 U507 ( .A1(n454), .A2(n514), .ZN(n559) );
  NOR2_X1 U508 ( .A1(n569), .A2(n559), .ZN(n457) );
  NOR2_X1 U509 ( .A1(n569), .A2(n573), .ZN(n458) );
  XNOR2_X1 U510 ( .A(KEYINPUT75), .B(n458), .ZN(n486) );
  NOR2_X1 U511 ( .A1(n557), .A2(n560), .ZN(n459) );
  XNOR2_X1 U512 ( .A(KEYINPUT16), .B(n459), .ZN(n473) );
  NAND2_X1 U513 ( .A1(n514), .A2(n511), .ZN(n460) );
  NAND2_X1 U514 ( .A1(n467), .A2(n460), .ZN(n461) );
  XOR2_X1 U515 ( .A(KEYINPUT25), .B(n461), .Z(n466) );
  XNOR2_X1 U516 ( .A(n511), .B(KEYINPUT27), .ZN(n523) );
  NOR2_X1 U517 ( .A1(n467), .A2(n514), .ZN(n462) );
  XNOR2_X1 U518 ( .A(n462), .B(KEYINPUT26), .ZN(n567) );
  NAND2_X1 U519 ( .A1(n523), .A2(n567), .ZN(n463) );
  XOR2_X1 U520 ( .A(KEYINPUT100), .B(n463), .Z(n464) );
  NOR2_X1 U521 ( .A1(n524), .A2(n464), .ZN(n465) );
  NAND2_X1 U522 ( .A1(n466), .A2(n465), .ZN(n471) );
  NOR2_X1 U523 ( .A1(n514), .A2(n522), .ZN(n468) );
  NAND2_X1 U524 ( .A1(n468), .A2(n523), .ZN(n469) );
  NAND2_X1 U525 ( .A1(n524), .A2(n469), .ZN(n470) );
  NAND2_X1 U526 ( .A1(n471), .A2(n470), .ZN(n472) );
  XNOR2_X1 U527 ( .A(KEYINPUT101), .B(n472), .ZN(n483) );
  NAND2_X1 U528 ( .A1(n473), .A2(n483), .ZN(n498) );
  NOR2_X1 U529 ( .A1(n486), .A2(n498), .ZN(n481) );
  NAND2_X1 U530 ( .A1(n481), .A2(n524), .ZN(n476) );
  XNOR2_X1 U531 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n474) );
  XNOR2_X1 U532 ( .A(n474), .B(KEYINPUT102), .ZN(n475) );
  XNOR2_X1 U533 ( .A(n476), .B(n475), .ZN(G1324GAT) );
  XOR2_X1 U534 ( .A(G8GAT), .B(KEYINPUT103), .Z(n478) );
  NAND2_X1 U535 ( .A1(n481), .A2(n511), .ZN(n477) );
  XNOR2_X1 U536 ( .A(n478), .B(n477), .ZN(G1325GAT) );
  XOR2_X1 U537 ( .A(G15GAT), .B(KEYINPUT35), .Z(n480) );
  NAND2_X1 U538 ( .A1(n481), .A2(n514), .ZN(n479) );
  XNOR2_X1 U539 ( .A(n480), .B(n479), .ZN(G1326GAT) );
  NAND2_X1 U540 ( .A1(n481), .A2(n522), .ZN(n482) );
  XNOR2_X1 U541 ( .A(n482), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U542 ( .A(G29GAT), .B(KEYINPUT39), .Z(n491) );
  NAND2_X1 U543 ( .A1(n580), .A2(n483), .ZN(n484) );
  NOR2_X1 U544 ( .A1(n577), .A2(n484), .ZN(n485) );
  XNOR2_X1 U545 ( .A(KEYINPUT37), .B(n485), .ZN(n509) );
  OR2_X1 U546 ( .A1(n486), .A2(n509), .ZN(n489) );
  XNOR2_X1 U547 ( .A(KEYINPUT104), .B(KEYINPUT105), .ZN(n487) );
  XNOR2_X1 U548 ( .A(n487), .B(KEYINPUT38), .ZN(n488) );
  XNOR2_X1 U549 ( .A(n489), .B(n488), .ZN(n495) );
  NAND2_X1 U550 ( .A1(n495), .A2(n524), .ZN(n490) );
  XNOR2_X1 U551 ( .A(n491), .B(n490), .ZN(G1328GAT) );
  NAND2_X1 U552 ( .A1(n495), .A2(n511), .ZN(n492) );
  XNOR2_X1 U553 ( .A(n492), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U554 ( .A1(n495), .A2(n514), .ZN(n493) );
  XNOR2_X1 U555 ( .A(n493), .B(KEYINPUT40), .ZN(n494) );
  XNOR2_X1 U556 ( .A(G43GAT), .B(n494), .ZN(G1330GAT) );
  NAND2_X1 U557 ( .A1(n495), .A2(n522), .ZN(n496) );
  XNOR2_X1 U558 ( .A(n496), .B(G50GAT), .ZN(G1331GAT) );
  NAND2_X1 U559 ( .A1(n569), .A2(n497), .ZN(n508) );
  NOR2_X1 U560 ( .A1(n508), .A2(n498), .ZN(n499) );
  XNOR2_X1 U561 ( .A(KEYINPUT106), .B(n499), .ZN(n505) );
  NAND2_X1 U562 ( .A1(n524), .A2(n505), .ZN(n500) );
  XNOR2_X1 U563 ( .A(KEYINPUT42), .B(n500), .ZN(n501) );
  XNOR2_X1 U564 ( .A(G57GAT), .B(n501), .ZN(G1332GAT) );
  XOR2_X1 U565 ( .A(G64GAT), .B(KEYINPUT107), .Z(n503) );
  NAND2_X1 U566 ( .A1(n511), .A2(n505), .ZN(n502) );
  XNOR2_X1 U567 ( .A(n503), .B(n502), .ZN(G1333GAT) );
  NAND2_X1 U568 ( .A1(n505), .A2(n514), .ZN(n504) );
  XNOR2_X1 U569 ( .A(n504), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U570 ( .A(G78GAT), .B(KEYINPUT43), .Z(n507) );
  NAND2_X1 U571 ( .A1(n522), .A2(n505), .ZN(n506) );
  XNOR2_X1 U572 ( .A(n507), .B(n506), .ZN(G1335GAT) );
  NOR2_X1 U573 ( .A1(n509), .A2(n508), .ZN(n516) );
  NAND2_X1 U574 ( .A1(n524), .A2(n516), .ZN(n510) );
  XNOR2_X1 U575 ( .A(G85GAT), .B(n510), .ZN(G1336GAT) );
  NAND2_X1 U576 ( .A1(n516), .A2(n511), .ZN(n512) );
  XNOR2_X1 U577 ( .A(n512), .B(KEYINPUT108), .ZN(n513) );
  XNOR2_X1 U578 ( .A(G92GAT), .B(n513), .ZN(G1337GAT) );
  NAND2_X1 U579 ( .A1(n516), .A2(n514), .ZN(n515) );
  XNOR2_X1 U580 ( .A(n515), .B(G99GAT), .ZN(G1338GAT) );
  XNOR2_X1 U581 ( .A(G106GAT), .B(KEYINPUT109), .ZN(n520) );
  XOR2_X1 U582 ( .A(KEYINPUT44), .B(KEYINPUT110), .Z(n518) );
  NAND2_X1 U583 ( .A1(n516), .A2(n522), .ZN(n517) );
  XNOR2_X1 U584 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X1 U585 ( .A(n520), .B(n519), .ZN(G1339GAT) );
  NOR2_X1 U586 ( .A1(n522), .A2(n521), .ZN(n528) );
  NAND2_X1 U587 ( .A1(n524), .A2(n523), .ZN(n525) );
  NOR2_X1 U588 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U589 ( .A(KEYINPUT112), .B(n527), .ZN(n541) );
  NAND2_X1 U590 ( .A1(n528), .A2(n541), .ZN(n537) );
  NOR2_X1 U591 ( .A1(n569), .A2(n537), .ZN(n530) );
  XNOR2_X1 U592 ( .A(G113GAT), .B(KEYINPUT113), .ZN(n529) );
  XNOR2_X1 U593 ( .A(n530), .B(n529), .ZN(G1340GAT) );
  NOR2_X1 U594 ( .A1(n553), .A2(n537), .ZN(n532) );
  XNOR2_X1 U595 ( .A(KEYINPUT114), .B(KEYINPUT49), .ZN(n531) );
  XNOR2_X1 U596 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U597 ( .A(G120GAT), .B(n533), .ZN(G1341GAT) );
  NOR2_X1 U598 ( .A1(n557), .A2(n537), .ZN(n535) );
  XNOR2_X1 U599 ( .A(KEYINPUT50), .B(KEYINPUT115), .ZN(n534) );
  XNOR2_X1 U600 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U601 ( .A(G127GAT), .B(n536), .ZN(G1342GAT) );
  XOR2_X1 U602 ( .A(G134GAT), .B(KEYINPUT51), .Z(n540) );
  INV_X1 U603 ( .A(n537), .ZN(n538) );
  NAND2_X1 U604 ( .A1(n538), .A2(n560), .ZN(n539) );
  XNOR2_X1 U605 ( .A(n540), .B(n539), .ZN(G1343GAT) );
  XNOR2_X1 U606 ( .A(KEYINPUT117), .B(KEYINPUT118), .ZN(n544) );
  NAND2_X1 U607 ( .A1(n541), .A2(n567), .ZN(n542) );
  XNOR2_X1 U608 ( .A(n542), .B(KEYINPUT116), .ZN(n550) );
  NOR2_X1 U609 ( .A1(n569), .A2(n550), .ZN(n543) );
  XNOR2_X1 U610 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U611 ( .A(G141GAT), .B(n545), .ZN(G1344GAT) );
  NOR2_X1 U612 ( .A1(n550), .A2(n553), .ZN(n547) );
  XNOR2_X1 U613 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n546) );
  XNOR2_X1 U614 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U615 ( .A(G148GAT), .B(n548), .ZN(G1345GAT) );
  NOR2_X1 U616 ( .A1(n550), .A2(n557), .ZN(n549) );
  XOR2_X1 U617 ( .A(G155GAT), .B(n549), .Z(G1346GAT) );
  NOR2_X1 U618 ( .A1(n551), .A2(n550), .ZN(n552) );
  XOR2_X1 U619 ( .A(G162GAT), .B(n552), .Z(G1347GAT) );
  NOR2_X1 U620 ( .A1(n553), .A2(n559), .ZN(n555) );
  XNOR2_X1 U621 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U623 ( .A(G176GAT), .B(n556), .ZN(G1349GAT) );
  NOR2_X1 U624 ( .A1(n557), .A2(n559), .ZN(n558) );
  XOR2_X1 U625 ( .A(G183GAT), .B(n558), .Z(G1350GAT) );
  XOR2_X1 U626 ( .A(KEYINPUT121), .B(KEYINPUT58), .Z(n563) );
  INV_X1 U627 ( .A(n559), .ZN(n561) );
  NAND2_X1 U628 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n563), .B(n562), .ZN(n564) );
  XNOR2_X1 U630 ( .A(G190GAT), .B(n564), .ZN(G1351GAT) );
  XOR2_X1 U631 ( .A(KEYINPUT60), .B(KEYINPUT122), .Z(n566) );
  XNOR2_X1 U632 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n565) );
  XNOR2_X1 U633 ( .A(n566), .B(n565), .ZN(n571) );
  NAND2_X1 U634 ( .A1(n568), .A2(n567), .ZN(n572) );
  NOR2_X1 U635 ( .A1(n569), .A2(n572), .ZN(n570) );
  XOR2_X1 U636 ( .A(n571), .B(n570), .Z(G1352GAT) );
  XOR2_X1 U637 ( .A(KEYINPUT123), .B(KEYINPUT61), .Z(n575) );
  INV_X1 U638 ( .A(n572), .ZN(n581) );
  NAND2_X1 U639 ( .A1(n581), .A2(n573), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(n576) );
  XOR2_X1 U641 ( .A(G204GAT), .B(n576), .Z(G1353GAT) );
  NAND2_X1 U642 ( .A1(n581), .A2(n577), .ZN(n578) );
  XNOR2_X1 U643 ( .A(n578), .B(KEYINPUT124), .ZN(n579) );
  XNOR2_X1 U644 ( .A(G211GAT), .B(n579), .ZN(G1354GAT) );
  XNOR2_X1 U645 ( .A(G218GAT), .B(KEYINPUT125), .ZN(n585) );
  XOR2_X1 U646 ( .A(KEYINPUT126), .B(KEYINPUT62), .Z(n583) );
  NAND2_X1 U647 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n585), .B(n584), .ZN(G1355GAT) );
endmodule

