//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 0 0 0 0 1 0 0 1 1 0 0 0 1 1 1 1 1 0 0 0 1 1 1 0 0 0 1 1 1 1 1 1 1 1 1 1 0 0 0 0 0 0 0 0 0 1 1 1 0 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:22 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n935, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007;
  XOR2_X1   g000(.A(KEYINPUT9), .B(G234), .Z(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  OAI21_X1  g002(.A(G221), .B1(new_n188), .B2(G902), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  XNOR2_X1  g004(.A(G110), .B(G140), .ZN(new_n191));
  INV_X1    g005(.A(G227), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n192), .A2(G953), .ZN(new_n193));
  XOR2_X1   g007(.A(new_n191), .B(new_n193), .Z(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT11), .ZN(new_n196));
  INV_X1    g010(.A(G134), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n196), .B1(new_n197), .B2(G137), .ZN(new_n198));
  INV_X1    g012(.A(G137), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n199), .A2(KEYINPUT11), .A3(G134), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n197), .A2(G137), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n198), .A2(new_n200), .A3(new_n201), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n202), .A2(KEYINPUT64), .A3(G131), .ZN(new_n203));
  NAND2_X1  g017(.A1(KEYINPUT64), .A2(G131), .ZN(new_n204));
  NAND4_X1  g018(.A1(new_n198), .A2(new_n200), .A3(new_n204), .A4(new_n201), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT73), .ZN(new_n208));
  INV_X1    g022(.A(G104), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT74), .ZN(new_n211));
  INV_X1    g025(.A(G107), .ZN(new_n212));
  NAND2_X1  g026(.A1(KEYINPUT73), .A2(G104), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n210), .A2(new_n211), .A3(new_n212), .A4(new_n213), .ZN(new_n214));
  OAI21_X1  g028(.A(KEYINPUT75), .B1(new_n212), .B2(G104), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT75), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n216), .A2(new_n209), .A3(G107), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n214), .A2(new_n215), .A3(new_n217), .ZN(new_n218));
  AND2_X1   g032(.A1(KEYINPUT73), .A2(G104), .ZN(new_n219));
  NOR2_X1   g033(.A1(KEYINPUT73), .A2(G104), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n211), .B1(new_n221), .B2(new_n212), .ZN(new_n222));
  OAI21_X1  g036(.A(G101), .B1(new_n218), .B2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G143), .ZN(new_n224));
  OAI21_X1  g038(.A(KEYINPUT1), .B1(new_n224), .B2(G146), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n224), .A2(G146), .ZN(new_n226));
  INV_X1    g040(.A(G146), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n227), .A2(G143), .ZN(new_n228));
  OAI211_X1 g042(.A(G128), .B(new_n225), .C1(new_n226), .C2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n227), .A2(G143), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n224), .A2(G146), .ZN(new_n231));
  INV_X1    g045(.A(G128), .ZN(new_n232));
  OAI211_X1 g046(.A(new_n230), .B(new_n231), .C1(KEYINPUT1), .C2(new_n232), .ZN(new_n233));
  AND2_X1   g047(.A1(new_n229), .A2(new_n233), .ZN(new_n234));
  OAI22_X1  g048(.A1(new_n219), .A2(new_n220), .B1(KEYINPUT3), .B2(G107), .ZN(new_n235));
  INV_X1    g049(.A(G101), .ZN(new_n236));
  NAND2_X1  g050(.A1(KEYINPUT3), .A2(G107), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT3), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n238), .A2(new_n212), .A3(G104), .ZN(new_n239));
  NAND4_X1  g053(.A1(new_n235), .A2(new_n236), .A3(new_n237), .A4(new_n239), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n223), .A2(KEYINPUT10), .A3(new_n234), .A4(new_n240), .ZN(new_n241));
  AOI22_X1  g055(.A1(new_n210), .A2(new_n213), .B1(new_n238), .B2(new_n212), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n239), .A2(new_n237), .ZN(new_n243));
  OAI21_X1  g057(.A(G101), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n244), .A2(KEYINPUT4), .A3(new_n240), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n230), .A2(new_n231), .A3(KEYINPUT0), .A4(G128), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n226), .A2(new_n228), .ZN(new_n247));
  XNOR2_X1  g061(.A(KEYINPUT0), .B(G128), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n246), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n251));
  OAI211_X1 g065(.A(new_n251), .B(G101), .C1(new_n242), .C2(new_n243), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n245), .A2(new_n250), .A3(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n241), .A2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT76), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n223), .A2(new_n234), .A3(new_n240), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT10), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n254), .B1(new_n255), .B2(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n256), .A2(KEYINPUT76), .A3(new_n257), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n207), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n258), .A2(new_n255), .ZN(new_n262));
  AND2_X1   g076(.A1(new_n241), .A2(new_n253), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n262), .A2(new_n263), .A3(new_n207), .A4(new_n260), .ZN(new_n264));
  INV_X1    g078(.A(new_n264), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n195), .B1(new_n261), .B2(new_n265), .ZN(new_n266));
  AND3_X1   g080(.A1(new_n223), .A2(new_n234), .A3(new_n240), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n234), .B1(new_n223), .B2(new_n240), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n206), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(KEYINPUT12), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n229), .A2(new_n233), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n215), .A2(new_n217), .ZN(new_n272));
  NOR3_X1   g086(.A1(new_n219), .A2(new_n220), .A3(G107), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n272), .B1(new_n273), .B2(new_n211), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n221), .A2(new_n212), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(KEYINPUT74), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n236), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n240), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n271), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(new_n256), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT12), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n280), .A2(new_n281), .A3(new_n206), .ZN(new_n282));
  NAND4_X1  g096(.A1(new_n264), .A2(new_n194), .A3(new_n270), .A4(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(KEYINPUT77), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n281), .B1(new_n280), .B2(new_n206), .ZN(new_n285));
  AOI211_X1 g099(.A(KEYINPUT12), .B(new_n207), .C1(new_n279), .C2(new_n256), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT77), .ZN(new_n288));
  NAND4_X1  g102(.A1(new_n287), .A2(new_n288), .A3(new_n194), .A4(new_n264), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n266), .A2(new_n284), .A3(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(G469), .ZN(new_n291));
  INV_X1    g105(.A(G902), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n290), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT78), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND4_X1  g109(.A1(new_n290), .A2(KEYINPUT78), .A3(new_n291), .A4(new_n292), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n287), .A2(new_n264), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(new_n195), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n262), .A2(new_n263), .A3(new_n260), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(new_n206), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(new_n264), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n299), .B1(new_n195), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(new_n292), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(G469), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n190), .B1(new_n297), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n249), .A2(G125), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n307), .B1(new_n234), .B2(G125), .ZN(new_n308));
  INV_X1    g122(.A(G224), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n309), .A2(G953), .ZN(new_n310));
  XNOR2_X1  g124(.A(new_n310), .B(KEYINPUT80), .ZN(new_n311));
  XNOR2_X1  g125(.A(new_n308), .B(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT67), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT66), .ZN(new_n314));
  INV_X1    g128(.A(G119), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n314), .B1(new_n315), .B2(G116), .ZN(new_n316));
  INV_X1    g130(.A(G116), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n317), .A2(KEYINPUT66), .A3(G119), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n317), .A2(G119), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  AND2_X1   g135(.A1(KEYINPUT2), .A2(G113), .ZN(new_n322));
  NOR2_X1   g136(.A1(KEYINPUT2), .A2(G113), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  AND3_X1   g138(.A1(new_n319), .A2(new_n321), .A3(new_n324), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n324), .B1(new_n319), .B2(new_n321), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n313), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  AND3_X1   g141(.A1(new_n317), .A2(KEYINPUT66), .A3(G119), .ZN(new_n328));
  AOI21_X1  g142(.A(KEYINPUT66), .B1(new_n317), .B2(G119), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n321), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(new_n324), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n320), .B1(new_n316), .B2(new_n318), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(new_n324), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n332), .A2(KEYINPUT67), .A3(new_n334), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n327), .A2(new_n335), .A3(new_n245), .A4(new_n252), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n333), .A2(KEYINPUT5), .ZN(new_n337));
  INV_X1    g151(.A(G113), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT5), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n338), .B1(new_n320), .B2(new_n339), .ZN(new_n340));
  AOI22_X1  g154(.A1(new_n337), .A2(new_n340), .B1(new_n333), .B2(new_n324), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n341), .A2(new_n240), .A3(new_n223), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n336), .A2(new_n342), .ZN(new_n343));
  XNOR2_X1  g157(.A(G110), .B(G122), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n336), .A2(new_n342), .A3(new_n344), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n346), .A2(KEYINPUT6), .A3(new_n347), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n344), .B1(new_n336), .B2(new_n342), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT79), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT6), .ZN(new_n351));
  AND3_X1   g165(.A1(new_n349), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n350), .B1(new_n349), .B2(new_n351), .ZN(new_n353));
  OAI211_X1 g167(.A(new_n312), .B(new_n348), .C1(new_n352), .C2(new_n353), .ZN(new_n354));
  XNOR2_X1  g168(.A(new_n344), .B(KEYINPUT8), .ZN(new_n355));
  INV_X1    g169(.A(new_n342), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n341), .B1(new_n240), .B2(new_n223), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n355), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT7), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n310), .A2(new_n359), .ZN(new_n360));
  XNOR2_X1  g174(.A(new_n308), .B(new_n360), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n358), .A2(new_n361), .A3(new_n347), .ZN(new_n362));
  AND2_X1   g176(.A1(new_n362), .A2(new_n292), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n354), .A2(new_n363), .ZN(new_n364));
  OAI21_X1  g178(.A(G210), .B1(G237), .B2(G902), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT81), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n354), .A2(new_n363), .A3(new_n365), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n367), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  OAI21_X1  g184(.A(G214), .B1(G237), .B2(G902), .ZN(new_n371));
  AND3_X1   g185(.A1(new_n354), .A2(new_n365), .A3(new_n363), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(KEYINPUT81), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n370), .A2(new_n371), .A3(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(G475), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT16), .ZN(new_n376));
  INV_X1    g190(.A(G140), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n376), .A2(new_n377), .A3(G125), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(G125), .ZN(new_n379));
  INV_X1    g193(.A(G125), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(G140), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n378), .B1(new_n382), .B2(new_n376), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(new_n227), .ZN(new_n384));
  NOR2_X1   g198(.A1(G237), .A2(G953), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(G214), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT82), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n386), .A2(new_n387), .A3(G143), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(G143), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n224), .A2(KEYINPUT82), .ZN(new_n390));
  NAND4_X1  g204(.A1(new_n389), .A2(new_n390), .A3(G214), .A4(new_n385), .ZN(new_n391));
  NAND4_X1  g205(.A1(new_n388), .A2(new_n391), .A3(KEYINPUT17), .A4(G131), .ZN(new_n392));
  OAI211_X1 g206(.A(G146), .B(new_n378), .C1(new_n382), .C2(new_n376), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n384), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT83), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n384), .A2(new_n392), .A3(KEYINPUT83), .A4(new_n393), .ZN(new_n397));
  AOI21_X1  g211(.A(G131), .B1(new_n388), .B2(new_n391), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT17), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n388), .A2(new_n391), .A3(G131), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n399), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n396), .A2(new_n397), .A3(new_n402), .ZN(new_n403));
  OAI21_X1  g217(.A(KEYINPUT69), .B1(new_n382), .B2(G146), .ZN(new_n404));
  XNOR2_X1  g218(.A(G125), .B(G140), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT69), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n405), .A2(new_n406), .A3(new_n227), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n408), .B1(new_n227), .B2(new_n405), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n388), .A2(new_n391), .A3(KEYINPUT18), .A4(G131), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n388), .A2(new_n391), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT18), .ZN(new_n412));
  INV_X1    g226(.A(G131), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n411), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n409), .A2(new_n410), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n403), .A2(new_n415), .ZN(new_n416));
  XNOR2_X1  g230(.A(G113), .B(G122), .ZN(new_n417));
  XNOR2_X1  g231(.A(new_n417), .B(new_n209), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n416), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n403), .A2(new_n418), .A3(new_n415), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n375), .B1(new_n422), .B2(new_n292), .ZN(new_n423));
  OR2_X1    g237(.A1(new_n382), .A2(KEYINPUT19), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n382), .A2(KEYINPUT19), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n424), .A2(new_n227), .A3(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(new_n401), .ZN(new_n427));
  OAI211_X1 g241(.A(new_n426), .B(new_n393), .C1(new_n427), .C2(new_n398), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n415), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(new_n419), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n421), .A2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT20), .ZN(new_n432));
  NOR2_X1   g246(.A1(G475), .A2(G902), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n431), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n432), .B1(new_n431), .B2(new_n433), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT84), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n434), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND4_X1  g251(.A1(new_n431), .A2(KEYINPUT84), .A3(new_n432), .A4(new_n433), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n423), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(G234), .A2(G237), .ZN(new_n440));
  INV_X1    g254(.A(G953), .ZN(new_n441));
  AND3_X1   g255(.A1(new_n440), .A2(G952), .A3(new_n441), .ZN(new_n442));
  XOR2_X1   g256(.A(KEYINPUT21), .B(G898), .Z(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  AND3_X1   g258(.A1(new_n440), .A2(G902), .A3(G953), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n442), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n224), .A2(KEYINPUT13), .A3(G128), .ZN(new_n448));
  AOI21_X1  g262(.A(KEYINPUT13), .B1(new_n224), .B2(G128), .ZN(new_n449));
  OAI221_X1 g263(.A(new_n448), .B1(G128), .B2(new_n224), .C1(new_n449), .C2(KEYINPUT85), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(KEYINPUT85), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  OAI21_X1  g266(.A(G134), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(G122), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(G116), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n317), .A2(G122), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(G107), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n455), .A2(new_n456), .A3(new_n212), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n232), .A2(G143), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n224), .A2(G128), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  AOI22_X1  g276(.A1(new_n458), .A2(new_n459), .B1(new_n462), .B2(new_n197), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n453), .A2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT86), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n453), .A2(KEYINPUT86), .A3(new_n463), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT14), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n468), .B1(new_n317), .B2(G122), .ZN(new_n469));
  OR2_X1    g283(.A1(new_n469), .A2(KEYINPUT87), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n469), .A2(KEYINPUT87), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n468), .A2(new_n317), .A3(G122), .ZN(new_n472));
  NAND4_X1  g286(.A1(new_n470), .A2(new_n471), .A3(new_n455), .A4(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(G107), .ZN(new_n474));
  INV_X1    g288(.A(new_n459), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n462), .A2(new_n197), .ZN(new_n476));
  OAI21_X1  g290(.A(G134), .B1(new_n460), .B2(new_n461), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n475), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n474), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n466), .A2(new_n467), .A3(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(G217), .ZN(new_n481));
  NOR3_X1   g295(.A1(new_n188), .A2(new_n481), .A3(G953), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  AOI22_X1  g298(.A1(new_n464), .A2(new_n465), .B1(new_n474), .B2(new_n478), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n482), .B1(new_n485), .B2(new_n467), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n292), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(G478), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n488), .A2(KEYINPUT15), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  OAI221_X1 g304(.A(new_n292), .B1(KEYINPUT15), .B2(new_n488), .C1(new_n484), .C2(new_n486), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n439), .A2(new_n447), .A3(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT88), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n439), .A2(KEYINPUT88), .A3(new_n447), .A4(new_n493), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n374), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  AND2_X1   g312(.A1(new_n306), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n384), .A2(new_n393), .ZN(new_n500));
  XOR2_X1   g314(.A(KEYINPUT24), .B(G110), .Z(new_n501));
  XNOR2_X1  g315(.A(G119), .B(G128), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT23), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n504), .B1(G119), .B2(new_n232), .ZN(new_n505));
  NOR3_X1   g319(.A1(new_n315), .A2(KEYINPUT23), .A3(G128), .ZN(new_n506));
  OAI22_X1  g320(.A1(new_n505), .A2(new_n506), .B1(G119), .B2(new_n232), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(G110), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n500), .A2(new_n503), .A3(new_n508), .ZN(new_n509));
  OAI22_X1  g323(.A1(new_n507), .A2(G110), .B1(new_n502), .B2(new_n501), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n510), .A2(new_n393), .A3(new_n408), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  XNOR2_X1  g326(.A(KEYINPUT22), .B(G137), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n441), .A2(G221), .A3(G234), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n513), .B(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n512), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n509), .A2(new_n511), .A3(new_n515), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n517), .A2(new_n292), .A3(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT70), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT25), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n481), .B1(G234), .B2(new_n292), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n519), .A2(new_n520), .A3(KEYINPUT25), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  AND2_X1   g340(.A1(new_n517), .A2(new_n518), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n524), .A2(G902), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n528), .B(KEYINPUT71), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n526), .A2(new_n530), .ZN(new_n531));
  XNOR2_X1  g345(.A(new_n531), .B(KEYINPUT72), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT32), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT31), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n327), .A2(new_n335), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n206), .A2(new_n250), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n202), .A2(new_n413), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n413), .B1(G134), .B2(new_n199), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(new_n201), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n234), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n535), .A2(new_n536), .A3(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n536), .A2(new_n541), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(KEYINPUT30), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT30), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT65), .ZN(new_n547));
  AOI22_X1  g361(.A1(new_n202), .A2(new_n413), .B1(new_n201), .B2(new_n538), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n234), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n540), .A2(KEYINPUT65), .ZN(new_n550));
  OAI211_X1 g364(.A(new_n546), .B(new_n536), .C1(new_n549), .C2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n545), .A2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n535), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n543), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n385), .A2(G210), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n555), .B(new_n236), .ZN(new_n556));
  XNOR2_X1  g370(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n556), .B(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n534), .B1(new_n554), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n540), .A2(KEYINPUT65), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n548), .A2(new_n547), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n561), .A2(new_n234), .A3(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n535), .B1(new_n563), .B2(new_n536), .ZN(new_n564));
  OAI21_X1  g378(.A(KEYINPUT28), .B1(new_n543), .B2(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n249), .B1(new_n203), .B2(new_n205), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n548), .A2(new_n271), .ZN(new_n567));
  OAI21_X1  g381(.A(KEYINPUT68), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT68), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n536), .A2(new_n541), .A3(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n568), .A2(new_n570), .A3(new_n535), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT28), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n559), .B1(new_n565), .B2(new_n573), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n535), .B1(new_n545), .B2(new_n551), .ZN(new_n575));
  NOR4_X1   g389(.A1(new_n575), .A2(new_n543), .A3(KEYINPUT31), .A4(new_n558), .ZN(new_n576));
  NOR3_X1   g390(.A1(new_n560), .A2(new_n574), .A3(new_n576), .ZN(new_n577));
  NOR2_X1   g391(.A1(G472), .A2(G902), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n533), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n554), .A2(new_n559), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(KEYINPUT31), .ZN(new_n582));
  INV_X1    g396(.A(new_n574), .ZN(new_n583));
  INV_X1    g397(.A(new_n576), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n585), .A2(KEYINPUT32), .A3(new_n578), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n565), .A2(new_n573), .A3(new_n559), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT29), .ZN(new_n588));
  OAI211_X1 g402(.A(new_n587), .B(new_n588), .C1(new_n559), .C2(new_n554), .ZN(new_n589));
  AND2_X1   g403(.A1(new_n571), .A2(new_n572), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n553), .A2(new_n544), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n572), .B1(new_n591), .B2(new_n542), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n558), .A2(new_n588), .ZN(new_n594));
  AOI21_X1  g408(.A(G902), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n589), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(G472), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n580), .A2(new_n586), .A3(new_n597), .ZN(new_n598));
  AND2_X1   g412(.A1(new_n532), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n499), .A2(new_n599), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n600), .B(G101), .ZN(G3));
  XOR2_X1   g415(.A(new_n531), .B(KEYINPUT72), .Z(new_n602));
  OAI21_X1  g416(.A(G472), .B1(new_n577), .B2(G902), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n603), .B1(new_n577), .B2(new_n579), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(new_n306), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n365), .B1(new_n354), .B2(new_n363), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n371), .B1(new_n372), .B2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT89), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT33), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n612), .B1(new_n484), .B2(new_n486), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n480), .A2(new_n483), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n485), .A2(new_n467), .A3(new_n482), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n614), .A2(KEYINPUT33), .A3(new_n615), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n488), .A2(G902), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n613), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n487), .A2(new_n488), .ZN(new_n619));
  AND2_X1   g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NOR3_X1   g434(.A1(new_n439), .A2(new_n446), .A3(new_n620), .ZN(new_n621));
  OAI211_X1 g435(.A(KEYINPUT89), .B(new_n371), .C1(new_n372), .C2(new_n608), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n611), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(KEYINPUT90), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT90), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n611), .A2(new_n621), .A3(new_n625), .A4(new_n622), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n607), .A2(new_n627), .ZN(new_n628));
  XOR2_X1   g442(.A(KEYINPUT34), .B(G104), .Z(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(G6));
  XOR2_X1   g444(.A(new_n446), .B(KEYINPUT91), .Z(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n423), .B1(new_n490), .B2(new_n491), .ZN(new_n633));
  INV_X1    g447(.A(new_n435), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(new_n434), .ZN(new_n635));
  AND2_X1   g449(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  AND4_X1   g450(.A1(new_n611), .A2(new_n622), .A3(new_n632), .A4(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n607), .A2(new_n637), .ZN(new_n638));
  XOR2_X1   g452(.A(KEYINPUT35), .B(G107), .Z(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G9));
  NOR2_X1   g454(.A1(new_n516), .A2(KEYINPUT36), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n512), .B(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(new_n529), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n526), .A2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n604), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n499), .A2(new_n646), .ZN(new_n647));
  XOR2_X1   g461(.A(KEYINPUT37), .B(G110), .Z(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G12));
  AND4_X1   g463(.A1(new_n598), .A2(new_n611), .A3(new_n622), .A4(new_n644), .ZN(new_n650));
  AND2_X1   g464(.A1(new_n650), .A2(new_n306), .ZN(new_n651));
  INV_X1    g465(.A(G900), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n442), .B1(new_n445), .B2(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  AND2_X1   g468(.A1(new_n636), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n651), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(G128), .ZN(G30));
  NOR2_X1   g471(.A1(new_n439), .A2(new_n493), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n658), .A2(new_n371), .A3(new_n645), .ZN(new_n659));
  XOR2_X1   g473(.A(new_n659), .B(KEYINPUT94), .Z(new_n660));
  AOI21_X1  g474(.A(new_n559), .B1(new_n591), .B2(new_n542), .ZN(new_n661));
  OR2_X1    g475(.A1(new_n661), .A2(KEYINPUT92), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n661), .A2(KEYINPUT92), .ZN(new_n663));
  AND3_X1   g477(.A1(new_n662), .A2(new_n581), .A3(new_n663), .ZN(new_n664));
  OAI21_X1  g478(.A(G472), .B1(new_n664), .B2(G902), .ZN(new_n665));
  AND3_X1   g479(.A1(new_n580), .A2(new_n586), .A3(new_n665), .ZN(new_n666));
  XOR2_X1   g480(.A(new_n666), .B(KEYINPUT93), .Z(new_n667));
  NAND2_X1  g481(.A1(new_n370), .A2(new_n373), .ZN(new_n668));
  XOR2_X1   g482(.A(new_n668), .B(KEYINPUT38), .Z(new_n669));
  NAND3_X1  g483(.A1(new_n660), .A2(new_n667), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(KEYINPUT95), .ZN(new_n671));
  XOR2_X1   g485(.A(new_n653), .B(KEYINPUT39), .Z(new_n672));
  NAND2_X1  g486(.A1(new_n306), .A2(new_n672), .ZN(new_n673));
  OR2_X1    g487(.A1(new_n673), .A2(KEYINPUT40), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n673), .A2(KEYINPUT40), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n671), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G143), .ZN(G45));
  NAND2_X1  g491(.A1(new_n437), .A2(new_n438), .ZN(new_n678));
  INV_X1    g492(.A(new_n423), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(new_n620), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n680), .A2(new_n681), .A3(new_n654), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n651), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G146), .ZN(G48));
  AOI21_X1  g499(.A(new_n291), .B1(new_n290), .B2(new_n292), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  AOI22_X1  g501(.A1(new_n302), .A2(new_n195), .B1(new_n283), .B2(KEYINPUT77), .ZN(new_n688));
  AOI21_X1  g502(.A(G902), .B1(new_n688), .B2(new_n289), .ZN(new_n689));
  AOI21_X1  g503(.A(KEYINPUT78), .B1(new_n689), .B2(new_n291), .ZN(new_n690));
  INV_X1    g504(.A(new_n296), .ZN(new_n691));
  OAI211_X1 g505(.A(new_n189), .B(new_n687), .C1(new_n690), .C2(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n532), .A2(new_n598), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n627), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(KEYINPUT41), .B(G113), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n695), .B(new_n696), .ZN(G15));
  NAND2_X1  g511(.A1(new_n694), .A2(new_n637), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G116), .ZN(G18));
  NAND2_X1  g513(.A1(new_n496), .A2(new_n497), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n700), .A2(new_n598), .A3(new_n644), .ZN(new_n701));
  AOI211_X1 g515(.A(new_n190), .B(new_n686), .C1(new_n295), .C2(new_n296), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT96), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n611), .A2(new_n622), .ZN(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n702), .A2(new_n703), .A3(new_n705), .ZN(new_n706));
  OAI21_X1  g520(.A(KEYINPUT96), .B1(new_n692), .B2(new_n704), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n701), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(new_n315), .ZN(G21));
  INV_X1    g523(.A(G472), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n710), .B1(new_n585), .B2(new_n292), .ZN(new_n711));
  XOR2_X1   g525(.A(new_n578), .B(KEYINPUT97), .Z(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n593), .A2(KEYINPUT98), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT98), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n715), .B1(new_n590), .B2(new_n592), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n714), .A2(new_n716), .A3(new_n558), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n560), .A2(new_n576), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n713), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NOR3_X1   g533(.A1(new_n711), .A2(new_n719), .A3(new_n531), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(new_n658), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n611), .A2(new_n622), .A3(new_n632), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(new_n702), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G122), .ZN(G24));
  NOR3_X1   g539(.A1(new_n711), .A2(new_n719), .A3(new_n645), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n620), .B1(new_n678), .B2(new_n679), .ZN(new_n727));
  AOI21_X1  g541(.A(KEYINPUT99), .B1(new_n727), .B2(new_n654), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT99), .ZN(new_n729));
  NOR4_X1   g543(.A1(new_n439), .A2(new_n620), .A3(new_n729), .A4(new_n653), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n726), .B1(new_n728), .B2(new_n730), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n731), .B1(new_n706), .B2(new_n707), .ZN(new_n732));
  XOR2_X1   g546(.A(KEYINPUT100), .B(G125), .Z(new_n733));
  XNOR2_X1  g547(.A(new_n732), .B(new_n733), .ZN(G27));
  NAND2_X1  g548(.A1(new_n682), .A2(new_n729), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n727), .A2(KEYINPUT99), .A3(new_n654), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(new_n531), .ZN(new_n738));
  AND3_X1   g552(.A1(new_n598), .A2(KEYINPUT101), .A3(new_n738), .ZN(new_n739));
  AOI21_X1  g553(.A(KEYINPUT101), .B1(new_n598), .B2(new_n738), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n737), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n668), .A2(new_n371), .ZN(new_n742));
  INV_X1    g556(.A(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n306), .A2(new_n743), .ZN(new_n744));
  OAI21_X1  g558(.A(KEYINPUT42), .B1(new_n741), .B2(new_n744), .ZN(new_n745));
  AOI22_X1  g559(.A1(new_n295), .A2(new_n296), .B1(G469), .B2(new_n304), .ZN(new_n746));
  NOR3_X1   g560(.A1(new_n746), .A2(new_n742), .A3(new_n190), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT42), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n747), .A2(new_n748), .A3(new_n599), .A4(new_n737), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n745), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(new_n413), .ZN(G33));
  NAND3_X1  g565(.A1(new_n747), .A2(new_n599), .A3(new_n655), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G134), .ZN(G36));
  NOR2_X1   g567(.A1(new_n291), .A2(new_n292), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT45), .ZN(new_n755));
  OR2_X1    g569(.A1(new_n303), .A2(new_n755), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n291), .B1(new_n303), .B2(new_n755), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n754), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(KEYINPUT46), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(new_n297), .ZN(new_n760));
  OAI22_X1  g574(.A1(new_n760), .A2(KEYINPUT102), .B1(KEYINPUT46), .B2(new_n758), .ZN(new_n761));
  AND2_X1   g575(.A1(new_n760), .A2(KEYINPUT102), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n189), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n439), .A2(new_n681), .ZN(new_n765));
  NAND2_X1  g579(.A1(KEYINPUT103), .A2(KEYINPUT43), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  XOR2_X1   g581(.A(KEYINPUT103), .B(KEYINPUT43), .Z(new_n768));
  OAI21_X1  g582(.A(new_n767), .B1(new_n765), .B2(new_n768), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n769), .A2(new_n604), .A3(new_n644), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT44), .ZN(new_n771));
  AND2_X1   g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n770), .A2(new_n771), .ZN(new_n773));
  NOR3_X1   g587(.A1(new_n772), .A2(new_n773), .A3(new_n742), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n764), .A2(new_n672), .A3(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(KEYINPUT104), .B(G137), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n775), .B(new_n776), .ZN(G39));
  INV_X1    g591(.A(KEYINPUT105), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n763), .B1(new_n778), .B2(KEYINPUT47), .ZN(new_n779));
  NOR4_X1   g593(.A1(new_n742), .A2(new_n532), .A3(new_n598), .A4(new_n682), .ZN(new_n780));
  XNOR2_X1  g594(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n781));
  OAI211_X1 g595(.A(new_n779), .B(new_n780), .C1(new_n763), .C2(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G140), .ZN(G42));
  INV_X1    g597(.A(KEYINPUT112), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n769), .A2(new_n442), .A3(new_n720), .ZN(new_n785));
  OR2_X1    g599(.A1(new_n785), .A2(new_n742), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n779), .B1(new_n763), .B2(new_n781), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n297), .A2(new_n687), .ZN(new_n788));
  XOR2_X1   g602(.A(new_n788), .B(KEYINPUT106), .Z(new_n789));
  NAND2_X1  g603(.A1(new_n789), .A2(new_n190), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n786), .B1(new_n787), .B2(new_n790), .ZN(new_n791));
  NOR4_X1   g605(.A1(new_n669), .A2(new_n785), .A3(new_n371), .A4(new_n692), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(KEYINPUT50), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n702), .A2(KEYINPUT113), .A3(new_n743), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(new_n442), .ZN(new_n795));
  AOI21_X1  g609(.A(KEYINPUT113), .B1(new_n702), .B2(new_n743), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n797), .A2(new_n726), .A3(new_n769), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n667), .A2(new_n602), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n797), .A2(new_n439), .A3(new_n620), .A4(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n793), .A2(new_n798), .A3(new_n800), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n784), .B1(new_n791), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n802), .A2(KEYINPUT51), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT51), .ZN(new_n804));
  OAI211_X1 g618(.A(new_n784), .B(new_n804), .C1(new_n791), .C2(new_n801), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n739), .A2(new_n740), .ZN(new_n806));
  INV_X1    g620(.A(new_n806), .ZN(new_n807));
  AND3_X1   g621(.A1(new_n797), .A2(new_n807), .A3(new_n769), .ZN(new_n808));
  XOR2_X1   g622(.A(KEYINPUT114), .B(KEYINPUT48), .Z(new_n809));
  OR2_X1    g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  AND3_X1   g624(.A1(new_n797), .A2(new_n727), .A3(new_n799), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n441), .A2(G952), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n785), .B1(new_n706), .B2(new_n707), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n811), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n808), .A2(new_n809), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n810), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT115), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  OR2_X1    g632(.A1(new_n816), .A2(new_n817), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n803), .A2(new_n805), .A3(new_n818), .A4(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT54), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n695), .A2(new_n698), .A3(new_n724), .ZN(new_n822));
  AND3_X1   g636(.A1(new_n370), .A2(new_n371), .A3(new_n373), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT107), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n823), .A2(new_n824), .A3(new_n727), .A4(new_n632), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n370), .A2(new_n371), .A3(new_n373), .A4(new_n632), .ZN(new_n826));
  INV_X1    g640(.A(new_n727), .ZN(new_n827));
  OAI21_X1  g641(.A(KEYINPUT107), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n825), .A2(new_n605), .A3(new_n306), .A4(new_n828), .ZN(new_n829));
  OAI211_X1 g643(.A(new_n306), .B(new_n498), .C1(new_n599), .C2(new_n646), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT108), .ZN(new_n831));
  AND3_X1   g645(.A1(new_n678), .A2(new_n633), .A3(new_n831), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n831), .B1(new_n678), .B2(new_n633), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n834), .A2(new_n826), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n306), .A2(new_n605), .A3(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n829), .A2(new_n830), .A3(new_n836), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n822), .A2(new_n837), .A3(new_n708), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n492), .A2(new_n423), .A3(new_n653), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n598), .A2(new_n635), .A3(new_n644), .A4(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n731), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n841), .A2(new_n747), .ZN(new_n842));
  AND4_X1   g656(.A1(new_n745), .A2(new_n749), .A3(new_n752), .A4(new_n842), .ZN(new_n843));
  AOI21_X1  g657(.A(KEYINPUT109), .B1(new_n838), .B2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(new_n731), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n703), .B1(new_n702), .B2(new_n705), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n692), .A2(KEYINPUT96), .A3(new_n704), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n845), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  OAI211_X1 g662(.A(new_n650), .B(new_n306), .C1(new_n655), .C2(new_n683), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n644), .A2(new_n653), .ZN(new_n850));
  XNOR2_X1  g664(.A(new_n850), .B(KEYINPUT110), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n851), .A2(new_n666), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n704), .A2(new_n439), .A3(new_n493), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n852), .A2(new_n853), .A3(new_n306), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n848), .A2(new_n849), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(KEYINPUT52), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT52), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n848), .A2(new_n857), .A3(new_n849), .A4(new_n854), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n844), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n838), .A2(KEYINPUT109), .A3(new_n843), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n860), .A2(KEYINPUT53), .A3(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(new_n849), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n732), .A2(new_n863), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n857), .B1(new_n864), .B2(new_n854), .ZN(new_n865));
  INV_X1    g679(.A(new_n858), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT109), .ZN(new_n868));
  AND3_X1   g682(.A1(new_n829), .A2(new_n830), .A3(new_n836), .ZN(new_n869));
  INV_X1    g683(.A(new_n701), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n870), .B1(new_n846), .B2(new_n847), .ZN(new_n871));
  AOI22_X1  g685(.A1(new_n627), .A2(new_n694), .B1(new_n723), .B2(new_n702), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n869), .A2(new_n698), .A3(new_n871), .A4(new_n872), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n745), .A2(new_n749), .A3(new_n752), .A4(new_n842), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n868), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n867), .A2(new_n875), .A3(new_n861), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT53), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n821), .B1(new_n862), .B2(new_n878), .ZN(new_n879));
  AOI21_X1  g693(.A(KEYINPUT53), .B1(new_n860), .B2(new_n861), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT111), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n881), .B1(new_n822), .B2(new_n708), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n877), .B1(new_n841), .B2(new_n747), .ZN(new_n883));
  AND4_X1   g697(.A1(new_n745), .A2(new_n883), .A3(new_n749), .A4(new_n752), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n871), .A2(new_n872), .A3(KEYINPUT111), .A4(new_n698), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n882), .A2(new_n884), .A3(new_n869), .A4(new_n885), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n886), .A2(new_n859), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n880), .A2(KEYINPUT54), .A3(new_n887), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n820), .A2(new_n879), .A3(new_n888), .ZN(new_n889));
  NOR2_X1   g703(.A1(G952), .A2(G953), .ZN(new_n890));
  INV_X1    g704(.A(new_n789), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n891), .A2(KEYINPUT49), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n891), .A2(KEYINPUT49), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n738), .A2(new_n189), .A3(new_n371), .ZN(new_n894));
  NOR4_X1   g708(.A1(new_n667), .A2(new_n669), .A3(new_n765), .A4(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  OAI22_X1  g710(.A1(new_n889), .A2(new_n890), .B1(new_n892), .B2(new_n896), .ZN(G75));
  INV_X1    g711(.A(KEYINPUT118), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n898), .A2(KEYINPUT56), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n348), .B1(new_n352), .B2(new_n353), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n900), .B(new_n312), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(KEYINPUT55), .ZN(new_n902));
  MUX2_X1   g716(.A(new_n898), .B(new_n899), .S(new_n902), .Z(new_n903));
  INV_X1    g717(.A(KEYINPUT117), .ZN(new_n904));
  INV_X1    g718(.A(new_n887), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n292), .B1(new_n878), .B2(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n904), .B1(new_n906), .B2(G210), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n887), .B1(new_n876), .B2(new_n877), .ZN(new_n908));
  INV_X1    g722(.A(G210), .ZN(new_n909));
  NOR4_X1   g723(.A1(new_n908), .A2(KEYINPUT117), .A3(new_n909), .A4(new_n292), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n903), .B1(new_n907), .B2(new_n910), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n441), .A2(G952), .ZN(new_n912));
  INV_X1    g726(.A(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  NOR3_X1   g728(.A1(new_n908), .A2(new_n909), .A3(new_n292), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT116), .ZN(new_n916));
  AOI21_X1  g730(.A(KEYINPUT56), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  OAI21_X1  g731(.A(G902), .B1(new_n880), .B2(new_n887), .ZN(new_n918));
  OAI21_X1  g732(.A(KEYINPUT116), .B1(new_n918), .B2(new_n909), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n902), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n914), .A2(new_n920), .ZN(G51));
  INV_X1    g735(.A(KEYINPUT119), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n922), .B1(new_n908), .B2(new_n821), .ZN(new_n923));
  OAI21_X1  g737(.A(KEYINPUT54), .B1(new_n880), .B2(new_n887), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  OAI211_X1 g739(.A(new_n922), .B(KEYINPUT54), .C1(new_n880), .C2(new_n887), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n754), .B(KEYINPUT57), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n925), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(new_n290), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n906), .A2(new_n756), .A3(new_n757), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n912), .B1(new_n929), .B2(new_n930), .ZN(G54));
  NAND2_X1  g745(.A1(KEYINPUT58), .A2(G475), .ZN(new_n932));
  XOR2_X1   g746(.A(new_n932), .B(KEYINPUT120), .Z(new_n933));
  NOR2_X1   g747(.A1(new_n918), .A2(new_n933), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n913), .B1(new_n934), .B2(new_n431), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n935), .B1(new_n431), .B2(new_n934), .ZN(G60));
  XNOR2_X1  g750(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n937));
  NAND2_X1  g751(.A1(G478), .A2(G902), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n937), .B(new_n938), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n939), .B1(new_n888), .B2(new_n879), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n613), .A2(new_n616), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n912), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(new_n941), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n925), .A2(new_n926), .A3(new_n943), .A4(new_n939), .ZN(new_n944));
  AND2_X1   g758(.A1(new_n942), .A2(new_n944), .ZN(G63));
  NAND2_X1  g759(.A1(G217), .A2(G902), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n946), .B(KEYINPUT60), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n908), .A2(new_n947), .ZN(new_n948));
  OR2_X1    g762(.A1(new_n948), .A2(new_n527), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n948), .A2(new_n642), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n949), .A2(new_n913), .A3(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT61), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n949), .A2(KEYINPUT61), .A3(new_n913), .A4(new_n950), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n953), .A2(new_n954), .ZN(G66));
  NOR2_X1   g769(.A1(new_n838), .A2(G953), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n956), .B(KEYINPUT122), .ZN(new_n957));
  OAI21_X1  g771(.A(G953), .B1(new_n444), .B2(new_n309), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n900), .B1(G898), .B2(new_n441), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n959), .B(new_n960), .ZN(G69));
  NAND2_X1  g775(.A1(new_n807), .A2(new_n853), .ZN(new_n962));
  INV_X1    g776(.A(new_n962), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n764), .A2(new_n672), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(KEYINPUT126), .ZN(new_n965));
  INV_X1    g779(.A(new_n750), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT126), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n764), .A2(new_n967), .A3(new_n672), .A4(new_n963), .ZN(new_n968));
  NAND4_X1  g782(.A1(new_n965), .A2(new_n966), .A3(new_n752), .A4(new_n968), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n864), .B(KEYINPUT124), .Z(new_n970));
  NAND3_X1  g784(.A1(new_n782), .A2(new_n970), .A3(new_n775), .ZN(new_n971));
  OR2_X1    g785(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n972), .A2(new_n441), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n424), .A2(new_n425), .ZN(new_n974));
  XOR2_X1   g788(.A(new_n974), .B(KEYINPUT123), .Z(new_n975));
  XNOR2_X1  g789(.A(new_n552), .B(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(new_n976), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n977), .B1(new_n652), .B2(G953), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n973), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n970), .A2(new_n676), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT62), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n981), .A2(KEYINPUT125), .ZN(new_n982));
  OR2_X1    g796(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n981), .A2(KEYINPUT125), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n982), .B1(new_n980), .B2(new_n984), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n742), .B1(new_n827), .B2(new_n834), .ZN(new_n986));
  NAND4_X1  g800(.A1(new_n986), .A2(new_n599), .A3(new_n306), .A4(new_n672), .ZN(new_n987));
  AND3_X1   g801(.A1(new_n782), .A2(new_n775), .A3(new_n987), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n983), .A2(new_n985), .A3(new_n988), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n989), .A2(new_n441), .A3(new_n977), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n979), .A2(new_n990), .ZN(new_n991));
  OAI21_X1  g805(.A(G953), .B1(new_n192), .B2(new_n652), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  INV_X1    g807(.A(new_n992), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n979), .A2(new_n990), .A3(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n993), .A2(new_n995), .ZN(G72));
  NAND2_X1  g810(.A1(G472), .A2(G902), .ZN(new_n997));
  XOR2_X1   g811(.A(new_n997), .B(KEYINPUT63), .Z(new_n998));
  OAI21_X1  g812(.A(new_n998), .B1(new_n972), .B2(new_n873), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n554), .A2(new_n558), .ZN(new_n1000));
  XOR2_X1   g814(.A(new_n1000), .B(KEYINPUT127), .Z(new_n1001));
  AND2_X1   g815(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n559), .B1(new_n575), .B2(new_n543), .ZN(new_n1003));
  NAND4_X1  g817(.A1(new_n983), .A2(new_n985), .A3(new_n838), .A4(new_n988), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n1003), .B1(new_n1004), .B2(new_n998), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n1000), .A2(new_n998), .A3(new_n1003), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n1006), .B1(new_n862), .B2(new_n878), .ZN(new_n1007));
  NOR4_X1   g821(.A1(new_n1002), .A2(new_n1005), .A3(new_n912), .A4(new_n1007), .ZN(G57));
endmodule


