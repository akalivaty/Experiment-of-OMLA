//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 0 0 1 0 0 0 0 1 1 0 0 0 0 0 0 1 0 1 0 1 1 1 1 1 1 1 1 0 0 1 0 1 0 0 1 0 1 0 1 1 0 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:11 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n546, new_n548, new_n549, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n562,
    new_n563, new_n564, new_n566, new_n567, new_n568, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n597, new_n598, new_n601, new_n602, new_n604, new_n605,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1152, new_n1153;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT65), .ZN(new_n437));
  INV_X1    g012(.A(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n437), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT66), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  XNOR2_X1  g037(.A(KEYINPUT3), .B(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G125), .ZN(new_n464));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  XNOR2_X1  g040(.A(new_n465), .B(KEYINPUT67), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(G101), .A2(G2104), .ZN(new_n469));
  INV_X1    g044(.A(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(KEYINPUT3), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT3), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(G137), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n469), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  AND2_X1   g053(.A1(new_n468), .A2(new_n478), .ZN(G160));
  OAI21_X1  g054(.A(KEYINPUT68), .B1(new_n474), .B2(new_n477), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT68), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n463), .A2(new_n481), .A3(G2105), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n474), .A2(G2105), .ZN(new_n484));
  AOI22_X1  g059(.A1(new_n483), .A2(G124), .B1(G136), .B2(new_n484), .ZN(new_n485));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n477), .ZN(new_n487));
  AND2_X1   g062(.A1(new_n485), .A2(new_n487), .ZN(G162));
  NOR2_X1   g063(.A1(new_n470), .A2(G2105), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G102), .ZN(new_n490));
  INV_X1    g065(.A(G114), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n491), .A2(new_n470), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n492), .B1(new_n463), .B2(G126), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n490), .B1(new_n493), .B2(new_n477), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n471), .A2(new_n473), .A3(G138), .A4(new_n477), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n463), .A2(KEYINPUT4), .A3(G138), .A4(new_n477), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n494), .A2(new_n499), .ZN(G164));
  XNOR2_X1  g075(.A(KEYINPUT69), .B(G651), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G75), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n501), .A2(KEYINPUT6), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT6), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G651), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(G50), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n503), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n502), .A2(G62), .ZN(new_n511));
  INV_X1    g086(.A(G88), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n511), .B1(new_n507), .B2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(KEYINPUT5), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT5), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G543), .ZN(new_n517));
  AND2_X1   g092(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n513), .A2(new_n518), .ZN(new_n519));
  AND2_X1   g094(.A1(new_n510), .A2(new_n519), .ZN(G166));
  NOR2_X1   g095(.A1(new_n507), .A2(new_n514), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G51), .ZN(new_n522));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  XNOR2_X1  g098(.A(new_n523), .B(KEYINPUT7), .ZN(new_n524));
  INV_X1    g099(.A(new_n507), .ZN(new_n525));
  AOI22_X1  g100(.A1(new_n525), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n515), .A2(new_n517), .ZN(new_n527));
  OAI211_X1 g102(.A(new_n522), .B(new_n524), .C1(new_n526), .C2(new_n527), .ZN(G286));
  INV_X1    g103(.A(G286), .ZN(G168));
  NAND2_X1  g104(.A1(G77), .A2(G543), .ZN(new_n530));
  INV_X1    g105(.A(G64), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n530), .B1(new_n527), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(new_n502), .ZN(new_n533));
  XOR2_X1   g108(.A(new_n533), .B(KEYINPUT70), .Z(new_n534));
  NOR2_X1   g109(.A1(new_n507), .A2(new_n527), .ZN(new_n535));
  AOI22_X1  g110(.A1(G52), .A2(new_n521), .B1(new_n535), .B2(G90), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n534), .A2(new_n536), .ZN(G301));
  INV_X1    g112(.A(G301), .ZN(G171));
  NAND2_X1  g113(.A1(new_n535), .A2(G81), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n521), .A2(G43), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n518), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n541));
  OR2_X1    g116(.A1(new_n541), .A2(new_n501), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n539), .A2(new_n540), .A3(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G860), .ZN(G153));
  AND3_X1   g120(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G36), .ZN(G176));
  NAND2_X1  g122(.A1(G1), .A2(G3), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT8), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n546), .A2(new_n549), .ZN(G188));
  NAND2_X1  g125(.A1(G78), .A2(G543), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT71), .ZN(new_n552));
  INV_X1    g127(.A(G65), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n552), .B1(new_n553), .B2(new_n527), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n535), .A2(G91), .B1(G651), .B2(new_n554), .ZN(new_n555));
  NAND4_X1  g130(.A1(new_n504), .A2(G53), .A3(G543), .A4(new_n506), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT9), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  OR2_X1    g133(.A1(new_n556), .A2(new_n557), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n555), .A2(new_n558), .A3(new_n559), .ZN(G299));
  NAND2_X1  g135(.A1(new_n510), .A2(new_n519), .ZN(G303));
  NAND2_X1  g136(.A1(new_n521), .A2(G49), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n535), .A2(G87), .ZN(new_n563));
  OAI21_X1  g138(.A(G651), .B1(new_n518), .B2(G74), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(G288));
  NAND4_X1  g140(.A1(new_n504), .A2(G86), .A3(new_n506), .A4(new_n518), .ZN(new_n566));
  NAND4_X1  g141(.A1(new_n504), .A2(G48), .A3(G543), .A4(new_n506), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n518), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n568));
  OAI211_X1 g143(.A(new_n566), .B(new_n567), .C1(new_n568), .C2(new_n501), .ZN(G305));
  AOI22_X1  g144(.A1(new_n518), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n570));
  NOR2_X1   g145(.A1(new_n570), .A2(new_n501), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n571), .B(KEYINPUT72), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n535), .A2(G85), .ZN(new_n574));
  INV_X1    g149(.A(G47), .ZN(new_n575));
  INV_X1    g150(.A(new_n521), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n574), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n573), .A2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(new_n578), .ZN(G290));
  INV_X1    g154(.A(KEYINPUT10), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT73), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n535), .A2(new_n581), .A3(G92), .ZN(new_n582));
  INV_X1    g157(.A(new_n582), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n581), .B1(new_n535), .B2(G92), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n580), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(new_n584), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n586), .A2(KEYINPUT10), .A3(new_n582), .ZN(new_n587));
  NAND2_X1  g162(.A1(G79), .A2(G543), .ZN(new_n588));
  INV_X1    g163(.A(G66), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n527), .B2(new_n589), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n521), .A2(G54), .B1(G651), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n585), .A2(new_n587), .A3(new_n591), .ZN(new_n592));
  XOR2_X1   g167(.A(new_n592), .B(KEYINPUT74), .Z(new_n593));
  NOR2_X1   g168(.A1(new_n593), .A2(G868), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n594), .B1(G868), .B2(G171), .ZN(G284));
  AOI21_X1  g170(.A(new_n594), .B1(G868), .B2(G171), .ZN(G321));
  NAND2_X1  g171(.A1(G286), .A2(G868), .ZN(new_n597));
  INV_X1    g172(.A(G299), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n598), .B2(G868), .ZN(G297));
  OAI21_X1  g174(.A(new_n597), .B1(new_n598), .B2(G868), .ZN(G280));
  XNOR2_X1  g175(.A(new_n592), .B(KEYINPUT74), .ZN(new_n601));
  INV_X1    g176(.A(G559), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n602), .B2(G860), .ZN(G148));
  NAND2_X1  g178(.A1(new_n601), .A2(new_n602), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n604), .A2(G868), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n605), .B1(G868), .B2(new_n544), .ZN(G323));
  XNOR2_X1  g181(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g182(.A(new_n483), .ZN(new_n608));
  INV_X1    g183(.A(G123), .ZN(new_n609));
  OR3_X1    g184(.A1(new_n608), .A2(KEYINPUT75), .A3(new_n609), .ZN(new_n610));
  OR2_X1    g185(.A1(G99), .A2(G2105), .ZN(new_n611));
  INV_X1    g186(.A(G111), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n470), .B1(new_n612), .B2(G2105), .ZN(new_n613));
  AOI22_X1  g188(.A1(new_n484), .A2(G135), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  OAI21_X1  g189(.A(KEYINPUT75), .B1(new_n608), .B2(new_n609), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n610), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  XOR2_X1   g191(.A(new_n616), .B(G2096), .Z(new_n617));
  NAND2_X1  g192(.A1(new_n463), .A2(new_n489), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT12), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT13), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(G2100), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n617), .A2(new_n621), .ZN(G156));
  XOR2_X1   g197(.A(KEYINPUT15), .B(G2435), .Z(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(G2438), .ZN(new_n624));
  XOR2_X1   g199(.A(G2427), .B(G2430), .Z(new_n625));
  NOR2_X1   g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  XOR2_X1   g201(.A(KEYINPUT76), .B(KEYINPUT14), .Z(new_n627));
  NOR2_X1   g202(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT77), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n624), .A2(new_n625), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(G2451), .B(G2454), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT16), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n631), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(G1341), .B(G1348), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(G2443), .B(G2446), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  AND2_X1   g213(.A1(new_n638), .A2(G14), .ZN(G401));
  XOR2_X1   g214(.A(G2072), .B(G2078), .Z(new_n640));
  XOR2_X1   g215(.A(G2067), .B(G2678), .Z(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(G2084), .B(G2090), .Z(new_n643));
  NAND2_X1  g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  AOI21_X1  g219(.A(new_n640), .B1(new_n644), .B2(KEYINPUT18), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2096), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(G2100), .Z(new_n647));
  AND2_X1   g222(.A1(new_n644), .A2(KEYINPUT17), .ZN(new_n648));
  OR2_X1    g223(.A1(new_n642), .A2(new_n643), .ZN(new_n649));
  AOI21_X1  g224(.A(KEYINPUT18), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n647), .B(new_n650), .ZN(G227));
  XOR2_X1   g226(.A(G1956), .B(G2474), .Z(new_n652));
  XOR2_X1   g227(.A(G1961), .B(G1966), .Z(new_n653));
  NOR2_X1   g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1971), .B(G1976), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT19), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n652), .A2(new_n653), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  INV_X1    g235(.A(KEYINPUT20), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n658), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n655), .A2(new_n657), .A3(new_n659), .ZN(new_n663));
  OAI211_X1 g238(.A(new_n662), .B(new_n663), .C1(new_n661), .C2(new_n660), .ZN(new_n664));
  XOR2_X1   g239(.A(KEYINPUT21), .B(G1986), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(G1991), .B(G1996), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(KEYINPUT22), .B(G1981), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n668), .B(new_n669), .Z(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(G229));
  OAI21_X1  g246(.A(KEYINPUT81), .B1(G4), .B2(G16), .ZN(new_n672));
  OR3_X1    g247(.A1(KEYINPUT81), .A2(G4), .A3(G16), .ZN(new_n673));
  INV_X1    g248(.A(G16), .ZN(new_n674));
  OAI211_X1 g249(.A(new_n672), .B(new_n673), .C1(new_n593), .C2(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(G1348), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT30), .B(G28), .ZN(new_n678));
  INV_X1    g253(.A(G29), .ZN(new_n679));
  OR2_X1    g254(.A1(KEYINPUT31), .A2(G11), .ZN(new_n680));
  NAND2_X1  g255(.A1(KEYINPUT31), .A2(G11), .ZN(new_n681));
  AOI22_X1  g256(.A1(new_n678), .A2(new_n679), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n682), .B1(new_n616), .B2(new_n679), .ZN(new_n683));
  XOR2_X1   g258(.A(new_n683), .B(KEYINPUT87), .Z(new_n684));
  NOR2_X1   g259(.A1(G16), .A2(G21), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n685), .B1(G168), .B2(G16), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n686), .A2(G1966), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT88), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n679), .A2(G27), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n689), .B1(G164), .B2(new_n679), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(G2078), .ZN(new_n691));
  NOR4_X1   g266(.A1(new_n677), .A2(new_n684), .A3(new_n688), .A4(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(G171), .A2(G16), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n693), .B1(G5), .B2(G16), .ZN(new_n694));
  INV_X1    g269(.A(G1961), .ZN(new_n695));
  OR2_X1    g270(.A1(G29), .A2(G32), .ZN(new_n696));
  NAND3_X1  g271(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT26), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n698), .B1(new_n483), .B2(G129), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n489), .A2(G105), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n484), .A2(G141), .ZN(new_n701));
  NAND3_X1  g276(.A1(new_n699), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n696), .B1(new_n702), .B2(new_n679), .ZN(new_n703));
  XNOR2_X1  g278(.A(KEYINPUT27), .B(G1996), .ZN(new_n704));
  OAI22_X1  g279(.A1(new_n694), .A2(new_n695), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  OAI21_X1  g280(.A(KEYINPUT83), .B1(G29), .B2(G33), .ZN(new_n706));
  OR3_X1    g281(.A1(KEYINPUT83), .A2(G29), .A3(G33), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n489), .A2(G103), .ZN(new_n708));
  INV_X1    g283(.A(KEYINPUT25), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n484), .A2(G139), .ZN(new_n711));
  AOI22_X1  g286(.A1(new_n463), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n712));
  OAI211_X1 g287(.A(new_n710), .B(new_n711), .C1(new_n477), .C2(new_n712), .ZN(new_n713));
  OAI211_X1 g288(.A(new_n706), .B(new_n707), .C1(new_n713), .C2(new_n679), .ZN(new_n714));
  XOR2_X1   g289(.A(new_n714), .B(G2072), .Z(new_n715));
  NAND2_X1  g290(.A1(KEYINPUT24), .A2(G34), .ZN(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g292(.A1(KEYINPUT24), .A2(G34), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n679), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n720), .A2(KEYINPUT84), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n468), .A2(new_n478), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n721), .B1(new_n722), .B2(new_n679), .ZN(new_n723));
  INV_X1    g298(.A(KEYINPUT84), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n723), .B1(new_n724), .B2(new_n719), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n715), .B1(G2084), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n703), .A2(new_n704), .ZN(new_n727));
  XOR2_X1   g302(.A(new_n727), .B(KEYINPUT85), .Z(new_n728));
  NAND2_X1  g303(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT86), .ZN(new_n730));
  AOI211_X1 g305(.A(new_n705), .B(new_n730), .C1(new_n695), .C2(new_n694), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n725), .A2(G2084), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(new_n686), .B2(G1966), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n674), .A2(G19), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(new_n544), .B2(new_n674), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(G1341), .Z(new_n736));
  NAND4_X1  g311(.A1(new_n692), .A2(new_n731), .A3(new_n733), .A4(new_n736), .ZN(new_n737));
  NOR2_X1   g312(.A1(G16), .A2(G23), .ZN(new_n738));
  INV_X1    g313(.A(G288), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n738), .B1(new_n739), .B2(G16), .ZN(new_n740));
  XNOR2_X1  g315(.A(KEYINPUT33), .B(G1976), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n674), .A2(G22), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(G166), .B2(new_n674), .ZN(new_n744));
  INV_X1    g319(.A(G1971), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n744), .B(new_n745), .ZN(new_n746));
  MUX2_X1   g321(.A(G6), .B(G305), .S(G16), .Z(new_n747));
  XOR2_X1   g322(.A(KEYINPUT32), .B(G1981), .Z(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n742), .A2(new_n746), .A3(new_n749), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(KEYINPUT34), .Z(new_n751));
  NOR2_X1   g326(.A1(G25), .A2(G29), .ZN(new_n752));
  AOI22_X1  g327(.A1(new_n483), .A2(G119), .B1(G131), .B2(new_n484), .ZN(new_n753));
  OR2_X1    g328(.A1(G95), .A2(G2105), .ZN(new_n754));
  OAI211_X1 g329(.A(new_n754), .B(G2104), .C1(G107), .C2(new_n477), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(KEYINPUT78), .Z(new_n757));
  INV_X1    g332(.A(new_n757), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n752), .B1(new_n758), .B2(G29), .ZN(new_n759));
  XNOR2_X1  g334(.A(KEYINPUT35), .B(G1991), .ZN(new_n760));
  INV_X1    g335(.A(new_n760), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n759), .B(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n674), .A2(G24), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(new_n578), .B2(new_n674), .ZN(new_n764));
  XNOR2_X1  g339(.A(KEYINPUT79), .B(G1986), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n764), .B(new_n765), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n751), .A2(new_n762), .A3(new_n766), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT80), .ZN(new_n768));
  INV_X1    g343(.A(KEYINPUT36), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  OR2_X1    g345(.A1(new_n767), .A2(KEYINPUT80), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n767), .A2(KEYINPUT80), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n771), .A2(KEYINPUT36), .A3(new_n772), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n737), .B1(new_n770), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n679), .A2(G35), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(G162), .B2(new_n679), .ZN(new_n776));
  MUX2_X1   g351(.A(new_n775), .B(new_n776), .S(KEYINPUT89), .Z(new_n777));
  XOR2_X1   g352(.A(KEYINPUT29), .B(G2090), .Z(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n679), .A2(G26), .ZN(new_n780));
  AOI22_X1  g355(.A1(new_n483), .A2(G128), .B1(G140), .B2(new_n484), .ZN(new_n781));
  OR2_X1    g356(.A1(G104), .A2(G2105), .ZN(new_n782));
  OAI211_X1 g357(.A(new_n782), .B(G2104), .C1(G116), .C2(new_n477), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  INV_X1    g359(.A(new_n784), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n780), .B1(new_n785), .B2(new_n679), .ZN(new_n786));
  MUX2_X1   g361(.A(new_n780), .B(new_n786), .S(KEYINPUT28), .Z(new_n787));
  XNOR2_X1  g362(.A(KEYINPUT82), .B(G2067), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NAND3_X1  g364(.A1(new_n674), .A2(KEYINPUT23), .A3(G20), .ZN(new_n790));
  INV_X1    g365(.A(KEYINPUT23), .ZN(new_n791));
  INV_X1    g366(.A(G20), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n791), .B1(new_n792), .B2(G16), .ZN(new_n793));
  OAI211_X1 g368(.A(new_n790), .B(new_n793), .C1(new_n598), .C2(new_n674), .ZN(new_n794));
  INV_X1    g369(.A(G1956), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NAND4_X1  g371(.A1(new_n774), .A2(new_n779), .A3(new_n789), .A4(new_n796), .ZN(G150));
  INV_X1    g372(.A(G150), .ZN(G311));
  NAND2_X1  g373(.A1(new_n535), .A2(G93), .ZN(new_n799));
  AOI22_X1  g374(.A1(new_n518), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n800));
  XOR2_X1   g375(.A(KEYINPUT90), .B(G55), .Z(new_n801));
  OAI221_X1 g376(.A(new_n799), .B1(new_n501), .B2(new_n800), .C1(new_n576), .C2(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n802), .A2(G860), .ZN(new_n803));
  XOR2_X1   g378(.A(new_n803), .B(KEYINPUT37), .Z(new_n804));
  NAND2_X1  g379(.A1(new_n601), .A2(G559), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT38), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT39), .ZN(new_n807));
  OR2_X1    g382(.A1(new_n802), .A2(KEYINPUT91), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n802), .A2(KEYINPUT91), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n808), .A2(new_n544), .A3(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(new_n810), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n544), .B1(new_n808), .B2(new_n809), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n807), .B(new_n813), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n804), .B1(new_n814), .B2(G860), .ZN(G145));
  NAND2_X1  g390(.A1(new_n483), .A2(G130), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n484), .A2(G142), .ZN(new_n817));
  OAI21_X1  g392(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n818));
  OR2_X1    g393(.A1(new_n818), .A2(KEYINPUT93), .ZN(new_n819));
  INV_X1    g394(.A(KEYINPUT92), .ZN(new_n820));
  OR3_X1    g395(.A1(new_n820), .A2(new_n477), .A3(G118), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n820), .B1(new_n477), .B2(G118), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n818), .A2(KEYINPUT93), .ZN(new_n823));
  NAND4_X1  g398(.A1(new_n819), .A2(new_n821), .A3(new_n822), .A4(new_n823), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n816), .A2(new_n817), .A3(new_n824), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n756), .B(new_n825), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT94), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n827), .B(new_n619), .Z(new_n828));
  INV_X1    g403(.A(KEYINPUT95), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n827), .B(new_n619), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n831), .A2(KEYINPUT95), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n784), .B(G164), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(new_n702), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(new_n713), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n830), .A2(new_n832), .A3(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT96), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n831), .B(new_n829), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n839), .A2(KEYINPUT96), .A3(new_n835), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n616), .B(G160), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(G162), .ZN(new_n843));
  INV_X1    g418(.A(new_n843), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n835), .B(KEYINPUT97), .Z(new_n845));
  OAI211_X1 g420(.A(new_n841), .B(new_n844), .C1(new_n828), .C2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(G37), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n839), .A2(new_n835), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n848), .B1(new_n838), .B2(new_n840), .ZN(new_n849));
  OAI211_X1 g424(.A(new_n846), .B(new_n847), .C1(new_n849), .C2(new_n844), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n850), .A2(KEYINPUT40), .ZN(new_n851));
  OR2_X1    g426(.A1(new_n849), .A2(new_n844), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT40), .ZN(new_n853));
  NAND4_X1  g428(.A1(new_n852), .A2(new_n853), .A3(new_n847), .A4(new_n846), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n851), .A2(new_n854), .ZN(G395));
  NOR2_X1   g430(.A1(new_n802), .A2(G868), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n604), .B(new_n813), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n592), .B(new_n598), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT98), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT41), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n858), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n858), .A2(new_n860), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n592), .B(G299), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n863), .A2(KEYINPUT41), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  OAI211_X1 g440(.A(new_n857), .B(new_n861), .C1(new_n859), .C2(new_n865), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n866), .B1(new_n863), .B2(new_n857), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT100), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(G288), .B(G303), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(G305), .ZN(new_n871));
  OR2_X1    g446(.A1(new_n871), .A2(G290), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(G290), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(KEYINPUT99), .B(KEYINPUT42), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n874), .B(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n869), .A2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n867), .B(new_n868), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n877), .B1(new_n878), .B2(new_n876), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n856), .B1(new_n879), .B2(G868), .ZN(G295));
  AOI21_X1  g455(.A(new_n856), .B1(new_n879), .B2(G868), .ZN(G331));
  INV_X1    g456(.A(KEYINPUT103), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n802), .B(KEYINPUT91), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n883), .A2(new_n543), .ZN(new_n884));
  XNOR2_X1  g459(.A(G168), .B(G301), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n884), .A2(new_n810), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n886), .A2(KEYINPUT101), .ZN(new_n887));
  INV_X1    g462(.A(new_n885), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n888), .B1(new_n811), .B2(new_n812), .ZN(new_n889));
  AND2_X1   g464(.A1(new_n889), .A2(new_n886), .ZN(new_n890));
  OAI211_X1 g465(.A(new_n858), .B(new_n887), .C1(new_n890), .C2(KEYINPUT101), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n889), .A2(new_n886), .ZN(new_n892));
  OAI211_X1 g467(.A(new_n861), .B(new_n892), .C1(new_n865), .C2(new_n859), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT102), .ZN(new_n895));
  INV_X1    g470(.A(new_n874), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT43), .ZN(new_n898));
  OAI211_X1 g473(.A(new_n891), .B(new_n893), .C1(KEYINPUT102), .C2(new_n874), .ZN(new_n899));
  NAND4_X1  g474(.A1(new_n897), .A2(new_n898), .A3(new_n899), .A4(new_n847), .ZN(new_n900));
  AND2_X1   g475(.A1(new_n900), .A2(KEYINPUT44), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n890), .A2(new_n858), .ZN(new_n902));
  INV_X1    g477(.A(new_n887), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT101), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n903), .B1(new_n904), .B2(new_n892), .ZN(new_n905));
  INV_X1    g480(.A(new_n865), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n902), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  AND2_X1   g482(.A1(new_n907), .A2(new_n896), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n891), .A2(new_n874), .A3(new_n893), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n909), .A2(new_n847), .ZN(new_n910));
  OAI21_X1  g485(.A(KEYINPUT43), .B1(new_n908), .B2(new_n910), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n882), .B1(new_n901), .B2(new_n911), .ZN(new_n912));
  AND4_X1   g487(.A1(new_n882), .A2(new_n911), .A3(KEYINPUT44), .A4(new_n900), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n897), .A2(new_n847), .A3(new_n899), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(KEYINPUT43), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n907), .A2(new_n896), .ZN(new_n916));
  NAND4_X1  g491(.A1(new_n916), .A2(new_n898), .A3(new_n847), .A4(new_n909), .ZN(new_n917));
  AND2_X1   g492(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  OAI22_X1  g493(.A1(new_n912), .A2(new_n913), .B1(new_n918), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g494(.A(G2067), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n784), .B(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(G1384), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n922), .B1(new_n494), .B2(new_n499), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT45), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  XNOR2_X1  g500(.A(KEYINPUT104), .B(G40), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n468), .A2(new_n478), .A3(new_n927), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n925), .A2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(new_n929), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n921), .A2(new_n930), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n931), .A2(KEYINPUT105), .ZN(new_n932));
  AND2_X1   g507(.A1(new_n931), .A2(KEYINPUT105), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n702), .B(G1996), .ZN(new_n934));
  AOI211_X1 g509(.A(new_n932), .B(new_n933), .C1(new_n929), .C2(new_n934), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n756), .B(new_n761), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n935), .B1(new_n930), .B2(new_n936), .ZN(new_n937));
  XOR2_X1   g512(.A(new_n578), .B(G1986), .Z(new_n938));
  AOI21_X1  g513(.A(new_n937), .B1(new_n929), .B2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT107), .ZN(new_n940));
  OAI211_X1 g515(.A(KEYINPUT45), .B(new_n922), .C1(new_n494), .C2(new_n499), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n941), .A2(G160), .A3(new_n927), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT106), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n925), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n923), .A2(KEYINPUT106), .A3(new_n924), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n942), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n940), .B1(new_n946), .B2(G1971), .ZN(new_n947));
  AND3_X1   g522(.A1(new_n941), .A2(G160), .A3(new_n927), .ZN(new_n948));
  INV_X1    g523(.A(new_n945), .ZN(new_n949));
  AOI21_X1  g524(.A(KEYINPUT106), .B1(new_n923), .B2(new_n924), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n948), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n951), .A2(KEYINPUT107), .A3(new_n745), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT108), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n923), .A2(new_n953), .ZN(new_n954));
  OAI211_X1 g529(.A(KEYINPUT108), .B(new_n922), .C1(new_n494), .C2(new_n499), .ZN(new_n955));
  AOI21_X1  g530(.A(KEYINPUT50), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(G2090), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n928), .B1(new_n923), .B2(KEYINPUT50), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n957), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n947), .A2(new_n952), .A3(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(KEYINPUT109), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT109), .ZN(new_n963));
  NAND4_X1  g538(.A1(new_n947), .A2(new_n952), .A3(new_n963), .A4(new_n960), .ZN(new_n964));
  NAND2_X1  g539(.A1(G303), .A2(G8), .ZN(new_n965));
  NAND2_X1  g540(.A1(KEYINPUT110), .A2(KEYINPUT55), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  XOR2_X1   g542(.A(KEYINPUT110), .B(KEYINPUT55), .Z(new_n968));
  OAI21_X1  g543(.A(new_n967), .B1(new_n965), .B2(new_n968), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n962), .A2(G8), .A3(new_n964), .A4(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(G8), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n954), .A2(new_n955), .ZN(new_n972));
  INV_X1    g547(.A(new_n928), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n971), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  AND2_X1   g549(.A1(G305), .A2(G1981), .ZN(new_n975));
  NOR2_X1   g550(.A1(G305), .A2(G1981), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT49), .ZN(new_n977));
  OR3_X1    g552(.A1(new_n975), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n977), .B1(new_n975), .B2(new_n976), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n974), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT112), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n974), .A2(new_n978), .A3(KEYINPUT112), .A4(new_n979), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT111), .ZN(new_n985));
  INV_X1    g560(.A(G1976), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n985), .B1(G288), .B2(new_n986), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n739), .A2(KEYINPUT111), .A3(G1976), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n974), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(KEYINPUT52), .ZN(new_n990));
  AOI21_X1  g565(.A(KEYINPUT52), .B1(G288), .B2(new_n986), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n974), .A2(new_n987), .A3(new_n988), .A4(new_n991), .ZN(new_n992));
  AND3_X1   g567(.A1(new_n984), .A2(new_n990), .A3(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT115), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n951), .A2(new_n745), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n954), .A2(KEYINPUT50), .A3(new_n955), .ZN(new_n996));
  INV_X1    g571(.A(new_n499), .ZN(new_n997));
  INV_X1    g572(.A(G126), .ZN(new_n998));
  OAI22_X1  g573(.A1(new_n474), .A2(new_n998), .B1(new_n491), .B2(new_n470), .ZN(new_n999));
  AOI22_X1  g574(.A1(new_n999), .A2(G2105), .B1(G102), .B2(new_n489), .ZN(new_n1000));
  AOI21_X1  g575(.A(G1384), .B1(new_n997), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT50), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n928), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n996), .A2(KEYINPUT114), .A3(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(new_n958), .ZN(new_n1005));
  AOI21_X1  g580(.A(KEYINPUT114), .B1(new_n996), .B2(new_n1003), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n995), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(G8), .ZN(new_n1008));
  INV_X1    g583(.A(new_n969), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n994), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  AOI211_X1 g585(.A(KEYINPUT115), .B(new_n969), .C1(new_n1007), .C2(G8), .ZN(new_n1011));
  OAI211_X1 g586(.A(new_n970), .B(new_n993), .C1(new_n1010), .C2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT51), .ZN(new_n1014));
  INV_X1    g589(.A(new_n959), .ZN(new_n1015));
  XNOR2_X1  g590(.A(KEYINPUT116), .B(G2084), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1016), .ZN(new_n1017));
  NOR3_X1   g592(.A1(new_n956), .A2(new_n1015), .A3(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n954), .A2(new_n924), .A3(new_n955), .ZN(new_n1019));
  AOI21_X1  g594(.A(G1966), .B1(new_n1019), .B2(new_n948), .ZN(new_n1020));
  NOR3_X1   g595(.A1(new_n1018), .A2(new_n1020), .A3(G286), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1014), .B1(new_n1021), .B2(new_n971), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1020), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n957), .A2(new_n959), .A3(new_n1016), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1023), .A2(new_n1024), .A3(G168), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1025), .A2(KEYINPUT51), .A3(G8), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1022), .A2(KEYINPUT124), .A3(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT124), .ZN(new_n1028));
  OAI211_X1 g603(.A(new_n1028), .B(new_n1014), .C1(new_n1021), .C2(new_n971), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n971), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(G286), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1027), .A2(new_n1029), .A3(new_n1031), .ZN(new_n1032));
  XNOR2_X1  g607(.A(KEYINPUT125), .B(KEYINPUT54), .ZN(new_n1033));
  INV_X1    g608(.A(G2078), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n946), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT53), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n957), .A2(new_n959), .ZN(new_n1037));
  AOI22_X1  g612(.A1(new_n1035), .A2(new_n1036), .B1(new_n1037), .B2(new_n695), .ZN(new_n1038));
  AND2_X1   g613(.A1(new_n941), .A2(G160), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1036), .A2(G2078), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1039), .A2(G40), .A3(new_n925), .A4(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1038), .A2(new_n1041), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1042), .A2(G171), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1019), .A2(new_n948), .A3(new_n1040), .ZN(new_n1044));
  AOI21_X1  g619(.A(G301), .B1(new_n1038), .B2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1033), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1038), .A2(G301), .A3(new_n1044), .ZN(new_n1047));
  OR2_X1    g622(.A1(new_n1047), .A2(KEYINPUT126), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1042), .A2(G171), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1047), .A2(KEYINPUT126), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1048), .A2(KEYINPUT54), .A3(new_n1049), .A4(new_n1050), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1013), .A2(new_n1032), .A3(new_n1046), .A4(new_n1051), .ZN(new_n1052));
  XNOR2_X1  g627(.A(KEYINPUT120), .B(KEYINPUT61), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n996), .A2(new_n1003), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(new_n795), .ZN(new_n1055));
  XNOR2_X1  g630(.A(KEYINPUT56), .B(G2072), .ZN(new_n1056));
  OAI211_X1 g631(.A(new_n948), .B(new_n1056), .C1(new_n949), .C2(new_n950), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1055), .A2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT57), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n555), .A2(new_n1060), .A3(new_n558), .A4(new_n559), .ZN(new_n1061));
  AND2_X1   g636(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1058), .A2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1055), .A2(new_n1062), .A3(new_n1057), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1053), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT121), .ZN(new_n1067));
  AOI22_X1  g642(.A1(new_n946), .A2(new_n1056), .B1(new_n1054), .B2(new_n795), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1067), .B1(new_n1068), .B2(new_n1062), .ZN(new_n1069));
  AND4_X1   g644(.A1(new_n1067), .A2(new_n1055), .A3(new_n1062), .A4(new_n1057), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  AND2_X1   g646(.A1(new_n1064), .A2(KEYINPUT61), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1066), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  XOR2_X1   g648(.A(KEYINPUT58), .B(G1341), .Z(new_n1074));
  INV_X1    g649(.A(KEYINPUT117), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1075), .B1(new_n972), .B2(new_n973), .ZN(new_n1076));
  AOI211_X1 g651(.A(KEYINPUT117), .B(new_n928), .C1(new_n954), .C2(new_n955), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1074), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(KEYINPUT119), .ZN(new_n1079));
  INV_X1    g654(.A(G1996), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n946), .A2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT119), .ZN(new_n1082));
  OAI211_X1 g657(.A(new_n1082), .B(new_n1074), .C1(new_n1076), .C2(new_n1077), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1079), .A2(new_n1081), .A3(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(new_n544), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT59), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1084), .A2(KEYINPUT59), .A3(new_n544), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1073), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT122), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1073), .A2(new_n1087), .A3(KEYINPUT122), .A4(new_n1088), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1076), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1077), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1093), .A2(new_n1094), .A3(new_n920), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1037), .A2(new_n676), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(new_n601), .ZN(new_n1098));
  XOR2_X1   g673(.A(KEYINPUT123), .B(KEYINPUT60), .Z(new_n1099));
  AND2_X1   g674(.A1(new_n1097), .A2(KEYINPUT60), .ZN(new_n1100));
  OAI211_X1 g675(.A(new_n1098), .B(new_n1099), .C1(new_n1100), .C2(new_n601), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1099), .ZN(new_n1102));
  AND2_X1   g677(.A1(new_n1097), .A2(new_n601), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n601), .B1(new_n1097), .B2(KEYINPUT60), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1102), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  AND2_X1   g680(.A1(new_n1101), .A2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1091), .A2(new_n1092), .A3(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1064), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1108), .B1(new_n1103), .B2(new_n1065), .ZN(new_n1109));
  XNOR2_X1  g684(.A(new_n1109), .B(KEYINPUT118), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1052), .B1(new_n1107), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT63), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1030), .A2(G168), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1112), .B1(new_n1012), .B2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n962), .A2(G8), .A3(new_n964), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1112), .B1(new_n1115), .B2(new_n1009), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1113), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1116), .A2(new_n970), .A3(new_n993), .A4(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1114), .A2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n739), .A2(new_n986), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1120), .B1(new_n982), .B2(new_n983), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n974), .B1(new_n1121), .B2(new_n976), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n984), .A2(new_n990), .A3(new_n992), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1122), .B1(new_n970), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT113), .ZN(new_n1125));
  XNOR2_X1  g700(.A(new_n1124), .B(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1032), .A2(KEYINPUT62), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT62), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1027), .A2(new_n1029), .A3(new_n1128), .A4(new_n1031), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1013), .A2(new_n1127), .A3(new_n1045), .A4(new_n1129), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1119), .A2(new_n1126), .A3(new_n1130), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n939), .B1(new_n1111), .B2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n935), .A2(new_n761), .A3(new_n758), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n785), .A2(new_n920), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n930), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  NOR3_X1   g710(.A1(G290), .A2(G1986), .A3(new_n930), .ZN(new_n1136));
  XNOR2_X1  g711(.A(new_n1136), .B(KEYINPUT48), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n937), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n929), .A2(new_n1080), .ZN(new_n1139));
  XNOR2_X1  g714(.A(new_n1139), .B(KEYINPUT46), .ZN(new_n1140));
  INV_X1    g715(.A(new_n921), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n929), .B1(new_n1141), .B2(new_n702), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1143));
  XOR2_X1   g718(.A(new_n1143), .B(KEYINPUT47), .Z(new_n1144));
  NOR3_X1   g719(.A1(new_n1135), .A2(new_n1138), .A3(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1132), .A2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(KEYINPUT127), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT127), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1132), .A2(new_n1148), .A3(new_n1145), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1147), .A2(new_n1149), .ZN(G329));
  assign    G231 = 1'b0;
  AOI21_X1  g725(.A(new_n461), .B1(new_n915), .B2(new_n917), .ZN(new_n1152));
  NOR2_X1   g726(.A1(G401), .A2(G227), .ZN(new_n1153));
  NAND4_X1  g727(.A1(new_n850), .A2(new_n1152), .A3(new_n670), .A4(new_n1153), .ZN(G225));
  INV_X1    g728(.A(G225), .ZN(G308));
endmodule


