//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 1 0 0 1 0 0 1 0 0 0 1 1 1 0 1 0 0 1 0 1 1 1 1 0 1 1 0 1 0 0 0 0 0 1 0 0 1 1 1 0 0 0 0 0 1 1 0 0 0 1 0 1 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:16 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n446, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n553, new_n554, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n575, new_n576,
    new_n577, new_n579, new_n580, new_n581, new_n582, new_n583, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n604, new_n605, new_n608, new_n609, new_n610, new_n612,
    new_n613, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1150, new_n1151, new_n1152, new_n1153;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XOR2_X1   g017(.A(new_n442), .B(KEYINPUT65), .Z(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  NAND2_X1  g020(.A1(G94), .A2(G452), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT66), .Z(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT67), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  AND2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  OAI211_X1 g037(.A(G137), .B(new_n460), .C1(new_n461), .C2(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT68), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT68), .ZN(new_n470));
  NAND4_X1  g045(.A1(new_n469), .A2(new_n470), .A3(G137), .A4(new_n460), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n464), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n466), .A2(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G101), .ZN(new_n474));
  AND2_X1   g049(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(G125), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n477), .B1(new_n467), .B2(new_n468), .ZN(new_n478));
  AND2_X1   g053(.A1(G113), .A2(G2104), .ZN(new_n479));
  OAI21_X1  g054(.A(G2105), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n476), .A2(new_n481), .ZN(G160));
  NOR2_X1   g057(.A1(new_n461), .A2(new_n462), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n483), .A2(new_n460), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  AOI21_X1  g060(.A(G2105), .B1(new_n467), .B2(new_n468), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G136), .ZN(new_n487));
  OR2_X1    g062(.A1(G100), .A2(G2105), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n488), .B(G2104), .C1(G112), .C2(new_n460), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n485), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  INV_X1    g066(.A(KEYINPUT70), .ZN(new_n492));
  OR2_X1    g067(.A1(new_n460), .A2(G114), .ZN(new_n493));
  OAI21_X1  g068(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  AND2_X1   g071(.A1(G126), .A2(G2105), .ZN(new_n497));
  INV_X1    g072(.A(G138), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n498), .A2(G2105), .ZN(new_n499));
  NAND2_X1  g074(.A1(KEYINPUT69), .A2(KEYINPUT4), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n497), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n496), .B1(new_n502), .B2(new_n483), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n501), .B1(new_n486), .B2(G138), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n492), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(G126), .A2(G2105), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n460), .A2(G138), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n506), .B1(new_n507), .B2(new_n500), .ZN(new_n508));
  AOI22_X1  g083(.A1(new_n508), .A2(new_n469), .B1(new_n493), .B2(new_n495), .ZN(new_n509));
  OAI211_X1 g084(.A(G138), .B(new_n460), .C1(new_n461), .C2(new_n462), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(new_n500), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n509), .A2(KEYINPUT70), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n505), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(new_n513), .ZN(G164));
  XNOR2_X1  g089(.A(KEYINPUT5), .B(G543), .ZN(new_n515));
  XNOR2_X1  g090(.A(KEYINPUT6), .B(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(G88), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n516), .A2(G543), .ZN(new_n519));
  INV_X1    g094(.A(G50), .ZN(new_n520));
  OAI22_X1  g095(.A1(new_n517), .A2(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n515), .A2(G62), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(KEYINPUT71), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT71), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n515), .A2(new_n524), .A3(G62), .ZN(new_n525));
  NAND2_X1  g100(.A1(G75), .A2(G543), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n523), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n521), .B1(new_n527), .B2(G651), .ZN(G166));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n529), .B(KEYINPUT7), .ZN(new_n530));
  INV_X1    g105(.A(G51), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n530), .B1(new_n519), .B2(new_n531), .ZN(new_n532));
  XOR2_X1   g107(.A(KEYINPUT5), .B(G543), .Z(new_n533));
  NAND2_X1  g108(.A1(new_n516), .A2(G89), .ZN(new_n534));
  NAND2_X1  g109(.A1(G63), .A2(G651), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n532), .A2(new_n536), .ZN(G168));
  INV_X1    g112(.A(G90), .ZN(new_n538));
  INV_X1    g113(.A(G52), .ZN(new_n539));
  OAI22_X1  g114(.A1(new_n517), .A2(new_n538), .B1(new_n519), .B2(new_n539), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n515), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n541));
  INV_X1    g116(.A(G651), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  OR2_X1    g118(.A1(new_n540), .A2(new_n543), .ZN(G301));
  INV_X1    g119(.A(G301), .ZN(G171));
  AND3_X1   g120(.A1(new_n515), .A2(new_n516), .A3(G81), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n515), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n547), .A2(new_n542), .ZN(new_n548));
  AND2_X1   g123(.A1(new_n516), .A2(G543), .ZN(new_n549));
  AOI211_X1 g124(.A(new_n546), .B(new_n548), .C1(G43), .C2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND4_X1  g129(.A1(G319), .A2(G483), .A3(G661), .A4(new_n554), .ZN(G188));
  NAND2_X1  g130(.A1(new_n517), .A2(KEYINPUT72), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT72), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n515), .A2(new_n516), .A3(new_n557), .ZN(new_n558));
  AND2_X1   g133(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n559), .A2(KEYINPUT73), .A3(G91), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT73), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n556), .A2(new_n558), .ZN(new_n562));
  INV_X1    g137(.A(G91), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n561), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n560), .A2(new_n564), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n515), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n566));
  NOR2_X1   g141(.A1(new_n566), .A2(new_n542), .ZN(new_n567));
  INV_X1    g142(.A(G53), .ZN(new_n568));
  OAI21_X1  g143(.A(KEYINPUT9), .B1(new_n519), .B2(new_n568), .ZN(new_n569));
  OR3_X1    g144(.A1(new_n519), .A2(KEYINPUT9), .A3(new_n568), .ZN(new_n570));
  AOI21_X1  g145(.A(new_n567), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n565), .A2(new_n571), .ZN(G299));
  INV_X1    g147(.A(G168), .ZN(G286));
  INV_X1    g148(.A(G166), .ZN(G303));
  OR2_X1    g149(.A1(new_n515), .A2(G74), .ZN(new_n575));
  AOI22_X1  g150(.A1(G651), .A2(new_n575), .B1(new_n549), .B2(G49), .ZN(new_n576));
  INV_X1    g151(.A(G87), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n576), .B1(new_n562), .B2(new_n577), .ZN(G288));
  NAND2_X1  g153(.A1(G73), .A2(G543), .ZN(new_n579));
  INV_X1    g154(.A(G61), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n579), .B1(new_n533), .B2(new_n580), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n581), .A2(G651), .B1(new_n549), .B2(G48), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n556), .A2(G86), .A3(new_n558), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(new_n583), .ZN(G305));
  INV_X1    g159(.A(G85), .ZN(new_n585));
  XNOR2_X1  g160(.A(KEYINPUT74), .B(G47), .ZN(new_n586));
  OAI22_X1  g161(.A1(new_n517), .A2(new_n585), .B1(new_n519), .B2(new_n586), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n515), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n588), .A2(new_n542), .ZN(new_n589));
  OR2_X1    g164(.A1(new_n587), .A2(new_n589), .ZN(G290));
  NAND2_X1  g165(.A1(G301), .A2(G868), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n559), .A2(G92), .ZN(new_n592));
  XNOR2_X1  g167(.A(KEYINPUT75), .B(KEYINPUT10), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(G79), .A2(G543), .ZN(new_n595));
  INV_X1    g170(.A(G66), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n533), .B2(new_n596), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n597), .A2(G651), .B1(new_n549), .B2(G54), .ZN(new_n598));
  AND2_X1   g173(.A1(new_n594), .A2(new_n598), .ZN(new_n599));
  OR2_X1    g174(.A1(new_n592), .A2(new_n593), .ZN(new_n600));
  AND2_X1   g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n591), .B1(new_n601), .B2(G868), .ZN(G284));
  OAI21_X1  g177(.A(new_n591), .B1(new_n601), .B2(G868), .ZN(G321));
  NAND2_X1  g178(.A1(G286), .A2(G868), .ZN(new_n604));
  INV_X1    g179(.A(G299), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n605), .B2(G868), .ZN(G297));
  OAI21_X1  g181(.A(new_n604), .B1(new_n605), .B2(G868), .ZN(G280));
  NAND2_X1  g182(.A1(new_n599), .A2(new_n600), .ZN(new_n608));
  INV_X1    g183(.A(G860), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n608), .B1(G559), .B2(new_n609), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT76), .ZN(G148));
  OR2_X1    g186(.A1(new_n608), .A2(G559), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(G868), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n613), .B1(G868), .B2(new_n550), .ZN(G323));
  XNOR2_X1  g189(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g190(.A1(new_n469), .A2(new_n473), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT12), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT13), .ZN(new_n618));
  INV_X1    g193(.A(G2100), .ZN(new_n619));
  OR2_X1    g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n618), .A2(new_n619), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n484), .A2(G123), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n486), .A2(G135), .ZN(new_n623));
  NOR2_X1   g198(.A1(new_n460), .A2(G111), .ZN(new_n624));
  OAI21_X1  g199(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n625));
  OAI211_X1 g200(.A(new_n622), .B(new_n623), .C1(new_n624), .C2(new_n625), .ZN(new_n626));
  INV_X1    g201(.A(G2096), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n620), .A2(new_n621), .A3(new_n628), .ZN(G156));
  XNOR2_X1  g204(.A(G2427), .B(G2438), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2430), .ZN(new_n631));
  XNOR2_X1  g206(.A(KEYINPUT15), .B(G2435), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n631), .A2(new_n632), .ZN(new_n634));
  NAND3_X1  g209(.A1(new_n633), .A2(KEYINPUT14), .A3(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2451), .B(G2454), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT16), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n635), .B(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(G2443), .B(G2446), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(G1341), .B(G1348), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT77), .ZN(new_n642));
  NOR2_X1   g217(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT78), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n640), .A2(new_n642), .ZN(new_n645));
  AND3_X1   g220(.A1(new_n644), .A2(G14), .A3(new_n645), .ZN(G401));
  INV_X1    g221(.A(KEYINPUT18), .ZN(new_n647));
  XOR2_X1   g222(.A(G2084), .B(G2090), .Z(new_n648));
  XNOR2_X1  g223(.A(G2067), .B(G2678), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n650), .A2(KEYINPUT17), .ZN(new_n651));
  NOR2_X1   g226(.A1(new_n648), .A2(new_n649), .ZN(new_n652));
  OAI21_X1  g227(.A(new_n647), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(new_n619), .ZN(new_n654));
  XOR2_X1   g229(.A(G2072), .B(G2078), .Z(new_n655));
  AOI21_X1  g230(.A(new_n655), .B1(new_n650), .B2(KEYINPUT18), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(new_n627), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n654), .B(new_n657), .ZN(G227));
  XOR2_X1   g233(.A(G1956), .B(G2474), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT79), .ZN(new_n660));
  XOR2_X1   g235(.A(G1961), .B(G1966), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT80), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1971), .B(G1976), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT19), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n666), .B(KEYINPUT20), .Z(new_n667));
  OR2_X1    g242(.A1(new_n660), .A2(new_n662), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n668), .A2(new_n665), .A3(new_n663), .ZN(new_n669));
  OAI211_X1 g244(.A(new_n667), .B(new_n669), .C1(new_n665), .C2(new_n668), .ZN(new_n670));
  XNOR2_X1  g245(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1991), .B(G1996), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1981), .B(G1986), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n674), .B(new_n675), .Z(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(G229));
  INV_X1    g252(.A(G29), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n678), .A2(G32), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n484), .A2(G129), .ZN(new_n680));
  INV_X1    g255(.A(KEYINPUT87), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n486), .A2(G141), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT86), .ZN(new_n684));
  XNOR2_X1  g259(.A(KEYINPUT88), .B(KEYINPUT26), .ZN(new_n685));
  NAND3_X1  g260(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  AOI21_X1  g262(.A(new_n687), .B1(G105), .B2(new_n473), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n682), .A2(new_n684), .A3(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n679), .B1(new_n690), .B2(new_n678), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT27), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(G1996), .ZN(new_n693));
  INV_X1    g268(.A(G16), .ZN(new_n694));
  NOR2_X1   g269(.A1(G171), .A2(new_n694), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n695), .B1(G5), .B2(new_n694), .ZN(new_n696));
  INV_X1    g271(.A(G1961), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n694), .A2(G21), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(G168), .B2(new_n694), .ZN(new_n700));
  OR2_X1    g275(.A1(new_n700), .A2(G1966), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n700), .A2(G1966), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n698), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  AND2_X1   g278(.A1(new_n678), .A2(G33), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n460), .A2(G103), .A3(G2104), .ZN(new_n705));
  XOR2_X1   g280(.A(new_n705), .B(KEYINPUT25), .Z(new_n706));
  NAND2_X1  g281(.A1(new_n486), .A2(G139), .ZN(new_n707));
  AOI22_X1  g282(.A1(new_n469), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n708));
  OAI211_X1 g283(.A(new_n706), .B(new_n707), .C1(new_n460), .C2(new_n708), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n704), .B1(new_n709), .B2(G29), .ZN(new_n710));
  INV_X1    g285(.A(G2072), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(new_n696), .B2(new_n697), .ZN(new_n713));
  XOR2_X1   g288(.A(KEYINPUT31), .B(G11), .Z(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT89), .ZN(new_n715));
  INV_X1    g290(.A(G28), .ZN(new_n716));
  OR2_X1    g291(.A1(new_n716), .A2(KEYINPUT30), .ZN(new_n717));
  AOI21_X1  g292(.A(G29), .B1(new_n716), .B2(KEYINPUT30), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n715), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  OAI221_X1 g294(.A(new_n719), .B1(new_n678), .B2(new_n626), .C1(new_n710), .C2(new_n711), .ZN(new_n720));
  NOR3_X1   g295(.A1(new_n703), .A2(new_n713), .A3(new_n720), .ZN(new_n721));
  NOR2_X1   g296(.A1(G27), .A2(G29), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(G164), .B2(G29), .ZN(new_n723));
  INV_X1    g298(.A(G2078), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n678), .B1(KEYINPUT24), .B2(G34), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(KEYINPUT24), .B2(G34), .ZN(new_n727));
  INV_X1    g302(.A(G160), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n727), .B1(new_n728), .B2(G29), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(G2084), .ZN(new_n730));
  NAND4_X1  g305(.A1(new_n693), .A2(new_n721), .A3(new_n725), .A4(new_n730), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n731), .A2(KEYINPUT90), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n731), .A2(KEYINPUT90), .ZN(new_n733));
  NOR2_X1   g308(.A1(G4), .A2(G16), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT84), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(new_n608), .B2(new_n694), .ZN(new_n736));
  INV_X1    g311(.A(G1348), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n678), .A2(G35), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(G162), .B2(new_n678), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT29), .ZN(new_n741));
  INV_X1    g316(.A(G2090), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n741), .B(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n678), .A2(G26), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT28), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n484), .A2(G128), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n486), .A2(G140), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n460), .A2(G116), .ZN(new_n748));
  OAI21_X1  g323(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n749));
  OAI211_X1 g324(.A(new_n746), .B(new_n747), .C1(new_n748), .C2(new_n749), .ZN(new_n750));
  AND3_X1   g325(.A1(new_n750), .A2(KEYINPUT85), .A3(G29), .ZN(new_n751));
  AOI21_X1  g326(.A(KEYINPUT85), .B1(new_n750), .B2(G29), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n745), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(G2067), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  XOR2_X1   g330(.A(KEYINPUT82), .B(G16), .Z(new_n756));
  NOR2_X1   g331(.A1(new_n756), .A2(G19), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(new_n550), .B2(new_n756), .ZN(new_n758));
  XOR2_X1   g333(.A(new_n758), .B(G1341), .Z(new_n759));
  NAND3_X1  g334(.A1(new_n743), .A2(new_n755), .A3(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(G20), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n756), .A2(new_n761), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(KEYINPUT23), .Z(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(new_n605), .B2(new_n694), .ZN(new_n764));
  XNOR2_X1  g339(.A(KEYINPUT91), .B(G1956), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n764), .B(new_n765), .ZN(new_n766));
  NOR3_X1   g341(.A1(new_n738), .A2(new_n760), .A3(new_n766), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n732), .A2(new_n733), .A3(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n694), .A2(G23), .ZN(new_n769));
  INV_X1    g344(.A(G288), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n769), .B1(new_n770), .B2(new_n694), .ZN(new_n771));
  XNOR2_X1  g346(.A(KEYINPUT33), .B(G1976), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  MUX2_X1   g348(.A(G6), .B(G305), .S(G16), .Z(new_n774));
  XOR2_X1   g349(.A(KEYINPUT32), .B(G1981), .Z(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n756), .A2(G22), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(G166), .B2(new_n756), .ZN(new_n778));
  INV_X1    g353(.A(G1971), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NAND3_X1  g355(.A1(new_n773), .A2(new_n776), .A3(new_n780), .ZN(new_n781));
  XOR2_X1   g356(.A(new_n781), .B(KEYINPUT83), .Z(new_n782));
  INV_X1    g357(.A(KEYINPUT34), .ZN(new_n783));
  OR2_X1    g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n782), .A2(new_n783), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n484), .A2(G119), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n486), .A2(G131), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n460), .A2(G107), .ZN(new_n788));
  OAI21_X1  g363(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n789));
  OAI211_X1 g364(.A(new_n786), .B(new_n787), .C1(new_n788), .C2(new_n789), .ZN(new_n790));
  MUX2_X1   g365(.A(G25), .B(new_n790), .S(G29), .Z(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT81), .ZN(new_n792));
  XOR2_X1   g367(.A(KEYINPUT35), .B(G1991), .Z(new_n793));
  INV_X1    g368(.A(new_n793), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n792), .B(new_n794), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n756), .A2(G24), .ZN(new_n796));
  INV_X1    g371(.A(G290), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n796), .B1(new_n797), .B2(new_n756), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(G1986), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n795), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n784), .A2(new_n785), .A3(new_n800), .ZN(new_n801));
  OR2_X1    g376(.A1(new_n801), .A2(KEYINPUT36), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n801), .A2(KEYINPUT36), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n768), .B1(new_n802), .B2(new_n803), .ZN(G311));
  INV_X1    g379(.A(KEYINPUT92), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n802), .A2(new_n803), .ZN(new_n806));
  INV_X1    g381(.A(new_n768), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n805), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  AOI211_X1 g383(.A(KEYINPUT92), .B(new_n768), .C1(new_n802), .C2(new_n803), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n808), .A2(new_n809), .ZN(G150));
  INV_X1    g385(.A(G93), .ZN(new_n811));
  XOR2_X1   g386(.A(KEYINPUT93), .B(G55), .Z(new_n812));
  OAI22_X1  g387(.A1(new_n517), .A2(new_n811), .B1(new_n519), .B2(new_n812), .ZN(new_n813));
  AOI22_X1  g388(.A1(new_n515), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n814), .A2(new_n542), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n816), .A2(new_n609), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT95), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(KEYINPUT37), .Z(new_n819));
  NAND2_X1  g394(.A1(new_n601), .A2(G559), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT38), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n550), .B(new_n816), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n821), .B(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT39), .ZN(new_n824));
  OR2_X1    g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT94), .ZN(new_n826));
  AOI21_X1  g401(.A(G860), .B1(new_n823), .B2(new_n824), .ZN(new_n827));
  AND3_X1   g402(.A1(new_n825), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n826), .B1(new_n825), .B2(new_n827), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n819), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT96), .ZN(G145));
  XNOR2_X1  g406(.A(new_n689), .B(new_n709), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n484), .A2(G130), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n486), .A2(G142), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n460), .A2(G118), .ZN(new_n835));
  OAI21_X1  g410(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n836));
  OAI211_X1 g411(.A(new_n833), .B(new_n834), .C1(new_n835), .C2(new_n836), .ZN(new_n837));
  XOR2_X1   g412(.A(new_n837), .B(new_n617), .Z(new_n838));
  XNOR2_X1  g413(.A(new_n832), .B(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n509), .A2(new_n511), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n750), .B(new_n840), .ZN(new_n841));
  XOR2_X1   g416(.A(new_n841), .B(new_n790), .Z(new_n842));
  XNOR2_X1  g417(.A(new_n839), .B(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n626), .B(new_n490), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(G160), .ZN(new_n845));
  XOR2_X1   g420(.A(KEYINPUT97), .B(KEYINPUT98), .Z(new_n846));
  XNOR2_X1  g421(.A(new_n845), .B(new_n846), .ZN(new_n847));
  AOI21_X1  g422(.A(G37), .B1(new_n843), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n848), .B1(new_n847), .B2(new_n843), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g425(.A(new_n612), .B(new_n822), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n608), .B(G299), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(KEYINPUT41), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n608), .B(new_n605), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT41), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT99), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n854), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n852), .A2(KEYINPUT99), .A3(KEYINPUT41), .ZN(new_n860));
  AND2_X1   g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n853), .B1(new_n861), .B2(new_n851), .ZN(new_n862));
  OR2_X1    g437(.A1(new_n862), .A2(KEYINPUT42), .ZN(new_n863));
  XOR2_X1   g438(.A(G290), .B(G305), .Z(new_n864));
  XNOR2_X1  g439(.A(G288), .B(G166), .ZN(new_n865));
  XOR2_X1   g440(.A(new_n864), .B(new_n865), .Z(new_n866));
  NAND2_X1  g441(.A1(new_n862), .A2(KEYINPUT42), .ZN(new_n867));
  AND3_X1   g442(.A1(new_n863), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n866), .B1(new_n863), .B2(new_n867), .ZN(new_n869));
  OAI21_X1  g444(.A(G868), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n870), .B1(G868), .B2(new_n816), .ZN(G295));
  OAI21_X1  g446(.A(new_n870), .B1(G868), .B2(new_n816), .ZN(G331));
  XNOR2_X1  g447(.A(KEYINPUT100), .B(KEYINPUT43), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(G301), .B(G286), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n822), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n822), .A2(new_n875), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(KEYINPUT101), .ZN(new_n878));
  OAI211_X1 g453(.A(new_n859), .B(new_n860), .C1(new_n876), .C2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n866), .ZN(new_n880));
  INV_X1    g455(.A(new_n876), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n855), .A2(new_n881), .A3(new_n877), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n879), .A2(new_n880), .A3(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(G37), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  XOR2_X1   g460(.A(new_n866), .B(KEYINPUT102), .Z(new_n886));
  AOI21_X1  g461(.A(new_n886), .B1(new_n879), .B2(new_n882), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n874), .B1(new_n885), .B2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT103), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n854), .A2(new_n857), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n881), .A2(new_n877), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n855), .A2(KEYINPUT103), .A3(new_n856), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n890), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  OR3_X1    g468(.A1(new_n878), .A2(new_n852), .A3(new_n876), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n886), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  NAND4_X1  g471(.A1(new_n896), .A2(new_n884), .A3(new_n883), .A4(new_n873), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n888), .A2(new_n897), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n898), .A2(KEYINPUT44), .ZN(new_n899));
  OAI21_X1  g474(.A(KEYINPUT104), .B1(new_n885), .B2(new_n895), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n900), .A2(KEYINPUT43), .ZN(new_n901));
  NOR3_X1   g476(.A1(new_n885), .A2(KEYINPUT104), .A3(new_n895), .ZN(new_n902));
  OR2_X1    g477(.A1(new_n885), .A2(new_n887), .ZN(new_n903));
  OAI22_X1  g478(.A1(new_n901), .A2(new_n902), .B1(new_n903), .B2(new_n874), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n899), .B1(new_n904), .B2(KEYINPUT44), .ZN(G397));
  XNOR2_X1  g480(.A(KEYINPUT105), .B(G1384), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n840), .A2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT106), .ZN(new_n909));
  AOI21_X1  g484(.A(KEYINPUT45), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n840), .A2(KEYINPUT106), .A3(new_n907), .ZN(new_n911));
  AND2_X1   g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND4_X1  g487(.A1(new_n472), .A2(G40), .A3(new_n480), .A4(new_n474), .ZN(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  AND2_X1   g489(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(G1996), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n917), .A2(new_n689), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n915), .B(KEYINPUT107), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n750), .B(new_n754), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n920), .B1(new_n690), .B2(new_n916), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n918), .B1(new_n919), .B2(new_n921), .ZN(new_n922));
  AND2_X1   g497(.A1(new_n790), .A2(new_n794), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n790), .A2(new_n794), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n919), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  AND2_X1   g500(.A1(new_n922), .A2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  XNOR2_X1  g502(.A(G290), .B(G1986), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n927), .B1(new_n915), .B2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT50), .ZN(new_n930));
  INV_X1    g505(.A(G1384), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n930), .B1(new_n513), .B2(new_n931), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n840), .A2(new_n930), .A3(new_n931), .ZN(new_n933));
  NAND4_X1  g508(.A1(new_n933), .A2(new_n475), .A3(G40), .A4(new_n480), .ZN(new_n934));
  OR3_X1    g509(.A1(new_n932), .A2(new_n934), .A3(G2084), .ZN(new_n935));
  AOI21_X1  g510(.A(G1384), .B1(new_n505), .B2(new_n512), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(KEYINPUT45), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT45), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n840), .A2(new_n931), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n913), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n937), .A2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(G1966), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n935), .A2(new_n943), .ZN(new_n944));
  OAI21_X1  g519(.A(G8), .B1(new_n944), .B2(G286), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT119), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n945), .A2(new_n946), .A3(KEYINPUT51), .ZN(new_n947));
  XNOR2_X1  g522(.A(KEYINPUT119), .B(KEYINPUT51), .ZN(new_n948));
  OAI211_X1 g523(.A(G8), .B(new_n948), .C1(new_n944), .C2(G286), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n944), .A2(G8), .A3(G286), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n947), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  OR2_X1    g526(.A1(new_n951), .A2(KEYINPUT62), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT55), .ZN(new_n953));
  INV_X1    g528(.A(G8), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n953), .B1(G166), .B2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT110), .ZN(new_n956));
  AOI22_X1  g531(.A1(new_n522), .A2(KEYINPUT71), .B1(G75), .B2(G543), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n542), .B1(new_n957), .B2(new_n525), .ZN(new_n958));
  OAI211_X1 g533(.A(KEYINPUT55), .B(G8), .C1(new_n958), .C2(new_n521), .ZN(new_n959));
  AND3_X1   g534(.A1(new_n955), .A2(new_n956), .A3(new_n959), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n956), .B1(new_n955), .B2(new_n959), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  AOI21_X1  g537(.A(KEYINPUT45), .B1(new_n513), .B2(new_n931), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n840), .A2(KEYINPUT45), .A3(new_n907), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n914), .A2(new_n964), .ZN(new_n965));
  OAI21_X1  g540(.A(KEYINPUT108), .B1(new_n963), .B2(new_n965), .ZN(new_n966));
  AOI211_X1 g541(.A(new_n938), .B(new_n906), .C1(new_n509), .C2(new_n511), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n967), .A2(new_n913), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT108), .ZN(new_n969));
  OAI211_X1 g544(.A(new_n968), .B(new_n969), .C1(KEYINPUT45), .C2(new_n936), .ZN(new_n970));
  AND3_X1   g545(.A1(new_n966), .A2(new_n779), .A3(new_n970), .ZN(new_n971));
  AOI211_X1 g546(.A(KEYINPUT50), .B(G1384), .C1(new_n509), .C2(new_n511), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n972), .A2(new_n913), .ZN(new_n973));
  OAI211_X1 g548(.A(new_n973), .B(new_n742), .C1(new_n930), .C2(new_n936), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(KEYINPUT109), .ZN(new_n975));
  INV_X1    g550(.A(new_n512), .ZN(new_n976));
  AOI21_X1  g551(.A(KEYINPUT70), .B1(new_n509), .B2(new_n511), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n931), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(KEYINPUT50), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT109), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n979), .A2(new_n980), .A3(new_n742), .A4(new_n973), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n975), .A2(new_n981), .ZN(new_n982));
  OAI211_X1 g557(.A(G8), .B(new_n962), .C1(new_n971), .C2(new_n982), .ZN(new_n983));
  AOI22_X1  g558(.A1(new_n515), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n984));
  INV_X1    g559(.A(G48), .ZN(new_n985));
  OAI22_X1  g560(.A1(new_n984), .A2(new_n542), .B1(new_n985), .B2(new_n519), .ZN(new_n986));
  AND3_X1   g561(.A1(new_n515), .A2(new_n516), .A3(G86), .ZN(new_n987));
  OAI21_X1  g562(.A(G1981), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n988), .B1(G305), .B2(G1981), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT49), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  OAI211_X1 g566(.A(new_n988), .B(KEYINPUT49), .C1(G305), .C2(G1981), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n913), .A2(new_n939), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n993), .A2(new_n954), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n991), .A2(new_n992), .A3(new_n994), .ZN(new_n995));
  OAI211_X1 g570(.A(new_n576), .B(G1976), .C1(new_n577), .C2(new_n562), .ZN(new_n996));
  OAI211_X1 g571(.A(new_n996), .B(G8), .C1(new_n913), .C2(new_n939), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(KEYINPUT52), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n995), .A2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(new_n997), .ZN(new_n1000));
  INV_X1    g575(.A(G1976), .ZN(new_n1001));
  AOI21_X1  g576(.A(KEYINPUT52), .B1(G288), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT111), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1000), .A2(KEYINPUT111), .A3(new_n1002), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n999), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n983), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n955), .A2(new_n959), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n966), .A2(new_n779), .A3(new_n970), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n913), .B1(KEYINPUT50), .B2(new_n939), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1011), .B1(new_n978), .B2(KEYINPUT50), .ZN(new_n1012));
  OR2_X1    g587(.A1(new_n1012), .A2(G2090), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1010), .A2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1009), .B1(new_n1014), .B2(G8), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1008), .A2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(G2078), .B1(new_n966), .B2(new_n970), .ZN(new_n1017));
  XOR2_X1   g592(.A(KEYINPUT121), .B(KEYINPUT53), .Z(new_n1018));
  NOR2_X1   g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT113), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1020), .B1(new_n932), .B2(new_n934), .ZN(new_n1021));
  OAI211_X1 g596(.A(new_n973), .B(KEYINPUT113), .C1(new_n930), .C2(new_n936), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1021), .A2(new_n697), .A3(new_n1022), .ZN(new_n1023));
  AND2_X1   g598(.A1(new_n724), .A2(KEYINPUT53), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n937), .A2(new_n940), .A3(new_n1024), .ZN(new_n1025));
  AOI21_X1  g600(.A(KEYINPUT120), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1023), .A2(new_n1025), .A3(KEYINPUT120), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1019), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1029), .A2(G301), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n951), .A2(KEYINPUT62), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n952), .A2(new_n1016), .A3(new_n1030), .A4(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT112), .ZN(new_n1033));
  INV_X1    g608(.A(new_n983), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(new_n1007), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n995), .A2(new_n1001), .A3(new_n770), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1036), .B1(G1981), .B2(G305), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(new_n994), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1035), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  AOI211_X1 g615(.A(new_n954), .B(G286), .C1(new_n935), .C2(new_n943), .ZN(new_n1041));
  AOI21_X1  g616(.A(KEYINPUT63), .B1(new_n1016), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1008), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n944), .A2(KEYINPUT63), .A3(G8), .A4(G168), .ZN(new_n1044));
  OAI21_X1  g619(.A(G8), .B1(new_n971), .B2(new_n982), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1009), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1044), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  AND2_X1   g622(.A1(new_n1043), .A2(new_n1047), .ZN(new_n1048));
  OAI211_X1 g623(.A(new_n1033), .B(new_n1040), .C1(new_n1042), .C2(new_n1048), .ZN(new_n1049));
  AND2_X1   g624(.A1(new_n1010), .A2(new_n1013), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1046), .B1(new_n1050), .B2(new_n954), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1051), .A2(new_n1007), .A3(new_n983), .A4(new_n1041), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT63), .ZN(new_n1053));
  AOI22_X1  g628(.A1(new_n1052), .A2(new_n1053), .B1(new_n1043), .B2(new_n1047), .ZN(new_n1054));
  OAI21_X1  g629(.A(KEYINPUT112), .B1(new_n1054), .B2(new_n1039), .ZN(new_n1055));
  OR2_X1    g630(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1056));
  AND3_X1   g631(.A1(new_n1023), .A2(KEYINPUT120), .A3(new_n1025), .ZN(new_n1057));
  OAI211_X1 g632(.A(new_n1056), .B(G301), .C1(new_n1057), .C2(new_n1026), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT54), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n478), .A2(new_n479), .ZN(new_n1060));
  OR2_X1    g635(.A1(new_n1060), .A2(KEYINPUT122), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(KEYINPUT122), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1061), .A2(new_n1062), .A3(G2105), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1063), .A2(G40), .A3(new_n475), .A4(new_n1024), .ZN(new_n1064));
  OR3_X1    g639(.A1(new_n912), .A2(new_n967), .A3(new_n1064), .ZN(new_n1065));
  OAI211_X1 g640(.A(new_n1065), .B(new_n1023), .C1(new_n1017), .C2(new_n1018), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1059), .B1(new_n1066), .B2(G171), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1058), .A2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1068), .A2(new_n1016), .A3(new_n951), .ZN(new_n1069));
  OR3_X1    g644(.A1(new_n1066), .A2(KEYINPUT123), .A3(G171), .ZN(new_n1070));
  OAI21_X1  g645(.A(KEYINPUT123), .B1(new_n1066), .B2(G171), .ZN(new_n1071));
  OAI211_X1 g646(.A(new_n1070), .B(new_n1071), .C1(G301), .C2(new_n1029), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1069), .B1(new_n1059), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(G1956), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1012), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT115), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n978), .A2(new_n938), .ZN(new_n1077));
  XNOR2_X1  g652(.A(KEYINPUT56), .B(G2072), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1077), .A2(new_n968), .A3(new_n1078), .ZN(new_n1079));
  AND3_X1   g654(.A1(new_n1075), .A2(new_n1076), .A3(new_n1079), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1076), .B1(new_n1075), .B2(new_n1079), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT57), .ZN(new_n1082));
  XNOR2_X1  g657(.A(G299), .B(new_n1082), .ZN(new_n1083));
  NOR3_X1   g658(.A1(new_n1080), .A2(new_n1081), .A3(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1021), .A2(new_n737), .A3(new_n1022), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n993), .A2(new_n754), .ZN(new_n1086));
  AND3_X1   g661(.A1(new_n1085), .A2(KEYINPUT114), .A3(new_n1086), .ZN(new_n1087));
  AOI21_X1  g662(.A(KEYINPUT114), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  XNOR2_X1  g664(.A(G299), .B(KEYINPUT57), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1075), .A2(new_n1079), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1092), .A2(new_n608), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1084), .B1(new_n1089), .B2(new_n1093), .ZN(new_n1094));
  OAI21_X1  g669(.A(KEYINPUT60), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(new_n601), .ZN(new_n1096));
  OAI211_X1 g671(.A(KEYINPUT60), .B(new_n608), .C1(new_n1087), .C2(new_n1088), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT60), .ZN(new_n1098));
  AOI22_X1  g673(.A1(new_n1096), .A2(new_n1097), .B1(new_n1098), .B2(new_n1089), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT118), .ZN(new_n1100));
  OAI21_X1  g675(.A(KEYINPUT61), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1100), .B1(new_n1084), .B2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n968), .B1(new_n936), .B2(KEYINPUT45), .ZN(new_n1103));
  OAI21_X1  g678(.A(KEYINPUT116), .B1(new_n1103), .B2(G1996), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT116), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1077), .A2(new_n1105), .A3(new_n916), .A4(new_n968), .ZN(new_n1106));
  XNOR2_X1  g681(.A(KEYINPUT58), .B(G1341), .ZN(new_n1107));
  OAI211_X1 g682(.A(new_n1104), .B(new_n1106), .C1(new_n993), .C2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(new_n550), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1109), .A2(KEYINPUT59), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT59), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1108), .A2(new_n1111), .A3(new_n550), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1113));
  XNOR2_X1  g688(.A(KEYINPUT117), .B(KEYINPUT61), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1091), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1115), .A2(new_n1083), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1114), .B1(new_n1116), .B2(new_n1092), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1091), .A2(KEYINPUT115), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1075), .A2(new_n1076), .A3(new_n1079), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1118), .A2(new_n1090), .A3(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT61), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1121), .B1(new_n1115), .B2(new_n1083), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1120), .A2(new_n1122), .A3(KEYINPUT118), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1102), .A2(new_n1113), .A3(new_n1117), .A4(new_n1123), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1094), .B1(new_n1099), .B2(new_n1124), .ZN(new_n1125));
  AOI22_X1  g700(.A1(new_n1049), .A2(new_n1055), .B1(new_n1073), .B2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT124), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1032), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1049), .A2(new_n1055), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1073), .A2(new_n1125), .ZN(new_n1130));
  AND3_X1   g705(.A1(new_n1129), .A2(new_n1130), .A3(new_n1127), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n929), .B1(new_n1128), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n690), .A2(new_n920), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n919), .A2(new_n1133), .ZN(new_n1134));
  XNOR2_X1  g709(.A(new_n1134), .B(KEYINPUT126), .ZN(new_n1135));
  XNOR2_X1  g710(.A(new_n917), .B(KEYINPUT46), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  XOR2_X1   g712(.A(KEYINPUT127), .B(KEYINPUT47), .Z(new_n1138));
  XNOR2_X1  g713(.A(new_n1137), .B(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(G1986), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n915), .A2(new_n1140), .A3(new_n797), .ZN(new_n1141));
  XOR2_X1   g716(.A(new_n1141), .B(KEYINPUT48), .Z(new_n1142));
  OAI21_X1  g717(.A(new_n1139), .B1(new_n927), .B2(new_n1142), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n750), .A2(G2067), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1144), .B1(new_n922), .B2(new_n924), .ZN(new_n1145));
  XOR2_X1   g720(.A(new_n1145), .B(KEYINPUT125), .Z(new_n1146));
  AOI21_X1  g721(.A(new_n1143), .B1(new_n919), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1132), .A2(new_n1147), .ZN(G329));
  assign    G231 = 1'b0;
  AND2_X1   g723(.A1(new_n888), .A2(new_n897), .ZN(new_n1150));
  INV_X1    g724(.A(G319), .ZN(new_n1151));
  NOR3_X1   g725(.A1(G401), .A2(new_n1151), .A3(G227), .ZN(new_n1152));
  NAND3_X1  g726(.A1(new_n676), .A2(new_n849), .A3(new_n1152), .ZN(new_n1153));
  NOR2_X1   g727(.A1(new_n1150), .A2(new_n1153), .ZN(G308));
  INV_X1    g728(.A(G308), .ZN(G225));
endmodule


