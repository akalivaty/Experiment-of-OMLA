//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 1 1 1 1 1 0 1 1 1 0 1 0 1 1 0 0 1 1 1 1 0 1 0 1 1 0 1 0 1 1 0 1 0 0 1 0 1 1 0 1 1 1 1 0 0 0 1 1 1 0 0 1 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:55 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1271, new_n1272,
    new_n1273, new_n1275, new_n1276, new_n1277, new_n1278, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1346, new_n1347,
    new_n1348, new_n1349, new_n1350;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  OAI21_X1  g0012(.A(G50), .B1(G58), .B2(G68), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT64), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n207), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n218));
  INV_X1    g0018(.A(G58), .ZN(new_n219));
  INV_X1    g0019(.A(G232), .ZN(new_n220));
  INV_X1    g0020(.A(G97), .ZN(new_n221));
  INV_X1    g0021(.A(G257), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n218), .B1(new_n219), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n209), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n212), .B(new_n217), .C1(KEYINPUT1), .C2(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XOR2_X1   g0029(.A(G238), .B(G244), .Z(new_n230));
  XNOR2_X1  g0030(.A(G226), .B(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XOR2_X1   g0038(.A(G58), .B(G77), .Z(new_n239));
  XNOR2_X1  g0039(.A(G50), .B(G68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G351));
  NAND3_X1  g0045(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n246));
  INV_X1    g0046(.A(new_n246), .ZN(new_n247));
  INV_X1    g0047(.A(G68), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(KEYINPUT12), .ZN(new_n250));
  NAND3_X1  g0050(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(new_n215), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n247), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n206), .A2(G20), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n253), .A2(G68), .A3(new_n254), .ZN(new_n255));
  NOR2_X1   g0055(.A1(G20), .A2(G33), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  OAI22_X1  g0057(.A1(new_n257), .A2(new_n202), .B1(new_n207), .B2(G68), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n207), .A2(G33), .ZN(new_n259));
  INV_X1    g0059(.A(G77), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n252), .B1(new_n258), .B2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT11), .ZN(new_n263));
  OAI211_X1 g0063(.A(new_n250), .B(new_n255), .C1(new_n262), .C2(new_n263), .ZN(new_n264));
  AND2_X1   g0064(.A1(new_n262), .A2(new_n263), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  XNOR2_X1  g0066(.A(new_n266), .B(KEYINPUT75), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT74), .ZN(new_n268));
  NAND2_X1  g0068(.A1(G33), .A2(G41), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n269), .A2(G1), .A3(G13), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n270), .A2(G238), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(G33), .A2(G97), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  NOR2_X1   g0074(.A1(G226), .A2(G1698), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n275), .B1(new_n220), .B2(G1698), .ZN(new_n276));
  XNOR2_X1  g0076(.A(KEYINPUT3), .B(G33), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n274), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n272), .B1(new_n278), .B2(new_n270), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT71), .ZN(new_n280));
  INV_X1    g0080(.A(G41), .ZN(new_n281));
  INV_X1    g0081(.A(G45), .ZN(new_n282));
  AOI21_X1  g0082(.A(G1), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  AND4_X1   g0083(.A1(new_n280), .A2(new_n283), .A3(new_n270), .A4(G274), .ZN(new_n284));
  INV_X1    g0084(.A(G274), .ZN(new_n285));
  AND2_X1   g0085(.A1(G1), .A2(G13), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n285), .B1(new_n286), .B2(new_n269), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n280), .B1(new_n287), .B2(new_n283), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n284), .A2(new_n288), .ZN(new_n289));
  OAI21_X1  g0089(.A(KEYINPUT13), .B1(new_n279), .B2(new_n289), .ZN(new_n290));
  AND3_X1   g0090(.A1(new_n270), .A2(G238), .A3(new_n271), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n220), .A2(G1698), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n292), .B1(G226), .B2(G1698), .ZN(new_n293));
  AND2_X1   g0093(.A1(KEYINPUT3), .A2(G33), .ZN(new_n294));
  NOR2_X1   g0094(.A1(KEYINPUT3), .A2(G33), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n273), .B1(new_n293), .B2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(new_n270), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n291), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT13), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n283), .A2(new_n270), .A3(G274), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(KEYINPUT71), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n287), .A2(new_n280), .A3(new_n283), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n299), .A2(new_n300), .A3(new_n304), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n290), .A2(G179), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(KEYINPUT73), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT73), .ZN(new_n308));
  NAND4_X1  g0108(.A1(new_n290), .A2(new_n308), .A3(G179), .A4(new_n305), .ZN(new_n309));
  AND2_X1   g0109(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  AND3_X1   g0110(.A1(new_n299), .A2(new_n300), .A3(new_n304), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n300), .B1(new_n299), .B2(new_n304), .ZN(new_n312));
  OAI21_X1  g0112(.A(G169), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(KEYINPUT14), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n290), .A2(new_n305), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT14), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n315), .A2(new_n316), .A3(G169), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n314), .A2(new_n317), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n268), .B1(new_n310), .B2(new_n318), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n316), .B1(new_n315), .B2(G169), .ZN(new_n320));
  INV_X1    g0120(.A(G169), .ZN(new_n321));
  AOI211_X1 g0121(.A(KEYINPUT14), .B(new_n321), .C1(new_n290), .C2(new_n305), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n307), .A2(new_n309), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n323), .A2(KEYINPUT74), .A3(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n267), .B1(new_n319), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n315), .A2(G200), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n290), .A2(G190), .A3(new_n305), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n327), .A2(new_n328), .A3(new_n266), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(KEYINPUT72), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT72), .ZN(new_n331));
  NAND4_X1  g0131(.A1(new_n327), .A2(new_n331), .A3(new_n328), .A4(new_n266), .ZN(new_n332));
  AND2_X1   g0132(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n326), .A2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT18), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n270), .A2(new_n271), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n301), .B1(new_n220), .B2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(G1698), .ZN(new_n338));
  OAI211_X1 g0138(.A(G223), .B(new_n338), .C1(new_n294), .C2(new_n295), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT76), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND4_X1  g0141(.A1(new_n277), .A2(KEYINPUT76), .A3(G223), .A4(new_n338), .ZN(new_n342));
  NAND2_X1  g0142(.A1(G33), .A2(G87), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n277), .A2(G226), .A3(G1698), .ZN(new_n344));
  NAND4_X1  g0144(.A1(new_n341), .A2(new_n342), .A3(new_n343), .A4(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n337), .B1(new_n345), .B2(new_n298), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n346), .A2(G169), .ZN(new_n347));
  AOI211_X1 g0147(.A(G179), .B(new_n337), .C1(new_n345), .C2(new_n298), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT16), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT7), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n351), .B1(new_n277), .B2(G20), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n296), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n248), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n219), .A2(new_n248), .ZN(new_n355));
  OAI21_X1  g0155(.A(G20), .B1(new_n355), .B2(new_n201), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n256), .A2(G159), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n350), .B1(new_n354), .B2(new_n358), .ZN(new_n359));
  AOI21_X1  g0159(.A(KEYINPUT7), .B1(new_n296), .B2(new_n207), .ZN(new_n360));
  NOR4_X1   g0160(.A1(new_n294), .A2(new_n295), .A3(new_n351), .A4(G20), .ZN(new_n361));
  OAI21_X1  g0161(.A(G68), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n358), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n362), .A2(KEYINPUT16), .A3(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n359), .A2(new_n364), .A3(new_n252), .ZN(new_n365));
  XNOR2_X1  g0165(.A(KEYINPUT8), .B(G58), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n366), .B1(new_n206), .B2(G20), .ZN(new_n367));
  AOI22_X1  g0167(.A1(new_n367), .A2(new_n253), .B1(new_n247), .B2(new_n366), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n365), .A2(new_n368), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n335), .B1(new_n349), .B2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n349), .A2(new_n335), .A3(new_n369), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT77), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n345), .A2(new_n298), .ZN(new_n375));
  INV_X1    g0175(.A(new_n337), .ZN(new_n376));
  AOI21_X1  g0176(.A(G200), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  AOI211_X1 g0177(.A(G190), .B(new_n337), .C1(new_n345), .C2(new_n298), .ZN(new_n378));
  OAI211_X1 g0178(.A(new_n365), .B(new_n368), .C1(new_n377), .C2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT17), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(new_n368), .ZN(new_n382));
  INV_X1    g0182(.A(new_n252), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n362), .A2(new_n363), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n383), .B1(new_n384), .B2(new_n350), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n382), .B1(new_n385), .B2(new_n364), .ZN(new_n386));
  INV_X1    g0186(.A(G190), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n375), .A2(new_n387), .A3(new_n376), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n388), .B1(G200), .B2(new_n346), .ZN(new_n389));
  AOI21_X1  g0189(.A(KEYINPUT17), .B1(new_n386), .B2(new_n389), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n374), .B1(new_n381), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n379), .A2(new_n380), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n386), .A2(KEYINPUT17), .A3(new_n389), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n392), .A2(new_n393), .A3(KEYINPUT77), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n373), .B1(new_n391), .B2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT70), .ZN(new_n396));
  INV_X1    g0196(.A(G226), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n301), .B1(new_n397), .B2(new_n336), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n277), .A2(G222), .A3(new_n338), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n277), .A2(G223), .A3(G1698), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n296), .A2(G77), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n399), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT66), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n270), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n399), .A2(new_n400), .A3(KEYINPUT66), .A4(new_n401), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n398), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(G200), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n396), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(KEYINPUT10), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n402), .A2(new_n403), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n410), .A2(new_n298), .A3(new_n405), .ZN(new_n411));
  INV_X1    g0211(.A(new_n398), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n413), .A2(new_n387), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT9), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n203), .A2(G20), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(KEYINPUT67), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT67), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n203), .A2(new_n419), .A3(G20), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(G150), .ZN(new_n422));
  OAI22_X1  g0222(.A1(new_n366), .A2(new_n259), .B1(new_n422), .B2(new_n257), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n383), .B1(new_n421), .B2(new_n424), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n202), .B1(new_n206), .B2(G20), .ZN(new_n426));
  AOI22_X1  g0226(.A1(new_n253), .A2(new_n426), .B1(new_n202), .B2(new_n247), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n416), .B1(new_n425), .B2(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n423), .B1(new_n420), .B2(new_n418), .ZN(new_n430));
  OAI211_X1 g0230(.A(KEYINPUT9), .B(new_n427), .C1(new_n430), .C2(new_n383), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n407), .B1(new_n411), .B2(new_n412), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n409), .A2(new_n415), .A3(new_n434), .ZN(new_n435));
  OAI211_X1 g0235(.A(new_n429), .B(new_n431), .C1(new_n406), .C2(new_n407), .ZN(new_n436));
  OAI211_X1 g0236(.A(KEYINPUT10), .B(new_n408), .C1(new_n436), .C2(new_n414), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n413), .A2(G179), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n427), .B1(new_n430), .B2(new_n383), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n440), .B1(new_n406), .B2(G169), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(G244), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n301), .B1(new_n444), .B2(new_n336), .ZN(new_n445));
  OR2_X1    g0245(.A1(KEYINPUT3), .A2(G33), .ZN(new_n446));
  NAND2_X1  g0246(.A1(KEYINPUT3), .A2(G33), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n338), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(G238), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n277), .A2(G232), .A3(new_n338), .ZN(new_n450));
  XNOR2_X1  g0250(.A(KEYINPUT68), .B(G107), .ZN(new_n451));
  OAI211_X1 g0251(.A(new_n449), .B(new_n450), .C1(new_n277), .C2(new_n451), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n445), .B1(new_n452), .B2(new_n298), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(G190), .ZN(new_n454));
  OR2_X1    g0254(.A1(new_n257), .A2(KEYINPUT69), .ZN(new_n455));
  INV_X1    g0255(.A(new_n366), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n257), .A2(KEYINPUT69), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n455), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  XNOR2_X1  g0258(.A(KEYINPUT15), .B(G87), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(new_n259), .ZN(new_n461));
  AOI22_X1  g0261(.A1(new_n460), .A2(new_n461), .B1(G20), .B2(G77), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n383), .B1(new_n458), .B2(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n253), .A2(G77), .A3(new_n254), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n464), .B1(G77), .B2(new_n246), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n454), .B(new_n466), .C1(new_n407), .C2(new_n453), .ZN(new_n467));
  OR2_X1    g0267(.A1(new_n453), .A2(G169), .ZN(new_n468));
  INV_X1    g0268(.A(new_n466), .ZN(new_n469));
  INV_X1    g0269(.A(G179), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n453), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n468), .A2(new_n469), .A3(new_n471), .ZN(new_n472));
  AND4_X1   g0272(.A1(new_n438), .A2(new_n443), .A3(new_n467), .A4(new_n472), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n334), .A2(new_n395), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n206), .A2(G33), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n246), .A2(new_n475), .A3(new_n215), .A4(new_n251), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT78), .ZN(new_n477));
  OR2_X1    g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n476), .A2(new_n477), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n478), .A2(G87), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n459), .A2(new_n247), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT19), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(KEYINPUT80), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT80), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(KEYINPUT19), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n483), .B(new_n485), .C1(new_n259), .C2(new_n221), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n207), .B(G68), .C1(new_n294), .C2(new_n295), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  XNOR2_X1  g0288(.A(KEYINPUT80), .B(KEYINPUT19), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n207), .B1(new_n489), .B2(new_n273), .ZN(new_n490));
  INV_X1    g0290(.A(G87), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n451), .A2(new_n491), .A3(new_n221), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n488), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n480), .B(new_n481), .C1(new_n493), .C2(new_n383), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n206), .A2(G45), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n270), .A2(G250), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n270), .A2(G274), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n496), .B1(new_n497), .B2(new_n495), .ZN(new_n498));
  OAI211_X1 g0298(.A(G244), .B(G1698), .C1(new_n294), .C2(new_n295), .ZN(new_n499));
  OAI211_X1 g0299(.A(G238), .B(new_n338), .C1(new_n294), .C2(new_n295), .ZN(new_n500));
  INV_X1    g0300(.A(G33), .ZN(new_n501));
  INV_X1    g0301(.A(G116), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n499), .B(new_n500), .C1(new_n501), .C2(new_n502), .ZN(new_n503));
  AOI211_X1 g0303(.A(new_n387), .B(new_n498), .C1(new_n298), .C2(new_n503), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n494), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n503), .A2(new_n298), .ZN(new_n506));
  INV_X1    g0306(.A(new_n498), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(G200), .ZN(new_n509));
  AOI211_X1 g0309(.A(G179), .B(new_n498), .C1(new_n298), .C2(new_n503), .ZN(new_n510));
  AOI21_X1  g0310(.A(G169), .B1(new_n506), .B2(new_n507), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n478), .A2(new_n460), .A3(new_n479), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n513), .B(new_n481), .C1(new_n493), .C2(new_n383), .ZN(new_n514));
  AOI22_X1  g0314(.A1(new_n505), .A2(new_n509), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g0315(.A1(KEYINPUT5), .A2(G41), .ZN(new_n516));
  INV_X1    g0316(.A(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(KEYINPUT5), .A2(G41), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n495), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(new_n287), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n282), .A2(G1), .ZN(new_n521));
  INV_X1    g0321(.A(new_n518), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n521), .B1(new_n522), .B2(new_n516), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(new_n270), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n520), .B1(new_n524), .B2(new_n222), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n277), .A2(KEYINPUT4), .A3(G244), .A4(new_n338), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT79), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n277), .A2(G244), .A3(new_n338), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT4), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  AOI22_X1  g0331(.A1(new_n448), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n444), .B1(new_n446), .B2(new_n447), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n533), .A2(KEYINPUT79), .A3(KEYINPUT4), .A4(new_n338), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n528), .A2(new_n531), .A3(new_n532), .A4(new_n534), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n525), .B1(new_n535), .B2(new_n298), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(G190), .ZN(new_n537));
  INV_X1    g0337(.A(new_n451), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n538), .B1(new_n360), .B2(new_n361), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT6), .ZN(new_n540));
  AND2_X1   g0340(.A1(G97), .A2(G107), .ZN(new_n541));
  NOR2_X1   g0341(.A1(G97), .A2(G107), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(G107), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n544), .A2(KEYINPUT6), .A3(G97), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  AOI22_X1  g0346(.A1(new_n546), .A2(G20), .B1(G77), .B2(new_n256), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n383), .B1(new_n539), .B2(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n478), .A2(G97), .A3(new_n479), .ZN(new_n549));
  INV_X1    g0349(.A(new_n549), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n246), .A2(G97), .ZN(new_n551));
  NOR3_X1   g0351(.A1(new_n548), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n537), .B(new_n552), .C1(new_n407), .C2(new_n536), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n536), .A2(new_n470), .ZN(new_n554));
  INV_X1    g0354(.A(new_n551), .ZN(new_n555));
  AND2_X1   g0355(.A1(new_n539), .A2(new_n547), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n549), .B(new_n555), .C1(new_n556), .C2(new_n383), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n554), .B(new_n557), .C1(G169), .C2(new_n536), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n515), .A2(new_n553), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n247), .A2(new_n544), .ZN(new_n560));
  XOR2_X1   g0360(.A(new_n560), .B(KEYINPUT25), .Z(new_n561));
  NAND3_X1  g0361(.A1(new_n478), .A2(G107), .A3(new_n479), .ZN(new_n562));
  AND2_X1   g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n544), .A2(KEYINPUT68), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT68), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(G107), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n564), .A2(new_n566), .A3(G20), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(KEYINPUT23), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(KEYINPUT84), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT83), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n491), .A2(G20), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT82), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT22), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n277), .A2(new_n570), .A3(new_n571), .A4(new_n574), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n571), .B(new_n570), .C1(new_n295), .C2(new_n294), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(new_n573), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n569), .A2(new_n575), .A3(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT84), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n567), .A2(new_n579), .A3(KEYINPUT23), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n571), .B1(new_n294), .B2(new_n295), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(new_n572), .ZN(new_n582));
  NOR3_X1   g0382(.A1(new_n501), .A2(new_n502), .A3(G20), .ZN(new_n583));
  NOR3_X1   g0383(.A1(new_n207), .A2(KEYINPUT23), .A3(G107), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n580), .A2(new_n582), .A3(new_n585), .ZN(new_n586));
  OAI21_X1  g0386(.A(KEYINPUT85), .B1(new_n578), .B2(new_n586), .ZN(new_n587));
  AND3_X1   g0387(.A1(new_n580), .A2(new_n582), .A3(new_n585), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT85), .ZN(new_n589));
  AOI22_X1  g0389(.A1(new_n568), .A2(KEYINPUT84), .B1(new_n576), .B2(new_n573), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n588), .A2(new_n589), .A3(new_n590), .A4(new_n575), .ZN(new_n591));
  AND3_X1   g0391(.A1(new_n587), .A2(new_n591), .A3(KEYINPUT24), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT24), .ZN(new_n593));
  OAI211_X1 g0393(.A(KEYINPUT85), .B(new_n593), .C1(new_n578), .C2(new_n586), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n252), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n563), .B1(new_n592), .B2(new_n595), .ZN(new_n596));
  OAI211_X1 g0396(.A(G257), .B(G1698), .C1(new_n294), .C2(new_n295), .ZN(new_n597));
  OAI211_X1 g0397(.A(G250), .B(new_n338), .C1(new_n294), .C2(new_n295), .ZN(new_n598));
  INV_X1    g0398(.A(G294), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n597), .B(new_n598), .C1(new_n501), .C2(new_n599), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n519), .A2(new_n298), .ZN(new_n601));
  AOI22_X1  g0401(.A1(new_n600), .A2(new_n298), .B1(new_n601), .B2(G264), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n602), .A2(G179), .A3(new_n520), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT86), .ZN(new_n604));
  OR2_X1    g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n321), .B1(new_n602), .B2(new_n520), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n603), .B1(new_n606), .B2(new_n604), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n596), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n523), .A2(G270), .A3(new_n270), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n520), .A2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(new_n611), .ZN(new_n612));
  OAI211_X1 g0412(.A(G264), .B(G1698), .C1(new_n294), .C2(new_n295), .ZN(new_n613));
  OAI211_X1 g0413(.A(G257), .B(new_n338), .C1(new_n294), .C2(new_n295), .ZN(new_n614));
  INV_X1    g0414(.A(G303), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n613), .B(new_n614), .C1(new_n615), .C2(new_n277), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(new_n298), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n612), .A2(new_n617), .ZN(new_n618));
  OR2_X1    g0418(.A1(new_n476), .A2(new_n502), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n247), .A2(new_n502), .ZN(new_n620));
  AOI22_X1  g0420(.A1(new_n251), .A2(new_n215), .B1(G20), .B2(new_n502), .ZN(new_n621));
  AOI21_X1  g0421(.A(G20), .B1(G33), .B2(G283), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n622), .B1(G33), .B2(new_n221), .ZN(new_n623));
  AND3_X1   g0423(.A1(new_n621), .A2(new_n623), .A3(KEYINPUT20), .ZN(new_n624));
  AOI21_X1  g0424(.A(KEYINPUT20), .B1(new_n621), .B2(new_n623), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n619), .B(new_n620), .C1(new_n624), .C2(new_n625), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n618), .A2(G169), .A3(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT21), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(KEYINPUT81), .ZN(new_n629));
  INV_X1    g0429(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n627), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n612), .A2(G190), .A3(new_n617), .ZN(new_n632));
  INV_X1    g0432(.A(new_n626), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n611), .B1(new_n298), .B2(new_n616), .ZN(new_n634));
  OAI211_X1 g0434(.A(new_n632), .B(new_n633), .C1(new_n634), .C2(new_n407), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n634), .A2(G179), .A3(new_n626), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n618), .A2(G169), .A3(new_n626), .A4(new_n629), .ZN(new_n637));
  AND4_X1   g0437(.A1(new_n631), .A2(new_n635), .A3(new_n636), .A4(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n600), .A2(new_n298), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n601), .A2(G264), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n639), .A2(new_n520), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(new_n407), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n642), .B1(G190), .B2(new_n641), .ZN(new_n643));
  OAI211_X1 g0443(.A(new_n563), .B(new_n643), .C1(new_n592), .C2(new_n595), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n609), .A2(new_n638), .A3(new_n644), .ZN(new_n645));
  NOR3_X1   g0445(.A1(new_n474), .A2(new_n559), .A3(new_n645), .ZN(G372));
  INV_X1    g0446(.A(new_n372), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n647), .A2(new_n370), .ZN(new_n648));
  INV_X1    g0448(.A(new_n267), .ZN(new_n649));
  AND4_X1   g0449(.A1(KEYINPUT74), .A2(new_n324), .A3(new_n314), .A4(new_n317), .ZN(new_n650));
  AOI21_X1  g0450(.A(KEYINPUT74), .B1(new_n323), .B2(new_n324), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n649), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n330), .A2(new_n332), .ZN(new_n653));
  INV_X1    g0453(.A(new_n472), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n652), .A2(KEYINPUT88), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n391), .A2(new_n394), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  AOI21_X1  g0458(.A(KEYINPUT88), .B1(new_n652), .B2(new_n655), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n648), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n442), .B1(new_n660), .B2(new_n438), .ZN(new_n661));
  AND3_X1   g0461(.A1(new_n334), .A2(new_n395), .A3(new_n473), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n644), .A2(new_n515), .A3(new_n553), .A4(new_n558), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n631), .A2(new_n636), .A3(new_n637), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n664), .B1(new_n596), .B2(new_n608), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n535), .A2(new_n298), .ZN(new_n667));
  INV_X1    g0467(.A(new_n525), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n548), .A2(new_n551), .ZN(new_n670));
  AOI22_X1  g0470(.A1(new_n321), .A2(new_n669), .B1(new_n670), .B2(new_n549), .ZN(new_n671));
  XOR2_X1   g0471(.A(KEYINPUT87), .B(KEYINPUT26), .Z(new_n672));
  NAND4_X1  g0472(.A1(new_n515), .A2(new_n554), .A3(new_n671), .A4(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n490), .A2(new_n492), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n674), .A2(new_n486), .A3(new_n487), .ZN(new_n675));
  AOI22_X1  g0475(.A1(new_n675), .A2(new_n252), .B1(new_n247), .B2(new_n459), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n498), .B1(new_n503), .B2(new_n298), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(G190), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n676), .A2(new_n509), .A3(new_n480), .A4(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n508), .A2(new_n321), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n677), .A2(new_n470), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n514), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(KEYINPUT26), .B1(new_n558), .B2(new_n683), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n673), .A2(new_n684), .A3(new_n682), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n662), .B1(new_n666), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n661), .A2(new_n686), .ZN(G369));
  NAND3_X1  g0487(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n688));
  OR2_X1    g0488(.A1(new_n688), .A2(KEYINPUT27), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(KEYINPUT27), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n689), .A2(G213), .A3(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(G343), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n587), .A2(new_n591), .A3(KEYINPUT24), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n694), .A2(new_n252), .A3(new_n594), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n693), .B1(new_n695), .B2(new_n563), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT89), .ZN(new_n697));
  OR2_X1    g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n644), .ZN(new_n699));
  AOI22_X1  g0499(.A1(new_n695), .A2(new_n563), .B1(new_n605), .B2(new_n607), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n696), .A2(new_n697), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n698), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n693), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n700), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n633), .A2(new_n693), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n664), .A2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n638), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n708), .B1(new_n709), .B2(new_n707), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(G330), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n706), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n700), .A2(new_n693), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n664), .A2(new_n693), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n698), .A2(new_n701), .A3(new_n702), .A4(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n713), .A2(new_n714), .A3(new_n717), .ZN(G399));
  INV_X1    g0518(.A(new_n210), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n719), .A2(G41), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n492), .A2(G116), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NOR3_X1   g0522(.A1(new_n720), .A2(new_n722), .A3(new_n206), .ZN(new_n723));
  INV_X1    g0523(.A(new_n213), .ZN(new_n724));
  AOI22_X1  g0524(.A1(new_n723), .A2(KEYINPUT90), .B1(new_n724), .B2(new_n720), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n725), .B1(KEYINPUT90), .B2(new_n723), .ZN(new_n726));
  XNOR2_X1  g0526(.A(new_n726), .B(KEYINPUT28), .ZN(new_n727));
  OAI211_X1 g0527(.A(KEYINPUT92), .B(new_n672), .C1(new_n558), .C2(new_n683), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n515), .A2(KEYINPUT26), .A3(new_n554), .A4(new_n671), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n671), .A2(new_n554), .A3(new_n682), .A4(new_n679), .ZN(new_n731));
  AOI21_X1  g0531(.A(KEYINPUT92), .B1(new_n731), .B2(new_n672), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n682), .B1(new_n663), .B2(new_n665), .ZN(new_n734));
  OAI211_X1 g0534(.A(KEYINPUT29), .B(new_n693), .C1(new_n733), .C2(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n693), .B1(new_n666), .B2(new_n685), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT29), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n735), .A2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT91), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n602), .A2(new_n677), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n612), .A2(G179), .A3(new_n617), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  AOI21_X1  g0543(.A(KEYINPUT30), .B1(new_n743), .B2(new_n536), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n618), .A2(new_n641), .A3(new_n470), .A4(new_n508), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(new_n536), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n740), .B1(new_n744), .B2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT30), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n634), .A2(G179), .A3(new_n677), .A4(new_n602), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n748), .B1(new_n749), .B2(new_n669), .ZN(new_n750));
  NOR3_X1   g0550(.A1(new_n634), .A2(G179), .A3(new_n677), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n751), .A2(new_n669), .A3(new_n641), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n750), .A2(new_n752), .A3(KEYINPUT91), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n743), .A2(KEYINPUT30), .A3(new_n536), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n747), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  AND2_X1   g0555(.A1(new_n704), .A2(KEYINPUT31), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n750), .A2(new_n754), .A3(new_n752), .ZN(new_n758));
  AOI21_X1  g0558(.A(KEYINPUT31), .B1(new_n758), .B2(new_n704), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n757), .A2(new_n760), .ZN(new_n761));
  NOR3_X1   g0561(.A1(new_n645), .A2(new_n559), .A3(new_n704), .ZN(new_n762));
  OAI21_X1  g0562(.A(G330), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  AND2_X1   g0563(.A1(new_n739), .A2(new_n763), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n727), .B1(new_n764), .B2(G1), .ZN(G364));
  AND2_X1   g0565(.A1(new_n207), .A2(G13), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(G45), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n206), .B1(new_n768), .B2(KEYINPUT93), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n769), .B1(KEYINPUT93), .B2(new_n768), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(new_n720), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n712), .A2(new_n771), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n772), .B1(G330), .B2(new_n710), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n719), .A2(new_n296), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(G355), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n775), .B1(G116), .B2(new_n210), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n719), .A2(new_n277), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n778), .B1(new_n214), .B2(new_n282), .ZN(new_n779));
  OR2_X1    g0579(.A1(new_n241), .A2(new_n282), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n776), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(G13), .A2(G33), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(G20), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n215), .B1(G20), .B2(new_n321), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n771), .B1(new_n781), .B2(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n207), .A2(new_n470), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(G200), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(G190), .ZN(new_n791));
  INV_X1    g0591(.A(G317), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(KEYINPUT33), .ZN(new_n793));
  OR2_X1    g0593(.A1(new_n792), .A2(KEYINPUT33), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n791), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  NOR3_X1   g0595(.A1(new_n387), .A2(G179), .A3(G200), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(new_n207), .ZN(new_n797));
  INV_X1    g0597(.A(G326), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n790), .A2(new_n387), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  OAI221_X1 g0600(.A(new_n795), .B1(new_n599), .B2(new_n797), .C1(new_n798), .C2(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n207), .A2(G190), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n802), .A2(G179), .A3(new_n407), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n802), .A2(new_n470), .A3(new_n407), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  AOI22_X1  g0606(.A1(new_n804), .A2(G311), .B1(new_n806), .B2(G329), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n789), .A2(G190), .A3(new_n407), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n277), .B1(new_n809), .B2(G322), .ZN(new_n810));
  NOR4_X1   g0610(.A1(new_n207), .A2(new_n387), .A3(new_n407), .A4(G179), .ZN(new_n811));
  NOR4_X1   g0611(.A1(new_n207), .A2(new_n407), .A3(G179), .A4(G190), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n811), .A2(G303), .B1(new_n812), .B2(G283), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n807), .A2(new_n810), .A3(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n801), .A2(new_n814), .ZN(new_n815));
  XOR2_X1   g0615(.A(new_n815), .B(KEYINPUT97), .Z(new_n816));
  NAND2_X1  g0616(.A1(new_n811), .A2(G87), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(new_n277), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n818), .B(KEYINPUT96), .ZN(new_n819));
  INV_X1    g0619(.A(new_n791), .ZN(new_n820));
  INV_X1    g0620(.A(new_n812), .ZN(new_n821));
  OAI22_X1  g0621(.A1(new_n820), .A2(new_n248), .B1(new_n544), .B2(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n800), .A2(new_n202), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n797), .A2(new_n221), .ZN(new_n824));
  NOR3_X1   g0624(.A1(new_n822), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(G159), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n805), .A2(new_n826), .ZN(new_n827));
  XNOR2_X1  g0627(.A(new_n827), .B(KEYINPUT32), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n819), .A2(new_n825), .A3(new_n828), .ZN(new_n829));
  XOR2_X1   g0629(.A(new_n808), .B(KEYINPUT94), .Z(new_n830));
  OAI22_X1  g0630(.A1(new_n830), .A2(new_n219), .B1(new_n260), .B2(new_n803), .ZN(new_n831));
  XNOR2_X1  g0631(.A(new_n831), .B(KEYINPUT95), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n816), .B1(new_n829), .B2(new_n832), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n788), .B1(new_n833), .B2(new_n785), .ZN(new_n834));
  INV_X1    g0634(.A(new_n784), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n834), .B1(new_n710), .B2(new_n835), .ZN(new_n836));
  AND2_X1   g0636(.A1(new_n773), .A2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(G396));
  NOR2_X1   g0638(.A1(new_n466), .A2(new_n693), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT100), .ZN(new_n840));
  XNOR2_X1  g0640(.A(new_n839), .B(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n472), .A2(KEYINPUT99), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT99), .ZN(new_n843));
  NAND4_X1  g0643(.A1(new_n468), .A2(new_n843), .A3(new_n469), .A4(new_n471), .ZN(new_n844));
  NAND4_X1  g0644(.A1(new_n841), .A2(new_n467), .A3(new_n842), .A4(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  OAI211_X1 g0646(.A(new_n693), .B(new_n846), .C1(new_n666), .C2(new_n685), .ZN(new_n847));
  INV_X1    g0647(.A(new_n736), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n654), .A2(new_n704), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n845), .A2(new_n849), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n847), .B1(new_n848), .B2(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n771), .B1(new_n851), .B2(new_n763), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n852), .B1(new_n763), .B2(new_n851), .ZN(new_n853));
  INV_X1    g0653(.A(new_n785), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(new_n783), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n771), .B1(G77), .B2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(G311), .ZN(new_n857));
  OAI22_X1  g0657(.A1(new_n821), .A2(new_n491), .B1(new_n857), .B2(new_n805), .ZN(new_n858));
  XOR2_X1   g0658(.A(new_n858), .B(KEYINPUT98), .Z(new_n859));
  OAI21_X1  g0659(.A(new_n296), .B1(new_n803), .B2(new_n502), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n860), .B1(G294), .B2(new_n809), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n824), .B1(G283), .B2(new_n791), .ZN(new_n862));
  AOI22_X1  g0662(.A1(new_n799), .A2(G303), .B1(G107), .B2(new_n811), .ZN(new_n863));
  NAND4_X1  g0663(.A1(new_n859), .A2(new_n861), .A3(new_n862), .A4(new_n863), .ZN(new_n864));
  AOI22_X1  g0664(.A1(new_n799), .A2(G137), .B1(new_n804), .B2(G159), .ZN(new_n865));
  INV_X1    g0665(.A(G143), .ZN(new_n866));
  OAI221_X1 g0666(.A(new_n865), .B1(new_n422), .B2(new_n820), .C1(new_n830), .C2(new_n866), .ZN(new_n867));
  XOR2_X1   g0667(.A(new_n867), .B(KEYINPUT34), .Z(new_n868));
  INV_X1    g0668(.A(G132), .ZN(new_n869));
  OAI221_X1 g0669(.A(new_n277), .B1(new_n805), .B2(new_n869), .C1(new_n797), .C2(new_n219), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n812), .A2(G68), .ZN(new_n871));
  INV_X1    g0671(.A(new_n811), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n871), .B1(new_n872), .B2(new_n202), .ZN(new_n873));
  OR2_X1    g0673(.A1(new_n870), .A2(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n864), .B1(new_n868), .B2(new_n874), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n856), .B1(new_n875), .B2(new_n785), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n876), .B1(new_n783), .B2(new_n850), .ZN(new_n877));
  AND2_X1   g0677(.A1(new_n853), .A2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(new_n878), .ZN(G384));
  OR2_X1    g0679(.A1(new_n546), .A2(KEYINPUT35), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n546), .A2(KEYINPUT35), .ZN(new_n881));
  NAND4_X1  g0681(.A1(new_n880), .A2(G116), .A3(new_n216), .A4(new_n881), .ZN(new_n882));
  XOR2_X1   g0682(.A(new_n882), .B(KEYINPUT36), .Z(new_n883));
  NOR3_X1   g0683(.A1(new_n355), .A2(new_n213), .A3(new_n260), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT101), .ZN(new_n885));
  OR2_X1    g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AOI22_X1  g0686(.A1(new_n884), .A2(new_n885), .B1(new_n202), .B2(G68), .ZN(new_n887));
  AOI211_X1 g0687(.A(new_n206), .B(G13), .C1(new_n886), .C2(new_n887), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n883), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n649), .A2(new_n704), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n652), .A2(new_n653), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n319), .A2(new_n325), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n649), .B(new_n704), .C1(new_n892), .C2(new_n333), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n842), .A2(new_n844), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(new_n693), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n847), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n894), .A2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT38), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n369), .A2(new_n692), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n901), .B1(new_n657), .B2(new_n648), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n691), .B1(new_n365), .B2(new_n368), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n903), .B1(new_n386), .B2(new_n389), .ZN(new_n904));
  INV_X1    g0704(.A(new_n347), .ZN(new_n905));
  INV_X1    g0705(.A(new_n348), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n369), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  OAI211_X1 g0707(.A(new_n904), .B(new_n907), .C1(KEYINPUT102), .C2(KEYINPUT37), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n907), .A2(new_n379), .A3(new_n901), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT37), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n901), .A2(KEYINPUT102), .A3(new_n379), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n909), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n908), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n900), .B1(new_n902), .B2(new_n913), .ZN(new_n914));
  AND2_X1   g0714(.A1(new_n908), .A2(new_n912), .ZN(new_n915));
  OAI211_X1 g0715(.A(new_n915), .B(KEYINPUT38), .C1(new_n395), .C2(new_n901), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  AOI22_X1  g0717(.A1(new_n899), .A2(new_n917), .B1(new_n373), .B2(new_n691), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n381), .A2(new_n390), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n901), .B1(new_n648), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n900), .B1(new_n920), .B2(new_n913), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n916), .A2(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT39), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n652), .A2(new_n704), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n914), .A2(KEYINPUT39), .A3(new_n916), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n924), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n918), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(KEYINPUT103), .B1(new_n739), .B2(new_n474), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT103), .ZN(new_n930));
  NAND4_X1  g0730(.A1(new_n662), .A2(new_n930), .A3(new_n738), .A4(new_n735), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(new_n661), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n928), .B(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(G330), .ZN(new_n935));
  INV_X1    g0735(.A(new_n850), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n936), .B1(new_n891), .B2(new_n893), .ZN(new_n937));
  INV_X1    g0737(.A(new_n559), .ZN(new_n938));
  NAND4_X1  g0738(.A1(new_n701), .A2(new_n938), .A3(new_n638), .A4(new_n693), .ZN(new_n939));
  AND3_X1   g0739(.A1(new_n758), .A2(KEYINPUT31), .A3(new_n704), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n940), .A2(new_n759), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n922), .A2(new_n937), .A3(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(KEYINPUT40), .ZN(new_n944));
  AOI221_X4 g0744(.A(new_n936), .B1(new_n939), .B2(new_n941), .C1(new_n891), .C2(new_n893), .ZN(new_n945));
  AOI21_X1  g0745(.A(KEYINPUT40), .B1(new_n914), .B2(new_n916), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n944), .A2(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n474), .B1(new_n939), .B2(new_n941), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n935), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(new_n949), .B2(new_n948), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n934), .A2(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n952), .B1(new_n206), .B2(new_n766), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n934), .A2(new_n951), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n889), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  XOR2_X1   g0755(.A(new_n955), .B(KEYINPUT104), .Z(G367));
  OAI211_X1 g0756(.A(new_n553), .B(new_n558), .C1(new_n552), .C2(new_n693), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n671), .A2(new_n554), .A3(new_n704), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  OR2_X1    g0760(.A1(new_n717), .A2(new_n960), .ZN(new_n961));
  OR2_X1    g0761(.A1(new_n961), .A2(KEYINPUT42), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n558), .B1(new_n957), .B2(new_n609), .ZN(new_n963));
  AOI22_X1  g0763(.A1(new_n961), .A2(KEYINPUT42), .B1(new_n693), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n494), .A2(new_n704), .ZN(new_n965));
  MUX2_X1   g0765(.A(new_n682), .B(new_n683), .S(new_n965), .Z(new_n966));
  XOR2_X1   g0766(.A(new_n966), .B(KEYINPUT105), .Z(new_n967));
  AOI22_X1  g0767(.A1(new_n962), .A2(new_n964), .B1(KEYINPUT43), .B2(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(KEYINPUT43), .B2(new_n967), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT43), .ZN(new_n970));
  INV_X1    g0770(.A(new_n967), .ZN(new_n971));
  NAND4_X1  g0771(.A1(new_n962), .A2(new_n964), .A3(new_n970), .A4(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n969), .A2(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(new_n713), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n974), .A2(new_n959), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n973), .B1(KEYINPUT106), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(KEYINPUT106), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n973), .A2(KEYINPUT106), .A3(new_n975), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n720), .B(KEYINPUT41), .Z(new_n980));
  NAND3_X1  g0780(.A1(new_n717), .A2(new_n714), .A3(new_n959), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT107), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND4_X1  g0783(.A1(new_n717), .A2(KEYINPUT107), .A3(new_n714), .A4(new_n959), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  XNOR2_X1  g0785(.A(KEYINPUT108), .B(KEYINPUT45), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n959), .B1(new_n717), .B2(new_n714), .ZN(new_n988));
  OR2_X1    g0788(.A1(new_n988), .A2(KEYINPUT44), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n988), .A2(KEYINPUT44), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(new_n986), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n983), .A2(new_n984), .A3(new_n992), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n987), .A2(new_n991), .A3(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(new_n974), .ZN(new_n995));
  AOI22_X1  g0795(.A1(new_n985), .A2(new_n986), .B1(new_n989), .B2(new_n990), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n996), .A2(new_n713), .A3(new_n993), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n703), .A2(new_n705), .A3(new_n715), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n998), .A2(new_n717), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(new_n712), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n1000), .A2(new_n764), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n995), .A2(new_n997), .A3(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n980), .B1(new_n1003), .B2(new_n764), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n978), .B(new_n979), .C1(new_n1004), .C2(new_n770), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n771), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n786), .B1(new_n210), .B2(new_n459), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1007), .B1(new_n777), .B2(new_n237), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(new_n791), .A2(G294), .B1(G97), .B2(new_n812), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n1009), .B1(new_n857), .B2(new_n800), .C1(new_n451), .C2(new_n797), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n811), .A2(G116), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n1011), .B(KEYINPUT46), .Z(new_n1012));
  NOR2_X1   g0812(.A1(new_n830), .A2(new_n615), .ZN(new_n1013));
  INV_X1    g0813(.A(G283), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n296), .B1(new_n805), .B2(new_n792), .C1(new_n1014), .C2(new_n803), .ZN(new_n1015));
  NOR4_X1   g0815(.A1(new_n1010), .A2(new_n1012), .A3(new_n1013), .A4(new_n1015), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n791), .A2(G159), .B1(G77), .B2(new_n812), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1017), .B1(new_n866), .B2(new_n800), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n277), .B1(new_n808), .B2(new_n422), .ZN(new_n1019));
  INV_X1    g0819(.A(G137), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n803), .A2(new_n202), .B1(new_n805), .B2(new_n1020), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n872), .A2(new_n219), .B1(new_n248), .B2(new_n797), .ZN(new_n1022));
  NOR4_X1   g0822(.A1(new_n1018), .A2(new_n1019), .A3(new_n1021), .A4(new_n1022), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n1016), .A2(new_n1023), .ZN(new_n1024));
  XOR2_X1   g0824(.A(new_n1024), .B(KEYINPUT47), .Z(new_n1025));
  AOI211_X1 g0825(.A(new_n1006), .B(new_n1008), .C1(new_n1025), .C2(new_n785), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1026), .B1(new_n967), .B2(new_n835), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1005), .A2(new_n1027), .ZN(G387));
  NOR2_X1   g0828(.A1(new_n1000), .A2(new_n764), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n720), .ZN(new_n1030));
  OR3_X1    g0830(.A1(new_n1002), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n703), .A2(new_n705), .A3(new_n784), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n778), .B1(new_n234), .B2(G45), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1033), .B1(new_n722), .B2(new_n774), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n282), .B1(new_n248), .B2(new_n260), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT50), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1036), .B1(new_n456), .B2(new_n202), .ZN(new_n1037));
  NOR3_X1   g0837(.A1(new_n366), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1038));
  NOR4_X1   g0838(.A1(new_n722), .A2(new_n1035), .A3(new_n1037), .A4(new_n1038), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n1034), .A2(new_n1039), .B1(G107), .B2(new_n210), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1006), .B1(new_n1040), .B2(new_n786), .ZN(new_n1041));
  XOR2_X1   g0841(.A(new_n1041), .B(KEYINPUT109), .Z(new_n1042));
  AOI22_X1  g0842(.A1(new_n791), .A2(G311), .B1(new_n804), .B2(G303), .ZN(new_n1043));
  INV_X1    g0843(.A(G322), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n1043), .B1(new_n1044), .B2(new_n800), .C1(new_n830), .C2(new_n792), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT48), .ZN(new_n1046));
  OR2_X1    g0846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n797), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n1049), .A2(G283), .B1(G294), .B2(new_n811), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1047), .A2(new_n1048), .A3(new_n1050), .ZN(new_n1051));
  INV_X1    g0851(.A(KEYINPUT49), .ZN(new_n1052));
  AND2_X1   g0852(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n296), .B1(new_n798), .B2(new_n805), .C1(new_n821), .C2(new_n502), .ZN(new_n1055));
  OR3_X1    g0855(.A1(new_n1053), .A2(new_n1054), .A3(new_n1055), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n791), .A2(new_n456), .B1(new_n804), .B2(G68), .ZN(new_n1057));
  XOR2_X1   g0857(.A(new_n1057), .B(KEYINPUT110), .Z(new_n1058));
  OAI221_X1 g0858(.A(new_n277), .B1(new_n805), .B2(new_n422), .C1(new_n808), .C2(new_n202), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n821), .A2(new_n221), .B1(new_n797), .B2(new_n459), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n800), .A2(new_n826), .B1(new_n260), .B2(new_n872), .ZN(new_n1061));
  OR4_X1    g0861(.A1(new_n1058), .A2(new_n1059), .A3(new_n1060), .A4(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n854), .B1(new_n1056), .B2(new_n1062), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n1042), .A2(new_n1063), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n1000), .A2(new_n770), .B1(new_n1032), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1031), .A2(new_n1065), .ZN(G393));
  NAND2_X1  g0866(.A1(new_n1003), .A2(new_n720), .ZN(new_n1067));
  AND2_X1   g0867(.A1(new_n995), .A2(new_n997), .ZN(new_n1068));
  OAI21_X1  g0868(.A(KEYINPUT111), .B1(new_n1068), .B2(new_n1002), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n995), .A2(new_n997), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT111), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1070), .A2(new_n1071), .A3(new_n1001), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1067), .B1(new_n1069), .B2(new_n1072), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n786), .B1(new_n221), .B2(new_n210), .C1(new_n778), .C2(new_n244), .ZN(new_n1074));
  AND2_X1   g0874(.A1(new_n1074), .A2(new_n771), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n797), .A2(new_n260), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n1076), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1077), .B1(new_n248), .B2(new_n872), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n820), .A2(new_n202), .B1(new_n491), .B2(new_n821), .ZN(new_n1079));
  OAI221_X1 g0879(.A(new_n277), .B1(new_n805), .B2(new_n866), .C1(new_n366), .C2(new_n803), .ZN(new_n1080));
  NOR3_X1   g0880(.A1(new_n1078), .A2(new_n1079), .A3(new_n1080), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n800), .A2(new_n422), .B1(new_n826), .B2(new_n808), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1082), .B(KEYINPUT51), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n800), .A2(new_n792), .B1(new_n857), .B2(new_n808), .ZN(new_n1084));
  XNOR2_X1  g0884(.A(new_n1084), .B(KEYINPUT52), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n820), .A2(new_n615), .B1(new_n544), .B2(new_n821), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n296), .B1(new_n805), .B2(new_n1044), .C1(new_n599), .C2(new_n803), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n872), .A2(new_n1014), .B1(new_n502), .B2(new_n797), .ZN(new_n1088));
  NOR3_X1   g0888(.A1(new_n1086), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n1081), .A2(new_n1083), .B1(new_n1085), .B2(new_n1089), .ZN(new_n1090));
  OAI221_X1 g0890(.A(new_n1075), .B1(new_n1090), .B2(new_n854), .C1(new_n959), .C2(new_n835), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n770), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1091), .B1(new_n1070), .B2(new_n1092), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n1073), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1094), .ZN(G390));
  AOI21_X1  g0895(.A(new_n935), .B1(new_n939), .B2(new_n941), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n662), .A2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n932), .A2(new_n661), .A3(new_n1097), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n894), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1096), .A2(new_n850), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n693), .B(new_n846), .C1(new_n733), .C2(new_n734), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1102), .A2(new_n896), .ZN(new_n1103));
  OAI211_X1 g0903(.A(G330), .B(new_n850), .C1(new_n761), .C2(new_n762), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1103), .B1(new_n1105), .B2(new_n894), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1104), .A2(new_n891), .A3(new_n893), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n894), .A2(new_n850), .A3(new_n1096), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n1101), .A2(new_n1106), .B1(new_n1109), .B2(new_n897), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n1098), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(KEYINPUT112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n924), .A2(new_n926), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n925), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n898), .A2(new_n1115), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n1102), .A2(new_n896), .B1(new_n891), .B2(new_n893), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n925), .B1(new_n916), .B2(new_n921), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n1114), .A2(new_n1116), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1105), .A2(new_n894), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1113), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  AND3_X1   g0922(.A1(new_n914), .A2(KEYINPUT39), .A3(new_n916), .ZN(new_n1123));
  AOI21_X1  g0923(.A(KEYINPUT39), .B1(new_n916), .B2(new_n921), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1116), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n1125), .A2(new_n1126), .A3(new_n1113), .A4(new_n1121), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1108), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n924), .A2(new_n926), .B1(new_n898), .B2(new_n1115), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1119), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n1130), .A2(new_n1117), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1128), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1127), .A2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1112), .B1(new_n1122), .B2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1125), .A2(new_n1126), .A3(new_n1121), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1135), .A2(KEYINPUT112), .ZN(new_n1136));
  NAND4_X1  g0936(.A1(new_n1111), .A2(new_n1136), .A3(new_n1132), .A4(new_n1127), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1134), .A2(new_n720), .A3(new_n1137), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n1133), .A2(new_n1122), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1114), .A2(new_n782), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n771), .B1(new_n456), .B2(new_n855), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n791), .A2(G137), .B1(G50), .B2(new_n812), .ZN(new_n1142));
  INV_X1    g0942(.A(G128), .ZN(new_n1143));
  OAI221_X1 g0943(.A(new_n1142), .B1(new_n1143), .B2(new_n800), .C1(new_n826), .C2(new_n797), .ZN(new_n1144));
  OR3_X1    g0944(.A1(new_n872), .A2(KEYINPUT53), .A3(new_n422), .ZN(new_n1145));
  OAI21_X1  g0945(.A(KEYINPUT53), .B1(new_n872), .B2(new_n422), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(KEYINPUT54), .B(G143), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n296), .B1(new_n804), .B2(new_n1148), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(G132), .A2(new_n809), .B1(new_n806), .B2(G125), .ZN(new_n1150));
  NAND4_X1  g0950(.A1(new_n1145), .A2(new_n1146), .A3(new_n1149), .A4(new_n1150), .ZN(new_n1151));
  OAI221_X1 g0951(.A(new_n1077), .B1(new_n820), .B2(new_n451), .C1(new_n1014), .C2(new_n800), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(G116), .A2(new_n809), .B1(new_n806), .B2(G294), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n277), .B1(new_n804), .B2(G97), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n1153), .A2(new_n817), .A3(new_n871), .A4(new_n1154), .ZN(new_n1155));
  OAI22_X1  g0955(.A1(new_n1144), .A2(new_n1151), .B1(new_n1152), .B2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1141), .B1(new_n1156), .B2(new_n785), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(new_n1139), .A2(new_n770), .B1(new_n1140), .B2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1138), .A2(new_n1158), .ZN(G378));
  XOR2_X1   g0959(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(KEYINPUT115), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n438), .A2(new_n443), .ZN(new_n1163));
  AND2_X1   g0963(.A1(new_n440), .A2(new_n692), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1164), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n438), .A2(new_n443), .A3(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1162), .B1(new_n1165), .B2(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1166), .B1(new_n438), .B2(new_n443), .ZN(new_n1169));
  AOI211_X1 g0969(.A(new_n442), .B(new_n1164), .C1(new_n435), .C2(new_n437), .ZN(new_n1170));
  NOR3_X1   g0970(.A1(new_n1169), .A2(new_n1170), .A3(KEYINPUT115), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1161), .B1(new_n1168), .B2(new_n1171), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1165), .A2(new_n1162), .A3(new_n1167), .ZN(new_n1173));
  OAI21_X1  g0973(.A(KEYINPUT115), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1173), .A2(new_n1174), .A3(new_n1160), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1172), .A2(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1177), .B1(new_n948), .B2(G330), .ZN(new_n1178));
  AOI211_X1 g0978(.A(new_n935), .B(new_n1176), .C1(new_n944), .C2(new_n947), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n928), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(new_n943), .A2(KEYINPUT40), .B1(new_n945), .B2(new_n946), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1176), .B1(new_n1181), .B2(new_n935), .ZN(new_n1182));
  INV_X1    g0982(.A(KEYINPUT40), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(new_n945), .B2(new_n922), .ZN(new_n1184));
  NOR3_X1   g0984(.A1(new_n902), .A2(new_n900), .A3(new_n913), .ZN(new_n1185));
  AND3_X1   g0985(.A1(new_n392), .A2(KEYINPUT77), .A3(new_n393), .ZN(new_n1186));
  AOI21_X1  g0986(.A(KEYINPUT77), .B1(new_n392), .B2(new_n393), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n648), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1188), .A2(new_n903), .ZN(new_n1189));
  AOI21_X1  g0989(.A(KEYINPUT38), .B1(new_n1189), .B2(new_n915), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1183), .B1(new_n1185), .B2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n937), .A2(new_n942), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  OAI211_X1 g0993(.A(G330), .B(new_n1177), .C1(new_n1184), .C2(new_n1193), .ZN(new_n1194));
  AND2_X1   g0994(.A1(new_n918), .A2(new_n927), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1182), .A2(new_n1194), .A3(new_n1195), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1180), .A2(KEYINPUT116), .A3(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1195), .B1(new_n1182), .B2(new_n1194), .ZN(new_n1198));
  INV_X1    g0998(.A(KEYINPUT116), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1197), .A2(new_n770), .A3(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1176), .A2(new_n782), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n771), .B1(G50), .B2(new_n855), .ZN(new_n1203));
  OAI22_X1  g1003(.A1(new_n808), .A2(new_n1143), .B1(new_n803), .B2(new_n1020), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n799), .A2(G125), .ZN(new_n1205));
  OAI221_X1 g1005(.A(new_n1205), .B1(new_n872), .B2(new_n1147), .C1(new_n820), .C2(new_n869), .ZN(new_n1206));
  AOI211_X1 g1006(.A(new_n1204), .B(new_n1206), .C1(G150), .C2(new_n1049), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT59), .ZN(new_n1208));
  OR2_X1    g1008(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n812), .A2(G159), .ZN(new_n1211));
  AOI211_X1 g1011(.A(G33), .B(G41), .C1(new_n806), .C2(G124), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n1209), .A2(new_n1210), .A3(new_n1211), .A4(new_n1212), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n791), .A2(G97), .B1(new_n804), .B2(new_n460), .ZN(new_n1214));
  XNOR2_X1  g1014(.A(new_n1214), .B(KEYINPUT114), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n296), .A2(new_n281), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1216), .B1(new_n806), .B2(G283), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n809), .A2(G107), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n872), .A2(new_n260), .B1(new_n248), .B2(new_n797), .ZN(new_n1220));
  OAI22_X1  g1020(.A1(new_n800), .A2(new_n502), .B1(new_n219), .B2(new_n821), .ZN(new_n1221));
  NOR4_X1   g1021(.A1(new_n1215), .A2(new_n1219), .A3(new_n1220), .A4(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1222), .A2(KEYINPUT58), .ZN(new_n1223));
  OR2_X1    g1023(.A1(new_n1222), .A2(KEYINPUT58), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n1216), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1225));
  XOR2_X1   g1025(.A(new_n1225), .B(KEYINPUT113), .Z(new_n1226));
  NAND4_X1  g1026(.A1(new_n1213), .A2(new_n1223), .A3(new_n1224), .A4(new_n1226), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1203), .B1(new_n1227), .B2(new_n785), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1202), .A2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1201), .A2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1098), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1137), .A2(new_n1232), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1233), .A2(new_n1197), .A3(new_n1200), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT57), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT117), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1098), .B1(new_n1139), .B2(new_n1111), .ZN(new_n1238));
  AND3_X1   g1038(.A1(new_n1182), .A2(new_n1194), .A3(new_n1195), .ZN(new_n1239));
  OAI21_X1  g1039(.A(KEYINPUT57), .B1(new_n1239), .B2(new_n1198), .ZN(new_n1240));
  OAI211_X1 g1040(.A(new_n1237), .B(new_n720), .C1(new_n1238), .C2(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1236), .A2(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1235), .B1(new_n1180), .B2(new_n1196), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1030), .B1(new_n1243), .B2(new_n1233), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1244), .A2(new_n1237), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1231), .B1(new_n1242), .B2(new_n1245), .ZN(G375));
  INV_X1    g1046(.A(new_n980), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1098), .A2(new_n1110), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1112), .A2(new_n1247), .A3(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1110), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1099), .A2(new_n782), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n771), .B1(G68), .B2(new_n855), .ZN(new_n1252));
  OAI22_X1  g1052(.A1(new_n800), .A2(new_n599), .B1(new_n221), .B2(new_n872), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1253), .B1(G116), .B2(new_n791), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n277), .B1(new_n804), .B2(new_n538), .ZN(new_n1255));
  AOI22_X1  g1055(.A1(G283), .A2(new_n809), .B1(new_n806), .B2(G303), .ZN(new_n1256));
  AOI22_X1  g1056(.A1(new_n1049), .A2(new_n460), .B1(G77), .B2(new_n812), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1254), .A2(new_n1255), .A3(new_n1256), .A4(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n799), .A2(G132), .ZN(new_n1259));
  XOR2_X1   g1059(.A(new_n1259), .B(KEYINPUT118), .Z(new_n1260));
  OAI21_X1  g1060(.A(new_n277), .B1(new_n803), .B2(new_n422), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1261), .B1(G128), .B2(new_n806), .ZN(new_n1262));
  OAI211_X1 g1062(.A(new_n1260), .B(new_n1262), .C1(new_n1020), .C2(new_n830), .ZN(new_n1263));
  AOI22_X1  g1063(.A1(new_n791), .A2(new_n1148), .B1(G159), .B2(new_n811), .ZN(new_n1264));
  OAI221_X1 g1064(.A(new_n1264), .B1(new_n202), .B2(new_n797), .C1(new_n219), .C2(new_n821), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1258), .B1(new_n1263), .B2(new_n1265), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1252), .B1(new_n1266), .B2(new_n785), .ZN(new_n1267));
  AOI22_X1  g1067(.A1(new_n1250), .A2(new_n770), .B1(new_n1251), .B2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1249), .A2(new_n1268), .ZN(new_n1269));
  XOR2_X1   g1069(.A(new_n1269), .B(KEYINPUT119), .Z(G381));
  XNOR2_X1  g1070(.A(G375), .B(KEYINPUT120), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1031), .A2(new_n837), .A3(new_n1065), .ZN(new_n1272));
  OR4_X1    g1072(.A1(G384), .A2(G390), .A3(G387), .A4(new_n1272), .ZN(new_n1273));
  OR4_X1    g1073(.A1(G378), .A2(new_n1271), .A3(G381), .A4(new_n1273), .ZN(G407));
  INV_X1    g1074(.A(G378), .ZN(new_n1275));
  INV_X1    g1075(.A(G213), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1276), .A2(G343), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1275), .A2(new_n1277), .ZN(new_n1278));
  OAI211_X1 g1078(.A(G407), .B(G213), .C1(new_n1271), .C2(new_n1278), .ZN(G409));
  INV_X1    g1079(.A(KEYINPUT123), .ZN(new_n1280));
  OAI211_X1 g1080(.A(G378), .B(new_n1231), .C1(new_n1242), .C2(new_n1245), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1180), .A2(new_n1196), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(new_n770), .ZN(new_n1283));
  OAI211_X1 g1083(.A(new_n1229), .B(new_n1283), .C1(new_n1234), .C2(new_n980), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1284), .A2(new_n1275), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1281), .A2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1277), .ZN(new_n1287));
  AND3_X1   g1087(.A1(new_n1248), .A2(KEYINPUT121), .A3(KEYINPUT60), .ZN(new_n1288));
  AOI21_X1  g1088(.A(KEYINPUT60), .B1(new_n1248), .B2(KEYINPUT121), .ZN(new_n1289));
  OAI211_X1 g1089(.A(new_n720), .B(new_n1112), .C1(new_n1288), .C2(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1290), .A2(new_n1268), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1291), .A2(new_n878), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1290), .A2(G384), .A3(new_n1268), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1294), .ZN(new_n1295));
  NAND4_X1  g1095(.A1(new_n1286), .A2(KEYINPUT122), .A3(new_n1287), .A4(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT63), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1277), .B1(new_n1281), .B2(new_n1285), .ZN(new_n1299));
  AOI21_X1  g1099(.A(KEYINPUT122), .B1(new_n1299), .B2(new_n1295), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1280), .B1(new_n1298), .B2(new_n1300), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1286), .A2(new_n1287), .A3(new_n1295), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT122), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1304));
  NAND4_X1  g1104(.A1(new_n1304), .A2(KEYINPUT123), .A3(new_n1297), .A4(new_n1296), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(G387), .A2(new_n1094), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT125), .ZN(new_n1307));
  OAI211_X1 g1107(.A(new_n1005), .B(new_n1027), .C1(new_n1073), .C2(new_n1093), .ZN(new_n1308));
  AND3_X1   g1108(.A1(new_n1306), .A2(new_n1307), .A3(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(G393), .A2(G396), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1310), .A2(new_n1272), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT124), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1310), .A2(KEYINPUT124), .A3(new_n1272), .ZN(new_n1314));
  OAI211_X1 g1114(.A(new_n1313), .B(new_n1314), .C1(new_n1308), .C2(new_n1307), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT126), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n1316), .B1(new_n1005), .B2(new_n1027), .ZN(new_n1317));
  AND2_X1   g1117(.A1(new_n1317), .A2(new_n1094), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1311), .B1(new_n1317), .B2(new_n1094), .ZN(new_n1319));
  OAI22_X1  g1119(.A1(new_n1309), .A2(new_n1315), .B1(new_n1318), .B2(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT61), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1277), .A2(G2897), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1292), .A2(new_n1293), .A3(new_n1322), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1323), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n1322), .B1(new_n1292), .B2(new_n1293), .ZN(new_n1325));
  OR2_X1    g1125(.A1(new_n1324), .A2(new_n1325), .ZN(new_n1326));
  OAI211_X1 g1126(.A(new_n1320), .B(new_n1321), .C1(new_n1299), .C2(new_n1326), .ZN(new_n1327));
  AND3_X1   g1127(.A1(new_n1299), .A2(KEYINPUT63), .A3(new_n1295), .ZN(new_n1328));
  NOR2_X1   g1128(.A1(new_n1327), .A2(new_n1328), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1301), .A2(new_n1305), .A3(new_n1329), .ZN(new_n1330));
  INV_X1    g1130(.A(new_n1320), .ZN(new_n1331));
  NOR2_X1   g1131(.A1(new_n1324), .A2(new_n1325), .ZN(new_n1332));
  AND2_X1   g1132(.A1(new_n1284), .A2(new_n1275), .ZN(new_n1333));
  AOI22_X1  g1133(.A1(new_n1244), .A2(new_n1237), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n720), .B1(new_n1238), .B2(new_n1240), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1335), .A2(KEYINPUT117), .ZN(new_n1336));
  AOI21_X1  g1136(.A(new_n1230), .B1(new_n1334), .B2(new_n1336), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n1333), .B1(new_n1337), .B2(G378), .ZN(new_n1338));
  OAI21_X1  g1138(.A(new_n1332), .B1(new_n1338), .B2(new_n1277), .ZN(new_n1339));
  AOI211_X1 g1139(.A(new_n1277), .B(new_n1294), .C1(new_n1281), .C2(new_n1285), .ZN(new_n1340));
  AOI21_X1  g1140(.A(new_n1303), .B1(KEYINPUT127), .B2(KEYINPUT62), .ZN(new_n1341));
  OAI211_X1 g1141(.A(new_n1339), .B(new_n1321), .C1(new_n1340), .C2(new_n1341), .ZN(new_n1342));
  AOI21_X1  g1142(.A(KEYINPUT62), .B1(new_n1296), .B2(KEYINPUT127), .ZN(new_n1343));
  OAI21_X1  g1143(.A(new_n1331), .B1(new_n1342), .B2(new_n1343), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1330), .A2(new_n1344), .ZN(G405));
  NOR2_X1   g1145(.A1(new_n1337), .A2(G378), .ZN(new_n1346));
  INV_X1    g1146(.A(new_n1281), .ZN(new_n1347));
  OR3_X1    g1147(.A1(new_n1346), .A2(new_n1347), .A3(new_n1295), .ZN(new_n1348));
  OAI21_X1  g1148(.A(new_n1295), .B1(new_n1346), .B2(new_n1347), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1348), .A2(new_n1349), .ZN(new_n1350));
  XNOR2_X1  g1150(.A(new_n1350), .B(new_n1331), .ZN(G402));
endmodule


