//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 0 0 0 1 1 1 0 1 0 1 0 1 0 1 0 0 0 0 1 1 1 1 0 1 1 1 0 0 0 1 1 1 0 0 1 0 1 1 1 1 1 1 1 1 0 1 0 0 0 1 0 1 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:30 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n775, new_n776, new_n777, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n789, new_n790,
    new_n791, new_n793, new_n794, new_n795, new_n796, new_n797, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n805, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n847, new_n848, new_n849, new_n850, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n918, new_n919,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n975, new_n976, new_n978, new_n979, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n992, new_n993, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1043, new_n1044,
    new_n1045, new_n1046;
  INV_X1    g000(.A(G169gat), .ZN(new_n202));
  INV_X1    g001(.A(G176gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT26), .ZN(new_n205));
  INV_X1    g004(.A(G183gat), .ZN(new_n206));
  INV_X1    g005(.A(G190gat), .ZN(new_n207));
  OAI22_X1  g006(.A1(new_n204), .A2(new_n205), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(G169gat), .A2(G176gat), .ZN(new_n209));
  NOR2_X1   g008(.A1(G169gat), .A2(G176gat), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n210), .A2(KEYINPUT26), .ZN(new_n211));
  AOI21_X1  g010(.A(new_n208), .B1(new_n209), .B2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n206), .A2(KEYINPUT27), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT27), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(G183gat), .ZN(new_n215));
  AND2_X1   g014(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n216), .A2(KEYINPUT28), .A3(new_n207), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n213), .A2(new_n215), .A3(new_n207), .ZN(new_n218));
  AND2_X1   g017(.A1(KEYINPUT67), .A2(KEYINPUT28), .ZN(new_n219));
  NOR2_X1   g018(.A1(KEYINPUT67), .A2(KEYINPUT28), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n218), .A2(KEYINPUT68), .A3(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n217), .A2(new_n222), .ZN(new_n223));
  AOI21_X1  g022(.A(KEYINPUT68), .B1(new_n218), .B2(new_n221), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n212), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n207), .A2(G183gat), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n206), .A2(G190gat), .ZN(new_n227));
  OAI21_X1  g026(.A(KEYINPUT24), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT23), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n229), .A2(G176gat), .ZN(new_n230));
  OR2_X1    g029(.A1(KEYINPUT64), .A2(G169gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(KEYINPUT64), .A2(G169gat), .ZN(new_n232));
  NAND4_X1  g031(.A1(new_n230), .A2(new_n231), .A3(KEYINPUT65), .A4(new_n232), .ZN(new_n233));
  NOR3_X1   g032(.A1(new_n206), .A2(new_n207), .A3(KEYINPUT24), .ZN(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  AND3_X1   g034(.A1(new_n228), .A2(new_n233), .A3(new_n235), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n210), .B1(KEYINPUT23), .B2(new_n209), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n230), .A2(new_n231), .A3(new_n232), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT65), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n237), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  AOI21_X1  g039(.A(KEYINPUT25), .B1(new_n236), .B2(new_n240), .ZN(new_n241));
  OAI21_X1  g040(.A(KEYINPUT25), .B1(new_n204), .B2(new_n229), .ZN(new_n242));
  OR2_X1    g041(.A1(new_n242), .A2(new_n237), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT66), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n228), .A2(new_n235), .A3(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT24), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n206), .A2(G190gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n207), .A2(G183gat), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n246), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  OAI21_X1  g048(.A(KEYINPUT66), .B1(new_n249), .B2(new_n234), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n243), .B1(new_n245), .B2(new_n250), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n225), .B1(new_n241), .B2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(G113gat), .ZN(new_n253));
  INV_X1    g052(.A(G120gat), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT1), .ZN(new_n256));
  NAND2_X1  g055(.A1(G113gat), .A2(G120gat), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n255), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  OR2_X1    g057(.A1(G127gat), .A2(G134gat), .ZN(new_n259));
  INV_X1    g058(.A(G127gat), .ZN(new_n260));
  XNOR2_X1  g059(.A(KEYINPUT69), .B(G134gat), .ZN(new_n261));
  OAI211_X1 g060(.A(new_n258), .B(new_n259), .C1(new_n260), .C2(new_n261), .ZN(new_n262));
  AOI21_X1  g061(.A(KEYINPUT1), .B1(new_n253), .B2(new_n254), .ZN(new_n263));
  XNOR2_X1  g062(.A(G127gat), .B(G134gat), .ZN(new_n264));
  XNOR2_X1  g063(.A(KEYINPUT70), .B(G113gat), .ZN(new_n265));
  OAI211_X1 g064(.A(new_n263), .B(new_n264), .C1(new_n265), .C2(new_n254), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n262), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(G227gat), .A2(G233gat), .ZN(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  OAI211_X1 g070(.A(new_n225), .B(new_n267), .C1(new_n241), .C2(new_n251), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n269), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(KEYINPUT32), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT33), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  XOR2_X1   g075(.A(G15gat), .B(G43gat), .Z(new_n277));
  XNOR2_X1  g076(.A(G71gat), .B(G99gat), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n277), .B(new_n278), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n274), .A2(new_n276), .A3(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n272), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT25), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n238), .A2(new_n239), .ZN(new_n283));
  INV_X1    g082(.A(new_n237), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n228), .A2(new_n233), .A3(new_n235), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n282), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n242), .A2(new_n237), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n244), .B1(new_n228), .B2(new_n235), .ZN(new_n289));
  NOR3_X1   g088(.A1(new_n249), .A2(KEYINPUT66), .A3(new_n234), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n288), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n287), .A2(new_n291), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n267), .B1(new_n292), .B2(new_n225), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n270), .B1(new_n281), .B2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT34), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n295), .B1(new_n270), .B2(KEYINPUT71), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n269), .A2(new_n272), .ZN(new_n298));
  INV_X1    g097(.A(new_n296), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n298), .A2(new_n270), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n279), .ZN(new_n302));
  OAI211_X1 g101(.A(new_n273), .B(KEYINPUT32), .C1(new_n275), .C2(new_n302), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n280), .A2(new_n301), .A3(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n301), .B1(new_n280), .B2(new_n303), .ZN(new_n306));
  NOR3_X1   g105(.A1(new_n305), .A2(new_n306), .A3(KEYINPUT36), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT72), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n301), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n280), .A2(new_n303), .ZN(new_n310));
  INV_X1    g109(.A(new_n301), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  OAI211_X1 g111(.A(new_n304), .B(new_n309), .C1(new_n312), .C2(new_n308), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n307), .B1(KEYINPUT36), .B2(new_n313), .ZN(new_n314));
  AND2_X1   g113(.A1(G155gat), .A2(G162gat), .ZN(new_n315));
  NOR2_X1   g114(.A1(G155gat), .A2(G162gat), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(G141gat), .B(G148gat), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT2), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n319), .B1(G155gat), .B2(G162gat), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n317), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(G141gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(G148gat), .ZN(new_n323));
  INV_X1    g122(.A(G148gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(G141gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(G155gat), .B(G162gat), .ZN(new_n327));
  INV_X1    g126(.A(G155gat), .ZN(new_n328));
  INV_X1    g127(.A(G162gat), .ZN(new_n329));
  OAI21_X1  g128(.A(KEYINPUT2), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n326), .A2(new_n327), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n321), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(KEYINPUT3), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT3), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n321), .A2(new_n331), .A3(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n333), .A2(new_n335), .A3(new_n267), .ZN(new_n336));
  NAND4_X1  g135(.A1(new_n262), .A2(new_n266), .A3(new_n321), .A4(new_n331), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(KEYINPUT4), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n337), .A2(KEYINPUT4), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n336), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(G225gat), .A2(G233gat), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n267), .A2(new_n332), .ZN(new_n345));
  AOI22_X1  g144(.A1(new_n262), .A2(new_n266), .B1(new_n321), .B2(new_n331), .ZN(new_n346));
  OR3_X1    g145(.A1(new_n345), .A2(new_n343), .A3(new_n346), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n344), .A2(KEYINPUT39), .A3(new_n347), .ZN(new_n348));
  XNOR2_X1  g147(.A(G1gat), .B(G29gat), .ZN(new_n349));
  XNOR2_X1  g148(.A(new_n349), .B(KEYINPUT0), .ZN(new_n350));
  XNOR2_X1  g149(.A(G57gat), .B(G85gat), .ZN(new_n351));
  XOR2_X1   g150(.A(new_n350), .B(new_n351), .Z(new_n352));
  INV_X1    g151(.A(KEYINPUT39), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n341), .A2(new_n353), .A3(new_n343), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n348), .A2(new_n352), .A3(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT40), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(new_n352), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n343), .B1(new_n345), .B2(new_n346), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(KEYINPUT5), .ZN(new_n360));
  AND2_X1   g159(.A1(new_n336), .A2(new_n342), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT77), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT4), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n345), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  OAI21_X1  g163(.A(KEYINPUT77), .B1(new_n337), .B2(KEYINPUT4), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n364), .A2(new_n365), .A3(new_n338), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n360), .B1(new_n361), .B2(new_n366), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n339), .A2(new_n340), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT5), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n336), .A2(new_n369), .A3(new_n342), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n358), .B1(new_n367), .B2(new_n371), .ZN(new_n372));
  NAND4_X1  g171(.A1(new_n348), .A2(KEYINPUT40), .A3(new_n352), .A4(new_n354), .ZN(new_n373));
  AND3_X1   g172(.A1(new_n357), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(G211gat), .A2(G218gat), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT22), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NOR2_X1   g176(.A1(G197gat), .A2(G204gat), .ZN(new_n378));
  AND2_X1   g177(.A1(G197gat), .A2(G204gat), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n377), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  XOR2_X1   g179(.A(G211gat), .B(G218gat), .Z(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  XNOR2_X1  g181(.A(G211gat), .B(G218gat), .ZN(new_n383));
  XNOR2_X1  g182(.A(G197gat), .B(G204gat), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n383), .A2(new_n384), .A3(new_n377), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n382), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(G226gat), .A2(G233gat), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT29), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n389), .B1(new_n252), .B2(new_n390), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n388), .B1(new_n292), .B2(new_n225), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n387), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  XOR2_X1   g192(.A(G8gat), .B(G36gat), .Z(new_n394));
  XNOR2_X1  g193(.A(new_n394), .B(KEYINPUT73), .ZN(new_n395));
  XNOR2_X1  g194(.A(G64gat), .B(G92gat), .ZN(new_n396));
  XNOR2_X1  g195(.A(new_n395), .B(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n218), .A2(new_n221), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT68), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n400), .A2(new_n217), .A3(new_n222), .ZN(new_n401));
  AOI22_X1  g200(.A1(new_n287), .A2(new_n291), .B1(new_n401), .B2(new_n212), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n388), .B1(new_n402), .B2(KEYINPUT29), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n252), .A2(new_n389), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n403), .A2(new_n386), .A3(new_n404), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n393), .A2(new_n397), .A3(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT76), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT30), .ZN(new_n408));
  AND3_X1   g207(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n407), .B1(new_n406), .B2(new_n408), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n397), .ZN(new_n412));
  NOR3_X1   g211(.A1(new_n391), .A2(new_n387), .A3(new_n392), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n386), .B1(new_n403), .B2(new_n404), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n412), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT74), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND4_X1  g216(.A1(new_n393), .A2(new_n405), .A3(KEYINPUT30), .A4(new_n397), .ZN(new_n418));
  OAI211_X1 g217(.A(KEYINPUT74), .B(new_n412), .C1(new_n413), .C2(new_n414), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n417), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n374), .B1(new_n411), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n366), .A2(new_n361), .ZN(new_n422));
  INV_X1    g221(.A(new_n360), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n371), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n424), .A2(new_n425), .A3(new_n352), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT6), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n426), .A2(new_n372), .A3(new_n427), .ZN(new_n428));
  OAI211_X1 g227(.A(KEYINPUT6), .B(new_n358), .C1(new_n367), .C2(new_n371), .ZN(new_n429));
  AND3_X1   g228(.A1(new_n428), .A2(new_n429), .A3(new_n406), .ZN(new_n430));
  OAI21_X1  g229(.A(KEYINPUT37), .B1(new_n413), .B2(new_n414), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT37), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n393), .A2(new_n432), .A3(new_n405), .ZN(new_n433));
  XOR2_X1   g232(.A(KEYINPUT82), .B(KEYINPUT38), .Z(new_n434));
  NAND4_X1  g233(.A1(new_n431), .A2(new_n412), .A3(new_n433), .A4(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n431), .A2(new_n412), .A3(new_n433), .ZN(new_n436));
  INV_X1    g235(.A(new_n434), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n430), .A2(new_n435), .A3(new_n438), .ZN(new_n439));
  AND2_X1   g238(.A1(new_n421), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(G228gat), .A2(G233gat), .ZN(new_n441));
  AND2_X1   g240(.A1(new_n321), .A2(new_n331), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n380), .A2(new_n381), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n383), .B1(new_n377), .B2(new_n384), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n390), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n442), .B1(new_n445), .B2(new_n334), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n386), .B1(new_n335), .B2(new_n390), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n441), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n335), .A2(new_n390), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(new_n387), .ZN(new_n450));
  AOI21_X1  g249(.A(KEYINPUT29), .B1(new_n382), .B2(new_n385), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n332), .B1(new_n451), .B2(KEYINPUT3), .ZN(new_n452));
  INV_X1    g251(.A(new_n441), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n450), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n448), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(G22gat), .ZN(new_n456));
  XNOR2_X1  g255(.A(G78gat), .B(G106gat), .ZN(new_n457));
  XNOR2_X1  g256(.A(KEYINPUT31), .B(G50gat), .ZN(new_n458));
  XOR2_X1   g257(.A(new_n457), .B(new_n458), .Z(new_n459));
  INV_X1    g258(.A(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(G22gat), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n448), .A2(new_n461), .A3(new_n454), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n456), .A2(new_n460), .A3(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT78), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n448), .A2(KEYINPUT78), .A3(new_n461), .A4(new_n454), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n465), .A2(new_n466), .A3(new_n456), .ZN(new_n467));
  AND3_X1   g266(.A1(new_n467), .A2(KEYINPUT79), .A3(new_n459), .ZN(new_n468));
  AOI21_X1  g267(.A(KEYINPUT79), .B1(new_n467), .B2(new_n459), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n463), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(KEYINPUT80), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT80), .ZN(new_n472));
  OAI211_X1 g271(.A(new_n472), .B(new_n463), .C1(new_n468), .C2(new_n469), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n314), .B1(new_n440), .B2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT81), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n467), .A2(new_n459), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT79), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n467), .A2(KEYINPUT79), .A3(new_n459), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n472), .B1(new_n481), .B2(new_n463), .ZN(new_n482));
  INV_X1    g281(.A(new_n473), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n476), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT75), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n419), .A2(new_n418), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n393), .A2(new_n405), .ZN(new_n487));
  AOI21_X1  g286(.A(KEYINPUT74), .B1(new_n487), .B2(new_n412), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n485), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n406), .A2(new_n408), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(KEYINPUT76), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n417), .A2(KEYINPUT75), .A3(new_n418), .A4(new_n419), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n428), .A2(new_n429), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n489), .A2(new_n493), .A3(new_n494), .A4(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n471), .A2(KEYINPUT81), .A3(new_n473), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n484), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n475), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n313), .B1(new_n482), .B2(new_n483), .ZN(new_n500));
  OAI21_X1  g299(.A(KEYINPUT35), .B1(new_n500), .B2(new_n496), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n486), .A2(new_n488), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n493), .A2(new_n502), .A3(new_n495), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT83), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n305), .A2(new_n306), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n506), .A2(KEYINPUT35), .ZN(new_n507));
  NAND4_X1  g306(.A1(new_n493), .A2(new_n502), .A3(KEYINPUT83), .A4(new_n495), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n505), .A2(new_n474), .A3(new_n507), .A4(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n501), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT84), .ZN(new_n511));
  AND3_X1   g310(.A1(new_n499), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n511), .B1(new_n499), .B2(new_n510), .ZN(new_n513));
  NAND2_X1  g312(.A1(G229gat), .A2(G233gat), .ZN(new_n514));
  OAI21_X1  g313(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT85), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  OAI211_X1 g316(.A(KEYINPUT85), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  OR2_X1    g318(.A1(new_n519), .A2(KEYINPUT86), .ZN(new_n520));
  NOR3_X1   g319(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n521), .B1(new_n519), .B2(KEYINPUT86), .ZN(new_n522));
  XNOR2_X1  g321(.A(KEYINPUT87), .B(G36gat), .ZN(new_n523));
  AOI22_X1  g322(.A1(new_n520), .A2(new_n522), .B1(G29gat), .B2(new_n523), .ZN(new_n524));
  XNOR2_X1  g323(.A(G43gat), .B(G50gat), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(KEYINPUT15), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n523), .A2(G29gat), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n521), .B1(new_n517), .B2(new_n518), .ZN(new_n529));
  OR2_X1    g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(KEYINPUT88), .B(G43gat), .ZN(new_n531));
  INV_X1    g330(.A(G50gat), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  XNOR2_X1  g332(.A(KEYINPUT89), .B(G50gat), .ZN(new_n534));
  INV_X1    g333(.A(G43gat), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(KEYINPUT15), .B1(new_n533), .B2(new_n536), .ZN(new_n537));
  OAI22_X1  g336(.A1(new_n524), .A2(new_n526), .B1(new_n530), .B2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT17), .ZN(new_n539));
  AOI21_X1  g338(.A(KEYINPUT91), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(G8gat), .ZN(new_n541));
  XNOR2_X1  g340(.A(G15gat), .B(G22gat), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT90), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n542), .B(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(G1gat), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  OR2_X1    g345(.A1(new_n542), .A2(new_n543), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n542), .A2(new_n543), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT16), .ZN(new_n549));
  OAI211_X1 g348(.A(new_n547), .B(new_n548), .C1(new_n549), .C2(G1gat), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n541), .B1(new_n546), .B2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n546), .A2(new_n550), .A3(new_n541), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n540), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT91), .ZN(new_n556));
  AND3_X1   g355(.A1(new_n546), .A2(new_n550), .A3(new_n541), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n556), .B1(new_n557), .B2(new_n551), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n538), .B1(new_n558), .B2(new_n539), .ZN(new_n559));
  OAI211_X1 g358(.A(KEYINPUT18), .B(new_n514), .C1(new_n555), .C2(new_n559), .ZN(new_n560));
  OR2_X1    g359(.A1(new_n538), .A2(KEYINPUT93), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n538), .A2(KEYINPUT93), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n561), .A2(new_n554), .A3(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n554), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n564), .A2(KEYINPUT93), .A3(new_n538), .ZN(new_n565));
  XOR2_X1   g364(.A(new_n514), .B(KEYINPUT13), .Z(new_n566));
  NAND3_X1  g365(.A1(new_n563), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  AND2_X1   g366(.A1(new_n560), .A2(new_n567), .ZN(new_n568));
  AOI21_X1  g367(.A(KEYINPUT17), .B1(new_n554), .B2(new_n556), .ZN(new_n569));
  OAI22_X1  g368(.A1(new_n569), .A2(new_n538), .B1(new_n540), .B2(new_n554), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n570), .A2(new_n514), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT18), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT92), .ZN(new_n574));
  XNOR2_X1  g373(.A(G113gat), .B(G141gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n575), .B(G197gat), .ZN(new_n576));
  XOR2_X1   g375(.A(KEYINPUT11), .B(G169gat), .Z(new_n577));
  XNOR2_X1  g376(.A(new_n576), .B(new_n577), .ZN(new_n578));
  XOR2_X1   g377(.A(new_n578), .B(KEYINPUT12), .Z(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  OAI211_X1 g379(.A(new_n568), .B(new_n573), .C1(new_n574), .C2(new_n580), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n560), .A2(new_n567), .A3(new_n574), .ZN(new_n582));
  AOI21_X1  g381(.A(KEYINPUT18), .B1(new_n570), .B2(new_n514), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n560), .A2(new_n567), .ZN(new_n584));
  OAI211_X1 g383(.A(new_n582), .B(new_n579), .C1(new_n583), .C2(new_n584), .ZN(new_n585));
  AND3_X1   g384(.A1(new_n581), .A2(KEYINPUT94), .A3(new_n585), .ZN(new_n586));
  AOI21_X1  g385(.A(KEYINPUT94), .B1(new_n581), .B2(new_n585), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  NOR3_X1   g388(.A1(new_n512), .A2(new_n513), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(G232gat), .A2(G233gat), .ZN(new_n591));
  XOR2_X1   g390(.A(new_n591), .B(KEYINPUT101), .Z(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n593), .A2(KEYINPUT41), .ZN(new_n594));
  XNOR2_X1  g393(.A(G134gat), .B(G162gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n594), .B(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n596), .B(KEYINPUT103), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT102), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n598), .A2(G85gat), .A3(G92gat), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT7), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(G99gat), .A2(G106gat), .ZN(new_n602));
  INV_X1    g401(.A(G85gat), .ZN(new_n603));
  INV_X1    g402(.A(G92gat), .ZN(new_n604));
  AOI22_X1  g403(.A1(KEYINPUT8), .A2(new_n602), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND4_X1  g404(.A1(new_n598), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n601), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  XOR2_X1   g406(.A(G99gat), .B(G106gat), .Z(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n609), .A2(new_n539), .ZN(new_n610));
  OR2_X1    g409(.A1(new_n538), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n593), .A2(KEYINPUT41), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n538), .A2(new_n610), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n611), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  XOR2_X1   g413(.A(G190gat), .B(G218gat), .Z(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n615), .ZN(new_n617));
  NAND4_X1  g416(.A1(new_n611), .A2(new_n612), .A3(new_n613), .A4(new_n617), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n597), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  AND2_X1   g418(.A1(new_n596), .A2(KEYINPUT103), .ZN(new_n620));
  AND2_X1   g419(.A1(new_n616), .A2(new_n618), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n619), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(G183gat), .B(G211gat), .ZN(new_n623));
  XOR2_X1   g422(.A(G57gat), .B(G64gat), .Z(new_n624));
  NAND2_X1  g423(.A1(new_n624), .A2(KEYINPUT9), .ZN(new_n625));
  XOR2_X1   g424(.A(G71gat), .B(G78gat), .Z(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT98), .ZN(new_n628));
  INV_X1    g427(.A(G57gat), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n629), .A2(KEYINPUT95), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT95), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n631), .A2(G57gat), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n630), .A2(new_n632), .A3(G64gat), .ZN(new_n633));
  OR2_X1    g432(.A1(new_n629), .A2(G64gat), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT96), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n633), .A2(KEYINPUT96), .A3(new_n634), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  AOI21_X1  g438(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n640));
  OR2_X1    g439(.A1(new_n640), .A2(KEYINPUT97), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(KEYINPUT97), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n626), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n628), .B1(new_n639), .B2(new_n643), .ZN(new_n644));
  AND3_X1   g443(.A1(new_n633), .A2(KEYINPUT96), .A3(new_n634), .ZN(new_n645));
  AOI21_X1  g444(.A(KEYINPUT96), .B1(new_n633), .B2(new_n634), .ZN(new_n646));
  OAI211_X1 g445(.A(new_n643), .B(new_n628), .C1(new_n645), .C2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n627), .B1(new_n644), .B2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT21), .ZN(new_n650));
  NAND2_X1  g449(.A1(G231gat), .A2(G233gat), .ZN(new_n651));
  AND3_X1   g450(.A1(new_n649), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n651), .B1(new_n649), .B2(new_n650), .ZN(new_n653));
  OAI21_X1  g452(.A(G127gat), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  NOR3_X1   g454(.A1(new_n652), .A2(new_n653), .A3(G127gat), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n623), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n656), .ZN(new_n658));
  INV_X1    g457(.A(new_n623), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n658), .A2(new_n659), .A3(new_n654), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n627), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n643), .B1(new_n645), .B2(new_n646), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n663), .A2(KEYINPUT98), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n662), .B1(new_n664), .B2(new_n647), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n665), .A2(KEYINPUT21), .ZN(new_n666));
  XNOR2_X1  g465(.A(KEYINPUT99), .B(KEYINPUT100), .ZN(new_n667));
  AND3_X1   g466(.A1(new_n666), .A2(new_n564), .A3(new_n667), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n667), .B1(new_n564), .B2(new_n666), .ZN(new_n669));
  XNOR2_X1  g468(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(new_n328), .ZN(new_n671));
  OR3_X1    g470(.A1(new_n668), .A2(new_n669), .A3(new_n671), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n671), .B1(new_n668), .B2(new_n669), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n661), .A2(new_n674), .ZN(new_n675));
  NAND4_X1  g474(.A1(new_n657), .A2(new_n660), .A3(new_n672), .A4(new_n673), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n622), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  XNOR2_X1  g477(.A(G120gat), .B(G148gat), .ZN(new_n679));
  XNOR2_X1  g478(.A(G176gat), .B(G204gat), .ZN(new_n680));
  XOR2_X1   g479(.A(new_n679), .B(new_n680), .Z(new_n681));
  NAND2_X1  g480(.A1(new_n649), .A2(new_n609), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT10), .ZN(new_n683));
  INV_X1    g482(.A(new_n609), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n665), .A2(new_n684), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n682), .A2(new_n683), .A3(new_n685), .ZN(new_n686));
  AOI211_X1 g485(.A(new_n662), .B(new_n609), .C1(new_n664), .C2(new_n647), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(KEYINPUT10), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(G230gat), .A2(G233gat), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n665), .A2(new_n684), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n692), .A2(new_n687), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n690), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n681), .B1(new_n691), .B2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT104), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n698), .B1(new_n689), .B2(new_n690), .ZN(new_n699));
  AOI211_X1 g498(.A(KEYINPUT104), .B(new_n695), .C1(new_n686), .C2(new_n688), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(new_n681), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n702), .B1(new_n694), .B2(new_n695), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n697), .B1(new_n701), .B2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  NOR3_X1   g504(.A1(new_n678), .A2(KEYINPUT105), .A3(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT105), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n707), .B1(new_n677), .B2(new_n704), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n590), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n710), .A2(new_n495), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n711), .B(new_n545), .ZN(G1324gat));
  INV_X1    g511(.A(new_n710), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n493), .A2(new_n502), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n541), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(new_n714), .ZN(new_n716));
  XNOR2_X1  g515(.A(KEYINPUT16), .B(G8gat), .ZN(new_n717));
  NOR3_X1   g516(.A1(new_n710), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  OAI21_X1  g517(.A(KEYINPUT42), .B1(new_n715), .B2(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n719), .B1(new_n718), .B2(KEYINPUT42), .ZN(G1325gat));
  OR3_X1    g519(.A1(new_n710), .A2(G15gat), .A3(new_n506), .ZN(new_n721));
  AND3_X1   g520(.A1(new_n310), .A2(new_n311), .A3(KEYINPUT72), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n304), .A2(new_n309), .ZN(new_n723));
  OAI21_X1  g522(.A(KEYINPUT36), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  OR3_X1    g523(.A1(new_n305), .A2(new_n306), .A3(KEYINPUT36), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  OAI21_X1  g525(.A(G15gat), .B1(new_n710), .B2(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n721), .A2(new_n727), .ZN(G1326gat));
  AND3_X1   g527(.A1(new_n471), .A2(KEYINPUT81), .A3(new_n473), .ZN(new_n729));
  AOI21_X1  g528(.A(KEYINPUT81), .B1(new_n471), .B2(new_n473), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(new_n731), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n710), .A2(new_n732), .ZN(new_n733));
  XOR2_X1   g532(.A(KEYINPUT43), .B(G22gat), .Z(new_n734));
  XNOR2_X1  g533(.A(new_n733), .B(new_n734), .ZN(G1327gat));
  INV_X1    g534(.A(new_n622), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT44), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(new_n738), .ZN(new_n739));
  NOR3_X1   g538(.A1(new_n512), .A2(new_n513), .A3(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT107), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n498), .A2(new_n741), .ZN(new_n742));
  NAND4_X1  g541(.A1(new_n484), .A2(KEYINPUT107), .A3(new_n496), .A4(new_n497), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n742), .A2(new_n475), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(new_n510), .ZN(new_n745));
  AOI21_X1  g544(.A(KEYINPUT44), .B1(new_n745), .B2(new_n622), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n740), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n675), .A2(new_n676), .ZN(new_n748));
  INV_X1    g547(.A(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(new_n704), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n581), .A2(new_n585), .ZN(new_n751));
  INV_X1    g550(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n747), .A2(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(G29gat), .B1(new_n754), .B2(new_n495), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n750), .A2(new_n736), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n590), .A2(new_n756), .ZN(new_n757));
  OR2_X1    g556(.A1(new_n495), .A2(G29gat), .ZN(new_n758));
  OR3_X1    g557(.A1(new_n757), .A2(KEYINPUT106), .A3(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT45), .ZN(new_n760));
  OAI21_X1  g559(.A(KEYINPUT106), .B1(new_n757), .B2(new_n758), .ZN(new_n761));
  AND3_X1   g560(.A1(new_n759), .A2(new_n760), .A3(new_n761), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n760), .B1(new_n759), .B2(new_n761), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n755), .B1(new_n762), .B2(new_n763), .ZN(G1328gat));
  OAI21_X1  g563(.A(new_n523), .B1(new_n754), .B2(new_n716), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n716), .A2(new_n523), .ZN(new_n766));
  INV_X1    g565(.A(new_n766), .ZN(new_n767));
  OR3_X1    g566(.A1(new_n757), .A2(KEYINPUT46), .A3(new_n767), .ZN(new_n768));
  OAI21_X1  g567(.A(KEYINPUT46), .B1(new_n757), .B2(new_n767), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n765), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(KEYINPUT108), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT108), .ZN(new_n772));
  NAND4_X1  g571(.A1(new_n765), .A2(new_n768), .A3(new_n772), .A4(new_n769), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n771), .A2(new_n773), .ZN(G1329gat));
  NOR2_X1   g573(.A1(new_n757), .A2(new_n506), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n314), .A2(new_n531), .ZN(new_n776));
  OAI22_X1  g575(.A1(new_n775), .A2(new_n531), .B1(new_n754), .B2(new_n776), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n777), .B(KEYINPUT47), .ZN(G1330gat));
  NOR3_X1   g577(.A1(new_n757), .A2(new_n732), .A3(new_n534), .ZN(new_n779));
  NOR4_X1   g578(.A1(new_n740), .A2(new_n746), .A3(new_n752), .A4(new_n750), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(new_n731), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n779), .B1(new_n781), .B2(new_n534), .ZN(new_n782));
  INV_X1    g581(.A(new_n534), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n482), .A2(new_n483), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n783), .B1(new_n780), .B2(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT48), .ZN(new_n786));
  OR2_X1    g585(.A1(new_n779), .A2(new_n786), .ZN(new_n787));
  OAI22_X1  g586(.A1(new_n782), .A2(KEYINPUT48), .B1(new_n785), .B2(new_n787), .ZN(G1331gat));
  NAND4_X1  g587(.A1(new_n745), .A2(new_n752), .A3(new_n677), .A4(new_n705), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n789), .A2(new_n495), .ZN(new_n790));
  AND2_X1   g589(.A1(new_n630), .A2(new_n632), .ZN(new_n791));
  XNOR2_X1  g590(.A(new_n790), .B(new_n791), .ZN(G1332gat));
  NOR2_X1   g591(.A1(new_n789), .A2(new_n716), .ZN(new_n793));
  NOR2_X1   g592(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n794));
  AND2_X1   g593(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n793), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n796), .B1(new_n793), .B2(new_n794), .ZN(new_n797));
  XNOR2_X1  g596(.A(new_n797), .B(KEYINPUT109), .ZN(G1333gat));
  XOR2_X1   g597(.A(new_n506), .B(KEYINPUT110), .Z(new_n799));
  INV_X1    g598(.A(new_n799), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n789), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n314), .A2(G71gat), .ZN(new_n802));
  OAI22_X1  g601(.A1(new_n801), .A2(G71gat), .B1(new_n789), .B2(new_n802), .ZN(new_n803));
  XNOR2_X1  g602(.A(new_n803), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g603(.A1(new_n789), .A2(new_n732), .ZN(new_n805));
  XOR2_X1   g604(.A(new_n805), .B(G78gat), .Z(G1335gat));
  NOR3_X1   g605(.A1(new_n748), .A2(new_n751), .A3(new_n704), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n747), .A2(new_n807), .ZN(new_n808));
  OAI21_X1  g607(.A(G85gat), .B1(new_n808), .B2(new_n495), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n748), .A2(new_n751), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n745), .A2(new_n622), .A3(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT51), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND4_X1  g612(.A1(new_n745), .A2(KEYINPUT51), .A3(new_n622), .A4(new_n810), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n704), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(new_n495), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n815), .A2(new_n603), .A3(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n809), .A2(new_n817), .ZN(G1336gat));
  NOR2_X1   g617(.A1(new_n716), .A2(G92gat), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n815), .A2(new_n819), .ZN(new_n820));
  AND2_X1   g619(.A1(new_n474), .A2(new_n507), .ZN(new_n821));
  AND2_X1   g620(.A1(new_n505), .A2(new_n508), .ZN(new_n822));
  INV_X1    g621(.A(new_n496), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n823), .A2(new_n474), .A3(new_n313), .ZN(new_n824));
  AOI22_X1  g623(.A1(new_n821), .A2(new_n822), .B1(new_n824), .B2(KEYINPUT35), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n421), .A2(new_n439), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n726), .B1(new_n784), .B2(new_n826), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n827), .B1(new_n741), .B2(new_n498), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n825), .B1(new_n828), .B2(new_n743), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n737), .B1(new_n829), .B2(new_n736), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n827), .B1(new_n496), .B2(new_n731), .ZN(new_n831));
  OAI21_X1  g630(.A(KEYINPUT84), .B1(new_n831), .B2(new_n825), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n499), .A2(new_n510), .A3(new_n511), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n832), .A2(new_n833), .A3(new_n738), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n830), .A2(new_n834), .A3(new_n714), .A4(new_n807), .ZN(new_n835));
  AND2_X1   g634(.A1(new_n835), .A2(G92gat), .ZN(new_n836));
  OAI21_X1  g635(.A(KEYINPUT52), .B1(new_n820), .B2(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT112), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n604), .B1(new_n835), .B2(new_n838), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n747), .A2(KEYINPUT112), .A3(new_n714), .A4(new_n807), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  XNOR2_X1  g640(.A(KEYINPUT111), .B(KEYINPUT52), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n842), .B1(new_n815), .B2(new_n819), .ZN(new_n843));
  AND3_X1   g642(.A1(new_n841), .A2(KEYINPUT113), .A3(new_n843), .ZN(new_n844));
  AOI21_X1  g643(.A(KEYINPUT113), .B1(new_n841), .B2(new_n843), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n837), .B1(new_n844), .B2(new_n845), .ZN(G1337gat));
  INV_X1    g645(.A(G99gat), .ZN(new_n847));
  NOR3_X1   g646(.A1(new_n808), .A2(new_n847), .A3(new_n726), .ZN(new_n848));
  INV_X1    g647(.A(new_n506), .ZN(new_n849));
  AOI21_X1  g648(.A(G99gat), .B1(new_n815), .B2(new_n849), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n848), .A2(new_n850), .ZN(G1338gat));
  OAI21_X1  g650(.A(G106gat), .B1(new_n808), .B2(new_n732), .ZN(new_n852));
  INV_X1    g651(.A(G106gat), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n815), .A2(new_n853), .A3(new_n784), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT114), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n852), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(KEYINPUT53), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT53), .ZN(new_n858));
  OAI211_X1 g657(.A(new_n858), .B(G106gat), .C1(new_n808), .C2(new_n474), .ZN(new_n859));
  OAI211_X1 g658(.A(new_n859), .B(new_n854), .C1(new_n855), .C2(new_n858), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n857), .A2(new_n860), .ZN(G1339gat));
  INV_X1    g660(.A(KEYINPUT55), .ZN(new_n862));
  OAI21_X1  g661(.A(KEYINPUT54), .B1(new_n689), .B2(new_n690), .ZN(new_n863));
  NOR3_X1   g662(.A1(new_n863), .A2(new_n699), .A3(new_n700), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n702), .B1(new_n691), .B2(KEYINPUT54), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n862), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n701), .A2(new_n703), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n691), .A2(KEYINPUT104), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT54), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n685), .A2(new_n683), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n870), .B1(new_n693), .B2(new_n683), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n869), .B1(new_n871), .B2(new_n695), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n689), .A2(new_n698), .A3(new_n690), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n868), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n871), .A2(new_n695), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n681), .B1(new_n875), .B2(new_n869), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n874), .A2(new_n876), .A3(KEYINPUT55), .ZN(new_n877));
  NAND4_X1  g676(.A1(new_n866), .A2(new_n751), .A3(new_n867), .A4(new_n877), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n570), .A2(new_n514), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n566), .B1(new_n563), .B2(new_n565), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n578), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n568), .A2(new_n573), .A3(new_n580), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n705), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT116), .ZN(new_n884));
  AND3_X1   g683(.A1(new_n878), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n884), .B1(new_n878), .B2(new_n883), .ZN(new_n886));
  NOR3_X1   g685(.A1(new_n885), .A2(new_n886), .A3(new_n622), .ZN(new_n887));
  AND2_X1   g686(.A1(new_n877), .A2(new_n867), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n882), .A2(new_n881), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n889), .A2(new_n736), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n888), .A2(new_n866), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(KEYINPUT115), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT115), .ZN(new_n893));
  NAND4_X1  g692(.A1(new_n888), .A2(new_n890), .A3(new_n893), .A4(new_n866), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n749), .B1(new_n887), .B2(new_n895), .ZN(new_n896));
  NOR3_X1   g695(.A1(new_n678), .A2(new_n751), .A3(new_n705), .ZN(new_n897));
  INV_X1    g696(.A(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n714), .A2(new_n495), .ZN(new_n900));
  AND2_X1   g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  INV_X1    g700(.A(new_n500), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(new_n903), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n904), .A2(new_n265), .A3(new_n751), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n731), .B1(new_n896), .B2(new_n898), .ZN(new_n906));
  NOR3_X1   g705(.A1(new_n714), .A2(new_n506), .A3(new_n495), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n906), .A2(new_n588), .A3(new_n907), .ZN(new_n908));
  AND3_X1   g707(.A1(new_n908), .A2(KEYINPUT117), .A3(G113gat), .ZN(new_n909));
  AOI21_X1  g708(.A(KEYINPUT117), .B1(new_n908), .B2(G113gat), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n905), .B1(new_n909), .B2(new_n910), .ZN(G1340gat));
  NAND2_X1  g710(.A1(new_n906), .A2(new_n907), .ZN(new_n912));
  NOR3_X1   g711(.A1(new_n912), .A2(new_n254), .A3(new_n704), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n904), .A2(new_n705), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n913), .B1(new_n914), .B2(new_n254), .ZN(G1341gat));
  NOR3_X1   g714(.A1(new_n912), .A2(new_n260), .A3(new_n749), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n903), .A2(new_n749), .ZN(new_n917));
  OR2_X1    g716(.A1(new_n917), .A2(KEYINPUT118), .ZN(new_n918));
  AOI21_X1  g717(.A(G127gat), .B1(new_n917), .B2(KEYINPUT118), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n916), .B1(new_n918), .B2(new_n919), .ZN(G1342gat));
  NAND4_X1  g719(.A1(new_n901), .A2(new_n261), .A3(new_n902), .A4(new_n622), .ZN(new_n921));
  OR2_X1    g720(.A1(new_n921), .A2(KEYINPUT56), .ZN(new_n922));
  OAI21_X1  g721(.A(G134gat), .B1(new_n912), .B2(new_n736), .ZN(new_n923));
  AND3_X1   g722(.A1(new_n921), .A2(KEYINPUT119), .A3(KEYINPUT56), .ZN(new_n924));
  AOI21_X1  g723(.A(KEYINPUT119), .B1(new_n921), .B2(KEYINPUT56), .ZN(new_n925));
  OAI211_X1 g724(.A(new_n922), .B(new_n923), .C1(new_n924), .C2(new_n925), .ZN(G1343gat));
  AND2_X1   g725(.A1(new_n892), .A2(new_n894), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n889), .A2(new_n704), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n877), .A2(new_n867), .ZN(new_n929));
  XNOR2_X1  g728(.A(KEYINPUT120), .B(KEYINPUT55), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n930), .B1(new_n874), .B2(new_n876), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n928), .B1(new_n588), .B2(new_n932), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n927), .B1(new_n622), .B2(new_n933), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n897), .B1(new_n934), .B2(new_n749), .ZN(new_n935));
  OAI21_X1  g734(.A(KEYINPUT57), .B1(new_n935), .B2(new_n732), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT57), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n899), .A2(new_n937), .A3(new_n784), .ZN(new_n938));
  AND2_X1   g737(.A1(new_n726), .A2(new_n900), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n936), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  OAI21_X1  g739(.A(G141gat), .B1(new_n940), .B2(new_n589), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT58), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n314), .A2(new_n474), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n589), .A2(G141gat), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n901), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n941), .A2(new_n942), .A3(new_n945), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n901), .A2(new_n943), .ZN(new_n947));
  INV_X1    g746(.A(new_n947), .ZN(new_n948));
  NAND4_X1  g747(.A1(new_n936), .A2(new_n751), .A3(new_n938), .A4(new_n939), .ZN(new_n949));
  AOI22_X1  g748(.A1(new_n948), .A2(new_n944), .B1(new_n949), .B2(G141gat), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n946), .B1(new_n942), .B2(new_n950), .ZN(G1344gat));
  INV_X1    g750(.A(KEYINPUT59), .ZN(new_n952));
  OAI211_X1 g751(.A(new_n952), .B(G148gat), .C1(new_n940), .C2(new_n704), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT121), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n878), .A2(new_n883), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n955), .A2(KEYINPUT116), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n878), .A2(new_n883), .A3(new_n884), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n956), .A2(new_n736), .A3(new_n957), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n748), .B1(new_n927), .B2(new_n958), .ZN(new_n959));
  NOR2_X1   g758(.A1(new_n959), .A2(new_n897), .ZN(new_n960));
  NOR2_X1   g759(.A1(new_n474), .A2(new_n937), .ZN(new_n961));
  INV_X1    g760(.A(new_n961), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n954), .B1(new_n960), .B2(new_n962), .ZN(new_n963));
  OAI211_X1 g762(.A(KEYINPUT121), .B(new_n961), .C1(new_n959), .C2(new_n897), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n891), .B1(new_n933), .B2(new_n622), .ZN(new_n965));
  AOI22_X1  g764(.A1(new_n965), .A2(new_n749), .B1(new_n709), .B2(new_n589), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n937), .B1(new_n966), .B2(new_n732), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n963), .A2(new_n964), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n939), .A2(new_n705), .ZN(new_n969));
  INV_X1    g768(.A(new_n969), .ZN(new_n970));
  AOI21_X1  g769(.A(new_n324), .B1(new_n968), .B2(new_n970), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n953), .B1(new_n971), .B2(new_n952), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n948), .A2(new_n324), .A3(new_n705), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n972), .A2(new_n973), .ZN(G1345gat));
  NAND3_X1  g773(.A1(new_n948), .A2(new_n328), .A3(new_n748), .ZN(new_n975));
  OAI21_X1  g774(.A(G155gat), .B1(new_n940), .B2(new_n749), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n975), .A2(new_n976), .ZN(G1346gat));
  AOI21_X1  g776(.A(G162gat), .B1(new_n948), .B2(new_n622), .ZN(new_n978));
  NOR3_X1   g777(.A1(new_n940), .A2(new_n329), .A3(new_n736), .ZN(new_n979));
  NOR2_X1   g778(.A1(new_n978), .A2(new_n979), .ZN(G1347gat));
  NOR2_X1   g779(.A1(new_n716), .A2(new_n816), .ZN(new_n981));
  INV_X1    g780(.A(new_n981), .ZN(new_n982));
  NOR2_X1   g781(.A1(new_n800), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n906), .A2(new_n983), .ZN(new_n984));
  OAI21_X1  g783(.A(G169gat), .B1(new_n984), .B2(new_n589), .ZN(new_n985));
  AND2_X1   g784(.A1(new_n985), .A2(KEYINPUT122), .ZN(new_n986));
  NOR2_X1   g785(.A1(new_n985), .A2(KEYINPUT122), .ZN(new_n987));
  NOR2_X1   g786(.A1(new_n960), .A2(new_n982), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n988), .A2(new_n902), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n751), .A2(new_n231), .A3(new_n232), .ZN(new_n990));
  OAI22_X1  g789(.A1(new_n986), .A2(new_n987), .B1(new_n989), .B2(new_n990), .ZN(G1348gat));
  OAI21_X1  g790(.A(G176gat), .B1(new_n984), .B2(new_n704), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n705), .A2(new_n203), .ZN(new_n993));
  OAI21_X1  g792(.A(new_n992), .B1(new_n989), .B2(new_n993), .ZN(G1349gat));
  NAND3_X1  g793(.A1(new_n906), .A2(new_n748), .A3(new_n983), .ZN(new_n995));
  INV_X1    g794(.A(KEYINPUT123), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND4_X1  g796(.A1(new_n906), .A2(KEYINPUT123), .A3(new_n748), .A4(new_n983), .ZN(new_n998));
  NAND3_X1  g797(.A1(new_n997), .A2(G183gat), .A3(new_n998), .ZN(new_n999));
  AND2_X1   g798(.A1(new_n748), .A2(new_n216), .ZN(new_n1000));
  NAND4_X1  g799(.A1(new_n899), .A2(new_n902), .A3(new_n981), .A4(new_n1000), .ZN(new_n1001));
  AND2_X1   g800(.A1(new_n1001), .A2(KEYINPUT124), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n999), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n1003), .A2(KEYINPUT60), .ZN(new_n1004));
  INV_X1    g803(.A(KEYINPUT60), .ZN(new_n1005));
  NAND3_X1  g804(.A1(new_n999), .A2(new_n1005), .A3(new_n1002), .ZN(new_n1006));
  NAND2_X1  g805(.A1(new_n1004), .A2(new_n1006), .ZN(G1350gat));
  NAND4_X1  g806(.A1(new_n988), .A2(new_n207), .A3(new_n902), .A4(new_n622), .ZN(new_n1008));
  INV_X1    g807(.A(KEYINPUT125), .ZN(new_n1009));
  XNOR2_X1  g808(.A(new_n1008), .B(new_n1009), .ZN(new_n1010));
  NAND3_X1  g809(.A1(new_n906), .A2(new_n622), .A3(new_n983), .ZN(new_n1011));
  AND2_X1   g810(.A1(new_n1011), .A2(G190gat), .ZN(new_n1012));
  NAND2_X1  g811(.A1(new_n1012), .A2(KEYINPUT61), .ZN(new_n1013));
  OR2_X1    g812(.A1(new_n1012), .A2(KEYINPUT61), .ZN(new_n1014));
  NAND3_X1  g813(.A1(new_n1010), .A2(new_n1013), .A3(new_n1014), .ZN(G1351gat));
  NAND3_X1  g814(.A1(new_n899), .A2(new_n943), .A3(new_n981), .ZN(new_n1016));
  INV_X1    g815(.A(new_n1016), .ZN(new_n1017));
  AOI21_X1  g816(.A(G197gat), .B1(new_n1017), .B2(new_n751), .ZN(new_n1018));
  NOR2_X1   g817(.A1(new_n982), .A2(new_n314), .ZN(new_n1019));
  AND2_X1   g818(.A1(new_n968), .A2(new_n1019), .ZN(new_n1020));
  AND2_X1   g819(.A1(new_n588), .A2(G197gat), .ZN(new_n1021));
  AOI21_X1  g820(.A(new_n1018), .B1(new_n1020), .B2(new_n1021), .ZN(G1352gat));
  INV_X1    g821(.A(KEYINPUT62), .ZN(new_n1023));
  NOR2_X1   g822(.A1(new_n704), .A2(G204gat), .ZN(new_n1024));
  INV_X1    g823(.A(new_n1024), .ZN(new_n1025));
  OAI21_X1  g824(.A(KEYINPUT126), .B1(new_n1016), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g825(.A(new_n1026), .ZN(new_n1027));
  NOR3_X1   g826(.A1(new_n1016), .A2(KEYINPUT126), .A3(new_n1025), .ZN(new_n1028));
  OAI21_X1  g827(.A(new_n1023), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g828(.A(new_n1028), .ZN(new_n1030));
  NAND3_X1  g829(.A1(new_n1030), .A2(KEYINPUT62), .A3(new_n1026), .ZN(new_n1031));
  AND3_X1   g830(.A1(new_n968), .A2(new_n705), .A3(new_n1019), .ZN(new_n1032));
  INV_X1    g831(.A(G204gat), .ZN(new_n1033));
  OAI211_X1 g832(.A(new_n1029), .B(new_n1031), .C1(new_n1032), .C2(new_n1033), .ZN(G1353gat));
  OR3_X1    g833(.A1(new_n1016), .A2(G211gat), .A3(new_n749), .ZN(new_n1035));
  AOI21_X1  g834(.A(new_n962), .B1(new_n896), .B2(new_n898), .ZN(new_n1036));
  OAI21_X1  g835(.A(new_n967), .B1(new_n1036), .B2(KEYINPUT121), .ZN(new_n1037));
  INV_X1    g836(.A(new_n964), .ZN(new_n1038));
  OAI211_X1 g837(.A(new_n748), .B(new_n1019), .C1(new_n1037), .C2(new_n1038), .ZN(new_n1039));
  AND3_X1   g838(.A1(new_n1039), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1040));
  AOI21_X1  g839(.A(KEYINPUT63), .B1(new_n1039), .B2(G211gat), .ZN(new_n1041));
  OAI21_X1  g840(.A(new_n1035), .B1(new_n1040), .B2(new_n1041), .ZN(G1354gat));
  INV_X1    g841(.A(G218gat), .ZN(new_n1043));
  OAI21_X1  g842(.A(new_n1043), .B1(new_n1016), .B2(new_n736), .ZN(new_n1044));
  XNOR2_X1  g843(.A(new_n1044), .B(KEYINPUT127), .ZN(new_n1045));
  NOR2_X1   g844(.A1(new_n736), .A2(new_n1043), .ZN(new_n1046));
  AOI21_X1  g845(.A(new_n1045), .B1(new_n1020), .B2(new_n1046), .ZN(G1355gat));
endmodule


