//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 0 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1 0 1 0 0 1 1 1 0 0 0 0 0 0 0 1 0 0 1 1 1 1 1 0 1 0 0 1 1 1 1 0 1 0 0 1 0 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:51 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n704, new_n705, new_n706,
    new_n707, new_n709, new_n710, new_n711, new_n713, new_n714, new_n715,
    new_n716, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n763, new_n764, new_n765, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n798, new_n799, new_n800, new_n801, new_n803, new_n804, new_n805,
    new_n806, new_n808, new_n809, new_n810, new_n811, new_n813, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n840, new_n841, new_n842, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n906, new_n907, new_n909, new_n910, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n972,
    new_n973, new_n975, new_n976, new_n977, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n989,
    new_n990, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1039, new_n1040, new_n1041, new_n1042, new_n1044,
    new_n1045;
  INV_X1    g000(.A(KEYINPUT94), .ZN(new_n202));
  INV_X1    g001(.A(G29gat), .ZN(new_n203));
  INV_X1    g002(.A(G36gat), .ZN(new_n204));
  NAND3_X1  g003(.A1(new_n203), .A2(new_n204), .A3(KEYINPUT14), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT14), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n206), .B1(G29gat), .B2(G36gat), .ZN(new_n207));
  OAI211_X1 g006(.A(new_n205), .B(new_n207), .C1(new_n203), .C2(new_n204), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT15), .ZN(new_n209));
  OR2_X1    g008(.A1(G43gat), .A2(G50gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(G43gat), .A2(G50gat), .ZN(new_n211));
  AOI21_X1  g010(.A(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n208), .A2(new_n212), .ZN(new_n213));
  AOI21_X1  g012(.A(KEYINPUT15), .B1(G43gat), .B2(G50gat), .ZN(new_n214));
  XOR2_X1   g013(.A(KEYINPUT88), .B(G50gat), .Z(new_n215));
  OAI21_X1  g014(.A(new_n214), .B1(new_n215), .B2(G43gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n213), .A2(new_n216), .ZN(new_n217));
  AOI21_X1  g016(.A(KEYINPUT87), .B1(new_n208), .B2(new_n212), .ZN(new_n218));
  AND3_X1   g017(.A1(new_n208), .A2(KEYINPUT87), .A3(new_n212), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n217), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT89), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT17), .ZN(new_n223));
  OAI211_X1 g022(.A(new_n217), .B(KEYINPUT89), .C1(new_n218), .C2(new_n219), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  XOR2_X1   g024(.A(G15gat), .B(G22gat), .Z(new_n226));
  INV_X1    g025(.A(G1gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  XNOR2_X1  g027(.A(G15gat), .B(G22gat), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT16), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n229), .B1(new_n230), .B2(G1gat), .ZN(new_n231));
  INV_X1    g030(.A(G8gat), .ZN(new_n232));
  OR2_X1    g031(.A1(new_n232), .A2(KEYINPUT90), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n228), .A2(new_n231), .A3(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n234), .A2(KEYINPUT90), .A3(new_n232), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n232), .A2(KEYINPUT90), .ZN(new_n236));
  NAND4_X1  g035(.A1(new_n228), .A2(new_n231), .A3(new_n236), .A4(new_n233), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  OAI211_X1 g037(.A(new_n217), .B(KEYINPUT17), .C1(new_n218), .C2(new_n219), .ZN(new_n239));
  AND2_X1   g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n225), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT91), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(G229gat), .A2(G233gat), .ZN(new_n244));
  INV_X1    g043(.A(new_n238), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n245), .A2(new_n222), .A3(new_n224), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n225), .A2(KEYINPUT91), .A3(new_n240), .ZN(new_n247));
  NAND4_X1  g046(.A1(new_n243), .A2(new_n244), .A3(new_n246), .A4(new_n247), .ZN(new_n248));
  XOR2_X1   g047(.A(KEYINPUT92), .B(KEYINPUT18), .Z(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  AND2_X1   g050(.A1(new_n247), .A2(new_n246), .ZN(new_n252));
  NAND4_X1  g051(.A1(new_n252), .A2(KEYINPUT18), .A3(new_n244), .A4(new_n243), .ZN(new_n253));
  XNOR2_X1  g052(.A(G113gat), .B(G141gat), .ZN(new_n254));
  XNOR2_X1  g053(.A(KEYINPUT85), .B(KEYINPUT11), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n254), .B(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(G169gat), .B(G197gat), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n256), .B(new_n257), .ZN(new_n258));
  XOR2_X1   g057(.A(KEYINPUT86), .B(KEYINPUT12), .Z(new_n259));
  XOR2_X1   g058(.A(new_n258), .B(new_n259), .Z(new_n260));
  XOR2_X1   g059(.A(new_n244), .B(KEYINPUT13), .Z(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n222), .A2(new_n224), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(new_n238), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n262), .B1(new_n264), .B2(new_n246), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  NAND4_X1  g065(.A1(new_n251), .A2(new_n253), .A3(new_n260), .A4(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT93), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n247), .A2(new_n246), .ZN(new_n270));
  INV_X1    g069(.A(new_n244), .ZN(new_n271));
  AOI21_X1  g070(.A(KEYINPUT91), .B1(new_n225), .B2(new_n240), .ZN(new_n272));
  NOR3_X1   g071(.A1(new_n270), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n265), .B1(new_n273), .B2(KEYINPUT18), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n260), .B1(new_n274), .B2(new_n251), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n269), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n251), .A2(new_n253), .A3(new_n266), .ZN(new_n277));
  INV_X1    g076(.A(new_n260), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n277), .A2(KEYINPUT93), .A3(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n202), .B1(new_n276), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n277), .A2(new_n278), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n282), .A2(new_n268), .A3(new_n267), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n283), .A2(KEYINPUT94), .A3(new_n279), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n281), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(G183gat), .A2(G190gat), .ZN(new_n286));
  INV_X1    g085(.A(G169gat), .ZN(new_n287));
  INV_X1    g086(.A(G176gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(KEYINPUT26), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT68), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n290), .B(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(G169gat), .A2(G176gat), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT69), .ZN(new_n294));
  OAI211_X1 g093(.A(new_n287), .B(new_n288), .C1(new_n294), .C2(KEYINPUT26), .ZN(new_n295));
  AND2_X1   g094(.A1(new_n294), .A2(KEYINPUT26), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n293), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n286), .B1(new_n292), .B2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(G183gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(KEYINPUT27), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT27), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(G183gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT28), .ZN(new_n304));
  NOR3_X1   g103(.A1(new_n303), .A2(new_n304), .A3(G190gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n303), .A2(KEYINPUT67), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT67), .ZN(new_n307));
  AOI21_X1  g106(.A(G190gat), .B1(new_n300), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n305), .B1(new_n309), .B2(new_n304), .ZN(new_n310));
  OR2_X1    g109(.A1(new_n298), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT25), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n286), .A2(KEYINPUT24), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  XNOR2_X1  g113(.A(G183gat), .B(G190gat), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT24), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n314), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT23), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n318), .A2(G169gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n288), .A2(KEYINPUT64), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT64), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(G176gat), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n319), .A2(new_n320), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n293), .A2(KEYINPUT23), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(new_n289), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n312), .B1(new_n317), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(KEYINPUT65), .ZN(new_n328));
  INV_X1    g127(.A(G190gat), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n329), .A2(G183gat), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n299), .A2(G190gat), .ZN(new_n331));
  OAI21_X1  g130(.A(KEYINPUT24), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND4_X1  g131(.A1(new_n332), .A2(new_n314), .A3(new_n323), .A4(new_n325), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT65), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n333), .A2(new_n334), .A3(new_n312), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n328), .A2(new_n335), .ZN(new_n336));
  OAI211_X1 g135(.A(new_n325), .B(KEYINPUT25), .C1(new_n318), .C2(new_n289), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n337), .A2(new_n317), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  AOI21_X1  g138(.A(KEYINPUT66), .B1(new_n336), .B2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT66), .ZN(new_n341));
  AOI211_X1 g140(.A(new_n341), .B(new_n338), .C1(new_n328), .C2(new_n335), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n311), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT70), .ZN(new_n344));
  INV_X1    g143(.A(G113gat), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n344), .B1(new_n345), .B2(G120gat), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(G120gat), .ZN(new_n347));
  INV_X1    g146(.A(G120gat), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n348), .A2(KEYINPUT70), .A3(G113gat), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n346), .A2(new_n347), .A3(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  XNOR2_X1  g150(.A(G127gat), .B(G134gat), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT1), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  OAI21_X1  g153(.A(KEYINPUT71), .B1(new_n351), .B2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT71), .ZN(new_n356));
  NAND4_X1  g155(.A1(new_n350), .A2(new_n356), .A3(new_n353), .A4(new_n352), .ZN(new_n357));
  INV_X1    g156(.A(new_n352), .ZN(new_n358));
  INV_X1    g157(.A(new_n347), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n345), .A2(G120gat), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n353), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  AOI22_X1  g160(.A1(new_n355), .A2(new_n357), .B1(new_n358), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n343), .A2(new_n362), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n298), .A2(new_n310), .ZN(new_n364));
  XNOR2_X1  g163(.A(KEYINPUT64), .B(G176gat), .ZN(new_n365));
  AOI22_X1  g164(.A1(new_n365), .A2(new_n319), .B1(new_n289), .B2(new_n324), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n299), .A2(G190gat), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n329), .A2(G183gat), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n313), .B1(new_n369), .B2(KEYINPUT24), .ZN(new_n370));
  AOI211_X1 g169(.A(KEYINPUT65), .B(KEYINPUT25), .C1(new_n366), .C2(new_n370), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n334), .B1(new_n333), .B2(new_n312), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n339), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(new_n341), .ZN(new_n374));
  OAI211_X1 g173(.A(KEYINPUT66), .B(new_n339), .C1(new_n371), .C2(new_n372), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n364), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(new_n362), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(G227gat), .A2(G233gat), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n363), .A2(new_n378), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(KEYINPUT32), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT33), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  XOR2_X1   g183(.A(G15gat), .B(G43gat), .Z(new_n385));
  XNOR2_X1  g184(.A(G71gat), .B(G99gat), .ZN(new_n386));
  XNOR2_X1  g185(.A(new_n385), .B(new_n386), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n382), .A2(new_n384), .A3(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(new_n387), .ZN(new_n389));
  OAI211_X1 g188(.A(new_n381), .B(KEYINPUT32), .C1(new_n383), .C2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT74), .ZN(new_n392));
  NAND2_X1  g191(.A1(KEYINPUT73), .A2(KEYINPUT34), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n374), .A2(new_n375), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n377), .B1(new_n394), .B2(new_n311), .ZN(new_n395));
  AOI211_X1 g194(.A(new_n362), .B(new_n364), .C1(new_n374), .C2(new_n375), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n393), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n363), .A2(new_n378), .A3(KEYINPUT73), .ZN(new_n398));
  AND3_X1   g197(.A1(new_n397), .A2(new_n398), .A3(new_n379), .ZN(new_n399));
  NAND2_X1  g198(.A1(KEYINPUT72), .A2(KEYINPUT34), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n380), .B1(new_n363), .B2(new_n378), .ZN(new_n401));
  NOR2_X1   g200(.A1(KEYINPUT72), .A2(KEYINPUT34), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n400), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n392), .B1(new_n399), .B2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(new_n400), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n379), .B1(new_n395), .B2(new_n396), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n406), .B1(new_n407), .B2(new_n402), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n397), .A2(new_n398), .A3(new_n379), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n408), .A2(KEYINPUT74), .A3(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n391), .B1(new_n405), .B2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(G22gat), .ZN(new_n412));
  XNOR2_X1  g211(.A(G197gat), .B(G204gat), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT22), .ZN(new_n414));
  INV_X1    g213(.A(G211gat), .ZN(new_n415));
  INV_X1    g214(.A(G218gat), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n414), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n413), .A2(new_n417), .ZN(new_n418));
  XNOR2_X1  g217(.A(G211gat), .B(G218gat), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n419), .A2(new_n413), .A3(new_n417), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT29), .ZN(new_n424));
  AOI21_X1  g223(.A(KEYINPUT3), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  XNOR2_X1  g224(.A(G155gat), .B(G162gat), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(G155gat), .ZN(new_n428));
  INV_X1    g227(.A(G162gat), .ZN(new_n429));
  OAI21_X1  g228(.A(KEYINPUT2), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  XNOR2_X1  g229(.A(G141gat), .B(G148gat), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n430), .B1(new_n431), .B2(KEYINPUT77), .ZN(new_n432));
  INV_X1    g231(.A(G148gat), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(G141gat), .ZN(new_n434));
  INV_X1    g233(.A(G141gat), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(G148gat), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT77), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n427), .B1(new_n432), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(KEYINPUT78), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n437), .A2(new_n438), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n431), .A2(KEYINPUT77), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n442), .A2(new_n443), .A3(new_n430), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT78), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n444), .A2(new_n445), .A3(new_n427), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n441), .A2(new_n446), .ZN(new_n447));
  XNOR2_X1  g246(.A(KEYINPUT79), .B(G141gat), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(G148gat), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(new_n434), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT2), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n451), .B1(G155gat), .B2(G162gat), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n427), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n450), .A2(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n425), .B1(new_n447), .B2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT3), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n452), .B1(new_n437), .B2(new_n438), .ZN(new_n457));
  AOI211_X1 g256(.A(KEYINPUT78), .B(new_n426), .C1(new_n457), .C2(new_n443), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n445), .B1(new_n444), .B2(new_n427), .ZN(new_n459));
  OAI211_X1 g258(.A(new_n456), .B(new_n454), .C1(new_n458), .C2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(new_n424), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT76), .ZN(new_n462));
  XNOR2_X1  g261(.A(new_n423), .B(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n455), .B1(new_n461), .B2(new_n464), .ZN(new_n465));
  AOI22_X1  g264(.A1(new_n441), .A2(new_n446), .B1(new_n450), .B2(new_n453), .ZN(new_n466));
  OAI21_X1  g265(.A(KEYINPUT81), .B1(new_n466), .B2(new_n425), .ZN(new_n467));
  NAND2_X1  g266(.A1(G228gat), .A2(G233gat), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n465), .A2(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n463), .B1(new_n460), .B2(new_n424), .ZN(new_n471));
  OAI211_X1 g270(.A(new_n468), .B(new_n467), .C1(new_n471), .C2(new_n455), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT82), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  XNOR2_X1  g274(.A(G78gat), .B(G106gat), .ZN(new_n476));
  XNOR2_X1  g275(.A(KEYINPUT31), .B(G50gat), .ZN(new_n477));
  XOR2_X1   g276(.A(new_n476), .B(new_n477), .Z(new_n478));
  AOI21_X1  g277(.A(new_n412), .B1(new_n475), .B2(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(KEYINPUT82), .B1(new_n470), .B2(new_n472), .ZN(new_n480));
  INV_X1    g279(.A(new_n478), .ZN(new_n481));
  NOR3_X1   g280(.A1(new_n480), .A2(G22gat), .A3(new_n481), .ZN(new_n482));
  OAI22_X1  g281(.A1(new_n479), .A2(new_n482), .B1(new_n474), .B2(new_n473), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n475), .A2(new_n412), .A3(new_n478), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n473), .A2(new_n474), .ZN(new_n485));
  OAI21_X1  g284(.A(G22gat), .B1(new_n480), .B2(new_n481), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n484), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n483), .A2(new_n487), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n411), .A2(new_n488), .ZN(new_n489));
  AND3_X1   g288(.A1(new_n408), .A2(KEYINPUT74), .A3(new_n409), .ZN(new_n490));
  AOI21_X1  g289(.A(KEYINPUT74), .B1(new_n408), .B2(new_n409), .ZN(new_n491));
  OAI21_X1  g290(.A(KEYINPUT75), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT75), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n405), .A2(new_n493), .A3(new_n410), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n492), .A2(new_n391), .A3(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT5), .ZN(new_n496));
  NAND2_X1  g295(.A1(G225gat), .A2(G233gat), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n454), .B1(new_n458), .B2(new_n459), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(new_n377), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n447), .A2(new_n454), .A3(new_n362), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n497), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT80), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n496), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n498), .A2(KEYINPUT3), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n504), .A2(new_n460), .A3(new_n377), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT4), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n500), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n466), .A2(KEYINPUT4), .A3(new_n362), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n505), .A2(new_n497), .A3(new_n507), .A4(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(new_n497), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n498), .A2(new_n377), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n362), .B1(new_n447), .B2(new_n454), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(KEYINPUT80), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n503), .A2(new_n509), .A3(new_n514), .ZN(new_n515));
  AND2_X1   g314(.A1(new_n507), .A2(new_n508), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n516), .A2(new_n496), .A3(new_n497), .A4(new_n505), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  XNOR2_X1  g317(.A(G1gat), .B(G29gat), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n519), .B(KEYINPUT0), .ZN(new_n520));
  XNOR2_X1  g319(.A(G57gat), .B(G85gat), .ZN(new_n521));
  XOR2_X1   g320(.A(new_n520), .B(new_n521), .Z(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n518), .A2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT6), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n515), .A2(new_n522), .A3(new_n517), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n524), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n518), .A2(KEYINPUT6), .A3(new_n523), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(G8gat), .B(G36gat), .ZN(new_n530));
  XNOR2_X1  g329(.A(G64gat), .B(G92gat), .ZN(new_n531));
  XOR2_X1   g330(.A(new_n530), .B(new_n531), .Z(new_n532));
  INV_X1    g331(.A(new_n532), .ZN(new_n533));
  AND2_X1   g332(.A1(G226gat), .A2(G233gat), .ZN(new_n534));
  AND3_X1   g333(.A1(new_n311), .A2(new_n373), .A3(new_n534), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n534), .A2(KEYINPUT29), .ZN(new_n536));
  AOI211_X1 g335(.A(new_n463), .B(new_n535), .C1(new_n343), .C2(new_n536), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n394), .A2(new_n311), .A3(new_n534), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n338), .B1(new_n328), .B2(new_n335), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n536), .B1(new_n539), .B2(new_n364), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n464), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n533), .B1(new_n537), .B2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(new_n535), .ZN(new_n543));
  INV_X1    g342(.A(new_n536), .ZN(new_n544));
  OAI211_X1 g343(.A(new_n543), .B(new_n464), .C1(new_n376), .C2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(new_n540), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n546), .B1(new_n376), .B2(new_n534), .ZN(new_n547));
  OAI211_X1 g346(.A(new_n545), .B(new_n532), .C1(new_n547), .C2(new_n464), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n542), .A2(KEYINPUT30), .A3(new_n548), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n537), .A2(new_n541), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT30), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n550), .A2(new_n551), .A3(new_n532), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  AND2_X1   g352(.A1(new_n529), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n489), .A2(new_n495), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n555), .A2(KEYINPUT35), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n405), .A2(new_n410), .ZN(new_n557));
  INV_X1    g356(.A(new_n391), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n405), .A2(new_n391), .A3(new_n410), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n528), .A2(KEYINPUT84), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n522), .B1(new_n515), .B2(new_n517), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT84), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n564), .A2(new_n565), .A3(KEYINPUT6), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n564), .A2(KEYINPUT6), .ZN(new_n567));
  AOI22_X1  g366(.A1(new_n563), .A2(new_n566), .B1(new_n567), .B2(new_n526), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT35), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n569), .ZN(new_n570));
  NOR3_X1   g369(.A1(new_n568), .A2(new_n488), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n562), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n572), .ZN(new_n573));
  AND3_X1   g372(.A1(new_n484), .A2(new_n485), .A3(new_n486), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n485), .B1(new_n484), .B2(new_n486), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT83), .ZN(new_n576));
  NOR3_X1   g375(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  AOI21_X1  g376(.A(KEYINPUT83), .B1(new_n483), .B2(new_n487), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n529), .A2(new_n553), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT40), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n377), .B1(new_n466), .B2(new_n456), .ZN(new_n582));
  INV_X1    g381(.A(new_n460), .ZN(new_n583));
  OAI211_X1 g382(.A(new_n507), .B(new_n508), .C1(new_n582), .C2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT39), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n584), .A2(new_n585), .A3(new_n510), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n586), .A2(new_n522), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n499), .A2(new_n500), .A3(new_n497), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n588), .A2(KEYINPUT39), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n589), .B1(new_n584), .B2(new_n510), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n581), .B1(new_n587), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n584), .A2(new_n510), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n592), .A2(KEYINPUT39), .A3(new_n588), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n593), .A2(KEYINPUT40), .A3(new_n522), .A4(new_n586), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n524), .A2(new_n591), .A3(new_n594), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n553), .A2(new_n595), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n596), .A2(new_n488), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n563), .A2(new_n566), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT37), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n532), .B1(new_n550), .B2(new_n599), .ZN(new_n600));
  OR2_X1    g399(.A1(new_n547), .A2(new_n463), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n535), .B1(new_n343), .B2(new_n536), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n599), .B1(new_n602), .B2(new_n463), .ZN(new_n603));
  AOI21_X1  g402(.A(KEYINPUT38), .B1(new_n601), .B2(new_n603), .ZN(new_n604));
  AOI22_X1  g403(.A1(new_n600), .A2(new_n604), .B1(new_n550), .B2(new_n532), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n550), .A2(new_n599), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n545), .B1(new_n547), .B2(new_n464), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n533), .B1(new_n607), .B2(KEYINPUT37), .ZN(new_n608));
  OAI21_X1  g407(.A(KEYINPUT38), .B1(new_n606), .B2(new_n608), .ZN(new_n609));
  NAND4_X1  g408(.A1(new_n598), .A2(new_n605), .A3(new_n527), .A4(new_n609), .ZN(new_n610));
  AOI22_X1  g409(.A1(new_n579), .A2(new_n580), .B1(new_n597), .B2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT36), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n612), .B1(new_n557), .B2(new_n558), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n495), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n560), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n612), .B1(new_n615), .B2(new_n411), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n611), .A2(new_n617), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n285), .B1(new_n573), .B2(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(G57gat), .B(G64gat), .ZN(new_n620));
  XOR2_X1   g419(.A(G71gat), .B(G78gat), .Z(new_n621));
  AOI21_X1  g420(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT96), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n622), .B(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT97), .ZN(new_n625));
  AOI211_X1 g424(.A(new_n620), .B(new_n621), .C1(new_n624), .C2(new_n625), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n626), .B1(new_n625), .B2(new_n624), .ZN(new_n627));
  XOR2_X1   g426(.A(new_n621), .B(KEYINPUT95), .Z(new_n628));
  OAI21_X1  g427(.A(new_n628), .B1(new_n624), .B2(new_n620), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT21), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(G231gat), .A2(G233gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(G127gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n634), .B(new_n635), .ZN(new_n636));
  AND2_X1   g435(.A1(new_n627), .A2(new_n629), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n245), .B1(new_n637), .B2(KEYINPUT21), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n634), .B(G127gat), .ZN(new_n640));
  INV_X1    g439(.A(new_n638), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n639), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n644), .B(new_n428), .ZN(new_n645));
  XNOR2_X1  g444(.A(G183gat), .B(G211gat), .ZN(new_n646));
  XOR2_X1   g445(.A(new_n645), .B(new_n646), .Z(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n643), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n639), .A2(new_n642), .A3(new_n647), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(G85gat), .A2(G92gat), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n652), .B(KEYINPUT7), .ZN(new_n653));
  NAND2_X1  g452(.A1(G99gat), .A2(G106gat), .ZN(new_n654));
  INV_X1    g453(.A(G85gat), .ZN(new_n655));
  INV_X1    g454(.A(G92gat), .ZN(new_n656));
  AOI22_X1  g455(.A1(KEYINPUT8), .A2(new_n654), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n653), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g457(.A(G99gat), .B(G106gat), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n658), .B(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT98), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n660), .B(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n239), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(new_n225), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n662), .A2(new_n222), .A3(new_n224), .ZN(new_n666));
  NAND3_X1  g465(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n665), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  XOR2_X1   g467(.A(G190gat), .B(G218gat), .Z(new_n669));
  XOR2_X1   g468(.A(new_n668), .B(new_n669), .Z(new_n670));
  XNOR2_X1  g469(.A(G134gat), .B(G162gat), .ZN(new_n671));
  AOI21_X1  g470(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n670), .B(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n660), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n630), .A2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT10), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n627), .A2(new_n629), .A3(new_n660), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n676), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n662), .A2(KEYINPUT10), .A3(new_n637), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(G230gat), .A2(G233gat), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n676), .A2(new_n678), .ZN(new_n684));
  INV_X1    g483(.A(new_n682), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g486(.A(G120gat), .B(G148gat), .ZN(new_n688));
  XNOR2_X1  g487(.A(G176gat), .B(G204gat), .ZN(new_n689));
  XOR2_X1   g488(.A(new_n688), .B(new_n689), .Z(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  NOR3_X1   g490(.A1(new_n687), .A2(KEYINPUT99), .A3(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  OAI21_X1  g492(.A(KEYINPUT99), .B1(new_n687), .B2(new_n691), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n687), .A2(new_n691), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n651), .A2(new_n674), .A3(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n619), .A2(new_n700), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n701), .A2(new_n529), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(new_n227), .ZN(G1324gat));
  NOR2_X1   g502(.A1(new_n701), .A2(new_n553), .ZN(new_n704));
  XOR2_X1   g503(.A(KEYINPUT16), .B(G8gat), .Z(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n706), .B1(new_n232), .B2(new_n704), .ZN(new_n707));
  MUX2_X1   g506(.A(new_n706), .B(new_n707), .S(KEYINPUT42), .Z(G1325gat));
  OAI21_X1  g507(.A(G15gat), .B1(new_n701), .B2(new_n617), .ZN(new_n709));
  OR2_X1    g508(.A1(new_n561), .A2(G15gat), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n709), .B1(new_n701), .B2(new_n710), .ZN(new_n711));
  XOR2_X1   g510(.A(new_n711), .B(KEYINPUT100), .Z(G1326gat));
  INV_X1    g511(.A(new_n579), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n701), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(KEYINPUT101), .ZN(new_n715));
  XNOR2_X1  g514(.A(KEYINPUT43), .B(G22gat), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n715), .B(new_n716), .ZN(G1327gat));
  INV_X1    g516(.A(new_n651), .ZN(new_n718));
  INV_X1    g517(.A(new_n674), .ZN(new_n719));
  NAND4_X1  g518(.A1(new_n619), .A2(new_n718), .A3(new_n719), .A4(new_n698), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n720), .A2(G29gat), .A3(new_n529), .ZN(new_n721));
  XOR2_X1   g520(.A(new_n721), .B(KEYINPUT45), .Z(new_n722));
  INV_X1    g521(.A(KEYINPUT102), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n723), .B1(new_n276), .B2(new_n280), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n283), .A2(KEYINPUT102), .A3(new_n279), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n718), .A2(new_n698), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(new_n729), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n674), .B1(new_n573), .B2(new_n618), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT44), .ZN(new_n732));
  OAI21_X1  g531(.A(KEYINPUT103), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  AOI22_X1  g532(.A1(new_n612), .A2(new_n561), .B1(new_n495), .B2(new_n613), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n574), .A2(new_n575), .ZN(new_n735));
  AND2_X1   g534(.A1(new_n524), .A2(new_n591), .ZN(new_n736));
  NAND4_X1  g535(.A1(new_n736), .A2(new_n552), .A3(new_n549), .A4(new_n594), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n605), .A2(new_n609), .ZN(new_n738));
  AND3_X1   g537(.A1(new_n564), .A2(new_n565), .A3(KEYINPUT6), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n565), .B1(new_n564), .B2(KEYINPUT6), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n527), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  OAI211_X1 g540(.A(new_n735), .B(new_n737), .C1(new_n738), .C2(new_n741), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n576), .B1(new_n574), .B2(new_n575), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n483), .A2(new_n487), .A3(KEYINPUT83), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n580), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n742), .A2(new_n745), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n734), .A2(new_n746), .ZN(new_n747));
  AOI22_X1  g546(.A1(new_n555), .A2(KEYINPUT35), .B1(new_n562), .B2(new_n571), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n719), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT103), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n749), .A2(new_n750), .A3(KEYINPUT44), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n733), .A2(new_n751), .ZN(new_n752));
  OAI211_X1 g551(.A(new_n732), .B(new_n719), .C1(new_n747), .C2(new_n748), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(KEYINPUT104), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n573), .A2(new_n618), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT104), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n755), .A2(new_n756), .A3(new_n732), .A4(new_n719), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n754), .A2(new_n757), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n730), .B1(new_n752), .B2(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(new_n759), .ZN(new_n760));
  OAI21_X1  g559(.A(G29gat), .B1(new_n760), .B2(new_n529), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n722), .A2(new_n761), .ZN(G1328gat));
  OAI21_X1  g561(.A(G36gat), .B1(new_n760), .B2(new_n553), .ZN(new_n763));
  NOR3_X1   g562(.A1(new_n720), .A2(G36gat), .A3(new_n553), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(KEYINPUT46), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n763), .A2(new_n765), .ZN(G1329gat));
  AOI211_X1 g565(.A(new_n617), .B(new_n730), .C1(new_n752), .C2(new_n758), .ZN(new_n767));
  INV_X1    g566(.A(G43gat), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n562), .A2(new_n768), .ZN(new_n769));
  OAI22_X1  g568(.A1(new_n767), .A2(new_n768), .B1(new_n720), .B2(new_n769), .ZN(new_n770));
  XNOR2_X1  g569(.A(KEYINPUT106), .B(KEYINPUT47), .ZN(new_n771));
  AND3_X1   g570(.A1(new_n770), .A2(KEYINPUT105), .A3(new_n771), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n771), .B1(new_n770), .B2(KEYINPUT105), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n772), .A2(new_n773), .ZN(G1330gat));
  INV_X1    g573(.A(KEYINPUT109), .ZN(new_n775));
  INV_X1    g574(.A(new_n215), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n776), .B1(new_n759), .B2(new_n488), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n579), .A2(new_n776), .ZN(new_n778));
  XOR2_X1   g577(.A(new_n778), .B(KEYINPUT107), .Z(new_n779));
  NOR2_X1   g578(.A1(new_n720), .A2(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT48), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(new_n782), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n775), .B1(new_n777), .B2(new_n783), .ZN(new_n784));
  AOI211_X1 g583(.A(new_n735), .B(new_n730), .C1(new_n752), .C2(new_n758), .ZN(new_n785));
  OAI211_X1 g584(.A(KEYINPUT109), .B(new_n782), .C1(new_n785), .C2(new_n776), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n752), .A2(new_n758), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n788), .A2(new_n579), .A3(new_n729), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n780), .B1(new_n789), .B2(new_n215), .ZN(new_n790));
  NOR3_X1   g589(.A1(new_n790), .A2(KEYINPUT108), .A3(KEYINPUT48), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT108), .ZN(new_n792));
  INV_X1    g591(.A(new_n780), .ZN(new_n793));
  AOI211_X1 g592(.A(new_n713), .B(new_n730), .C1(new_n752), .C2(new_n758), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n793), .B1(new_n794), .B2(new_n776), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n792), .B1(new_n795), .B2(new_n781), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n787), .B1(new_n791), .B2(new_n796), .ZN(G1331gat));
  NOR4_X1   g596(.A1(new_n726), .A2(new_n718), .A3(new_n719), .A4(new_n698), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n755), .A2(new_n798), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n799), .A2(new_n529), .ZN(new_n800));
  XNOR2_X1  g599(.A(KEYINPUT110), .B(G57gat), .ZN(new_n801));
  XNOR2_X1  g600(.A(new_n800), .B(new_n801), .ZN(G1332gat));
  NOR2_X1   g601(.A1(new_n799), .A2(new_n553), .ZN(new_n803));
  NOR2_X1   g602(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n804));
  AND2_X1   g603(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n803), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n806), .B1(new_n803), .B2(new_n804), .ZN(G1333gat));
  OAI21_X1  g606(.A(G71gat), .B1(new_n799), .B2(new_n617), .ZN(new_n808));
  OR2_X1    g607(.A1(new_n561), .A2(G71gat), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n808), .B1(new_n799), .B2(new_n809), .ZN(new_n810));
  XOR2_X1   g609(.A(KEYINPUT111), .B(KEYINPUT50), .Z(new_n811));
  XNOR2_X1  g610(.A(new_n810), .B(new_n811), .ZN(G1334gat));
  NOR2_X1   g611(.A1(new_n799), .A2(new_n713), .ZN(new_n813));
  XOR2_X1   g612(.A(new_n813), .B(G78gat), .Z(G1335gat));
  NOR2_X1   g613(.A1(new_n726), .A2(new_n651), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(new_n697), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n816), .B1(new_n752), .B2(new_n758), .ZN(new_n817));
  INV_X1    g616(.A(new_n817), .ZN(new_n818));
  OAI21_X1  g617(.A(G85gat), .B1(new_n818), .B2(new_n529), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n755), .A2(new_n719), .A3(new_n815), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT51), .ZN(new_n821));
  XNOR2_X1  g620(.A(new_n820), .B(new_n821), .ZN(new_n822));
  AND2_X1   g621(.A1(new_n822), .A2(new_n697), .ZN(new_n823));
  INV_X1    g622(.A(new_n529), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n823), .A2(new_n655), .A3(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n819), .A2(new_n825), .ZN(G1336gat));
  INV_X1    g625(.A(new_n553), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n697), .A2(new_n827), .A3(new_n656), .ZN(new_n828));
  XOR2_X1   g627(.A(new_n828), .B(KEYINPUT112), .Z(new_n829));
  AND2_X1   g628(.A1(new_n822), .A2(new_n829), .ZN(new_n830));
  XNOR2_X1  g629(.A(KEYINPUT113), .B(KEYINPUT52), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  AOI211_X1 g631(.A(new_n553), .B(new_n816), .C1(new_n752), .C2(new_n758), .ZN(new_n833));
  AND2_X1   g632(.A1(new_n833), .A2(KEYINPUT114), .ZN(new_n834));
  OAI21_X1  g633(.A(G92gat), .B1(new_n833), .B2(KEYINPUT114), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n832), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n833), .A2(new_n656), .ZN(new_n837));
  OAI21_X1  g636(.A(KEYINPUT52), .B1(new_n837), .B2(new_n830), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n836), .A2(new_n838), .ZN(G1337gat));
  OAI21_X1  g638(.A(G99gat), .B1(new_n818), .B2(new_n617), .ZN(new_n840));
  INV_X1    g639(.A(G99gat), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n823), .A2(new_n841), .A3(new_n562), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n840), .A2(new_n842), .ZN(G1338gat));
  NOR2_X1   g642(.A1(new_n735), .A2(G106gat), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n822), .A2(new_n697), .A3(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT115), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND4_X1  g646(.A1(new_n822), .A2(KEYINPUT115), .A3(new_n697), .A4(new_n844), .ZN(new_n848));
  AOI21_X1  g647(.A(KEYINPUT53), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  AOI211_X1 g648(.A(new_n735), .B(new_n816), .C1(new_n752), .C2(new_n758), .ZN(new_n850));
  OAI21_X1  g649(.A(G106gat), .B1(new_n850), .B2(KEYINPUT116), .ZN(new_n851));
  AND2_X1   g650(.A1(new_n850), .A2(KEYINPUT116), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n849), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(G106gat), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n854), .B1(new_n817), .B2(new_n579), .ZN(new_n855));
  INV_X1    g654(.A(new_n845), .ZN(new_n856));
  OAI21_X1  g655(.A(KEYINPUT53), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n853), .A2(new_n857), .ZN(G1339gat));
  INV_X1    g657(.A(KEYINPUT99), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n685), .B1(new_n679), .B2(new_n680), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n860), .B1(new_n685), .B2(new_n684), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n859), .B1(new_n861), .B2(new_n690), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT55), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n679), .A2(new_n680), .A3(new_n685), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n683), .A2(KEYINPUT54), .A3(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT54), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n690), .B1(new_n860), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  OAI22_X1  g667(.A1(new_n862), .A2(new_n692), .B1(new_n863), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n863), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT117), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n868), .A2(KEYINPUT117), .A3(new_n863), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n869), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  AND3_X1   g673(.A1(new_n283), .A2(KEYINPUT102), .A3(new_n279), .ZN(new_n875));
  AOI21_X1  g674(.A(KEYINPUT102), .B1(new_n283), .B2(new_n279), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n874), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n264), .A2(new_n246), .A3(new_n262), .ZN(new_n878));
  XNOR2_X1  g677(.A(new_n878), .B(KEYINPUT118), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n244), .B1(new_n252), .B2(new_n243), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n258), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  AND2_X1   g680(.A1(new_n881), .A2(new_n267), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n697), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n719), .B1(new_n877), .B2(new_n883), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n719), .A2(new_n874), .A3(new_n882), .ZN(new_n885));
  INV_X1    g684(.A(new_n885), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n718), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n699), .A2(new_n726), .ZN(new_n888));
  INV_X1    g687(.A(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n579), .A2(new_n561), .ZN(new_n891));
  AND2_X1   g690(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n827), .A2(new_n529), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NOR3_X1   g693(.A1(new_n894), .A2(new_n345), .A3(new_n285), .ZN(new_n895));
  AND2_X1   g694(.A1(new_n697), .A2(new_n882), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n896), .B1(new_n726), .B2(new_n874), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n885), .B1(new_n897), .B2(new_n719), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n888), .B1(new_n898), .B2(new_n718), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n899), .A2(new_n529), .ZN(new_n900));
  AND2_X1   g699(.A1(new_n489), .A2(new_n495), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n900), .A2(new_n553), .A3(new_n901), .ZN(new_n902));
  INV_X1    g701(.A(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(new_n726), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n895), .B1(new_n345), .B2(new_n904), .ZN(G1340gat));
  NOR3_X1   g704(.A1(new_n894), .A2(new_n348), .A3(new_n698), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n903), .A2(new_n697), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n906), .B1(new_n348), .B2(new_n907), .ZN(G1341gat));
  OAI21_X1  g707(.A(G127gat), .B1(new_n894), .B2(new_n718), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n651), .A2(new_n635), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n909), .B1(new_n902), .B2(new_n910), .ZN(G1342gat));
  NOR3_X1   g710(.A1(new_n674), .A2(G134gat), .A3(new_n827), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n900), .A2(new_n901), .A3(new_n912), .ZN(new_n913));
  OR2_X1    g712(.A1(new_n913), .A2(KEYINPUT56), .ZN(new_n914));
  OAI21_X1  g713(.A(G134gat), .B1(new_n894), .B2(new_n674), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n913), .A2(KEYINPUT56), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n914), .A2(new_n915), .A3(new_n916), .ZN(G1343gat));
  NAND2_X1  g716(.A1(new_n900), .A2(KEYINPUT120), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n734), .A2(new_n735), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n900), .A2(KEYINPUT120), .ZN(new_n921));
  OAI21_X1  g720(.A(KEYINPUT121), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(new_n921), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT121), .ZN(new_n924));
  NAND4_X1  g723(.A1(new_n923), .A2(new_n924), .A3(new_n919), .A4(new_n918), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n285), .A2(G141gat), .ZN(new_n926));
  NAND4_X1  g725(.A1(new_n922), .A2(new_n925), .A3(new_n553), .A4(new_n926), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT58), .ZN(new_n928));
  AND2_X1   g727(.A1(new_n617), .A2(new_n893), .ZN(new_n929));
  INV_X1    g728(.A(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT57), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n713), .A2(new_n931), .ZN(new_n932));
  INV_X1    g731(.A(new_n869), .ZN(new_n933));
  NAND4_X1  g732(.A1(new_n281), .A2(new_n284), .A3(new_n933), .A4(new_n870), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n719), .B1(new_n934), .B2(new_n883), .ZN(new_n935));
  INV_X1    g734(.A(new_n935), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n651), .B1(new_n936), .B2(new_n885), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n937), .A2(KEYINPUT119), .ZN(new_n938));
  OAI211_X1 g737(.A(KEYINPUT119), .B(new_n718), .C1(new_n935), .C2(new_n886), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n939), .A2(new_n889), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n932), .B1(new_n938), .B2(new_n940), .ZN(new_n941));
  AOI21_X1  g740(.A(KEYINPUT57), .B1(new_n890), .B2(new_n488), .ZN(new_n942));
  INV_X1    g741(.A(new_n942), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n930), .B1(new_n941), .B2(new_n943), .ZN(new_n944));
  INV_X1    g743(.A(new_n944), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n945), .A2(new_n285), .ZN(new_n946));
  OAI211_X1 g745(.A(new_n927), .B(new_n928), .C1(new_n448), .C2(new_n946), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n448), .B1(new_n944), .B2(new_n726), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n926), .A2(new_n553), .ZN(new_n949));
  NOR3_X1   g748(.A1(new_n920), .A2(new_n921), .A3(new_n949), .ZN(new_n950));
  OAI21_X1  g749(.A(KEYINPUT58), .B1(new_n948), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n947), .A2(new_n951), .ZN(G1344gat));
  OAI21_X1  g751(.A(KEYINPUT57), .B1(new_n899), .B2(new_n735), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n699), .B1(new_n284), .B2(new_n281), .ZN(new_n954));
  OAI211_X1 g753(.A(new_n931), .B(new_n579), .C1(new_n937), .C2(new_n954), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n698), .B1(new_n930), .B2(KEYINPUT123), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n957), .B1(KEYINPUT123), .B2(new_n930), .ZN(new_n958));
  OAI21_X1  g757(.A(G148gat), .B1(new_n956), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n959), .A2(KEYINPUT59), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n944), .A2(new_n697), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n433), .A2(KEYINPUT59), .ZN(new_n962));
  AOI21_X1  g761(.A(KEYINPUT122), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT122), .ZN(new_n964));
  INV_X1    g763(.A(new_n962), .ZN(new_n965));
  AOI211_X1 g764(.A(new_n964), .B(new_n965), .C1(new_n944), .C2(new_n697), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n960), .B1(new_n963), .B2(new_n966), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n922), .A2(new_n925), .A3(new_n553), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n697), .A2(new_n433), .ZN(new_n969));
  OR2_X1    g768(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n967), .A2(new_n970), .ZN(G1345gat));
  OAI21_X1  g770(.A(G155gat), .B1(new_n945), .B2(new_n718), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n651), .A2(new_n428), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n972), .B1(new_n968), .B2(new_n973), .ZN(G1346gat));
  OAI21_X1  g773(.A(G162gat), .B1(new_n945), .B2(new_n674), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n922), .A2(new_n925), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n719), .A2(new_n429), .A3(new_n553), .ZN(new_n977));
  OAI21_X1  g776(.A(new_n975), .B1(new_n976), .B2(new_n977), .ZN(G1347gat));
  NOR2_X1   g777(.A1(new_n824), .A2(new_n553), .ZN(new_n979));
  AND3_X1   g778(.A1(new_n890), .A2(new_n891), .A3(new_n979), .ZN(new_n980));
  INV_X1    g779(.A(new_n980), .ZN(new_n981));
  NOR3_X1   g780(.A1(new_n981), .A2(new_n287), .A3(new_n285), .ZN(new_n982));
  OAI21_X1  g781(.A(KEYINPUT124), .B1(new_n899), .B2(new_n824), .ZN(new_n983));
  INV_X1    g782(.A(KEYINPUT124), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n890), .A2(new_n984), .A3(new_n529), .ZN(new_n985));
  AOI21_X1  g784(.A(new_n553), .B1(new_n983), .B2(new_n985), .ZN(new_n986));
  NAND3_X1  g785(.A1(new_n986), .A2(new_n901), .A3(new_n726), .ZN(new_n987));
  AOI21_X1  g786(.A(new_n982), .B1(new_n987), .B2(new_n287), .ZN(G1348gat));
  NOR3_X1   g787(.A1(new_n981), .A2(new_n365), .A3(new_n698), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n986), .A2(new_n901), .A3(new_n697), .ZN(new_n990));
  AOI21_X1  g789(.A(new_n989), .B1(new_n990), .B2(new_n288), .ZN(G1349gat));
  INV_X1    g790(.A(KEYINPUT126), .ZN(new_n992));
  AOI21_X1  g791(.A(new_n299), .B1(new_n980), .B2(new_n651), .ZN(new_n993));
  NOR3_X1   g792(.A1(new_n718), .A2(new_n303), .A3(new_n553), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n994), .A2(new_n901), .ZN(new_n995));
  INV_X1    g794(.A(new_n995), .ZN(new_n996));
  AOI21_X1  g795(.A(new_n984), .B1(new_n890), .B2(new_n529), .ZN(new_n997));
  AOI211_X1 g796(.A(KEYINPUT124), .B(new_n824), .C1(new_n887), .C2(new_n889), .ZN(new_n998));
  OAI21_X1  g797(.A(new_n996), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  INV_X1    g798(.A(KEYINPUT125), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g800(.A1(new_n983), .A2(new_n985), .ZN(new_n1002));
  NAND3_X1  g801(.A1(new_n1002), .A2(KEYINPUT125), .A3(new_n996), .ZN(new_n1003));
  AOI21_X1  g802(.A(new_n993), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g803(.A(KEYINPUT60), .ZN(new_n1005));
  OAI21_X1  g804(.A(new_n992), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g805(.A(new_n993), .ZN(new_n1007));
  AOI21_X1  g806(.A(KEYINPUT125), .B1(new_n1002), .B2(new_n996), .ZN(new_n1008));
  AOI211_X1 g807(.A(new_n1000), .B(new_n995), .C1(new_n983), .C2(new_n985), .ZN(new_n1009));
  OAI21_X1  g808(.A(new_n1007), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g809(.A1(new_n1010), .A2(KEYINPUT126), .A3(KEYINPUT60), .ZN(new_n1011));
  NAND2_X1  g810(.A1(new_n1006), .A2(new_n1011), .ZN(new_n1012));
  OAI211_X1 g811(.A(new_n1005), .B(new_n1007), .C1(new_n1008), .C2(new_n1009), .ZN(new_n1013));
  INV_X1    g812(.A(KEYINPUT127), .ZN(new_n1014));
  NAND2_X1  g813(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g814(.A1(new_n1004), .A2(KEYINPUT127), .A3(new_n1005), .ZN(new_n1016));
  NAND2_X1  g815(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g816(.A1(new_n1012), .A2(new_n1017), .ZN(G1350gat));
  OAI21_X1  g817(.A(G190gat), .B1(new_n981), .B2(new_n674), .ZN(new_n1019));
  AND2_X1   g818(.A1(new_n1019), .A2(KEYINPUT61), .ZN(new_n1020));
  NOR2_X1   g819(.A1(new_n1019), .A2(KEYINPUT61), .ZN(new_n1021));
  NAND2_X1  g820(.A1(new_n986), .A2(new_n901), .ZN(new_n1022));
  NAND2_X1  g821(.A1(new_n719), .A2(new_n329), .ZN(new_n1023));
  OAI22_X1  g822(.A1(new_n1020), .A2(new_n1021), .B1(new_n1022), .B2(new_n1023), .ZN(G1351gat));
  NAND2_X1  g823(.A1(new_n986), .A2(new_n919), .ZN(new_n1025));
  INV_X1    g824(.A(new_n1025), .ZN(new_n1026));
  AOI21_X1  g825(.A(G197gat), .B1(new_n1026), .B2(new_n726), .ZN(new_n1027));
  NAND2_X1  g826(.A1(new_n617), .A2(new_n979), .ZN(new_n1028));
  OR2_X1    g827(.A1(new_n956), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g828(.A(G197gat), .ZN(new_n1030));
  NOR3_X1   g829(.A1(new_n1029), .A2(new_n1030), .A3(new_n285), .ZN(new_n1031));
  NOR2_X1   g830(.A1(new_n1027), .A2(new_n1031), .ZN(G1352gat));
  NOR2_X1   g831(.A1(new_n698), .A2(G204gat), .ZN(new_n1033));
  INV_X1    g832(.A(new_n1033), .ZN(new_n1034));
  OR3_X1    g833(.A1(new_n1025), .A2(KEYINPUT62), .A3(new_n1034), .ZN(new_n1035));
  OAI21_X1  g834(.A(G204gat), .B1(new_n1029), .B2(new_n698), .ZN(new_n1036));
  OAI21_X1  g835(.A(KEYINPUT62), .B1(new_n1025), .B2(new_n1034), .ZN(new_n1037));
  NAND3_X1  g836(.A1(new_n1035), .A2(new_n1036), .A3(new_n1037), .ZN(G1353gat));
  NAND3_X1  g837(.A1(new_n1026), .A2(new_n415), .A3(new_n651), .ZN(new_n1039));
  OR3_X1    g838(.A1(new_n956), .A2(new_n718), .A3(new_n1028), .ZN(new_n1040));
  AND3_X1   g839(.A1(new_n1040), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1041));
  AOI21_X1  g840(.A(KEYINPUT63), .B1(new_n1040), .B2(G211gat), .ZN(new_n1042));
  OAI21_X1  g841(.A(new_n1039), .B1(new_n1041), .B2(new_n1042), .ZN(G1354gat));
  NAND3_X1  g842(.A1(new_n1026), .A2(new_n416), .A3(new_n719), .ZN(new_n1044));
  OAI21_X1  g843(.A(G218gat), .B1(new_n1029), .B2(new_n674), .ZN(new_n1045));
  NAND2_X1  g844(.A1(new_n1044), .A2(new_n1045), .ZN(G1355gat));
endmodule


