//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 1 0 1 0 1 0 0 1 1 0 1 0 1 0 0 1 0 1 0 1 0 0 1 0 0 1 1 0 0 0 0 0 1 1 1 0 0 0 1 1 0 0 0 1 1 0 0 0 1 0 0 1 0 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:56 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n210, new_n211, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1297, new_n1298, new_n1299, new_n1300, new_n1301, new_n1303,
    new_n1304, new_n1305, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1358, new_n1359,
    new_n1360, new_n1361, new_n1362, new_n1363, new_n1364, new_n1365,
    new_n1366, new_n1367, new_n1368, new_n1369, new_n1370;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G50), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G77), .ZN(G353));
  NOR2_X1   g0009(.A1(G97), .A2(G107), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n211), .A2(G87), .ZN(G355));
  NAND2_X1  g0012(.A1(G1), .A2(G20), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT65), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(G13), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n215), .B(G250), .C1(G257), .C2(G264), .ZN(new_n216));
  XOR2_X1   g0016(.A(new_n216), .B(KEYINPUT0), .Z(new_n217));
  NAND2_X1  g0017(.A1(G1), .A2(G13), .ZN(new_n218));
  INV_X1    g0018(.A(G20), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n206), .A2(new_n207), .ZN(new_n221));
  AOI21_X1  g0021(.A(new_n217), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n223));
  XOR2_X1   g0023(.A(new_n223), .B(KEYINPUT66), .Z(new_n224));
  AOI22_X1  g0024(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G97), .A2(G257), .B1(G107), .B2(G264), .ZN(new_n227));
  NAND3_X1  g0027(.A1(new_n225), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n214), .B1(new_n224), .B2(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT67), .ZN(new_n230));
  INV_X1    g0030(.A(KEYINPUT1), .ZN(new_n231));
  OR2_X1    g0031(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n230), .A2(new_n231), .ZN(new_n233));
  AND3_X1   g0033(.A1(new_n222), .A2(new_n232), .A3(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n238), .B(new_n241), .Z(G358));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n207), .A2(G68), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n203), .A2(G50), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G58), .B(G77), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n245), .B(new_n250), .ZN(G351));
  NAND3_X1  g0051(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n252));
  AND2_X1   g0052(.A1(new_n252), .A2(new_n218), .ZN(new_n253));
  AOI21_X1  g0053(.A(new_n219), .B1(new_n206), .B2(new_n207), .ZN(new_n254));
  OR2_X1    g0054(.A1(new_n254), .A2(KEYINPUT70), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(KEYINPUT70), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NOR2_X1   g0057(.A1(KEYINPUT8), .A2(G58), .ZN(new_n258));
  XNOR2_X1  g0058(.A(KEYINPUT69), .B(G58), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n258), .B1(new_n259), .B2(KEYINPUT8), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n219), .A2(G33), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  NOR2_X1   g0062(.A1(G20), .A2(G33), .ZN(new_n263));
  AOI22_X1  g0063(.A1(new_n260), .A2(new_n262), .B1(G150), .B2(new_n263), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n253), .B1(new_n257), .B2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G1), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n266), .A2(G13), .A3(G20), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n267), .A2(G50), .ZN(new_n268));
  OAI211_X1 g0068(.A(new_n252), .B(new_n218), .C1(G1), .C2(new_n219), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n268), .B1(new_n270), .B2(G50), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  OR3_X1    g0072(.A1(new_n265), .A2(KEYINPUT9), .A3(new_n272), .ZN(new_n273));
  OAI21_X1  g0073(.A(KEYINPUT9), .B1(new_n265), .B2(new_n272), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT10), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n218), .B1(G33), .B2(G41), .ZN(new_n277));
  XNOR2_X1  g0077(.A(KEYINPUT3), .B(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G1698), .ZN(new_n279));
  XOR2_X1   g0079(.A(KEYINPUT68), .B(G223), .Z(new_n280));
  INV_X1    g0080(.A(G77), .ZN(new_n281));
  OAI22_X1  g0081(.A1(new_n279), .A2(new_n280), .B1(new_n281), .B2(new_n278), .ZN(new_n282));
  INV_X1    g0082(.A(G1698), .ZN(new_n283));
  AND3_X1   g0083(.A1(new_n278), .A2(G222), .A3(new_n283), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n277), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n266), .B1(G41), .B2(G45), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G33), .ZN(new_n288));
  INV_X1    g0088(.A(G41), .ZN(new_n289));
  OAI211_X1 g0089(.A(G1), .B(G13), .C1(new_n288), .C2(new_n289), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n287), .A2(new_n290), .A3(G274), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n277), .A2(new_n287), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n292), .B1(G226), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n285), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n296), .A2(KEYINPUT72), .A3(G190), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT72), .ZN(new_n298));
  INV_X1    g0098(.A(G190), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n298), .B1(new_n295), .B2(new_n299), .ZN(new_n300));
  AOI22_X1  g0100(.A1(new_n297), .A2(new_n300), .B1(G200), .B2(new_n295), .ZN(new_n301));
  AND3_X1   g0101(.A1(new_n275), .A2(new_n276), .A3(new_n301), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n276), .B1(new_n275), .B2(new_n301), .ZN(new_n303));
  OR2_X1    g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n265), .A2(new_n272), .ZN(new_n305));
  INV_X1    g0105(.A(G169), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n305), .B1(new_n306), .B2(new_n295), .ZN(new_n307));
  INV_X1    g0107(.A(G179), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n296), .A2(new_n308), .ZN(new_n309));
  AND2_X1   g0109(.A1(new_n309), .A2(KEYINPUT71), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n309), .A2(KEYINPUT71), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n307), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT12), .ZN(new_n313));
  INV_X1    g0113(.A(new_n267), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n313), .B1(new_n314), .B2(new_n203), .ZN(new_n315));
  NOR3_X1   g0115(.A1(new_n267), .A2(KEYINPUT12), .A3(G68), .ZN(new_n316));
  OAI22_X1  g0116(.A1(new_n315), .A2(new_n316), .B1(new_n269), .B2(new_n203), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT11), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n252), .A2(new_n218), .ZN(new_n319));
  INV_X1    g0119(.A(new_n263), .ZN(new_n320));
  OAI22_X1  g0120(.A1(new_n320), .A2(new_n207), .B1(new_n219), .B2(G68), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n261), .A2(new_n281), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n319), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n317), .B1(new_n318), .B2(new_n323), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n324), .B1(new_n318), .B2(new_n323), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n292), .B1(G238), .B2(new_n293), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n278), .A2(G232), .A3(G1698), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n278), .A2(G226), .A3(new_n283), .ZN(new_n328));
  NAND2_X1  g0128(.A1(G33), .A2(G97), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n327), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(new_n277), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n326), .A2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT13), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n326), .A2(KEYINPUT13), .A3(new_n331), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n334), .A2(G169), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(KEYINPUT14), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT73), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n335), .A2(new_n338), .ZN(new_n339));
  AOI22_X1  g0139(.A1(new_n326), .A2(new_n331), .B1(KEYINPUT73), .B2(KEYINPUT13), .ZN(new_n340));
  OAI21_X1  g0140(.A(G179), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n337), .A2(new_n341), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n336), .A2(KEYINPUT14), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n325), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  AND2_X1   g0144(.A1(new_n334), .A2(new_n335), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n325), .B1(new_n345), .B2(G200), .ZN(new_n346));
  OAI21_X1  g0146(.A(G190), .B1(new_n339), .B2(new_n340), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n344), .A2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  XOR2_X1   g0150(.A(KEYINPUT8), .B(G58), .Z(new_n351));
  AOI22_X1  g0151(.A1(new_n351), .A2(new_n263), .B1(G20), .B2(G77), .ZN(new_n352));
  XNOR2_X1  g0152(.A(KEYINPUT15), .B(G87), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n352), .B1(new_n261), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(new_n319), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n270), .A2(G77), .ZN(new_n356));
  OAI211_X1 g0156(.A(new_n355), .B(new_n356), .C1(G77), .C2(new_n267), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n278), .A2(G232), .A3(new_n283), .ZN(new_n358));
  INV_X1    g0158(.A(G107), .ZN(new_n359));
  INV_X1    g0159(.A(G238), .ZN(new_n360));
  OAI221_X1 g0160(.A(new_n358), .B1(new_n359), .B2(new_n278), .C1(new_n279), .C2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(new_n277), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n292), .B1(G244), .B2(new_n293), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n357), .B1(G200), .B2(new_n364), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n365), .B1(new_n299), .B2(new_n364), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n364), .A2(new_n306), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n362), .A2(new_n308), .A3(new_n363), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n367), .A2(new_n368), .A3(new_n357), .ZN(new_n369));
  AND2_X1   g0169(.A1(new_n366), .A2(new_n369), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n304), .A2(new_n312), .A3(new_n350), .A4(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT16), .ZN(new_n372));
  OR2_X1    g0172(.A1(KEYINPUT69), .A2(G58), .ZN(new_n373));
  NAND2_X1  g0173(.A1(KEYINPUT69), .A2(G58), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n203), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  OAI21_X1  g0175(.A(G20), .B1(new_n375), .B2(new_n206), .ZN(new_n376));
  INV_X1    g0176(.A(G159), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n376), .B1(new_n377), .B2(new_n320), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT7), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n379), .B1(new_n278), .B2(G20), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n288), .A2(KEYINPUT3), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT3), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(G33), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n384), .A2(KEYINPUT7), .A3(new_n219), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n203), .B1(new_n380), .B2(new_n385), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n372), .B1(new_n378), .B2(new_n386), .ZN(new_n387));
  NOR3_X1   g0187(.A1(new_n278), .A2(new_n379), .A3(G20), .ZN(new_n388));
  AOI21_X1  g0188(.A(KEYINPUT7), .B1(new_n384), .B2(new_n219), .ZN(new_n389));
  OAI21_X1  g0189(.A(G68), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  AND2_X1   g0190(.A1(KEYINPUT69), .A2(G58), .ZN(new_n391));
  NOR2_X1   g0191(.A1(KEYINPUT69), .A2(G58), .ZN(new_n392));
  OAI21_X1  g0192(.A(G68), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n393), .A2(new_n204), .A3(new_n205), .ZN(new_n394));
  AOI22_X1  g0194(.A1(new_n394), .A2(G20), .B1(G159), .B2(new_n263), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n390), .A2(new_n395), .A3(KEYINPUT16), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n387), .A2(new_n396), .A3(new_n319), .ZN(new_n397));
  INV_X1    g0197(.A(new_n258), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n391), .A2(new_n392), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT8), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n398), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(new_n267), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n260), .A2(new_n269), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT74), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n402), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(new_n405), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n404), .B1(new_n402), .B2(new_n403), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n290), .A2(G232), .A3(new_n286), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n291), .A2(new_n409), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n381), .A2(new_n383), .A3(G226), .A4(G1698), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n381), .A2(new_n383), .A3(G223), .A4(new_n283), .ZN(new_n412));
  NAND2_X1  g0212(.A1(G33), .A2(G87), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n410), .B1(new_n414), .B2(new_n277), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(G190), .ZN(new_n416));
  INV_X1    g0216(.A(G200), .ZN(new_n417));
  OR2_X1    g0217(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n397), .A2(new_n408), .A3(new_n416), .A4(new_n418), .ZN(new_n419));
  XNOR2_X1  g0219(.A(new_n419), .B(KEYINPUT17), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n414), .A2(new_n277), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n421), .A2(new_n308), .A3(new_n291), .A4(new_n409), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n422), .B1(new_n415), .B2(G169), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n423), .B1(new_n397), .B2(new_n408), .ZN(new_n424));
  AOI21_X1  g0224(.A(KEYINPUT75), .B1(new_n424), .B2(KEYINPUT18), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n424), .A2(KEYINPUT18), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NOR3_X1   g0227(.A1(new_n424), .A2(KEYINPUT75), .A3(KEYINPUT18), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n420), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n371), .A2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  XNOR2_X1  g0231(.A(KEYINPUT5), .B(G41), .ZN(new_n432));
  INV_X1    g0232(.A(G45), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n433), .A2(G1), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n435), .A2(G270), .A3(new_n290), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n432), .A2(new_n290), .A3(G274), .A4(new_n434), .ZN(new_n437));
  AND2_X1   g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n278), .A2(G264), .A3(G1698), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n278), .A2(G257), .A3(new_n283), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n384), .A2(G303), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n439), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(new_n277), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n438), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT20), .ZN(new_n445));
  INV_X1    g0245(.A(G97), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n219), .B1(new_n446), .B2(G33), .ZN(new_n447));
  NAND2_X1  g0247(.A1(G33), .A2(G283), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(KEYINPUT76), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT76), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n450), .A2(G33), .A3(G283), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n447), .B1(new_n449), .B2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(G116), .ZN(new_n453));
  AOI22_X1  g0253(.A1(new_n252), .A2(new_n218), .B1(G20), .B2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n445), .B1(new_n452), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n449), .A2(new_n451), .ZN(new_n457));
  INV_X1    g0257(.A(new_n447), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n459), .A2(KEYINPUT20), .A3(new_n454), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n456), .A2(new_n460), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n267), .A2(G116), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n266), .A2(G33), .ZN(new_n463));
  AND3_X1   g0263(.A1(new_n253), .A2(new_n267), .A3(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n462), .B1(new_n464), .B2(G116), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n461), .A2(new_n465), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n444), .A2(new_n466), .A3(KEYINPUT21), .A4(G169), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n436), .A2(new_n437), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n468), .B1(new_n277), .B2(new_n442), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n469), .A2(new_n466), .A3(G179), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n306), .B1(new_n438), .B2(new_n443), .ZN(new_n472));
  AOI21_X1  g0272(.A(KEYINPUT21), .B1(new_n472), .B2(new_n466), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  AND2_X1   g0274(.A1(new_n461), .A2(new_n465), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n438), .A2(new_n443), .A3(G190), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n475), .B(new_n476), .C1(new_n469), .C2(new_n417), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n474), .A2(KEYINPUT79), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n472), .A2(new_n466), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT21), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n481), .A2(new_n477), .A3(new_n470), .A4(new_n467), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT79), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n478), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n435), .A2(G264), .A3(new_n290), .ZN(new_n486));
  AND2_X1   g0286(.A1(new_n486), .A2(new_n437), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n278), .A2(G257), .A3(G1698), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n278), .A2(G250), .A3(new_n283), .ZN(new_n489));
  NAND2_X1  g0289(.A1(G33), .A2(G294), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n488), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(new_n277), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n487), .A2(new_n492), .A3(G179), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n486), .A2(new_n437), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n494), .B1(new_n277), .B2(new_n491), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n493), .B1(new_n495), .B2(new_n306), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(KEYINPUT82), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT82), .ZN(new_n498));
  OAI211_X1 g0298(.A(new_n493), .B(new_n498), .C1(new_n495), .C2(new_n306), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n381), .A2(new_n383), .A3(new_n219), .A4(G87), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(KEYINPUT22), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT22), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n278), .A2(new_n502), .A3(new_n219), .A4(G87), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  XNOR2_X1  g0304(.A(KEYINPUT80), .B(KEYINPUT24), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT23), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n506), .B1(new_n219), .B2(G107), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n359), .A2(KEYINPUT23), .A3(G20), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n288), .A2(new_n453), .ZN(new_n509));
  AOI22_X1  g0309(.A1(new_n507), .A2(new_n508), .B1(new_n509), .B2(new_n219), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n504), .A2(new_n505), .A3(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n505), .B1(new_n504), .B2(new_n510), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n319), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT81), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT25), .ZN(new_n516));
  AOI211_X1 g0316(.A(G107), .B(new_n267), .C1(new_n515), .C2(new_n516), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n515), .A2(new_n516), .ZN(new_n518));
  OR2_X1    g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n517), .A2(new_n518), .ZN(new_n520));
  AOI22_X1  g0320(.A1(new_n519), .A2(new_n520), .B1(G107), .B2(new_n464), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n514), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n497), .A2(new_n499), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n487), .A2(new_n492), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(G200), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n487), .A2(new_n492), .A3(G190), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n514), .A2(new_n525), .A3(new_n521), .A4(new_n526), .ZN(new_n527));
  AND2_X1   g0327(.A1(new_n523), .A2(new_n527), .ZN(new_n528));
  OAI21_X1  g0328(.A(G107), .B1(new_n388), .B2(new_n389), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n359), .A2(KEYINPUT6), .A3(G97), .ZN(new_n530));
  AND2_X1   g0330(.A1(G97), .A2(G107), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n531), .A2(new_n210), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n530), .B1(new_n532), .B2(KEYINPUT6), .ZN(new_n533));
  AOI22_X1  g0333(.A1(new_n533), .A2(G20), .B1(G77), .B2(new_n263), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n529), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n319), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n267), .A2(G97), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n253), .A2(new_n267), .A3(new_n463), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n538), .B1(new_n539), .B2(new_n446), .ZN(new_n540));
  INV_X1    g0340(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n536), .A2(new_n541), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n381), .A2(new_n383), .A3(G244), .A4(new_n283), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT4), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n278), .A2(KEYINPUT4), .A3(G244), .A4(new_n283), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n278), .A2(G250), .A3(G1698), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n545), .A2(new_n546), .A3(new_n457), .A4(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n277), .ZN(new_n549));
  AND3_X1   g0349(.A1(new_n435), .A2(G257), .A3(new_n290), .ZN(new_n550));
  INV_X1    g0350(.A(new_n550), .ZN(new_n551));
  AND4_X1   g0351(.A1(G179), .A2(new_n549), .A3(new_n437), .A4(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n550), .B1(new_n548), .B2(new_n277), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n306), .B1(new_n553), .B2(new_n437), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n542), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n553), .A2(G190), .A3(new_n437), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n540), .B1(new_n535), .B2(new_n319), .ZN(new_n557));
  INV_X1    g0357(.A(new_n437), .ZN(new_n558));
  AOI211_X1 g0358(.A(new_n558), .B(new_n550), .C1(new_n277), .C2(new_n548), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n556), .B(new_n557), .C1(new_n559), .C2(new_n417), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n555), .A2(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(new_n561), .ZN(new_n562));
  AND3_X1   g0362(.A1(new_n290), .A2(G274), .A3(new_n434), .ZN(new_n563));
  INV_X1    g0363(.A(new_n509), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n360), .A2(new_n283), .ZN(new_n565));
  INV_X1    g0365(.A(G244), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(G1698), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n564), .B1(new_n384), .B2(new_n568), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n563), .B1(new_n569), .B2(new_n277), .ZN(new_n570));
  OAI21_X1  g0370(.A(G250), .B1(new_n433), .B2(G1), .ZN(new_n571));
  OAI21_X1  g0371(.A(KEYINPUT77), .B1(new_n277), .B2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(new_n571), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT77), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n573), .A2(new_n290), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n570), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n306), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT19), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n219), .B1(new_n329), .B2(new_n579), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n580), .B1(G87), .B2(new_n211), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n381), .A2(new_n383), .A3(new_n219), .A4(G68), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n579), .B1(new_n261), .B2(new_n446), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n319), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n353), .A2(new_n314), .ZN(new_n586));
  OAI211_X1 g0386(.A(new_n585), .B(new_n586), .C1(new_n353), .C2(new_n539), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n570), .A2(new_n308), .A3(new_n576), .ZN(new_n588));
  AND3_X1   g0388(.A1(new_n578), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n464), .A2(G87), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n585), .A2(new_n586), .A3(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(new_n591), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n570), .A2(KEYINPUT78), .A3(G190), .A4(new_n576), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n569), .A2(new_n277), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n290), .A2(G274), .A3(new_n434), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n594), .A2(new_n576), .A3(G190), .A4(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT78), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n417), .B1(new_n570), .B2(new_n576), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n593), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n589), .B1(new_n592), .B2(new_n600), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n485), .A2(new_n528), .A3(new_n562), .A4(new_n601), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n431), .A2(new_n602), .ZN(G372));
  INV_X1    g0403(.A(KEYINPUT18), .ZN(new_n604));
  AOI211_X1 g0404(.A(new_n604), .B(new_n423), .C1(new_n397), .C2(new_n408), .ZN(new_n605));
  OR2_X1    g0405(.A1(new_n426), .A2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT89), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n369), .A2(new_n608), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n367), .A2(KEYINPUT89), .A3(new_n357), .A4(new_n368), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n348), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n344), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n607), .B1(new_n612), .B2(new_n420), .ZN(new_n613));
  INV_X1    g0413(.A(new_n304), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n312), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT84), .ZN(new_n617));
  NOR2_X1   g0417(.A1(G238), .A2(G1698), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n618), .B1(new_n566), .B2(G1698), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n509), .B1(new_n619), .B2(new_n278), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n595), .B1(new_n620), .B2(new_n290), .ZN(new_n621));
  AND2_X1   g0421(.A1(new_n572), .A2(new_n575), .ZN(new_n622));
  OAI21_X1  g0422(.A(G200), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n623), .A2(new_n597), .A3(new_n596), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n591), .A2(KEYINPUT83), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT83), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n585), .A2(new_n626), .A3(new_n586), .A4(new_n590), .ZN(new_n627));
  AOI22_X1  g0427(.A1(new_n624), .A2(new_n593), .B1(new_n625), .B2(new_n627), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n617), .B1(new_n628), .B2(new_n589), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n625), .A2(new_n627), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n600), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n578), .A2(new_n587), .A3(new_n588), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n631), .A2(KEYINPUT84), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n629), .A2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n513), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n253), .B1(new_n635), .B2(new_n511), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n519), .A2(new_n520), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n464), .A2(G107), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n496), .B1(new_n636), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(KEYINPUT85), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT85), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n522), .A2(new_n642), .A3(new_n496), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n641), .A2(new_n474), .A3(new_n643), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n555), .A2(new_n527), .A3(new_n560), .ZN(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n634), .A2(new_n644), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(KEYINPUT86), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n645), .B1(new_n629), .B2(new_n633), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT86), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n649), .A2(new_n650), .A3(new_n644), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n589), .B1(new_n648), .B2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT88), .ZN(new_n653));
  OAI21_X1  g0453(.A(KEYINPUT87), .B1(new_n552), .B2(new_n554), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n553), .A2(G179), .A3(new_n437), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT87), .ZN(new_n656));
  OAI211_X1 g0456(.A(new_n655), .B(new_n656), .C1(new_n559), .C2(new_n306), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n654), .A2(new_n542), .A3(new_n657), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n658), .B1(new_n629), .B2(new_n633), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n653), .B1(new_n659), .B2(KEYINPUT26), .ZN(new_n660));
  AND3_X1   g0460(.A1(new_n654), .A2(new_n542), .A3(new_n657), .ZN(new_n661));
  NOR3_X1   g0461(.A1(new_n628), .A2(new_n589), .A3(new_n617), .ZN(new_n662));
  AOI21_X1  g0462(.A(KEYINPUT84), .B1(new_n631), .B2(new_n632), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n661), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT26), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n664), .A2(KEYINPUT88), .A3(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n554), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n557), .B1(new_n667), .B2(new_n655), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n601), .A2(KEYINPUT26), .A3(new_n668), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n660), .A2(new_n666), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n652), .A2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n616), .B1(new_n431), .B2(new_n672), .ZN(G369));
  NAND3_X1  g0473(.A1(new_n266), .A2(new_n219), .A3(G13), .ZN(new_n674));
  XNOR2_X1  g0474(.A(new_n674), .B(KEYINPUT90), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT27), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(G213), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n675), .A2(new_n676), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(G343), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n684), .A2(new_n475), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT91), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n685), .B1(new_n485), .B2(new_n686), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n687), .B1(new_n686), .B2(new_n485), .ZN(new_n688));
  INV_X1    g0488(.A(new_n474), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(new_n685), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n522), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n528), .B1(new_n692), .B2(new_n684), .ZN(new_n693));
  OR2_X1    g0493(.A1(new_n523), .A2(new_n684), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n691), .A2(G330), .A3(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n474), .A2(new_n683), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n528), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n641), .A2(new_n643), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(new_n684), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n696), .A2(new_n702), .ZN(G399));
  INV_X1    g0503(.A(new_n215), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n704), .A2(G41), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NOR3_X1   g0506(.A1(new_n211), .A2(G87), .A3(G116), .ZN(new_n707));
  AND3_X1   g0507(.A1(new_n706), .A2(G1), .A3(new_n707), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n708), .B1(new_n221), .B2(new_n705), .ZN(new_n709));
  XOR2_X1   g0509(.A(new_n709), .B(KEYINPUT28), .Z(new_n710));
  AND3_X1   g0510(.A1(new_n660), .A2(new_n666), .A3(new_n669), .ZN(new_n711));
  AND4_X1   g0511(.A1(new_n650), .A2(new_n634), .A3(new_n644), .A4(new_n646), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n650), .B1(new_n649), .B2(new_n644), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n632), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n684), .B1(new_n711), .B2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT29), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n715), .A2(KEYINPUT93), .A3(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT93), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n683), .B1(new_n652), .B2(new_n670), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n718), .B1(new_n719), .B2(KEYINPUT29), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n717), .A2(new_n720), .ZN(new_n721));
  OR2_X1    g0521(.A1(new_n561), .A2(KEYINPUT95), .ZN(new_n722));
  INV_X1    g0522(.A(new_n527), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n723), .B1(new_n523), .B2(new_n474), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n561), .A2(KEYINPUT95), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n722), .A2(new_n724), .A3(new_n634), .A4(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n600), .A2(new_n592), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n668), .A2(new_n665), .A3(new_n727), .A4(new_n632), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(new_n632), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n729), .B1(new_n664), .B2(KEYINPUT26), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT94), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n726), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  OAI211_X1 g0532(.A(new_n632), .B(new_n728), .C1(new_n659), .C2(new_n665), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n733), .A2(KEYINPUT94), .ZN(new_n734));
  OAI211_X1 g0534(.A(KEYINPUT29), .B(new_n684), .C1(new_n732), .C2(new_n734), .ZN(new_n735));
  AND2_X1   g0535(.A1(new_n721), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n444), .A2(new_n308), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n524), .A2(new_n577), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n737), .A2(new_n738), .A3(new_n553), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT30), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n444), .A2(new_n524), .A3(new_n308), .A4(new_n577), .ZN(new_n741));
  OAI22_X1  g0541(.A1(new_n739), .A2(new_n740), .B1(new_n559), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n739), .A2(new_n740), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT92), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n739), .A2(KEYINPUT92), .A3(new_n740), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n742), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT31), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  AOI22_X1  g0549(.A1(new_n602), .A2(KEYINPUT31), .B1(new_n749), .B2(new_n683), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n684), .A2(new_n748), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n742), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n752), .B1(new_n753), .B2(new_n743), .ZN(new_n754));
  OAI21_X1  g0554(.A(G330), .B1(new_n750), .B2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n736), .A2(new_n756), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n710), .B1(new_n757), .B2(G1), .ZN(G364));
  NAND2_X1  g0558(.A1(new_n308), .A2(G200), .ZN(new_n759));
  INV_X1    g0559(.A(KEYINPUT98), .ZN(new_n760));
  XNOR2_X1  g0560(.A(new_n759), .B(new_n760), .ZN(new_n761));
  NOR3_X1   g0561(.A1(new_n761), .A2(new_n219), .A3(new_n299), .ZN(new_n762));
  OR2_X1    g0562(.A1(new_n762), .A2(KEYINPUT99), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n762), .A2(KEYINPUT99), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(G87), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n219), .A2(G190), .ZN(new_n768));
  NOR2_X1   g0568(.A1(G179), .A2(G200), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(G159), .ZN(new_n772));
  XNOR2_X1  g0572(.A(new_n772), .B(KEYINPUT32), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n219), .B1(new_n769), .B2(G190), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n773), .B1(G97), .B2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n219), .A2(new_n308), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR3_X1   g0578(.A1(new_n778), .A2(G190), .A3(G200), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NOR3_X1   g0580(.A1(new_n778), .A2(new_n299), .A3(G200), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  OAI221_X1 g0582(.A(new_n278), .B1(new_n780), .B2(new_n281), .C1(new_n399), .C2(new_n782), .ZN(new_n783));
  NOR3_X1   g0583(.A1(new_n761), .A2(new_n219), .A3(G190), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n783), .B1(G107), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n777), .A2(G200), .ZN(new_n786));
  INV_X1    g0586(.A(KEYINPUT97), .ZN(new_n787));
  XNOR2_X1  g0587(.A(new_n786), .B(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n788), .A2(new_n299), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n788), .A2(G190), .ZN(new_n790));
  AOI22_X1  g0590(.A1(G50), .A2(new_n789), .B1(new_n790), .B2(G68), .ZN(new_n791));
  NAND4_X1  g0591(.A1(new_n767), .A2(new_n776), .A3(new_n785), .A4(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(G294), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n774), .A2(new_n793), .ZN(new_n794));
  AOI22_X1  g0594(.A1(new_n779), .A2(G311), .B1(G329), .B2(new_n771), .ZN(new_n795));
  INV_X1    g0595(.A(G322), .ZN(new_n796));
  OAI211_X1 g0596(.A(new_n795), .B(new_n384), .C1(new_n796), .C2(new_n782), .ZN(new_n797));
  AOI211_X1 g0597(.A(new_n794), .B(new_n797), .C1(G283), .C2(new_n784), .ZN(new_n798));
  INV_X1    g0598(.A(G303), .ZN(new_n799));
  INV_X1    g0599(.A(new_n790), .ZN(new_n800));
  XOR2_X1   g0600(.A(KEYINPUT33), .B(G317), .Z(new_n801));
  OAI221_X1 g0601(.A(new_n798), .B1(new_n799), .B2(new_n765), .C1(new_n800), .C2(new_n801), .ZN(new_n802));
  XNOR2_X1  g0602(.A(new_n789), .B(KEYINPUT100), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  AND2_X1   g0604(.A1(new_n804), .A2(G326), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n792), .B1(new_n802), .B2(new_n805), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n806), .B(KEYINPUT101), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n218), .B1(G20), .B2(new_n306), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  AND2_X1   g0609(.A1(new_n219), .A2(G13), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n266), .B1(new_n810), .B2(G45), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n705), .A2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n215), .A2(new_n278), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n815), .B1(G87), .B2(new_n211), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n250), .A2(new_n433), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n704), .A2(new_n278), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  AOI211_X1 g0619(.A(new_n817), .B(new_n819), .C1(new_n433), .C2(new_n221), .ZN(new_n820));
  AOI211_X1 g0620(.A(new_n816), .B(new_n820), .C1(new_n453), .C2(new_n704), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n822), .A2(KEYINPUT96), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(G13), .A2(G33), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n826), .A2(G20), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n827), .A2(new_n808), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n829), .B1(new_n822), .B2(KEYINPUT96), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n814), .B1(new_n824), .B2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n827), .ZN(new_n832));
  OAI211_X1 g0632(.A(new_n809), .B(new_n831), .C1(new_n691), .C2(new_n832), .ZN(new_n833));
  AND2_X1   g0633(.A1(new_n688), .A2(new_n690), .ZN(new_n834));
  INV_X1    g0634(.A(G330), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n836), .A2(new_n813), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n691), .A2(G330), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n833), .B1(new_n838), .B2(new_n839), .ZN(G396));
  AND2_X1   g0640(.A1(new_n370), .A2(new_n684), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n841), .B1(new_n711), .B2(new_n714), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n683), .A2(new_n357), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n366), .A2(new_n369), .A3(new_n843), .ZN(new_n844));
  NAND4_X1  g0644(.A1(new_n609), .A2(new_n357), .A3(new_n610), .A4(new_n683), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n842), .B1(new_n719), .B2(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n813), .B1(new_n847), .B2(new_n755), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n848), .B1(new_n755), .B2(new_n847), .ZN(new_n849));
  OR2_X1    g0649(.A1(new_n808), .A2(new_n825), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n813), .B1(G77), .B2(new_n850), .ZN(new_n851));
  AOI22_X1  g0651(.A1(G143), .A2(new_n781), .B1(new_n779), .B2(G159), .ZN(new_n852));
  INV_X1    g0652(.A(new_n789), .ZN(new_n853));
  INV_X1    g0653(.A(G137), .ZN(new_n854));
  INV_X1    g0654(.A(G150), .ZN(new_n855));
  OAI221_X1 g0655(.A(new_n852), .B1(new_n853), .B2(new_n854), .C1(new_n855), .C2(new_n800), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT34), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(G132), .ZN(new_n859));
  OAI221_X1 g0659(.A(new_n278), .B1(new_n770), .B2(new_n859), .C1(new_n399), .C2(new_n774), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n860), .B1(new_n784), .B2(G68), .ZN(new_n861));
  OAI211_X1 g0661(.A(new_n858), .B(new_n861), .C1(new_n207), .C2(new_n765), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n856), .A2(new_n857), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n784), .A2(G87), .ZN(new_n864));
  INV_X1    g0664(.A(G311), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n864), .B1(new_n865), .B2(new_n770), .ZN(new_n866));
  XOR2_X1   g0666(.A(new_n866), .B(KEYINPUT103), .Z(new_n867));
  OAI221_X1 g0667(.A(new_n384), .B1(new_n774), .B2(new_n446), .C1(new_n782), .C2(new_n793), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n868), .B1(new_n789), .B2(G303), .ZN(new_n869));
  OAI211_X1 g0669(.A(new_n867), .B(new_n869), .C1(new_n359), .C2(new_n765), .ZN(new_n870));
  AOI22_X1  g0670(.A1(new_n790), .A2(G283), .B1(G116), .B2(new_n779), .ZN(new_n871));
  XOR2_X1   g0671(.A(new_n871), .B(KEYINPUT102), .Z(new_n872));
  OAI22_X1  g0672(.A1(new_n862), .A2(new_n863), .B1(new_n870), .B2(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n851), .B1(new_n873), .B2(new_n808), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n874), .B1(new_n846), .B2(new_n826), .ZN(new_n875));
  AND3_X1   g0675(.A1(new_n849), .A2(KEYINPUT104), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g0676(.A(KEYINPUT104), .B1(new_n849), .B2(new_n875), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(new_n878), .ZN(G384));
  OR2_X1    g0679(.A1(new_n533), .A2(KEYINPUT35), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n533), .A2(KEYINPUT35), .ZN(new_n881));
  NAND4_X1  g0681(.A1(new_n880), .A2(G116), .A3(new_n220), .A4(new_n881), .ZN(new_n882));
  XOR2_X1   g0682(.A(new_n882), .B(KEYINPUT36), .Z(new_n883));
  NAND3_X1  g0683(.A1(new_n221), .A2(G77), .A3(new_n393), .ZN(new_n884));
  AOI211_X1 g0684(.A(new_n266), .B(G13), .C1(new_n884), .C2(new_n246), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n735), .A2(new_n430), .ZN(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(KEYINPUT93), .B1(new_n715), .B2(new_n716), .ZN(new_n889));
  NOR3_X1   g0689(.A1(new_n719), .A2(new_n718), .A3(KEYINPUT29), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n888), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(KEYINPUT107), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT107), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n721), .A2(new_n893), .A3(new_n888), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(new_n616), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n683), .A2(new_n325), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n344), .A2(new_n348), .A3(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n897), .B1(new_n344), .B2(new_n348), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n369), .A2(new_n683), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n901), .B1(new_n842), .B2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT38), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n397), .A2(new_n408), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(new_n680), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n402), .A2(new_n403), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(KEYINPUT74), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(new_n405), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n390), .A2(new_n395), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n253), .B1(new_n911), .B2(new_n372), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n910), .B1(new_n912), .B2(new_n396), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n604), .B1(new_n913), .B2(new_n423), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n914), .B1(new_n605), .B2(KEYINPUT75), .ZN(new_n915));
  INV_X1    g0715(.A(new_n428), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n907), .B1(new_n917), .B2(new_n420), .ZN(new_n918));
  INV_X1    g0718(.A(new_n424), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n919), .A2(new_n907), .A3(new_n419), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n681), .B1(new_n397), .B2(new_n408), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT105), .ZN(new_n922));
  OAI21_X1  g0722(.A(KEYINPUT37), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n920), .B(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n905), .B1(new_n918), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n429), .A2(new_n921), .ZN(new_n926));
  INV_X1    g0726(.A(new_n923), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n927), .B(new_n920), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n926), .A2(KEYINPUT38), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n925), .A2(new_n929), .ZN(new_n930));
  AOI22_X1  g0730(.A1(new_n904), .A2(new_n930), .B1(new_n607), .B2(new_n681), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT39), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT37), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n920), .B(new_n933), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n907), .B1(new_n606), .B2(new_n420), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n905), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  AND3_X1   g0736(.A1(new_n929), .A2(new_n932), .A3(new_n936), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n932), .B1(new_n925), .B2(new_n929), .ZN(new_n938));
  OAI21_X1  g0738(.A(KEYINPUT106), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NOR3_X1   g0739(.A1(new_n918), .A2(new_n924), .A3(new_n905), .ZN(new_n940));
  AOI21_X1  g0740(.A(KEYINPUT38), .B1(new_n926), .B2(new_n928), .ZN(new_n941));
  OAI21_X1  g0741(.A(KEYINPUT39), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT106), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n929), .A2(new_n932), .A3(new_n936), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n942), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n344), .A2(new_n683), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n939), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n931), .A2(new_n947), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n896), .B(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n929), .A2(new_n936), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(new_n846), .ZN(new_n952));
  INV_X1    g0752(.A(new_n900), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n952), .B1(new_n953), .B2(new_n898), .ZN(new_n954));
  OAI21_X1  g0754(.A(KEYINPUT108), .B1(new_n747), .B2(new_n752), .ZN(new_n955));
  INV_X1    g0755(.A(new_n746), .ZN(new_n956));
  AOI21_X1  g0756(.A(KEYINPUT92), .B1(new_n739), .B2(new_n740), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n753), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT108), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n958), .A2(new_n959), .A3(new_n751), .ZN(new_n960));
  AND2_X1   g0760(.A1(new_n955), .A2(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n954), .B1(new_n961), .B2(new_n750), .ZN(new_n962));
  OAI21_X1  g0762(.A(KEYINPUT40), .B1(new_n951), .B2(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n846), .B1(new_n899), .B2(new_n900), .ZN(new_n964));
  AND2_X1   g0764(.A1(new_n478), .A2(new_n484), .ZN(new_n965));
  NAND4_X1  g0765(.A1(new_n562), .A2(new_n601), .A3(new_n527), .A4(new_n523), .ZN(new_n966));
  OAI21_X1  g0766(.A(KEYINPUT31), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(new_n749), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n967), .B1(new_n968), .B2(new_n684), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n955), .A2(new_n960), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n964), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  AOI21_X1  g0771(.A(KEYINPUT40), .B1(new_n925), .B2(new_n929), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n963), .A2(new_n973), .ZN(new_n974));
  OAI211_X1 g0774(.A(new_n974), .B(new_n430), .C1(new_n750), .C2(new_n961), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n971), .A2(new_n950), .ZN(new_n976));
  AOI22_X1  g0776(.A1(new_n976), .A2(KEYINPUT40), .B1(new_n971), .B2(new_n972), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n961), .A2(new_n750), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n977), .B1(new_n431), .B2(new_n978), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n975), .A2(G330), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n949), .A2(new_n980), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n981), .B1(new_n266), .B2(new_n810), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n949), .A2(new_n980), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n886), .B1(new_n982), .B2(new_n983), .ZN(G367));
  NAND2_X1  g0784(.A1(new_n818), .A2(new_n241), .ZN(new_n985));
  INV_X1    g0785(.A(new_n353), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n829), .B1(new_n704), .B2(new_n986), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n814), .B1(new_n985), .B2(new_n987), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n684), .A2(new_n630), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n989), .B1(new_n629), .B2(new_n633), .ZN(new_n990));
  NOR3_X1   g0790(.A1(new_n630), .A2(new_n632), .A3(new_n684), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n766), .A2(G116), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT46), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(KEYINPUT112), .ZN(new_n997));
  INV_X1    g0797(.A(new_n784), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n998), .A2(new_n446), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n278), .B1(new_n779), .B2(G283), .ZN(new_n1000));
  XOR2_X1   g0800(.A(KEYINPUT113), .B(G317), .Z(new_n1001));
  OAI221_X1 g0801(.A(new_n1000), .B1(new_n782), .B2(new_n799), .C1(new_n770), .C2(new_n1001), .ZN(new_n1002));
  AOI211_X1 g0802(.A(new_n999), .B(new_n1002), .C1(G107), .C2(new_n775), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n1003), .B1(new_n793), .B2(new_n800), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n994), .A2(new_n995), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  OAI211_X1 g0806(.A(new_n997), .B(new_n1006), .C1(new_n865), .C2(new_n803), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(KEYINPUT114), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n765), .A2(new_n399), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n782), .A2(new_n855), .B1(new_n780), .B2(new_n207), .ZN(new_n1010));
  AOI211_X1 g0810(.A(new_n384), .B(new_n1010), .C1(G137), .C2(new_n771), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n790), .A2(G159), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n784), .A2(G77), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n774), .A2(new_n203), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n1014), .ZN(new_n1015));
  NAND4_X1  g0815(.A1(new_n1011), .A2(new_n1012), .A3(new_n1013), .A4(new_n1015), .ZN(new_n1016));
  AOI211_X1 g0816(.A(new_n1009), .B(new_n1016), .C1(G143), .C2(new_n804), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n1008), .A2(new_n1017), .ZN(new_n1018));
  AND2_X1   g0818(.A1(new_n1018), .A2(KEYINPUT47), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n808), .B1(new_n1018), .B2(KEYINPUT47), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n988), .B1(new_n993), .B2(new_n832), .C1(new_n1019), .C2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n683), .A2(new_n542), .ZN(new_n1022));
  AND3_X1   g0822(.A1(new_n722), .A2(new_n725), .A3(new_n1022), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n1023), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n658), .A2(new_n684), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n1025), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1024), .A2(new_n701), .A3(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT44), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1030), .A2(KEYINPUT44), .A3(new_n701), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT45), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n1030), .B2(new_n701), .ZN(new_n1034));
  OAI211_X1 g0834(.A(new_n702), .B(KEYINPUT45), .C1(new_n1023), .C2(new_n1025), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1032), .A2(new_n696), .A3(new_n1036), .ZN(new_n1037));
  INV_X1    g0837(.A(KEYINPUT111), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n696), .B1(new_n1032), .B2(new_n1036), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1040), .A2(new_n1038), .A3(new_n1037), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n698), .B1(new_n695), .B2(new_n697), .ZN(new_n1045));
  XOR2_X1   g0845(.A(new_n836), .B(new_n1045), .Z(new_n1046));
  OAI21_X1  g0846(.A(new_n757), .B1(new_n1044), .B2(new_n1046), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(KEYINPUT110), .B(KEYINPUT41), .ZN(new_n1048));
  XOR2_X1   g0848(.A(new_n705), .B(new_n1048), .Z(new_n1049));
  AOI21_X1  g0849(.A(new_n812), .B1(new_n1047), .B2(new_n1049), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n1030), .A2(new_n698), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT42), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n993), .A2(KEYINPUT43), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n555), .B1(new_n1030), .B2(new_n523), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1054), .A2(new_n684), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1052), .A2(new_n1053), .A3(new_n1055), .ZN(new_n1056));
  INV_X1    g0856(.A(KEYINPUT109), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  NAND4_X1  g0858(.A1(new_n1052), .A2(new_n1055), .A3(KEYINPUT109), .A4(new_n1053), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1052), .A2(new_n1055), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n992), .B(KEYINPUT43), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1060), .A2(new_n1063), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n696), .A2(new_n1030), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1064), .A2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1060), .A2(new_n1065), .A3(new_n1063), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1021), .B1(new_n1050), .B2(new_n1069), .ZN(G387));
  NAND2_X1  g0870(.A1(new_n351), .A2(new_n207), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT50), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n433), .B1(new_n203), .B2(new_n281), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1073), .B1(new_n707), .B2(KEYINPUT115), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1074), .B1(KEYINPUT115), .B2(new_n707), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n818), .B1(new_n1072), .B2(new_n1075), .C1(new_n238), .C2(new_n433), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n1076), .B1(G107), .B2(new_n215), .C1(new_n707), .C2(new_n815), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1077), .A2(new_n828), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1078), .A2(new_n813), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n695), .A2(new_n832), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n781), .A2(G50), .B1(G150), .B2(new_n771), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n1081), .B(new_n278), .C1(new_n203), .C2(new_n780), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n774), .A2(new_n353), .ZN(new_n1083));
  NOR3_X1   g0883(.A1(new_n999), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(G159), .A2(new_n789), .B1(new_n790), .B2(new_n260), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n1084), .B(new_n1085), .C1(new_n281), .C2(new_n765), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n782), .A2(new_n1001), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n780), .A2(new_n799), .ZN(new_n1088));
  AOI211_X1 g0888(.A(new_n1087), .B(new_n1088), .C1(G311), .C2(new_n790), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1089), .B1(new_n803), .B2(new_n796), .ZN(new_n1090));
  INV_X1    g0890(.A(KEYINPUT48), .ZN(new_n1091));
  OR2_X1    g0891(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(G283), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n765), .A2(new_n793), .B1(new_n1093), .B2(new_n774), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1094), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1092), .A2(KEYINPUT49), .A3(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n278), .B1(new_n771), .B2(G326), .ZN(new_n1097));
  OAI211_X1 g0897(.A(new_n1096), .B(new_n1097), .C1(new_n453), .C2(new_n998), .ZN(new_n1098));
  AOI21_X1  g0898(.A(KEYINPUT49), .B1(new_n1092), .B2(new_n1095), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1086), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  AOI211_X1 g0900(.A(new_n1079), .B(new_n1080), .C1(new_n1100), .C2(new_n808), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1046), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1101), .B1(new_n1102), .B2(new_n812), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n757), .A2(new_n1102), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(new_n705), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n757), .A2(new_n1102), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1103), .B1(new_n1105), .B2(new_n1106), .ZN(G393));
  AND2_X1   g0907(.A1(new_n1041), .A2(new_n1037), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1030), .A2(new_n827), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n819), .A2(new_n245), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n828), .B1(new_n215), .B2(new_n446), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n813), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n774), .A2(new_n453), .ZN(new_n1113));
  OAI221_X1 g0913(.A(new_n384), .B1(new_n796), .B2(new_n770), .C1(new_n780), .C2(new_n793), .ZN(new_n1114));
  AOI211_X1 g0914(.A(new_n1113), .B(new_n1114), .C1(G107), .C2(new_n784), .ZN(new_n1115));
  OAI221_X1 g0915(.A(new_n1115), .B1(new_n1093), .B2(new_n765), .C1(new_n799), .C2(new_n800), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n789), .A2(G317), .B1(G311), .B2(new_n781), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(new_n1117), .B(KEYINPUT52), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n384), .B1(new_n779), .B2(new_n351), .ZN(new_n1119));
  INV_X1    g0919(.A(G143), .ZN(new_n1120));
  OAI221_X1 g0920(.A(new_n1119), .B1(new_n281), .B2(new_n774), .C1(new_n1120), .C2(new_n770), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1121), .B1(G87), .B2(new_n784), .ZN(new_n1122));
  OAI221_X1 g0922(.A(new_n1122), .B1(new_n207), .B2(new_n800), .C1(new_n203), .C2(new_n765), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n789), .A2(G150), .B1(G159), .B2(new_n781), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(new_n1124), .B(KEYINPUT51), .ZN(new_n1125));
  OAI22_X1  g0925(.A1(new_n1116), .A2(new_n1118), .B1(new_n1123), .B2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1112), .B1(new_n1126), .B2(new_n808), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(new_n1108), .A2(new_n812), .B1(new_n1109), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  NOR3_X1   g0929(.A1(new_n1046), .A2(new_n736), .A3(new_n756), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1044), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n706), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1108), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1104), .A2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1129), .B1(new_n1132), .B2(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(G390));
  OAI21_X1  g0936(.A(KEYINPUT116), .B1(new_n904), .B2(new_n946), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n939), .A2(new_n945), .ZN(new_n1138));
  INV_X1    g0938(.A(KEYINPUT116), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n946), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n902), .B1(new_n671), .B2(new_n841), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n1139), .B(new_n1140), .C1(new_n1141), .C2(new_n901), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1137), .A2(new_n1138), .A3(new_n1142), .ZN(new_n1143));
  AND2_X1   g0943(.A1(new_n722), .A2(new_n725), .ZN(new_n1144));
  AND2_X1   g0944(.A1(new_n724), .A2(new_n634), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(new_n733), .A2(KEYINPUT94), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n730), .A2(new_n731), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n683), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n902), .B1(new_n1148), .B2(new_n846), .ZN(new_n1149));
  OAI211_X1 g0949(.A(new_n1140), .B(new_n950), .C1(new_n1149), .C2(new_n901), .ZN(new_n1150));
  OAI211_X1 g0950(.A(G330), .B(new_n846), .C1(new_n750), .C2(new_n754), .ZN(new_n1151));
  OR2_X1    g0951(.A1(new_n1151), .A2(new_n901), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1143), .A2(new_n1150), .A3(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n950), .A2(new_n1140), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1148), .A2(new_n846), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1155), .A2(new_n903), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n901), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1154), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1140), .B1(new_n1141), .B2(new_n901), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n1159), .A2(KEYINPUT116), .B1(new_n939), .B2(new_n945), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1158), .B1(new_n1160), .B2(new_n1142), .ZN(new_n1161));
  OAI21_X1  g0961(.A(G330), .B1(new_n961), .B2(new_n750), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1163), .A2(new_n954), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1153), .B1(new_n1161), .B2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1163), .A2(new_n430), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n901), .B1(new_n1162), .B2(new_n952), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1152), .A2(new_n1167), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n1163), .A2(new_n954), .B1(new_n901), .B2(new_n1151), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n1168), .A2(new_n1156), .B1(new_n1169), .B2(new_n1141), .ZN(new_n1170));
  NAND4_X1  g0970(.A1(new_n895), .A2(new_n616), .A3(new_n1166), .A4(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n706), .B1(new_n1165), .B2(new_n1171), .ZN(new_n1172));
  AOI211_X1 g0972(.A(KEYINPUT107), .B(new_n887), .C1(new_n720), .C2(new_n717), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n893), .B1(new_n721), .B2(new_n888), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n616), .B(new_n1166), .C1(new_n1173), .C2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1170), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1143), .A2(new_n1150), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1178), .A2(new_n954), .A3(new_n1163), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1177), .A2(new_n1153), .A3(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1172), .A2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1179), .A2(new_n812), .A3(new_n1153), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n813), .B1(new_n260), .B2(new_n850), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n784), .A2(G68), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(new_n781), .A2(G116), .B1(G294), .B2(new_n771), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n1185), .B(new_n384), .C1(new_n446), .C2(new_n780), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1186), .B1(G77), .B2(new_n775), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(G107), .A2(new_n790), .B1(new_n789), .B2(G283), .ZN(new_n1188));
  NAND4_X1  g0988(.A1(new_n767), .A2(new_n1184), .A3(new_n1187), .A4(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n766), .A2(G150), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(new_n1190), .B(KEYINPUT53), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(KEYINPUT54), .B(G143), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n790), .A2(G137), .B1(new_n779), .B2(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT117), .ZN(new_n1195));
  OR2_X1    g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n774), .A2(new_n377), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n771), .A2(G125), .ZN(new_n1199));
  OAI211_X1 g0999(.A(new_n278), .B(new_n1199), .C1(new_n782), .C2(new_n859), .ZN(new_n1200));
  AOI211_X1 g1000(.A(new_n1198), .B(new_n1200), .C1(G50), .C2(new_n784), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n789), .A2(G128), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n1196), .A2(new_n1197), .A3(new_n1201), .A4(new_n1202), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1189), .B1(new_n1191), .B2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1183), .B1(new_n1204), .B2(new_n808), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1138), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1205), .B1(new_n1206), .B2(new_n826), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1181), .A2(new_n1182), .A3(new_n1207), .ZN(G378));
  INV_X1    g1008(.A(KEYINPUT57), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n312), .B1(new_n302), .B2(new_n303), .ZN(new_n1210));
  XOR2_X1   g1010(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1211));
  NAND2_X1  g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n305), .A2(new_n681), .ZN(new_n1213));
  XNOR2_X1  g1013(.A(new_n1213), .B(KEYINPUT121), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1211), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n312), .B(new_n1215), .C1(new_n302), .C2(new_n303), .ZN(new_n1216));
  AND3_X1   g1016(.A1(new_n1212), .A2(new_n1214), .A3(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1214), .B1(new_n1212), .B2(new_n1216), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1220), .B1(new_n974), .B2(G330), .ZN(new_n1221));
  AOI211_X1 g1021(.A(new_n835), .B(new_n1219), .C1(new_n963), .C2(new_n973), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n948), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1219), .B1(new_n977), .B2(new_n835), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n973), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT40), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1226), .B1(new_n971), .B2(new_n950), .ZN(new_n1227));
  OAI211_X1 g1027(.A(new_n1220), .B(G330), .C1(new_n1225), .C2(new_n1227), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1224), .A2(new_n947), .A3(new_n1228), .A4(new_n931), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1209), .B1(new_n1223), .B2(new_n1229), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1165), .A2(new_n1171), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT123), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1175), .A2(new_n1232), .ZN(new_n1233));
  NAND4_X1  g1033(.A1(new_n895), .A2(KEYINPUT123), .A3(new_n616), .A4(new_n1166), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1230), .B1(new_n1231), .B2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(new_n705), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1223), .A2(new_n1229), .A3(KEYINPUT122), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT122), .ZN(new_n1239));
  OAI211_X1 g1039(.A(new_n1239), .B(new_n948), .C1(new_n1221), .C2(new_n1222), .ZN(new_n1240));
  AND2_X1   g1040(.A1(new_n1238), .A2(new_n1240), .ZN(new_n1241));
  OAI211_X1 g1041(.A(new_n1233), .B(new_n1234), .C1(new_n1165), .C2(new_n1171), .ZN(new_n1242));
  AOI21_X1  g1042(.A(KEYINPUT57), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1243));
  OR2_X1    g1043(.A1(new_n1237), .A2(new_n1243), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n813), .B1(G50), .B2(new_n850), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n1220), .A2(new_n826), .ZN(new_n1246));
  AOI211_X1 g1046(.A(G33), .B(G41), .C1(new_n771), .C2(G124), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1247), .B1(new_n998), .B2(new_n377), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(new_n789), .A2(G125), .B1(G150), .B2(new_n775), .ZN(new_n1249));
  XOR2_X1   g1049(.A(new_n1249), .B(KEYINPUT119), .Z(new_n1250));
  OAI21_X1  g1050(.A(KEYINPUT118), .B1(new_n765), .B2(new_n1192), .ZN(new_n1251));
  OR3_X1    g1051(.A1(new_n765), .A2(KEYINPUT118), .A3(new_n1192), .ZN(new_n1252));
  INV_X1    g1052(.A(G128), .ZN(new_n1253));
  OAI22_X1  g1053(.A1(new_n782), .A2(new_n1253), .B1(new_n780), .B2(new_n854), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1254), .B1(new_n790), .B2(G132), .ZN(new_n1255));
  AND4_X1   g1055(.A1(new_n1250), .A2(new_n1251), .A3(new_n1252), .A4(new_n1255), .ZN(new_n1256));
  XOR2_X1   g1056(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n1257));
  AOI21_X1  g1057(.A(new_n1248), .B1(new_n1256), .B2(new_n1257), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1258), .B1(new_n1256), .B2(new_n1257), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n784), .A2(new_n259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n384), .A2(new_n289), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1261), .B1(new_n781), .B2(G107), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(new_n779), .A2(new_n986), .B1(G283), .B2(new_n771), .ZN(new_n1263));
  AND4_X1   g1063(.A1(new_n1015), .A2(new_n1260), .A3(new_n1262), .A4(new_n1263), .ZN(new_n1264));
  AOI22_X1  g1064(.A1(G97), .A2(new_n790), .B1(new_n789), .B2(G116), .ZN(new_n1265));
  OAI211_X1 g1065(.A(new_n1264), .B(new_n1265), .C1(new_n281), .C2(new_n765), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT58), .ZN(new_n1267));
  OR2_X1    g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  OAI211_X1 g1068(.A(new_n1261), .B(new_n207), .C1(G33), .C2(G41), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1259), .A2(new_n1268), .A3(new_n1269), .A4(new_n1270), .ZN(new_n1271));
  AOI211_X1 g1071(.A(new_n1245), .B(new_n1246), .C1(new_n808), .C2(new_n1271), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1272), .B1(new_n1241), .B2(new_n812), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1244), .A2(new_n1273), .ZN(G375));
  NAND2_X1  g1074(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1275), .A2(new_n1171), .A3(new_n1049), .ZN(new_n1276));
  XOR2_X1   g1076(.A(new_n1276), .B(KEYINPUT124), .Z(new_n1277));
  NAND2_X1  g1077(.A1(new_n901), .A2(new_n825), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n813), .B1(G68), .B2(new_n850), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n766), .A2(G97), .ZN(new_n1280));
  AOI22_X1  g1080(.A1(G116), .A2(new_n790), .B1(new_n789), .B2(G294), .ZN(new_n1281));
  OAI22_X1  g1081(.A1(new_n782), .A2(new_n1093), .B1(new_n770), .B2(new_n799), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n384), .B1(new_n780), .B2(new_n359), .ZN(new_n1283));
  NOR3_X1   g1083(.A1(new_n1282), .A2(new_n1283), .A3(new_n1083), .ZN(new_n1284));
  NAND4_X1  g1084(.A1(new_n1280), .A2(new_n1281), .A3(new_n1013), .A4(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1260), .A2(new_n278), .ZN(new_n1286));
  XOR2_X1   g1086(.A(new_n1286), .B(KEYINPUT125), .Z(new_n1287));
  OAI21_X1  g1087(.A(new_n1287), .B1(new_n377), .B2(new_n765), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n774), .A2(new_n207), .ZN(new_n1289));
  OAI22_X1  g1089(.A1(new_n780), .A2(new_n855), .B1(new_n770), .B2(new_n1253), .ZN(new_n1290));
  AOI211_X1 g1090(.A(new_n1289), .B(new_n1290), .C1(G137), .C2(new_n781), .ZN(new_n1291));
  OAI221_X1 g1091(.A(new_n1291), .B1(new_n859), .B2(new_n853), .C1(new_n800), .C2(new_n1192), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1285), .B1(new_n1288), .B2(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1279), .B1(new_n1293), .B2(new_n808), .ZN(new_n1294));
  AOI22_X1  g1094(.A1(new_n1170), .A2(new_n812), .B1(new_n1278), .B2(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1277), .A2(new_n1295), .ZN(G381));
  NAND2_X1  g1096(.A1(new_n1135), .A2(new_n878), .ZN(new_n1297));
  NOR4_X1   g1097(.A1(new_n1297), .A2(G387), .A3(G396), .A4(G393), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1182), .A2(new_n1207), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1299), .B1(new_n1180), .B2(new_n1172), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1298), .A2(new_n1300), .ZN(new_n1301));
  OR3_X1    g1101(.A1(new_n1301), .A2(G375), .A3(G381), .ZN(G407));
  NAND2_X1  g1102(.A1(new_n682), .A2(G213), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1300), .A2(new_n1304), .ZN(new_n1305));
  OAI211_X1 g1105(.A(G407), .B(G213), .C1(G375), .C2(new_n1305), .ZN(G409));
  XNOR2_X1  g1106(.A(G393), .B(G396), .ZN(new_n1307));
  AND2_X1   g1107(.A1(G387), .A2(new_n1135), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(G387), .A2(new_n1135), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1307), .B1(new_n1308), .B2(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(G396), .ZN(new_n1311));
  XNOR2_X1  g1111(.A(G393), .B(new_n1311), .ZN(new_n1312));
  OR2_X1    g1112(.A1(new_n1050), .A2(new_n1069), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1313), .A2(G390), .A3(new_n1021), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(G387), .A2(new_n1135), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1312), .A2(new_n1314), .A3(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1310), .A2(new_n1316), .ZN(new_n1317));
  OAI211_X1 g1117(.A(G378), .B(new_n1273), .C1(new_n1237), .C2(new_n1243), .ZN(new_n1318));
  AND3_X1   g1118(.A1(new_n1241), .A2(new_n1242), .A3(new_n1049), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n811), .B1(new_n1223), .B2(new_n1229), .ZN(new_n1320));
  OR2_X1    g1120(.A1(new_n1320), .A2(new_n1272), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n1300), .B1(new_n1319), .B2(new_n1321), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1304), .B1(new_n1318), .B2(new_n1322), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1175), .A2(KEYINPUT60), .A3(new_n1176), .ZN(new_n1324));
  AND2_X1   g1124(.A1(new_n1324), .A2(new_n705), .ZN(new_n1325));
  OAI21_X1  g1125(.A(KEYINPUT60), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1326), .A2(new_n1275), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1325), .A2(new_n1327), .ZN(new_n1328));
  AOI21_X1  g1128(.A(G384), .B1(new_n1328), .B2(new_n1295), .ZN(new_n1329));
  INV_X1    g1129(.A(new_n1295), .ZN(new_n1330));
  AOI211_X1 g1130(.A(new_n878), .B(new_n1330), .C1(new_n1325), .C2(new_n1327), .ZN(new_n1331));
  NOR2_X1   g1131(.A1(new_n1329), .A2(new_n1331), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1323), .A2(new_n1332), .ZN(new_n1333));
  INV_X1    g1133(.A(KEYINPUT63), .ZN(new_n1334));
  AOI21_X1  g1134(.A(new_n1317), .B1(new_n1333), .B2(new_n1334), .ZN(new_n1335));
  INV_X1    g1135(.A(new_n1323), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1304), .A2(G2897), .ZN(new_n1337));
  INV_X1    g1137(.A(new_n1337), .ZN(new_n1338));
  OAI21_X1  g1138(.A(new_n1338), .B1(new_n1329), .B2(new_n1331), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1324), .A2(new_n705), .ZN(new_n1340));
  AOI21_X1  g1140(.A(new_n1340), .B1(new_n1275), .B2(new_n1326), .ZN(new_n1341));
  OAI21_X1  g1141(.A(new_n878), .B1(new_n1341), .B2(new_n1330), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1328), .A2(G384), .A3(new_n1295), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1342), .A2(new_n1343), .A3(new_n1337), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1339), .A2(new_n1344), .ZN(new_n1345));
  INV_X1    g1145(.A(new_n1345), .ZN(new_n1346));
  AOI21_X1  g1146(.A(KEYINPUT61), .B1(new_n1336), .B2(new_n1346), .ZN(new_n1347));
  NAND3_X1  g1147(.A1(new_n1323), .A2(KEYINPUT63), .A3(new_n1332), .ZN(new_n1348));
  NAND3_X1  g1148(.A1(new_n1335), .A2(new_n1347), .A3(new_n1348), .ZN(new_n1349));
  INV_X1    g1149(.A(KEYINPUT62), .ZN(new_n1350));
  AND3_X1   g1150(.A1(new_n1323), .A2(new_n1350), .A3(new_n1332), .ZN(new_n1351));
  INV_X1    g1151(.A(KEYINPUT61), .ZN(new_n1352));
  OAI21_X1  g1152(.A(new_n1352), .B1(new_n1323), .B2(new_n1345), .ZN(new_n1353));
  AOI21_X1  g1153(.A(new_n1350), .B1(new_n1323), .B2(new_n1332), .ZN(new_n1354));
  NOR3_X1   g1154(.A1(new_n1351), .A2(new_n1353), .A3(new_n1354), .ZN(new_n1355));
  AND2_X1   g1155(.A1(new_n1310), .A2(new_n1316), .ZN(new_n1356));
  OAI21_X1  g1156(.A(new_n1349), .B1(new_n1355), .B2(new_n1356), .ZN(G405));
  NAND2_X1  g1157(.A1(new_n1332), .A2(KEYINPUT126), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1358), .A2(KEYINPUT127), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1359), .A2(new_n1356), .ZN(new_n1360));
  NAND3_X1  g1160(.A1(new_n1317), .A2(KEYINPUT127), .A3(new_n1358), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(new_n1360), .A2(new_n1361), .ZN(new_n1362));
  AOI21_X1  g1162(.A(G378), .B1(new_n1244), .B2(new_n1273), .ZN(new_n1363));
  INV_X1    g1163(.A(new_n1318), .ZN(new_n1364));
  NOR2_X1   g1164(.A1(new_n1363), .A2(new_n1364), .ZN(new_n1365));
  INV_X1    g1165(.A(KEYINPUT127), .ZN(new_n1366));
  NAND2_X1  g1166(.A1(new_n1332), .A2(new_n1366), .ZN(new_n1367));
  NAND2_X1  g1167(.A1(new_n1365), .A2(new_n1367), .ZN(new_n1368));
  NAND2_X1  g1168(.A1(new_n1362), .A2(new_n1368), .ZN(new_n1369));
  NAND4_X1  g1169(.A1(new_n1360), .A2(new_n1367), .A3(new_n1365), .A4(new_n1361), .ZN(new_n1370));
  AND2_X1   g1170(.A1(new_n1369), .A2(new_n1370), .ZN(G402));
endmodule


