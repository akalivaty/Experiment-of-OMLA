//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 1 1 1 0 0 0 0 0 1 1 0 0 0 0 0 0 0 1 1 1 0 0 1 1 1 1 1 1 1 0 1 1 1 1 1 0 1 1 1 0 0 0 0 0 0 0 1 0 1 1 0 0 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:19 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n689,
    new_n690, new_n691, new_n692, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n769, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT75), .ZN(new_n190));
  XNOR2_X1  g004(.A(G125), .B(G140), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(KEYINPUT16), .ZN(new_n192));
  INV_X1    g006(.A(G125), .ZN(new_n193));
  OR3_X1    g007(.A1(new_n193), .A2(KEYINPUT16), .A3(G140), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G146), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n192), .A2(G146), .A3(new_n194), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G128), .ZN(new_n200));
  OAI211_X1 g014(.A(new_n200), .B(G119), .C1(KEYINPUT74), .C2(KEYINPUT23), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT23), .ZN(new_n202));
  INV_X1    g016(.A(G119), .ZN(new_n203));
  AOI21_X1  g017(.A(new_n202), .B1(new_n203), .B2(G128), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT74), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n205), .B1(new_n203), .B2(G128), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n201), .B1(new_n204), .B2(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G110), .ZN(new_n208));
  XOR2_X1   g022(.A(KEYINPUT24), .B(G110), .Z(new_n209));
  XNOR2_X1  g023(.A(G119), .B(G128), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n199), .A2(new_n208), .A3(new_n211), .ZN(new_n212));
  OAI22_X1  g026(.A1(new_n207), .A2(G110), .B1(new_n210), .B2(new_n209), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n191), .A2(new_n196), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n213), .A2(new_n198), .A3(new_n214), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n190), .B1(new_n212), .B2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(new_n216), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n212), .A2(new_n190), .A3(new_n215), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  XNOR2_X1  g033(.A(KEYINPUT22), .B(G137), .ZN(new_n220));
  INV_X1    g034(.A(G953), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n221), .A2(G221), .A3(G234), .ZN(new_n222));
  XNOR2_X1  g036(.A(new_n220), .B(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n219), .A2(new_n224), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n224), .B1(new_n212), .B2(new_n215), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  AOI21_X1  g042(.A(KEYINPUT25), .B1(new_n228), .B2(new_n188), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n226), .B1(new_n219), .B2(new_n224), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT25), .ZN(new_n231));
  NOR3_X1   g045(.A1(new_n230), .A2(new_n231), .A3(G902), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n189), .B1(new_n229), .B2(new_n232), .ZN(new_n233));
  NOR3_X1   g047(.A1(new_n230), .A2(G902), .A3(new_n189), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  AND2_X1   g049(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  OR2_X1    g051(.A1(KEYINPUT66), .A2(KEYINPUT1), .ZN(new_n238));
  NAND2_X1  g052(.A1(KEYINPUT66), .A2(KEYINPUT1), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n238), .A2(G128), .A3(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n196), .A2(G143), .ZN(new_n241));
  INV_X1    g055(.A(G143), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(G146), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  OAI21_X1  g058(.A(KEYINPUT67), .B1(new_n240), .B2(new_n244), .ZN(new_n245));
  AND2_X1   g059(.A1(KEYINPUT66), .A2(KEYINPUT1), .ZN(new_n246));
  NOR2_X1   g060(.A1(KEYINPUT66), .A2(KEYINPUT1), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  XNOR2_X1  g062(.A(G143), .B(G146), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT67), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n248), .A2(new_n249), .A3(new_n250), .A4(G128), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n245), .A2(new_n251), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n241), .B1(new_n246), .B2(new_n247), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G128), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(new_n244), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n252), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(G134), .ZN(new_n257));
  OAI21_X1  g071(.A(KEYINPUT11), .B1(new_n257), .B2(G137), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT11), .ZN(new_n259));
  INV_X1    g073(.A(G137), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n259), .A2(new_n260), .A3(G134), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n258), .A2(new_n261), .ZN(new_n262));
  AND2_X1   g076(.A1(KEYINPUT64), .A2(G131), .ZN(new_n263));
  NOR2_X1   g077(.A1(KEYINPUT64), .A2(G131), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n257), .A2(G137), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n262), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT65), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n268), .B1(new_n260), .B2(G134), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n260), .A2(G134), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n257), .A2(KEYINPUT65), .A3(G137), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n269), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(G131), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n267), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(KEYINPUT71), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT71), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n267), .A2(new_n273), .A3(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n256), .A2(new_n275), .A3(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT69), .ZN(new_n279));
  INV_X1    g093(.A(G116), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(KEYINPUT69), .A2(G116), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n281), .A2(G119), .A3(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n203), .A2(G116), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  XNOR2_X1  g099(.A(KEYINPUT2), .B(G113), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(new_n286), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n288), .A2(new_n283), .A3(new_n284), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(KEYINPUT0), .A2(G128), .ZN(new_n292));
  OR2_X1    g106(.A1(KEYINPUT0), .A2(G128), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n244), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n249), .A2(KEYINPUT0), .A3(G128), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(G131), .ZN(new_n298));
  AOI22_X1  g112(.A1(new_n258), .A2(new_n261), .B1(new_n257), .B2(G137), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n267), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT70), .ZN(new_n301));
  AND3_X1   g115(.A1(new_n297), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n301), .B1(new_n297), .B2(new_n300), .ZN(new_n303));
  OAI211_X1 g117(.A(new_n278), .B(new_n291), .C1(new_n302), .C2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT72), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n297), .A2(new_n300), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(KEYINPUT70), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n297), .A2(new_n300), .A3(new_n301), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND4_X1  g124(.A1(new_n310), .A2(KEYINPUT72), .A3(new_n291), .A4(new_n278), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n306), .A2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(new_n274), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n256), .A2(KEYINPUT68), .A3(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT68), .ZN(new_n315));
  AOI22_X1  g129(.A1(new_n245), .A2(new_n251), .B1(new_n254), .B2(new_n244), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n315), .B1(new_n316), .B2(new_n274), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n314), .A2(new_n317), .A3(new_n307), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT30), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  OAI211_X1 g134(.A(new_n278), .B(KEYINPUT30), .C1(new_n302), .C2(new_n303), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n320), .A2(new_n290), .A3(new_n321), .ZN(new_n322));
  NOR2_X1   g136(.A1(G237), .A2(G953), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G210), .ZN(new_n324));
  XOR2_X1   g138(.A(new_n324), .B(KEYINPUT27), .Z(new_n325));
  XNOR2_X1  g139(.A(KEYINPUT26), .B(G101), .ZN(new_n326));
  XOR2_X1   g140(.A(new_n325), .B(new_n326), .Z(new_n327));
  NAND3_X1  g141(.A1(new_n312), .A2(new_n322), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(KEYINPUT31), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT31), .ZN(new_n330));
  NAND4_X1  g144(.A1(new_n312), .A2(new_n322), .A3(new_n330), .A4(new_n327), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n290), .B1(new_n300), .B2(new_n297), .ZN(new_n332));
  AOI21_X1  g146(.A(KEYINPUT28), .B1(new_n278), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n318), .A2(new_n290), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n312), .A2(new_n334), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n333), .B1(new_n335), .B2(KEYINPUT28), .ZN(new_n336));
  OAI211_X1 g150(.A(new_n329), .B(new_n331), .C1(new_n336), .C2(new_n327), .ZN(new_n337));
  NOR2_X1   g151(.A1(G472), .A2(G902), .ZN(new_n338));
  AOI211_X1 g152(.A(KEYINPUT73), .B(KEYINPUT32), .C1(new_n337), .C2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT73), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n335), .A2(KEYINPUT28), .ZN(new_n341));
  INV_X1    g155(.A(new_n333), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n327), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n329), .A2(new_n331), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n338), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT32), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n340), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n339), .A2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(new_n338), .ZN(new_n349));
  AND2_X1   g163(.A1(new_n329), .A2(new_n331), .ZN(new_n350));
  INV_X1    g164(.A(new_n327), .ZN(new_n351));
  AOI22_X1  g165(.A1(new_n306), .A2(new_n311), .B1(new_n290), .B2(new_n318), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT28), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n351), .B1(new_n354), .B2(new_n333), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n349), .B1(new_n350), .B2(new_n355), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n342), .B(new_n327), .C1(new_n352), .C2(new_n353), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n327), .B1(new_n312), .B2(new_n322), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT29), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n357), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n310), .A2(new_n278), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(new_n290), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n312), .A2(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n333), .B1(new_n364), .B2(KEYINPUT28), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n351), .A2(new_n360), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n361), .A2(new_n367), .A3(new_n188), .ZN(new_n368));
  AOI22_X1  g182(.A1(new_n356), .A2(KEYINPUT32), .B1(new_n368), .B2(G472), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n237), .B1(new_n348), .B2(new_n369), .ZN(new_n370));
  XNOR2_X1  g184(.A(KEYINPUT9), .B(G234), .ZN(new_n371));
  NOR3_X1   g185(.A1(new_n371), .A2(new_n187), .A3(G953), .ZN(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT89), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n374), .B1(new_n200), .B2(G143), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n242), .A2(KEYINPUT89), .A3(G128), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n377), .B1(G128), .B2(new_n242), .ZN(new_n378));
  XNOR2_X1  g192(.A(new_n378), .B(G134), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n281), .A2(G122), .A3(new_n282), .ZN(new_n380));
  INV_X1    g194(.A(G122), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(KEYINPUT88), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT88), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(G122), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  AOI22_X1  g199(.A1(new_n380), .A2(KEYINPUT14), .B1(new_n385), .B2(G116), .ZN(new_n386));
  OR2_X1    g200(.A1(new_n380), .A2(KEYINPUT14), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(G107), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n385), .A2(G116), .ZN(new_n390));
  INV_X1    g204(.A(G107), .ZN(new_n391));
  AND3_X1   g205(.A1(new_n390), .A2(new_n391), .A3(new_n380), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n379), .A2(new_n389), .A3(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n391), .B1(new_n390), .B2(new_n380), .ZN(new_n396));
  OAI22_X1  g210(.A1(new_n392), .A2(new_n396), .B1(G134), .B2(new_n378), .ZN(new_n397));
  AOI21_X1  g211(.A(KEYINPUT13), .B1(new_n375), .B2(new_n376), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT90), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n242), .A2(G128), .ZN(new_n400));
  OR3_X1    g214(.A1(new_n398), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n399), .B1(new_n398), .B2(new_n400), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n375), .A2(KEYINPUT13), .A3(new_n376), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT91), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  OR2_X1    g219(.A1(new_n403), .A2(new_n404), .ZN(new_n406));
  NAND4_X1  g220(.A1(new_n401), .A2(new_n402), .A3(new_n405), .A4(new_n406), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n397), .B1(new_n407), .B2(G134), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n373), .B1(new_n395), .B2(new_n408), .ZN(new_n409));
  AND2_X1   g223(.A1(new_n407), .A2(G134), .ZN(new_n410));
  OAI211_X1 g224(.A(new_n394), .B(new_n372), .C1(new_n410), .C2(new_n397), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n409), .A2(new_n411), .A3(KEYINPUT92), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT92), .ZN(new_n413));
  OAI211_X1 g227(.A(new_n413), .B(new_n373), .C1(new_n395), .C2(new_n408), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n412), .A2(new_n188), .A3(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(G478), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n416), .A2(KEYINPUT15), .ZN(new_n417));
  XNOR2_X1  g231(.A(new_n415), .B(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(G237), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n419), .A2(new_n221), .A3(G214), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(new_n242), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n323), .A2(G143), .A3(G214), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n265), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n423), .A2(KEYINPUT17), .A3(new_n424), .ZN(new_n425));
  AND3_X1   g239(.A1(new_n197), .A2(new_n425), .A3(new_n198), .ZN(new_n426));
  OAI21_X1  g240(.A(KEYINPUT85), .B1(new_n423), .B2(new_n424), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT17), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n423), .A2(new_n424), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT85), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n421), .A2(new_n430), .A3(new_n265), .A4(new_n422), .ZN(new_n431));
  NAND4_X1  g245(.A1(new_n427), .A2(new_n428), .A3(new_n429), .A4(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n426), .A2(new_n432), .ZN(new_n433));
  XNOR2_X1  g247(.A(G113), .B(G122), .ZN(new_n434));
  XNOR2_X1  g248(.A(new_n434), .B(G104), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n423), .A2(KEYINPUT18), .A3(G131), .ZN(new_n437));
  XNOR2_X1  g251(.A(new_n191), .B(new_n196), .ZN(new_n438));
  NAND2_X1  g252(.A1(KEYINPUT18), .A2(G131), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n421), .A2(new_n422), .A3(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n437), .A2(new_n438), .A3(new_n440), .ZN(new_n441));
  AND3_X1   g255(.A1(new_n433), .A2(new_n436), .A3(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n436), .B1(new_n433), .B2(new_n441), .ZN(new_n443));
  OR2_X1    g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(new_n188), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(G475), .ZN(new_n446));
  NOR2_X1   g260(.A1(G475), .A2(G902), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n427), .A2(new_n429), .A3(new_n431), .ZN(new_n449));
  NAND2_X1  g263(.A1(KEYINPUT86), .A2(KEYINPUT19), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n191), .A2(new_n450), .ZN(new_n451));
  XOR2_X1   g265(.A(KEYINPUT86), .B(KEYINPUT19), .Z(new_n452));
  OAI21_X1  g266(.A(new_n451), .B1(new_n191), .B2(new_n452), .ZN(new_n453));
  OR2_X1    g267(.A1(new_n453), .A2(G146), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n449), .A2(new_n454), .A3(new_n198), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(new_n441), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(new_n435), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n433), .A2(new_n436), .A3(new_n441), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n448), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT20), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n459), .A2(KEYINPUT87), .A3(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n436), .B1(new_n455), .B2(new_n441), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n447), .B1(new_n442), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(KEYINPUT20), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g279(.A(KEYINPUT87), .B1(new_n459), .B2(new_n460), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n446), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n221), .A2(G952), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n468), .B1(G234), .B2(G237), .ZN(new_n469));
  AOI211_X1 g283(.A(new_n188), .B(new_n221), .C1(G234), .C2(G237), .ZN(new_n470));
  XNOR2_X1  g284(.A(KEYINPUT21), .B(G898), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n469), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NOR3_X1   g286(.A1(new_n418), .A2(new_n467), .A3(new_n472), .ZN(new_n473));
  OAI21_X1  g287(.A(G210), .B1(G237), .B2(G902), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT81), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n283), .A2(KEYINPUT5), .A3(new_n284), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n284), .A2(KEYINPUT5), .ZN(new_n477));
  INV_X1    g291(.A(G113), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n476), .A2(new_n479), .ZN(new_n480));
  AND2_X1   g294(.A1(new_n480), .A2(new_n289), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT3), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(KEYINPUT78), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n482), .A2(KEYINPUT78), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n391), .A2(G104), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(G101), .ZN(new_n487));
  INV_X1    g301(.A(G104), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(G107), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n482), .A2(new_n391), .A3(KEYINPUT78), .A4(G104), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n486), .A2(new_n487), .A3(new_n489), .A4(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT79), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n487), .B1(new_n485), .B2(new_n489), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  AND3_X1   g308(.A1(new_n491), .A2(new_n492), .A3(new_n494), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n492), .B1(new_n491), .B2(new_n494), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n481), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  XNOR2_X1  g311(.A(G110), .B(G122), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT78), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n499), .A2(KEYINPUT3), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n488), .A2(G107), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n499), .A2(KEYINPUT3), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n490), .A2(new_n489), .ZN(new_n504));
  OAI21_X1  g318(.A(G101), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n505), .A2(KEYINPUT4), .A3(new_n491), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT4), .ZN(new_n507));
  OAI211_X1 g321(.A(new_n507), .B(G101), .C1(new_n503), .C2(new_n504), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n506), .A2(new_n290), .A3(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n497), .A2(new_n498), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(KEYINPUT6), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n498), .B1(new_n497), .B2(new_n509), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n475), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n497), .A2(new_n509), .ZN(new_n514));
  INV_X1    g328(.A(new_n498), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n516), .A2(KEYINPUT81), .A3(KEYINPUT6), .A4(new_n510), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n513), .A2(new_n517), .ZN(new_n518));
  XOR2_X1   g332(.A(KEYINPUT82), .B(KEYINPUT6), .Z(new_n519));
  NOR2_X1   g333(.A1(new_n516), .A2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n316), .A2(new_n193), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n296), .A2(G125), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(G224), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n525), .A2(G953), .ZN(new_n526));
  XNOR2_X1  g340(.A(new_n524), .B(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n518), .A2(new_n521), .A3(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT83), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n520), .B1(new_n513), .B2(new_n517), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n531), .A2(KEYINPUT83), .A3(new_n527), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  OAI21_X1  g347(.A(KEYINPUT7), .B1(new_n525), .B2(G953), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n524), .A2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n534), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n522), .A2(new_n523), .A3(new_n536), .ZN(new_n537));
  AND2_X1   g351(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n480), .A2(new_n289), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n491), .A2(new_n494), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n497), .A2(new_n541), .ZN(new_n542));
  XOR2_X1   g356(.A(new_n498), .B(KEYINPUT8), .Z(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n538), .A2(KEYINPUT84), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(new_n510), .ZN(new_n547));
  AOI21_X1  g361(.A(KEYINPUT84), .B1(new_n538), .B2(new_n545), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n188), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n474), .B1(new_n533), .B2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(new_n474), .ZN(new_n552));
  AOI211_X1 g366(.A(new_n552), .B(new_n549), .C1(new_n530), .C2(new_n532), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  OAI21_X1  g368(.A(G214), .B1(G237), .B2(G902), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(G469), .ZN(new_n557));
  NOR3_X1   g371(.A1(new_n503), .A2(new_n504), .A3(G101), .ZN(new_n558));
  OAI21_X1  g372(.A(KEYINPUT79), .B1(new_n558), .B2(new_n493), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n491), .A2(new_n492), .A3(new_n494), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n561), .A2(KEYINPUT10), .A3(new_n256), .ZN(new_n562));
  INV_X1    g376(.A(new_n300), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT10), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT1), .ZN(new_n565));
  OAI22_X1  g379(.A1(new_n249), .A2(G128), .B1(new_n565), .B2(new_n243), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n566), .B1(new_n245), .B2(new_n251), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n564), .B1(new_n567), .B2(new_n540), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n506), .A2(new_n297), .A3(new_n508), .ZN(new_n569));
  NAND4_X1  g383(.A1(new_n562), .A2(new_n563), .A3(new_n568), .A4(new_n569), .ZN(new_n570));
  XNOR2_X1  g384(.A(G110), .B(G140), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n571), .B(KEYINPUT77), .ZN(new_n572));
  AND2_X1   g386(.A1(new_n221), .A2(G227), .ZN(new_n573));
  XOR2_X1   g387(.A(new_n572), .B(new_n573), .Z(new_n574));
  NAND2_X1  g388(.A1(new_n570), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n559), .A2(new_n316), .A3(new_n560), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(KEYINPUT80), .ZN(new_n577));
  OR2_X1    g391(.A1(new_n567), .A2(new_n540), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT80), .ZN(new_n579));
  NAND4_X1  g393(.A1(new_n559), .A2(new_n579), .A3(new_n316), .A4(new_n560), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n577), .A2(new_n578), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(new_n300), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT12), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n581), .A2(KEYINPUT12), .A3(new_n300), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n575), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n562), .A2(new_n568), .A3(new_n569), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(new_n300), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n574), .B1(new_n588), .B2(new_n570), .ZN(new_n589));
  OAI211_X1 g403(.A(new_n557), .B(new_n188), .C1(new_n586), .C2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n575), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(new_n588), .ZN(new_n592));
  INV_X1    g406(.A(new_n570), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n593), .B1(new_n584), .B2(new_n585), .ZN(new_n594));
  OAI211_X1 g408(.A(G469), .B(new_n592), .C1(new_n594), .C2(new_n574), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n557), .A2(new_n188), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n590), .A2(new_n595), .A3(new_n597), .ZN(new_n598));
  OAI21_X1  g412(.A(G221), .B1(new_n371), .B2(G902), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n599), .B(KEYINPUT76), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  NOR3_X1   g416(.A1(new_n554), .A2(new_n556), .A3(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n370), .A2(new_n473), .A3(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(KEYINPUT93), .B(G101), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n604), .B(new_n605), .ZN(G3));
  INV_X1    g420(.A(new_n602), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n337), .A2(new_n188), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n356), .B1(G472), .B2(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n607), .A2(new_n609), .A3(new_n236), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n610), .B(KEYINPUT94), .ZN(new_n611));
  INV_X1    g425(.A(new_n472), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT33), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n412), .A2(new_n613), .A3(new_n414), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n409), .A2(new_n411), .A3(KEYINPUT33), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n416), .A2(G902), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  XOR2_X1   g431(.A(KEYINPUT96), .B(G478), .Z(new_n618));
  NAND2_X1  g432(.A1(new_n415), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(new_n467), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT97), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n621), .B(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT95), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n556), .B1(new_n553), .B2(new_n624), .ZN(new_n625));
  AND4_X1   g439(.A1(KEYINPUT83), .A2(new_n518), .A3(new_n521), .A4(new_n527), .ZN(new_n626));
  AOI21_X1  g440(.A(KEYINPUT83), .B1(new_n531), .B2(new_n527), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n550), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(new_n552), .ZN(new_n629));
  OAI211_X1 g443(.A(new_n550), .B(new_n474), .C1(new_n626), .C2(new_n627), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n629), .A2(KEYINPUT95), .A3(new_n630), .ZN(new_n631));
  AND4_X1   g445(.A1(new_n612), .A2(new_n623), .A3(new_n625), .A4(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n611), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g448(.A(KEYINPUT34), .B(G104), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G6));
  NAND2_X1  g450(.A1(new_n459), .A2(new_n460), .ZN(new_n637));
  AOI22_X1  g451(.A1(new_n637), .A2(new_n464), .B1(new_n445), .B2(G475), .ZN(new_n638));
  AND2_X1   g452(.A1(new_n418), .A2(new_n638), .ZN(new_n639));
  AND4_X1   g453(.A1(new_n612), .A2(new_n625), .A3(new_n631), .A4(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n611), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(KEYINPUT35), .B(G107), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G9));
  OR2_X1    g458(.A1(new_n224), .A2(KEYINPUT36), .ZN(new_n645));
  OR2_X1    g459(.A1(new_n645), .A2(KEYINPUT98), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(KEYINPUT98), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n219), .A2(new_n648), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n189), .A2(G902), .ZN(new_n650));
  NAND4_X1  g464(.A1(new_n217), .A2(new_n218), .A3(new_n647), .A4(new_n646), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n649), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(KEYINPUT99), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n233), .A2(new_n653), .ZN(new_n654));
  AND2_X1   g468(.A1(new_n473), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n603), .A2(new_n609), .A3(new_n655), .ZN(new_n656));
  XOR2_X1   g470(.A(KEYINPUT37), .B(G110), .Z(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(G12));
  AOI21_X1  g472(.A(new_n602), .B1(new_n348), .B2(new_n369), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n555), .B1(new_n630), .B2(KEYINPUT95), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n660), .B1(new_n554), .B2(KEYINPUT95), .ZN(new_n661));
  INV_X1    g475(.A(G900), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n469), .B1(new_n470), .B2(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n418), .A2(new_n638), .A3(new_n664), .ZN(new_n665));
  OR2_X1    g479(.A1(new_n665), .A2(KEYINPUT100), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n665), .A2(KEYINPUT100), .ZN(new_n667));
  AND3_X1   g481(.A1(new_n666), .A2(new_n654), .A3(new_n667), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n659), .A2(new_n661), .A3(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(G128), .ZN(G30));
  XOR2_X1   g484(.A(KEYINPUT101), .B(KEYINPUT39), .Z(new_n671));
  XNOR2_X1  g485(.A(new_n663), .B(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n607), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g487(.A(new_n673), .B(KEYINPUT40), .Z(new_n674));
  INV_X1    g488(.A(G472), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n364), .A2(new_n327), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n676), .A2(G902), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n312), .A2(new_n322), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(new_n327), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n675), .B1(new_n677), .B2(new_n679), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n680), .B1(new_n356), .B2(KEYINPUT32), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n654), .B1(new_n348), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n629), .A2(new_n630), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(KEYINPUT38), .ZN(new_n684));
  AND2_X1   g498(.A1(new_n418), .A2(new_n467), .ZN(new_n685));
  AND2_X1   g499(.A1(new_n685), .A2(new_n555), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n674), .A2(new_n682), .A3(new_n684), .A4(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G143), .ZN(G45));
  NAND3_X1  g502(.A1(new_n620), .A2(new_n467), .A3(new_n664), .ZN(new_n689));
  INV_X1    g503(.A(new_n689), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n659), .A2(new_n661), .A3(new_n654), .A4(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(KEYINPUT102), .B(G146), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(G48));
  OR2_X1    g507(.A1(new_n586), .A2(new_n589), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n557), .B1(new_n694), .B2(new_n188), .ZN(new_n695));
  INV_X1    g509(.A(new_n590), .ZN(new_n696));
  NOR3_X1   g510(.A1(new_n695), .A2(new_n696), .A3(new_n600), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n632), .A2(new_n370), .A3(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(KEYINPUT41), .B(G113), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n698), .B(new_n699), .ZN(G15));
  NAND3_X1  g514(.A1(new_n640), .A2(new_n370), .A3(new_n697), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G116), .ZN(G18));
  OAI21_X1  g516(.A(KEYINPUT73), .B1(new_n356), .B2(KEYINPUT32), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n345), .A2(new_n340), .A3(new_n346), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n369), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  AND2_X1   g519(.A1(new_n705), .A2(new_n655), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n625), .A2(new_n631), .A3(new_n697), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G119), .ZN(G21));
  AND3_X1   g524(.A1(new_n625), .A2(new_n631), .A3(new_n685), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT103), .ZN(new_n712));
  OAI211_X1 g526(.A(new_n329), .B(new_n331), .C1(new_n365), .C2(new_n327), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(new_n338), .ZN(new_n714));
  AOI21_X1  g528(.A(G902), .B1(new_n350), .B2(new_n355), .ZN(new_n715));
  OAI211_X1 g529(.A(new_n236), .B(new_n714), .C1(new_n675), .C2(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n694), .A2(new_n188), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(G469), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n718), .A2(new_n612), .A3(new_n601), .A4(new_n590), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n716), .A2(new_n719), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n711), .A2(new_n712), .A3(new_n720), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n625), .A2(new_n631), .A3(new_n685), .ZN(new_n722));
  AOI22_X1  g536(.A1(new_n608), .A2(G472), .B1(new_n338), .B2(new_n713), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n697), .A2(new_n723), .A3(new_n236), .A4(new_n612), .ZN(new_n724));
  OAI21_X1  g538(.A(KEYINPUT103), .B1(new_n722), .B2(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n721), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G122), .ZN(G24));
  INV_X1    g541(.A(KEYINPUT104), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n689), .A2(new_n728), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n620), .A2(new_n467), .A3(KEYINPUT104), .A4(new_n664), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  OAI211_X1 g545(.A(new_n654), .B(new_n714), .C1(new_n715), .C2(new_n675), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT105), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n661), .A2(new_n733), .A3(new_n734), .A4(new_n697), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n723), .A2(new_n654), .A3(new_n729), .A4(new_n730), .ZN(new_n736));
  OAI21_X1  g550(.A(KEYINPUT105), .B1(new_n707), .B2(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G125), .ZN(G27));
  INV_X1    g553(.A(KEYINPUT108), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n629), .A2(new_n555), .A3(new_n630), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(KEYINPUT107), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT106), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n598), .A2(new_n743), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n590), .A2(new_n595), .A3(KEYINPUT106), .A4(new_n597), .ZN(new_n745));
  AND3_X1   g559(.A1(new_n744), .A2(new_n601), .A3(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT107), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n629), .A2(new_n747), .A3(new_n555), .A4(new_n630), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n742), .A2(new_n746), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n705), .A2(new_n236), .ZN(new_n750));
  NOR3_X1   g564(.A1(new_n749), .A2(new_n750), .A3(new_n731), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n740), .B1(new_n751), .B2(KEYINPUT42), .ZN(new_n752));
  AND2_X1   g566(.A1(new_n742), .A2(new_n748), .ZN(new_n753));
  INV_X1    g567(.A(new_n731), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n753), .A2(new_n370), .A3(new_n754), .A4(new_n746), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT42), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n755), .A2(KEYINPUT108), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n752), .A2(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(new_n749), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT109), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n345), .A2(new_n760), .A3(new_n346), .ZN(new_n761));
  OAI21_X1  g575(.A(KEYINPUT109), .B1(new_n356), .B2(KEYINPUT32), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n761), .A2(new_n369), .A3(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n763), .A2(new_n236), .ZN(new_n764));
  INV_X1    g578(.A(new_n764), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n759), .A2(new_n765), .A3(KEYINPUT42), .A4(new_n754), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n758), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G131), .ZN(G33));
  NAND4_X1  g582(.A1(new_n759), .A2(new_n370), .A3(new_n666), .A4(new_n667), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G134), .ZN(G36));
  NAND2_X1  g584(.A1(new_n584), .A2(new_n585), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(new_n570), .ZN(new_n772));
  INV_X1    g586(.A(new_n574), .ZN(new_n773));
  AOI22_X1  g587(.A1(new_n772), .A2(new_n773), .B1(new_n588), .B2(new_n591), .ZN(new_n774));
  OAI21_X1  g588(.A(G469), .B1(new_n774), .B2(KEYINPUT45), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n775), .B1(KEYINPUT45), .B2(new_n774), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n776), .A2(new_n596), .ZN(new_n777));
  OR3_X1    g591(.A1(new_n777), .A2(KEYINPUT110), .A3(KEYINPUT46), .ZN(new_n778));
  OAI21_X1  g592(.A(KEYINPUT110), .B1(new_n777), .B2(KEYINPUT46), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n696), .B1(new_n777), .B2(KEYINPUT46), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n778), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n781), .A2(new_n601), .A3(new_n672), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n742), .A2(new_n748), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n467), .B1(new_n617), .B2(new_n619), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n784), .B1(KEYINPUT111), .B2(KEYINPUT43), .ZN(new_n785));
  XOR2_X1   g599(.A(KEYINPUT111), .B(KEYINPUT43), .Z(new_n786));
  OAI21_X1  g600(.A(new_n785), .B1(new_n784), .B2(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(new_n609), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n787), .A2(new_n788), .A3(new_n654), .ZN(new_n789));
  INV_X1    g603(.A(new_n789), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n783), .B1(new_n790), .B2(KEYINPUT44), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n791), .B1(KEYINPUT44), .B2(new_n790), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n782), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(new_n260), .ZN(G39));
  NAND2_X1  g608(.A1(new_n781), .A2(new_n601), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n795), .A2(KEYINPUT112), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT112), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n781), .A2(new_n797), .A3(new_n601), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT113), .ZN(new_n799));
  OR2_X1    g613(.A1(new_n799), .A2(KEYINPUT47), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n796), .A2(new_n798), .A3(new_n800), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n799), .A2(KEYINPUT47), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n801), .B(new_n802), .ZN(new_n803));
  NOR4_X1   g617(.A1(new_n783), .A2(new_n705), .A3(new_n236), .A4(new_n689), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(G140), .ZN(G42));
  INV_X1    g620(.A(KEYINPUT54), .ZN(new_n807));
  MUX2_X1   g621(.A(new_n418), .B(new_n620), .S(new_n467), .Z(new_n808));
  NAND4_X1  g622(.A1(new_n683), .A2(new_n808), .A3(new_n612), .A4(new_n555), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n604), .B(new_n656), .C1(new_n611), .C2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT53), .ZN(new_n811));
  OR2_X1    g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  AND2_X1   g626(.A1(new_n738), .A2(new_n669), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT52), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  AND2_X1   g629(.A1(new_n721), .A2(new_n725), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n698), .A2(new_n701), .A3(new_n709), .ZN(new_n817));
  NOR4_X1   g631(.A1(new_n812), .A2(new_n815), .A3(new_n816), .A4(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n654), .A2(new_n638), .A3(new_n664), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n819), .A2(new_n602), .A3(new_n418), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n753), .A2(new_n705), .A3(new_n820), .ZN(new_n821));
  OAI211_X1 g635(.A(new_n769), .B(new_n821), .C1(new_n736), .C2(new_n749), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n822), .B1(new_n758), .B2(new_n766), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n682), .A2(new_n711), .A3(new_n664), .A4(new_n746), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n738), .A2(new_n669), .A3(new_n691), .A4(new_n824), .ZN(new_n825));
  XNOR2_X1  g639(.A(new_n825), .B(new_n814), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n818), .A2(new_n823), .A3(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT115), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n828), .B1(new_n817), .B2(new_n816), .ZN(new_n829));
  INV_X1    g643(.A(new_n697), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n750), .A2(new_n830), .ZN(new_n831));
  AOI22_X1  g645(.A1(new_n831), .A2(new_n632), .B1(new_n708), .B2(new_n706), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n832), .A2(KEYINPUT115), .A3(new_n701), .A4(new_n726), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n810), .B1(new_n829), .B2(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n826), .A2(new_n834), .A3(new_n823), .ZN(new_n835));
  AND3_X1   g649(.A1(new_n835), .A2(KEYINPUT116), .A3(new_n811), .ZN(new_n836));
  AOI21_X1  g650(.A(KEYINPUT116), .B1(new_n835), .B2(new_n811), .ZN(new_n837));
  OAI211_X1 g651(.A(new_n807), .B(new_n827), .C1(new_n836), .C2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT117), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n835), .A2(new_n811), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n811), .B1(new_n813), .B2(new_n814), .ZN(new_n841));
  INV_X1    g655(.A(new_n841), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n840), .B1(new_n835), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n843), .A2(KEYINPUT54), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n838), .A2(new_n839), .A3(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n838), .A2(new_n844), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n846), .A2(KEYINPUT117), .ZN(new_n847));
  INV_X1    g661(.A(new_n684), .ZN(new_n848));
  AND4_X1   g662(.A1(new_n236), .A2(new_n787), .A3(new_n469), .A4(new_n723), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n848), .A2(new_n556), .A3(new_n697), .A4(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n850), .A2(KEYINPUT118), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT50), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n783), .A2(new_n830), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n854), .A2(new_n469), .A3(new_n787), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n853), .B1(new_n732), .B2(new_n855), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n348), .A2(new_n681), .ZN(new_n857));
  AND4_X1   g671(.A1(new_n236), .A2(new_n854), .A3(new_n469), .A4(new_n857), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n620), .A2(new_n467), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n860), .B1(new_n852), .B2(new_n851), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n856), .A2(new_n861), .ZN(new_n862));
  XOR2_X1   g676(.A(new_n862), .B(KEYINPUT119), .Z(new_n863));
  NAND2_X1  g677(.A1(new_n718), .A2(new_n590), .ZN(new_n864));
  XNOR2_X1  g678(.A(new_n864), .B(KEYINPUT114), .ZN(new_n865));
  INV_X1    g679(.A(new_n865), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n866), .A2(new_n601), .ZN(new_n867));
  OAI211_X1 g681(.A(new_n753), .B(new_n849), .C1(new_n803), .C2(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n863), .A2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT51), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n855), .A2(new_n764), .ZN(new_n872));
  XOR2_X1   g686(.A(new_n872), .B(KEYINPUT48), .Z(new_n873));
  NAND2_X1  g687(.A1(new_n858), .A2(new_n623), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n468), .B1(new_n849), .B2(new_n708), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n873), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  NOR3_X1   g690(.A1(new_n856), .A2(new_n870), .A3(new_n861), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n876), .B1(new_n868), .B2(new_n877), .ZN(new_n878));
  AND4_X1   g692(.A1(new_n845), .A2(new_n847), .A3(new_n871), .A4(new_n878), .ZN(new_n879));
  NOR2_X1   g693(.A1(G952), .A2(G953), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n236), .A2(new_n555), .A3(new_n601), .A4(new_n784), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n881), .B1(new_n866), .B2(KEYINPUT49), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n882), .B1(KEYINPUT49), .B2(new_n866), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n848), .A2(new_n857), .ZN(new_n884));
  OAI22_X1  g698(.A1(new_n879), .A2(new_n880), .B1(new_n883), .B2(new_n884), .ZN(G75));
  OAI21_X1  g699(.A(new_n827), .B1(new_n836), .B2(new_n837), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n886), .A2(G210), .A3(G902), .ZN(new_n887));
  OR2_X1    g701(.A1(new_n887), .A2(KEYINPUT120), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n887), .A2(KEYINPUT120), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n531), .B(new_n527), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n890), .B(KEYINPUT55), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n891), .A2(KEYINPUT56), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n888), .A2(new_n889), .A3(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(new_n887), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n891), .B1(new_n894), .B2(KEYINPUT56), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n221), .A2(G952), .ZN(new_n896));
  INV_X1    g710(.A(new_n896), .ZN(new_n897));
  AND3_X1   g711(.A1(new_n893), .A2(new_n895), .A3(new_n897), .ZN(G51));
  NAND2_X1  g712(.A1(new_n886), .A2(KEYINPUT54), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT121), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n899), .A2(new_n900), .A3(new_n838), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n886), .A2(KEYINPUT121), .A3(KEYINPUT54), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n596), .B(KEYINPUT57), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n901), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(new_n694), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT116), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n840), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n835), .A2(KEYINPUT116), .A3(new_n811), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n188), .B1(new_n909), .B2(new_n827), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(new_n776), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n896), .B1(new_n905), .B2(new_n911), .ZN(G54));
  NAND2_X1  g726(.A1(new_n457), .A2(new_n458), .ZN(new_n913));
  NAND2_X1  g727(.A1(KEYINPUT58), .A2(G475), .ZN(new_n914));
  XOR2_X1   g728(.A(new_n914), .B(KEYINPUT122), .Z(new_n915));
  AND3_X1   g729(.A1(new_n910), .A2(new_n913), .A3(new_n915), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n913), .B1(new_n910), .B2(new_n915), .ZN(new_n917));
  NOR3_X1   g731(.A1(new_n916), .A2(new_n917), .A3(new_n896), .ZN(G60));
  NAND2_X1  g732(.A1(new_n847), .A2(new_n845), .ZN(new_n919));
  NAND2_X1  g733(.A1(G478), .A2(G902), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n920), .B(KEYINPUT59), .Z(new_n921));
  INV_X1    g735(.A(new_n921), .ZN(new_n922));
  AOI22_X1  g736(.A1(new_n919), .A2(new_n922), .B1(new_n614), .B2(new_n615), .ZN(new_n923));
  AND3_X1   g737(.A1(new_n614), .A2(new_n615), .A3(new_n922), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n901), .A2(new_n902), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n925), .A2(new_n897), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n923), .A2(new_n926), .ZN(G63));
  XNOR2_X1  g741(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n187), .A2(new_n188), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n928), .B(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n886), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n896), .B1(new_n931), .B2(new_n230), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT124), .ZN(new_n933));
  INV_X1    g747(.A(new_n930), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n934), .B1(new_n909), .B2(new_n827), .ZN(new_n935));
  AND2_X1   g749(.A1(new_n649), .A2(new_n651), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n933), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  AND4_X1   g751(.A1(new_n933), .A2(new_n886), .A3(new_n936), .A4(new_n930), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n932), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT61), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  OAI211_X1 g755(.A(KEYINPUT61), .B(new_n932), .C1(new_n937), .C2(new_n938), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n941), .A2(new_n942), .ZN(G66));
  OAI21_X1  g757(.A(G953), .B1(new_n471), .B2(new_n525), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(KEYINPUT125), .ZN(new_n945));
  INV_X1    g759(.A(new_n834), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n946), .A2(new_n221), .ZN(new_n947));
  MUX2_X1   g761(.A(KEYINPUT125), .B(new_n945), .S(new_n947), .Z(new_n948));
  INV_X1    g762(.A(new_n531), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n949), .B1(G898), .B2(new_n221), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n948), .B(new_n950), .ZN(G69));
  AOI21_X1  g765(.A(new_n221), .B1(G227), .B2(G900), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n320), .A2(new_n321), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n953), .B(new_n453), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n813), .A2(new_n687), .A3(new_n691), .ZN(new_n955));
  XOR2_X1   g769(.A(new_n955), .B(KEYINPUT62), .Z(new_n956));
  XOR2_X1   g770(.A(new_n808), .B(KEYINPUT126), .Z(new_n957));
  NOR3_X1   g771(.A1(new_n957), .A2(new_n750), .A3(new_n673), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n793), .B1(new_n753), .B2(new_n958), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n805), .A2(new_n956), .A3(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n954), .B1(new_n960), .B2(new_n221), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(KEYINPUT127), .ZN(new_n962));
  INV_X1    g776(.A(new_n962), .ZN(new_n963));
  NOR3_X1   g777(.A1(new_n782), .A2(new_n722), .A3(new_n764), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n769), .B1(new_n782), .B2(new_n792), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n813), .A2(new_n691), .ZN(new_n966));
  NOR3_X1   g780(.A1(new_n964), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n805), .A2(new_n221), .A3(new_n767), .A4(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(G900), .A2(G953), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n968), .A2(new_n954), .A3(new_n969), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n970), .B1(new_n961), .B2(KEYINPUT127), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n952), .B1(new_n963), .B2(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(KEYINPUT127), .ZN(new_n973));
  AND2_X1   g787(.A1(new_n960), .A2(new_n221), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n973), .B1(new_n974), .B2(new_n954), .ZN(new_n975));
  INV_X1    g789(.A(new_n952), .ZN(new_n976));
  NAND4_X1  g790(.A1(new_n975), .A2(new_n976), .A3(new_n962), .A4(new_n970), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n972), .A2(new_n977), .ZN(G72));
  NAND2_X1  g792(.A1(G472), .A2(G902), .ZN(new_n979));
  XOR2_X1   g793(.A(new_n979), .B(KEYINPUT63), .Z(new_n980));
  INV_X1    g794(.A(new_n980), .ZN(new_n981));
  AND3_X1   g795(.A1(new_n805), .A2(new_n767), .A3(new_n967), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n981), .B1(new_n982), .B2(new_n834), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n312), .A2(new_n351), .A3(new_n322), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n897), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  OR2_X1    g799(.A1(new_n960), .A2(new_n946), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n679), .B1(new_n986), .B2(new_n980), .ZN(new_n987));
  INV_X1    g801(.A(new_n843), .ZN(new_n988));
  AOI211_X1 g802(.A(new_n981), .B(new_n988), .C1(new_n328), .C2(new_n359), .ZN(new_n989));
  NOR3_X1   g803(.A1(new_n985), .A2(new_n987), .A3(new_n989), .ZN(G57));
endmodule


