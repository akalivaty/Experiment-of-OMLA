//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 1 0 1 0 0 0 0 1 1 0 1 0 1 1 1 0 1 1 0 0 1 0 1 0 1 0 1 0 1 0 0 0 1 0 0 1 1 0 0 1 0 1 1 0 1 1 1 1 0 0 1 0 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:30 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n555, new_n556, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n613, new_n614, new_n615, new_n616,
    new_n619, new_n620, new_n622, new_n623, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT64), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XNOR2_X1  g012(.A(KEYINPUT65), .B(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g018(.A(KEYINPUT66), .B(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  OR4_X1    g024(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(new_n452), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n456), .A2(G2106), .ZN(new_n457));
  INV_X1    g032(.A(new_n453), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n458), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT68), .ZN(new_n463));
  XNOR2_X1  g038(.A(KEYINPUT3), .B(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n463), .B1(new_n464), .B2(G125), .ZN(new_n465));
  AND2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  OAI211_X1 g042(.A(new_n463), .B(G125), .C1(new_n466), .C2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(new_n468), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n462), .B1(new_n465), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n472), .A2(G101), .A3(G2104), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n466), .A2(new_n467), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n472), .A2(G137), .ZN(new_n476));
  OAI21_X1  g051(.A(KEYINPUT69), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT69), .ZN(new_n478));
  NAND4_X1  g053(.A1(new_n464), .A2(new_n478), .A3(G137), .A4(new_n472), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n474), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n471), .A2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G160));
  OAI21_X1  g057(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n484), .B1(G112), .B2(new_n472), .ZN(new_n485));
  XNOR2_X1  g060(.A(new_n485), .B(KEYINPUT70), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n475), .A2(G2105), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n475), .A2(new_n472), .ZN(new_n489));
  AOI22_X1  g064(.A1(new_n488), .A2(G136), .B1(G124), .B2(new_n489), .ZN(new_n490));
  AND2_X1   g065(.A1(new_n487), .A2(new_n490), .ZN(G162));
  OAI211_X1 g066(.A(G126), .B(G2105), .C1(new_n466), .C2(new_n467), .ZN(new_n492));
  INV_X1    g067(.A(G114), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(G2105), .ZN(new_n494));
  OAI211_X1 g069(.A(new_n494), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n492), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(G138), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n497), .A2(G2105), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n498), .B1(new_n466), .B2(new_n467), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(KEYINPUT4), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n501));
  OAI211_X1 g076(.A(new_n498), .B(new_n501), .C1(new_n467), .C2(new_n466), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n496), .B1(new_n500), .B2(new_n502), .ZN(G164));
  OR2_X1    g078(.A1(KEYINPUT6), .A2(G651), .ZN(new_n504));
  NAND2_X1  g079(.A1(KEYINPUT6), .A2(G651), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT5), .ZN(new_n506));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(KEYINPUT5), .A2(G543), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n504), .A2(new_n505), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n507), .B1(new_n504), .B2(new_n505), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n510), .A2(G88), .B1(new_n511), .B2(G50), .ZN(new_n512));
  INV_X1    g087(.A(G651), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n508), .A2(new_n509), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n514), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n512), .B1(new_n513), .B2(new_n515), .ZN(G303));
  INV_X1    g091(.A(G303), .ZN(G166));
  NAND3_X1  g092(.A1(new_n514), .A2(G63), .A3(G651), .ZN(new_n518));
  XNOR2_X1  g093(.A(KEYINPUT6), .B(G651), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G543), .ZN(new_n520));
  INV_X1    g095(.A(G51), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n518), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(KEYINPUT71), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT71), .ZN(new_n524));
  OAI211_X1 g099(.A(new_n518), .B(new_n524), .C1(new_n521), .C2(new_n520), .ZN(new_n525));
  XNOR2_X1  g100(.A(KEYINPUT72), .B(KEYINPUT7), .ZN(new_n526));
  AND3_X1   g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  OR2_X1    g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n526), .A2(new_n527), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n528), .A2(new_n529), .B1(G89), .B2(new_n510), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n523), .A2(new_n525), .A3(new_n530), .ZN(G286));
  INV_X1    g106(.A(G286), .ZN(G168));
  NAND2_X1  g107(.A1(new_n514), .A2(G64), .ZN(new_n533));
  NAND2_X1  g108(.A1(G77), .A2(G543), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n513), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT73), .ZN(new_n536));
  AND2_X1   g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  XOR2_X1   g112(.A(KEYINPUT74), .B(G90), .Z(new_n538));
  AOI22_X1  g113(.A1(new_n510), .A2(new_n538), .B1(new_n511), .B2(G52), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n539), .B1(new_n535), .B2(new_n536), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n537), .A2(new_n540), .ZN(G171));
  AOI22_X1  g116(.A1(new_n514), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n542), .A2(new_n513), .ZN(new_n543));
  INV_X1    g118(.A(G43), .ZN(new_n544));
  NOR2_X1   g119(.A1(KEYINPUT5), .A2(G543), .ZN(new_n545));
  AND2_X1   g120(.A1(KEYINPUT5), .A2(G543), .ZN(new_n546));
  AND2_X1   g121(.A1(KEYINPUT6), .A2(G651), .ZN(new_n547));
  NOR2_X1   g122(.A1(KEYINPUT6), .A2(G651), .ZN(new_n548));
  OAI22_X1  g123(.A1(new_n545), .A2(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(G81), .ZN(new_n550));
  OAI22_X1  g125(.A1(new_n520), .A2(new_n544), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n543), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  NAND4_X1  g128(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND4_X1  g131(.A1(G319), .A2(G483), .A3(G661), .A4(new_n556), .ZN(G188));
  AND2_X1   g132(.A1(G53), .A2(G543), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n558), .B1(new_n547), .B2(new_n548), .ZN(new_n559));
  XNOR2_X1  g134(.A(KEYINPUT76), .B(KEYINPUT9), .ZN(new_n560));
  OAI21_X1  g135(.A(KEYINPUT77), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT9), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(KEYINPUT76), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT76), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(KEYINPUT9), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT77), .ZN(new_n567));
  NAND4_X1  g142(.A1(new_n566), .A2(new_n519), .A3(new_n567), .A4(new_n558), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n561), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n559), .A2(KEYINPUT75), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT75), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n519), .A2(new_n571), .A3(new_n558), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n570), .A2(new_n572), .A3(KEYINPUT9), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n569), .A2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT78), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n569), .A2(new_n573), .A3(KEYINPUT78), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(G78), .A2(G543), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n546), .A2(new_n545), .ZN(new_n580));
  INV_X1    g155(.A(G65), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n579), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n582), .A2(G651), .B1(new_n510), .B2(G91), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n578), .A2(new_n583), .ZN(G299));
  INV_X1    g159(.A(G171), .ZN(G301));
  NAND2_X1  g160(.A1(new_n510), .A2(G87), .ZN(new_n586));
  OAI21_X1  g161(.A(G651), .B1(new_n514), .B2(G74), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n511), .A2(G49), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(G288));
  OAI211_X1 g164(.A(G48), .B(G543), .C1(new_n547), .C2(new_n548), .ZN(new_n590));
  INV_X1    g165(.A(G86), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n549), .B2(new_n591), .ZN(new_n592));
  OAI21_X1  g167(.A(G61), .B1(new_n546), .B2(new_n545), .ZN(new_n593));
  NAND2_X1  g168(.A1(G73), .A2(G543), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n513), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(G305));
  AOI22_X1  g172(.A1(new_n514), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n598));
  OR2_X1    g173(.A1(new_n598), .A2(new_n513), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n510), .A2(G85), .B1(new_n511), .B2(G47), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(G290));
  AND3_X1   g176(.A1(new_n514), .A2(new_n519), .A3(G92), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n602), .B(KEYINPUT10), .ZN(new_n603));
  NAND2_X1  g178(.A1(G79), .A2(G543), .ZN(new_n604));
  INV_X1    g179(.A(G66), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n580), .B2(new_n605), .ZN(new_n606));
  AOI22_X1  g181(.A1(new_n606), .A2(G651), .B1(G54), .B2(new_n511), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n603), .A2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(G868), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n610), .B1(G171), .B2(new_n609), .ZN(G284));
  OAI21_X1  g186(.A(new_n610), .B1(G171), .B2(new_n609), .ZN(G321));
  NAND2_X1  g187(.A1(G286), .A2(G868), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT79), .ZN(new_n614));
  INV_X1    g189(.A(new_n583), .ZN(new_n615));
  AOI21_X1  g190(.A(new_n615), .B1(new_n576), .B2(new_n577), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n614), .B1(G868), .B2(new_n616), .ZN(G297));
  OAI21_X1  g192(.A(new_n614), .B1(G868), .B2(new_n616), .ZN(G280));
  INV_X1    g193(.A(new_n608), .ZN(new_n619));
  INV_X1    g194(.A(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n620), .B2(G860), .ZN(G148));
  NAND2_X1  g196(.A1(new_n619), .A2(new_n620), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n622), .A2(G868), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n623), .B1(G868), .B2(new_n552), .ZN(G323));
  XNOR2_X1  g199(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g200(.A1(new_n488), .A2(G135), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n489), .A2(G123), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n472), .A2(G111), .ZN(new_n628));
  OAI21_X1  g203(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n629));
  OAI211_X1 g204(.A(new_n626), .B(new_n627), .C1(new_n628), .C2(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT82), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(G2096), .Z(new_n632));
  NAND3_X1  g207(.A1(new_n472), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT81), .ZN(new_n634));
  XNOR2_X1  g209(.A(KEYINPUT80), .B(KEYINPUT12), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(KEYINPUT13), .Z(new_n637));
  INV_X1    g212(.A(G2100), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n637), .A2(new_n638), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n632), .A2(new_n639), .A3(new_n640), .ZN(G156));
  XNOR2_X1  g216(.A(G2427), .B(G2438), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G2430), .ZN(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT15), .B(G2435), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n643), .A2(new_n644), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n645), .A2(KEYINPUT14), .A3(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2451), .B(G2454), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT16), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n647), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2443), .B(G2446), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G1341), .B(G1348), .ZN(new_n653));
  OAI21_X1  g228(.A(G14), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n652), .A2(new_n653), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n655), .A2(KEYINPUT83), .ZN(new_n656));
  INV_X1    g231(.A(KEYINPUT83), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n652), .A2(new_n657), .A3(new_n653), .ZN(new_n658));
  AOI21_X1  g233(.A(new_n654), .B1(new_n656), .B2(new_n658), .ZN(G401));
  XNOR2_X1  g234(.A(G2084), .B(G2090), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT84), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2067), .B(G2678), .ZN(new_n662));
  AND2_X1   g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2072), .B(G2078), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n665), .B(KEYINPUT18), .Z(new_n666));
  NOR2_X1   g241(.A1(new_n661), .A2(new_n662), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n664), .B(KEYINPUT85), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n664), .B(KEYINPUT17), .ZN(new_n670));
  OR3_X1    g245(.A1(new_n663), .A2(new_n667), .A3(new_n670), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n666), .A2(new_n669), .A3(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(G2096), .B(G2100), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(G227));
  XOR2_X1   g249(.A(G1971), .B(G1976), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT19), .ZN(new_n676));
  XOR2_X1   g251(.A(G1956), .B(G2474), .Z(new_n677));
  XOR2_X1   g252(.A(G1961), .B(G1966), .Z(new_n678));
  AND2_X1   g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT20), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n677), .A2(new_n678), .ZN(new_n682));
  NOR3_X1   g257(.A1(new_n676), .A2(new_n679), .A3(new_n682), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n683), .B1(new_n676), .B2(new_n682), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(G1981), .ZN(new_n686));
  XOR2_X1   g261(.A(KEYINPUT86), .B(KEYINPUT87), .Z(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n686), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1991), .B(G1996), .ZN(new_n691));
  INV_X1    g266(.A(G1986), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n690), .B(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(G229));
  NOR2_X1   g270(.A1(G29), .A2(G35), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(G162), .B2(G29), .ZN(new_n697));
  XOR2_X1   g272(.A(new_n697), .B(KEYINPUT29), .Z(new_n698));
  INV_X1    g273(.A(G2090), .ZN(new_n699));
  INV_X1    g274(.A(G1961), .ZN(new_n700));
  INV_X1    g275(.A(G16), .ZN(new_n701));
  NOR2_X1   g276(.A1(G171), .A2(new_n701), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n702), .B1(G5), .B2(new_n701), .ZN(new_n703));
  OAI22_X1  g278(.A1(new_n698), .A2(new_n699), .B1(new_n700), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n489), .A2(G129), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT97), .ZN(new_n706));
  NAND3_X1  g281(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT26), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n472), .A2(G105), .A3(G2104), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT98), .ZN(new_n710));
  AOI211_X1 g285(.A(new_n708), .B(new_n710), .C1(G141), .C2(new_n488), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n706), .A2(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(G29), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n715), .B1(new_n714), .B2(G32), .ZN(new_n716));
  XNOR2_X1  g291(.A(KEYINPUT27), .B(G1996), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n714), .A2(G27), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT101), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(G164), .B2(new_n714), .ZN(new_n721));
  INV_X1    g296(.A(G2078), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n718), .A2(new_n723), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n716), .A2(new_n717), .ZN(new_n725));
  NOR2_X1   g300(.A1(G286), .A2(new_n701), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n726), .A2(KEYINPUT99), .ZN(new_n727));
  INV_X1    g302(.A(KEYINPUT99), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(G16), .B2(G21), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n727), .B1(new_n726), .B2(new_n729), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(G1966), .ZN(new_n731));
  NOR4_X1   g306(.A1(new_n704), .A2(new_n724), .A3(new_n725), .A4(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n698), .A2(new_n699), .ZN(new_n733));
  AND2_X1   g308(.A1(new_n714), .A2(G33), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n472), .A2(G103), .A3(G2104), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(KEYINPUT25), .Z(new_n736));
  INV_X1    g311(.A(new_n488), .ZN(new_n737));
  INV_X1    g312(.A(G139), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n736), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  AND2_X1   g314(.A1(new_n464), .A2(G127), .ZN(new_n740));
  AND2_X1   g315(.A1(G115), .A2(G2104), .ZN(new_n741));
  OAI21_X1  g316(.A(G2105), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n739), .B1(KEYINPUT96), .B2(new_n742), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(KEYINPUT96), .B2(new_n742), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n734), .B1(new_n744), .B2(G29), .ZN(new_n745));
  INV_X1    g320(.A(G2072), .ZN(new_n746));
  OR2_X1    g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n745), .A2(new_n746), .ZN(new_n748));
  XNOR2_X1  g323(.A(KEYINPUT30), .B(G28), .ZN(new_n749));
  OR2_X1    g324(.A1(KEYINPUT31), .A2(G11), .ZN(new_n750));
  NAND2_X1  g325(.A1(KEYINPUT31), .A2(G11), .ZN(new_n751));
  AOI22_X1  g326(.A1(new_n749), .A2(new_n714), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(new_n631), .B2(new_n714), .ZN(new_n753));
  INV_X1    g328(.A(KEYINPUT100), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND4_X1  g330(.A1(new_n733), .A2(new_n747), .A3(new_n748), .A4(new_n755), .ZN(new_n756));
  AND2_X1   g331(.A1(KEYINPUT24), .A2(G34), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n714), .B1(KEYINPUT24), .B2(G34), .ZN(new_n758));
  OAI22_X1  g333(.A1(G160), .A2(new_n714), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  AOI22_X1  g334(.A1(new_n703), .A2(new_n700), .B1(G2084), .B2(new_n759), .ZN(new_n760));
  OAI221_X1 g335(.A(new_n760), .B1(new_n754), .B2(new_n753), .C1(G2084), .C2(new_n759), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n756), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n701), .A2(G20), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT23), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(new_n616), .B2(new_n701), .ZN(new_n765));
  INV_X1    g340(.A(G1956), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n732), .A2(new_n762), .A3(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n488), .A2(G140), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n489), .A2(G128), .ZN(new_n770));
  OR2_X1    g345(.A1(G104), .A2(G2105), .ZN(new_n771));
  OAI211_X1 g346(.A(new_n771), .B(G2104), .C1(G116), .C2(new_n472), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n769), .A2(new_n770), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n773), .A2(G29), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(KEYINPUT94), .Z(new_n775));
  NAND2_X1  g350(.A1(new_n714), .A2(G26), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT28), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(G2067), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n701), .A2(G19), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(new_n552), .B2(new_n701), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(G1341), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n619), .A2(G16), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(G4), .B2(G16), .ZN(new_n785));
  INV_X1    g360(.A(G1348), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n783), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  OAI211_X1 g362(.A(new_n780), .B(new_n787), .C1(new_n786), .C2(new_n785), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT95), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n768), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n701), .A2(G23), .ZN(new_n791));
  INV_X1    g366(.A(G288), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n791), .B1(new_n792), .B2(new_n701), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT93), .ZN(new_n794));
  XOR2_X1   g369(.A(KEYINPUT33), .B(G1976), .Z(new_n795));
  OR2_X1    g370(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n794), .A2(new_n795), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n701), .A2(G22), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(G166), .B2(new_n701), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(G1971), .Z(new_n800));
  NOR2_X1   g375(.A1(G6), .A2(G16), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(new_n596), .B2(G16), .ZN(new_n802));
  XOR2_X1   g377(.A(KEYINPUT32), .B(G1981), .Z(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NAND4_X1  g379(.A1(new_n796), .A2(new_n797), .A3(new_n800), .A4(new_n804), .ZN(new_n805));
  OR2_X1    g380(.A1(new_n805), .A2(KEYINPUT34), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n701), .A2(G24), .ZN(new_n807));
  XOR2_X1   g382(.A(new_n807), .B(KEYINPUT91), .Z(new_n808));
  AOI21_X1  g383(.A(new_n808), .B1(G290), .B2(G16), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT92), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(G1986), .ZN(new_n811));
  AND2_X1   g386(.A1(new_n714), .A2(G25), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n488), .A2(G131), .ZN(new_n813));
  NOR2_X1   g388(.A1(G95), .A2(G2105), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT89), .ZN(new_n815));
  OAI21_X1  g390(.A(G2104), .B1(new_n472), .B2(G107), .ZN(new_n816));
  AND3_X1   g391(.A1(new_n489), .A2(KEYINPUT88), .A3(G119), .ZN(new_n817));
  AOI21_X1  g392(.A(KEYINPUT88), .B1(new_n489), .B2(G119), .ZN(new_n818));
  OAI221_X1 g393(.A(new_n813), .B1(new_n815), .B2(new_n816), .C1(new_n817), .C2(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(KEYINPUT90), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n812), .B1(new_n821), .B2(G29), .ZN(new_n822));
  XOR2_X1   g397(.A(KEYINPUT35), .B(G1991), .Z(new_n823));
  AND2_X1   g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n822), .A2(new_n823), .ZN(new_n825));
  NOR3_X1   g400(.A1(new_n811), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n805), .A2(KEYINPUT34), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n806), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(KEYINPUT36), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n790), .A2(new_n829), .ZN(G150));
  INV_X1    g405(.A(G150), .ZN(G311));
  NAND2_X1  g406(.A1(new_n619), .A2(G559), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT38), .ZN(new_n833));
  INV_X1    g408(.A(G67), .ZN(new_n834));
  INV_X1    g409(.A(G80), .ZN(new_n835));
  OAI22_X1  g410(.A1(new_n580), .A2(new_n834), .B1(new_n835), .B2(new_n507), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n836), .A2(KEYINPUT102), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT102), .ZN(new_n838));
  OAI221_X1 g413(.A(new_n838), .B1(new_n835), .B2(new_n507), .C1(new_n580), .C2(new_n834), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n837), .A2(G651), .A3(new_n839), .ZN(new_n840));
  XOR2_X1   g415(.A(KEYINPUT103), .B(G93), .Z(new_n841));
  AOI22_X1  g416(.A1(new_n510), .A2(new_n841), .B1(new_n511), .B2(G55), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  OR2_X1    g418(.A1(new_n543), .A2(new_n551), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n552), .A2(new_n840), .A3(new_n842), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n833), .B(new_n847), .Z(new_n848));
  OR2_X1    g423(.A1(new_n848), .A2(KEYINPUT39), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(KEYINPUT39), .ZN(new_n850));
  XOR2_X1   g425(.A(KEYINPUT104), .B(G860), .Z(new_n851));
  NAND3_X1  g426(.A1(new_n849), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n851), .B1(new_n840), .B2(new_n842), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(KEYINPUT37), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n852), .A2(new_n854), .ZN(G145));
  NAND2_X1  g430(.A1(new_n488), .A2(G142), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n489), .A2(G130), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n472), .A2(G118), .ZN(new_n858));
  OAI21_X1  g433(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n859));
  OAI211_X1 g434(.A(new_n856), .B(new_n857), .C1(new_n858), .C2(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n636), .B(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(new_n819), .ZN(new_n862));
  INV_X1    g437(.A(new_n773), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n862), .B(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n744), .B(new_n712), .ZN(new_n865));
  INV_X1    g440(.A(new_n502), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n501), .B1(new_n464), .B2(new_n498), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  OAI21_X1  g443(.A(KEYINPUT106), .B1(new_n868), .B2(new_n496), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n500), .A2(new_n502), .ZN(new_n870));
  AND2_X1   g445(.A1(new_n492), .A2(new_n495), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT106), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n870), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n869), .A2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n865), .B(new_n875), .ZN(new_n876));
  OR2_X1    g451(.A1(new_n864), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n864), .A2(new_n876), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n631), .B(KEYINPUT105), .ZN(new_n880));
  OR2_X1    g455(.A1(new_n880), .A2(new_n481), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n481), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(G162), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n881), .A2(new_n882), .A3(G162), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n879), .A2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(G37), .ZN(new_n889));
  NAND4_X1  g464(.A1(new_n877), .A2(new_n878), .A3(new_n886), .A4(new_n885), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n888), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  XOR2_X1   g466(.A(KEYINPUT107), .B(KEYINPUT40), .Z(new_n892));
  XNOR2_X1  g467(.A(new_n891), .B(new_n892), .ZN(G395));
  NAND2_X1  g468(.A1(new_n843), .A2(new_n609), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT108), .ZN(new_n895));
  NAND3_X1  g470(.A1(G299), .A2(new_n895), .A3(new_n619), .ZN(new_n896));
  OAI21_X1  g471(.A(KEYINPUT108), .B1(new_n616), .B2(new_n608), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n616), .A2(new_n608), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n622), .B(new_n847), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  OR2_X1    g477(.A1(new_n902), .A2(KEYINPUT109), .ZN(new_n903));
  NAND2_X1  g478(.A1(G299), .A2(new_n619), .ZN(new_n904));
  AOI21_X1  g479(.A(KEYINPUT41), .B1(new_n904), .B2(new_n899), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n899), .A2(KEYINPUT41), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n905), .B1(new_n898), .B2(new_n907), .ZN(new_n908));
  OR2_X1    g483(.A1(new_n908), .A2(new_n901), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n902), .A2(KEYINPUT109), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n903), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(G290), .B(new_n596), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n792), .B(G303), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n912), .B(new_n913), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n914), .B(KEYINPUT42), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n911), .A2(new_n916), .ZN(new_n917));
  NAND4_X1  g492(.A1(new_n903), .A2(new_n909), .A3(new_n910), .A4(new_n915), .ZN(new_n918));
  AND2_X1   g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n894), .B1(new_n919), .B2(new_n609), .ZN(G295));
  INV_X1    g495(.A(KEYINPUT110), .ZN(new_n921));
  OAI211_X1 g496(.A(new_n921), .B(new_n894), .C1(new_n919), .C2(new_n609), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n609), .B1(new_n917), .B2(new_n918), .ZN(new_n923));
  INV_X1    g498(.A(new_n894), .ZN(new_n924));
  OAI21_X1  g499(.A(KEYINPUT110), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n922), .A2(new_n925), .ZN(G331));
  AND3_X1   g501(.A1(new_n845), .A2(G286), .A3(new_n846), .ZN(new_n927));
  AOI21_X1  g502(.A(G286), .B1(new_n845), .B2(new_n846), .ZN(new_n928));
  OAI21_X1  g503(.A(G301), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n847), .A2(G168), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n845), .A2(G286), .A3(new_n846), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n930), .A2(G171), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n929), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(new_n900), .ZN(new_n934));
  OAI211_X1 g509(.A(new_n934), .B(new_n914), .C1(new_n908), .C2(new_n933), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(new_n889), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n906), .B1(new_n897), .B2(new_n896), .ZN(new_n937));
  OAI211_X1 g512(.A(new_n932), .B(new_n929), .C1(new_n937), .C2(new_n905), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n914), .B1(new_n938), .B2(new_n934), .ZN(new_n939));
  OAI21_X1  g514(.A(KEYINPUT43), .B1(new_n936), .B2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT111), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  OAI211_X1 g517(.A(KEYINPUT111), .B(KEYINPUT43), .C1(new_n936), .C2(new_n939), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n934), .A2(KEYINPUT112), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT112), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n933), .A2(new_n900), .A3(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT41), .ZN(new_n947));
  AOI22_X1  g522(.A1(new_n900), .A2(new_n947), .B1(new_n904), .B2(new_n907), .ZN(new_n948));
  OAI211_X1 g523(.A(new_n944), .B(new_n946), .C1(new_n933), .C2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(new_n914), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT43), .ZN(new_n952));
  INV_X1    g527(.A(new_n936), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n951), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n942), .A2(new_n943), .A3(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT44), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n951), .A2(KEYINPUT43), .A3(new_n953), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n952), .B1(new_n936), .B2(new_n939), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n960), .A2(KEYINPUT44), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n957), .A2(new_n961), .ZN(G397));
  INV_X1    g537(.A(KEYINPUT45), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n963), .B1(new_n874), .B2(G1384), .ZN(new_n964));
  INV_X1    g539(.A(new_n462), .ZN(new_n965));
  INV_X1    g540(.A(G125), .ZN(new_n966));
  OAI21_X1  g541(.A(KEYINPUT68), .B1(new_n475), .B2(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n965), .B1(new_n967), .B2(new_n468), .ZN(new_n968));
  OAI211_X1 g543(.A(new_n480), .B(G40), .C1(new_n968), .C2(new_n472), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n964), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(G1996), .ZN(new_n971));
  AOI21_X1  g546(.A(KEYINPUT114), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT114), .ZN(new_n973));
  NOR4_X1   g548(.A1(new_n964), .A2(new_n973), .A3(G1996), .A4(new_n969), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n713), .B1(new_n972), .B2(new_n974), .ZN(new_n975));
  XNOR2_X1  g550(.A(new_n773), .B(new_n779), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n976), .B1(new_n713), .B2(new_n971), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n970), .A2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(new_n970), .ZN(new_n979));
  XNOR2_X1  g554(.A(new_n819), .B(new_n823), .ZN(new_n980));
  OAI211_X1 g555(.A(new_n975), .B(new_n978), .C1(new_n979), .C2(new_n980), .ZN(new_n981));
  NOR2_X1   g556(.A1(G290), .A2(G1986), .ZN(new_n982));
  XOR2_X1   g557(.A(new_n982), .B(KEYINPUT113), .Z(new_n983));
  NAND2_X1  g558(.A1(G290), .A2(G1986), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n979), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n981), .A2(new_n985), .ZN(new_n986));
  AND3_X1   g561(.A1(new_n569), .A2(KEYINPUT78), .A3(new_n573), .ZN(new_n987));
  AOI21_X1  g562(.A(KEYINPUT78), .B1(new_n569), .B2(new_n573), .ZN(new_n988));
  OAI211_X1 g563(.A(KEYINPUT57), .B(new_n583), .C1(new_n987), .C2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT119), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n574), .A2(new_n583), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT57), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n990), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n989), .A2(new_n993), .ZN(new_n994));
  NAND4_X1  g569(.A1(new_n578), .A2(new_n990), .A3(KEYINPUT57), .A4(new_n583), .ZN(new_n995));
  INV_X1    g570(.A(G40), .ZN(new_n996));
  AOI211_X1 g571(.A(new_n996), .B(new_n474), .C1(new_n477), .C2(new_n479), .ZN(new_n997));
  AOI21_X1  g572(.A(G1384), .B1(new_n870), .B2(new_n871), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT50), .ZN(new_n999));
  OAI211_X1 g574(.A(new_n471), .B(new_n997), .C1(new_n998), .C2(new_n999), .ZN(new_n1000));
  NOR3_X1   g575(.A1(G164), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n766), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n963), .A2(G1384), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n869), .A2(new_n873), .A3(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n967), .A2(new_n468), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n472), .B1(new_n1005), .B2(new_n462), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n477), .A2(new_n479), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1007), .A2(G40), .A3(new_n473), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n963), .B1(G164), .B2(G1384), .ZN(new_n1010));
  XNOR2_X1  g585(.A(KEYINPUT56), .B(G2072), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n1004), .A2(new_n1009), .A3(new_n1010), .A4(new_n1011), .ZN(new_n1012));
  AOI22_X1  g587(.A1(new_n994), .A2(new_n995), .B1(new_n1002), .B2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g588(.A(KEYINPUT61), .B1(new_n1013), .B2(KEYINPUT121), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n994), .A2(new_n995), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1002), .A2(new_n1012), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT121), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n994), .A2(new_n995), .A3(new_n1002), .A4(new_n1012), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1017), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1014), .A2(new_n1020), .ZN(new_n1021));
  AND3_X1   g596(.A1(new_n994), .A2(new_n995), .A3(KEYINPUT120), .ZN(new_n1022));
  AOI21_X1  g597(.A(KEYINPUT120), .B1(new_n994), .B2(new_n995), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1016), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  AND2_X1   g599(.A1(new_n1019), .A2(KEYINPUT61), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n998), .A2(new_n999), .ZN(new_n1027));
  OAI21_X1  g602(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1009), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n471), .A2(new_n997), .A3(new_n998), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1030), .ZN(new_n1031));
  AOI22_X1  g606(.A1(new_n1029), .A2(new_n786), .B1(new_n1031), .B2(new_n779), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n608), .A2(KEYINPUT60), .ZN(new_n1033));
  AND2_X1   g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1004), .A2(new_n971), .A3(new_n1009), .A4(new_n1010), .ZN(new_n1035));
  XOR2_X1   g610(.A(KEYINPUT58), .B(G1341), .Z(new_n1036));
  NAND2_X1  g611(.A1(new_n1030), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1035), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(new_n552), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(KEYINPUT59), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT59), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1038), .A2(new_n1041), .A3(new_n552), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1034), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1043));
  AND2_X1   g618(.A1(new_n1032), .A2(new_n608), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n1032), .A2(new_n608), .ZN(new_n1045));
  OAI21_X1  g620(.A(KEYINPUT60), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1021), .A2(new_n1026), .A3(new_n1043), .A4(new_n1046), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1024), .B1(new_n608), .B2(new_n1032), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(new_n1019), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1047), .A2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n870), .A2(new_n871), .ZN(new_n1051));
  INV_X1    g626(.A(G1384), .ZN(new_n1052));
  AOI21_X1  g627(.A(KEYINPUT45), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1053), .A2(new_n969), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1051), .A2(new_n1003), .ZN(new_n1055));
  AOI21_X1  g630(.A(G1966), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  NOR3_X1   g631(.A1(new_n1000), .A2(G2084), .A3(new_n1001), .ZN(new_n1057));
  OAI211_X1 g632(.A(KEYINPUT122), .B(G8), .C1(new_n1056), .C2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(G8), .ZN(new_n1059));
  NOR2_X1   g634(.A1(G168), .A2(new_n1059), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1060), .A2(KEYINPUT51), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1058), .A2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1009), .A2(new_n1055), .A3(new_n1010), .ZN(new_n1063));
  INV_X1    g638(.A(G1966), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(G2084), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1009), .A2(new_n1027), .A3(new_n1028), .A4(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1065), .A2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(KEYINPUT122), .B1(new_n1068), .B2(G8), .ZN(new_n1069));
  OAI21_X1  g644(.A(KEYINPUT123), .B1(new_n1062), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT122), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1072));
  AOI22_X1  g647(.A1(new_n1072), .A2(new_n1066), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1071), .B1(new_n1073), .B2(new_n1059), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT123), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1074), .A2(new_n1075), .A3(new_n1058), .A4(new_n1061), .ZN(new_n1076));
  OAI211_X1 g651(.A(KEYINPUT51), .B(G8), .C1(new_n1068), .C2(G286), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1070), .A2(new_n1076), .A3(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1068), .A2(new_n1060), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1004), .A2(new_n722), .A3(new_n1009), .A4(new_n1010), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT53), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1081), .A2(KEYINPUT124), .A3(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(KEYINPUT124), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1029), .A2(new_n700), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1082), .A2(G2078), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1088), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1087), .B1(new_n1063), .B2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g665(.A(G171), .B1(new_n1086), .B2(new_n1090), .ZN(new_n1091));
  OR2_X1    g666(.A1(new_n968), .A2(KEYINPUT125), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n472), .B1(new_n968), .B2(KEYINPUT125), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1008), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n964), .A2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT126), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n964), .A2(KEYINPUT126), .A3(new_n1094), .ZN(new_n1098));
  AND3_X1   g673(.A1(new_n870), .A2(new_n872), .A3(new_n871), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n872), .B1(new_n870), .B2(new_n871), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1003), .ZN(new_n1101));
  NOR3_X1   g676(.A1(new_n1099), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1102), .A2(new_n1089), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1097), .A2(new_n1098), .A3(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT124), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(new_n1083), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1104), .A2(new_n1108), .A3(G301), .A4(new_n1087), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1091), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT54), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n515), .A2(new_n513), .ZN(new_n1114));
  INV_X1    g689(.A(G50), .ZN(new_n1115));
  INV_X1    g690(.A(G88), .ZN(new_n1116));
  OAI22_X1  g691(.A1(new_n520), .A2(new_n1115), .B1(new_n549), .B2(new_n1116), .ZN(new_n1117));
  OAI211_X1 g692(.A(KEYINPUT55), .B(G8), .C1(new_n1114), .C2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1118), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1113), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1120), .ZN(new_n1121));
  XOR2_X1   g696(.A(KEYINPUT115), .B(G1971), .Z(new_n1122));
  OAI211_X1 g697(.A(new_n471), .B(new_n997), .C1(new_n998), .C2(KEYINPUT45), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1122), .B1(new_n1102), .B2(new_n1123), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1009), .A2(new_n1027), .A3(new_n1028), .A4(new_n699), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1121), .B1(new_n1126), .B2(G8), .ZN(new_n1127));
  AOI211_X1 g702(.A(new_n1059), .B(new_n1120), .C1(new_n1124), .C2(new_n1125), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(G1976), .ZN(new_n1130));
  AOI21_X1  g705(.A(KEYINPUT52), .B1(G288), .B2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n792), .A2(G1976), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1030), .A2(new_n1131), .A3(G8), .A4(new_n1132), .ZN(new_n1133));
  OAI21_X1  g708(.A(G1981), .B1(new_n592), .B2(new_n595), .ZN(new_n1134));
  INV_X1    g709(.A(G61), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1135), .B1(new_n508), .B2(new_n509), .ZN(new_n1136));
  INV_X1    g711(.A(new_n594), .ZN(new_n1137));
  OAI21_X1  g712(.A(G651), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(G1981), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n514), .A2(new_n519), .A3(G86), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1138), .A2(new_n1139), .A3(new_n1140), .A4(new_n590), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1134), .A2(KEYINPUT49), .A3(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1142), .A2(KEYINPUT117), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT117), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1134), .A2(new_n1141), .A3(new_n1144), .A4(KEYINPUT49), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1143), .A2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT49), .ZN(new_n1147));
  AOI22_X1  g722(.A1(new_n510), .A2(G86), .B1(new_n511), .B2(G48), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1139), .B1(new_n1148), .B2(new_n1138), .ZN(new_n1149));
  NOR3_X1   g724(.A1(new_n592), .A2(new_n595), .A3(G1981), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1147), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1151), .A2(new_n1030), .A3(G8), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1133), .B1(new_n1146), .B2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1030), .A2(G8), .A3(new_n1132), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1154), .A2(KEYINPUT52), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1155), .A2(KEYINPUT116), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT116), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1154), .A2(new_n1157), .A3(KEYINPUT52), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1153), .B1(new_n1156), .B2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1129), .A2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1104), .A2(new_n1108), .A3(new_n1087), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1161), .A2(G171), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1090), .B1(new_n1107), .B2(new_n1083), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1111), .B1(new_n1163), .B2(G301), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1160), .B1(new_n1162), .B2(new_n1164), .ZN(new_n1165));
  NAND4_X1  g740(.A1(new_n1050), .A2(new_n1080), .A3(new_n1112), .A4(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(new_n1122), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1167), .B1(new_n1054), .B2(new_n1004), .ZN(new_n1168));
  INV_X1    g743(.A(new_n1125), .ZN(new_n1169));
  OAI21_X1  g744(.A(G8), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1170), .A2(new_n1120), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1126), .A2(G8), .A3(new_n1121), .ZN(new_n1172));
  AOI211_X1 g747(.A(new_n1059), .B(G286), .C1(new_n1065), .C2(new_n1067), .ZN(new_n1173));
  NAND4_X1  g748(.A1(new_n1159), .A2(new_n1171), .A3(new_n1172), .A4(new_n1173), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT63), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  NAND4_X1  g751(.A1(new_n1129), .A2(KEYINPUT63), .A3(new_n1159), .A4(new_n1173), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT118), .ZN(new_n1179));
  OR2_X1    g754(.A1(new_n1146), .A2(new_n1152), .ZN(new_n1180));
  NOR2_X1   g755(.A1(G288), .A2(G1976), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1182), .A2(new_n1141), .ZN(new_n1183));
  NOR2_X1   g758(.A1(new_n1031), .A2(new_n1059), .ZN(new_n1184));
  AOI22_X1  g759(.A1(new_n1183), .A2(new_n1184), .B1(new_n1159), .B2(new_n1128), .ZN(new_n1185));
  AND3_X1   g760(.A1(new_n1178), .A2(new_n1179), .A3(new_n1185), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1179), .B1(new_n1178), .B2(new_n1185), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1166), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1080), .A2(KEYINPUT62), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT62), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1078), .A2(new_n1190), .A3(new_n1079), .ZN(new_n1191));
  NOR2_X1   g766(.A1(new_n1160), .A2(new_n1091), .ZN(new_n1192));
  AND3_X1   g767(.A1(new_n1189), .A2(new_n1191), .A3(new_n1192), .ZN(new_n1193));
  OAI21_X1  g768(.A(new_n986), .B1(new_n1188), .B2(new_n1193), .ZN(new_n1194));
  INV_X1    g769(.A(new_n821), .ZN(new_n1195));
  NAND4_X1  g770(.A1(new_n975), .A2(new_n1195), .A3(new_n823), .A4(new_n978), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n863), .A2(new_n779), .ZN(new_n1197));
  AOI21_X1  g772(.A(new_n979), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  NOR2_X1   g773(.A1(new_n979), .A2(new_n983), .ZN(new_n1199));
  XNOR2_X1  g774(.A(new_n1199), .B(KEYINPUT48), .ZN(new_n1200));
  NOR2_X1   g775(.A1(new_n1200), .A2(new_n981), .ZN(new_n1201));
  AOI21_X1  g776(.A(new_n979), .B1(new_n713), .B2(new_n976), .ZN(new_n1202));
  INV_X1    g777(.A(KEYINPUT46), .ZN(new_n1203));
  OR3_X1    g778(.A1(new_n972), .A2(new_n1203), .A3(new_n974), .ZN(new_n1204));
  OAI21_X1  g779(.A(new_n1203), .B1(new_n972), .B2(new_n974), .ZN(new_n1205));
  AOI21_X1  g780(.A(new_n1202), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  INV_X1    g781(.A(KEYINPUT47), .ZN(new_n1207));
  OR2_X1    g782(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1209));
  AOI211_X1 g784(.A(new_n1198), .B(new_n1201), .C1(new_n1208), .C2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1194), .A2(new_n1210), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g786(.A1(G227), .A2(new_n460), .ZN(new_n1213));
  AND2_X1   g787(.A1(new_n656), .A2(new_n658), .ZN(new_n1214));
  OAI211_X1 g788(.A(KEYINPUT127), .B(new_n1213), .C1(new_n1214), .C2(new_n654), .ZN(new_n1215));
  INV_X1    g789(.A(KEYINPUT127), .ZN(new_n1216));
  INV_X1    g790(.A(new_n1213), .ZN(new_n1217));
  OAI21_X1  g791(.A(new_n1216), .B1(G401), .B2(new_n1217), .ZN(new_n1218));
  AND3_X1   g792(.A1(new_n1215), .A2(new_n694), .A3(new_n1218), .ZN(new_n1219));
  AND3_X1   g793(.A1(new_n1219), .A2(new_n955), .A3(new_n891), .ZN(G308));
  NAND3_X1  g794(.A1(new_n1219), .A2(new_n955), .A3(new_n891), .ZN(G225));
endmodule


