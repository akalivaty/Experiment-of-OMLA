//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 1 1 1 0 1 1 1 0 0 1 0 0 0 1 0 1 1 0 0 0 1 1 0 1 1 1 0 1 0 0 1 0 0 1 1 1 1 0 1 0 0 1 1 1 1 1 1 0 0 0 1 0 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:42 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n449, new_n450, new_n452, new_n455,
    new_n456, new_n457, new_n458, new_n459, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n551,
    new_n552, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n571, new_n573, new_n574, new_n575,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n613, new_n614, new_n616, new_n617, new_n618, new_n620,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1210, new_n1211, new_n1212, new_n1213;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT64), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g023(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n449));
  NAND2_X1  g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n449), .B(new_n450), .ZN(G223));
  INV_X1    g026(.A(new_n450), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n452), .A2(G567), .ZN(G234));
  NAND2_X1  g028(.A1(new_n452), .A2(G2106), .ZN(G217));
  NOR4_X1   g029(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT2), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR4_X1   g032(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n457), .A2(new_n459), .ZN(G325));
  INV_X1    g035(.A(G325), .ZN(G261));
  AOI22_X1  g036(.A1(new_n457), .A2(G2106), .B1(G567), .B2(new_n459), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  AND2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  OAI21_X1  g040(.A(G125), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n463), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  OAI211_X1 g043(.A(G137), .B(new_n463), .C1(new_n464), .C2(new_n465), .ZN(new_n469));
  INV_X1    g044(.A(G2104), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G101), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n468), .A2(new_n473), .ZN(G160));
  OAI21_X1  g049(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n475));
  INV_X1    g050(.A(G112), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n475), .B1(new_n476), .B2(G2105), .ZN(new_n477));
  OR2_X1    g052(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n463), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n481), .B(KEYINPUT66), .ZN(new_n482));
  XNOR2_X1  g057(.A(KEYINPUT3), .B(G2104), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(new_n463), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  AOI211_X1 g060(.A(new_n477), .B(new_n482), .C1(G136), .C2(new_n485), .ZN(G162));
  OAI21_X1  g061(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(G114), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G2105), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n488), .A2(KEYINPUT67), .A3(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT67), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n463), .A2(G114), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n492), .B1(new_n493), .B2(new_n487), .ZN(new_n494));
  AOI22_X1  g069(.A1(new_n491), .A2(new_n494), .B1(new_n480), .B2(G126), .ZN(new_n495));
  INV_X1    g070(.A(G138), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n496), .A2(G2105), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n497), .B1(new_n464), .B2(new_n465), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT4), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n500));
  OAI211_X1 g075(.A(new_n497), .B(new_n500), .C1(new_n465), .C2(new_n464), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n495), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(G164));
  XNOR2_X1  g079(.A(KEYINPUT6), .B(G651), .ZN(new_n505));
  XNOR2_X1  g080(.A(KEYINPUT5), .B(G543), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT69), .ZN(new_n507));
  AND3_X1   g082(.A1(new_n505), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n507), .B1(new_n505), .B2(new_n506), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  XNOR2_X1  g085(.A(KEYINPUT70), .B(G88), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n505), .A2(G50), .A3(G543), .ZN(new_n513));
  XNOR2_X1  g088(.A(new_n513), .B(KEYINPUT68), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n506), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  OR2_X1    g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n512), .A2(new_n514), .A3(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(new_n518), .ZN(G166));
  XOR2_X1   g094(.A(KEYINPUT72), .B(G89), .Z(new_n520));
  NAND2_X1  g095(.A1(new_n510), .A2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(new_n521), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n506), .A2(G63), .A3(G651), .ZN(new_n523));
  XNOR2_X1  g098(.A(new_n523), .B(KEYINPUT71), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n505), .A2(G543), .ZN(new_n525));
  INV_X1    g100(.A(new_n525), .ZN(new_n526));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(KEYINPUT7), .ZN(new_n528));
  OR2_X1    g103(.A1(new_n527), .A2(KEYINPUT7), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n526), .A2(G51), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n524), .A2(new_n530), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n522), .A2(new_n531), .ZN(G168));
  XNOR2_X1  g107(.A(KEYINPUT73), .B(G90), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n510), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(G77), .A2(G543), .ZN(new_n535));
  XOR2_X1   g110(.A(KEYINPUT5), .B(G543), .Z(new_n536));
  INV_X1    g111(.A(G64), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n535), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n538), .A2(G651), .B1(new_n526), .B2(G52), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n534), .A2(new_n539), .ZN(G301));
  INV_X1    g115(.A(G301), .ZN(G171));
  NAND2_X1  g116(.A1(new_n510), .A2(G81), .ZN(new_n542));
  NAND2_X1  g117(.A1(G68), .A2(G543), .ZN(new_n543));
  INV_X1    g118(.A(G56), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n543), .B1(new_n536), .B2(new_n544), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n545), .A2(G651), .B1(new_n526), .B2(G43), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n542), .A2(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  NAND4_X1  g124(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT8), .ZN(new_n552));
  NAND4_X1  g127(.A1(G319), .A2(G483), .A3(G661), .A4(new_n552), .ZN(G188));
  INV_X1    g128(.A(KEYINPUT9), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n526), .A2(new_n554), .A3(G53), .ZN(new_n555));
  INV_X1    g130(.A(G53), .ZN(new_n556));
  OAI21_X1  g131(.A(KEYINPUT9), .B1(new_n525), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n506), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n559));
  OR2_X1    g134(.A1(new_n559), .A2(new_n516), .ZN(new_n560));
  AND2_X1   g135(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT74), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n562), .B1(new_n508), .B2(new_n509), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n505), .A2(new_n506), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(KEYINPUT69), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n505), .A2(new_n506), .A3(new_n507), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n565), .A2(KEYINPUT74), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n563), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G91), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n561), .A2(new_n569), .ZN(G299));
  INV_X1    g145(.A(new_n531), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(new_n521), .ZN(G286));
  INV_X1    g147(.A(KEYINPUT75), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n518), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g149(.A1(new_n512), .A2(KEYINPUT75), .A3(new_n514), .A4(new_n517), .ZN(new_n575));
  AND2_X1   g150(.A1(new_n574), .A2(new_n575), .ZN(G303));
  NAND2_X1  g151(.A1(new_n568), .A2(G87), .ZN(new_n577));
  OR2_X1    g152(.A1(new_n506), .A2(G74), .ZN(new_n578));
  AOI22_X1  g153(.A1(G49), .A2(new_n526), .B1(new_n578), .B2(G651), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n577), .A2(new_n579), .ZN(G288));
  INV_X1    g155(.A(G86), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n581), .B1(new_n563), .B2(new_n567), .ZN(new_n582));
  NAND2_X1  g157(.A1(G73), .A2(G543), .ZN(new_n583));
  INV_X1    g158(.A(G61), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n536), .B2(new_n584), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n585), .A2(G651), .B1(new_n526), .B2(G48), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n582), .A2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(G305));
  NAND2_X1  g164(.A1(new_n526), .A2(G47), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n506), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n565), .A2(new_n566), .ZN(new_n592));
  INV_X1    g167(.A(G85), .ZN(new_n593));
  OAI221_X1 g168(.A(new_n590), .B1(new_n516), .B2(new_n591), .C1(new_n592), .C2(new_n593), .ZN(G290));
  NAND2_X1  g169(.A1(G301), .A2(G868), .ZN(new_n595));
  XOR2_X1   g170(.A(KEYINPUT76), .B(G66), .Z(new_n596));
  AOI22_X1  g171(.A1(new_n596), .A2(new_n506), .B1(G79), .B2(G543), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n598), .A2(G651), .B1(new_n526), .B2(G54), .ZN(new_n599));
  AND3_X1   g174(.A1(new_n568), .A2(KEYINPUT10), .A3(G92), .ZN(new_n600));
  AOI21_X1  g175(.A(KEYINPUT10), .B1(new_n568), .B2(G92), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n599), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(new_n602), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n595), .B1(new_n603), .B2(G868), .ZN(G284));
  OAI21_X1  g179(.A(new_n595), .B1(new_n603), .B2(G868), .ZN(G321));
  INV_X1    g180(.A(G868), .ZN(new_n606));
  NOR2_X1   g181(.A1(G168), .A2(new_n606), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n607), .B(KEYINPUT77), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n558), .A2(new_n560), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n609), .B1(new_n568), .B2(G91), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n608), .B1(G868), .B2(new_n610), .ZN(G297));
  OAI21_X1  g186(.A(new_n608), .B1(G868), .B2(new_n610), .ZN(G280));
  INV_X1    g187(.A(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n603), .B1(new_n613), .B2(G860), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT78), .ZN(G148));
  NOR2_X1   g190(.A1(new_n548), .A2(G868), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n603), .A2(new_n613), .ZN(new_n617));
  AOI21_X1  g192(.A(new_n616), .B1(new_n617), .B2(G868), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT79), .ZN(G323));
  XOR2_X1   g194(.A(KEYINPUT80), .B(KEYINPUT11), .Z(new_n620));
  XNOR2_X1  g195(.A(G323), .B(new_n620), .ZN(G282));
  NAND2_X1  g196(.A1(new_n483), .A2(new_n471), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT12), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT13), .ZN(new_n624));
  INV_X1    g199(.A(G2100), .ZN(new_n625));
  OR2_X1    g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n624), .A2(new_n625), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n480), .A2(G123), .ZN(new_n628));
  NOR2_X1   g203(.A1(new_n463), .A2(G111), .ZN(new_n629));
  OAI21_X1  g204(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n630));
  INV_X1    g205(.A(G135), .ZN(new_n631));
  OAI221_X1 g206(.A(new_n628), .B1(new_n629), .B2(new_n630), .C1(new_n631), .C2(new_n484), .ZN(new_n632));
  XOR2_X1   g207(.A(new_n632), .B(G2096), .Z(new_n633));
  NAND3_X1  g208(.A1(new_n626), .A2(new_n627), .A3(new_n633), .ZN(G156));
  XOR2_X1   g209(.A(G2451), .B(G2454), .Z(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT16), .ZN(new_n636));
  XNOR2_X1  g211(.A(G1341), .B(G1348), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  INV_X1    g213(.A(KEYINPUT14), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2427), .B(G2438), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2430), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT15), .B(G2435), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n639), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n643), .B1(new_n642), .B2(new_n641), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n638), .B(new_n644), .Z(new_n645));
  XNOR2_X1  g220(.A(G2443), .B(G2446), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n645), .A2(new_n646), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n647), .A2(new_n648), .A3(G14), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT81), .ZN(G401));
  XNOR2_X1  g225(.A(G2067), .B(G2678), .ZN(new_n651));
  NOR2_X1   g226(.A1(G2072), .A2(G2078), .ZN(new_n652));
  NOR2_X1   g227(.A1(new_n444), .A2(new_n652), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  AOI21_X1  g229(.A(new_n651), .B1(new_n654), .B2(KEYINPUT82), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n655), .B1(KEYINPUT82), .B2(new_n654), .ZN(new_n656));
  XOR2_X1   g231(.A(G2084), .B(G2090), .Z(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n653), .B(KEYINPUT17), .ZN(new_n659));
  INV_X1    g234(.A(new_n651), .ZN(new_n660));
  OAI211_X1 g235(.A(new_n656), .B(new_n658), .C1(new_n659), .C2(new_n660), .ZN(new_n661));
  NOR3_X1   g236(.A1(new_n658), .A2(new_n653), .A3(new_n660), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT18), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n659), .A2(new_n660), .A3(new_n657), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n661), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(G2096), .B(G2100), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(G227));
  XOR2_X1   g242(.A(G1971), .B(G1976), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT19), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1956), .B(G2474), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1961), .B(G1966), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT20), .ZN(new_n674));
  AND2_X1   g249(.A1(new_n670), .A2(new_n671), .ZN(new_n675));
  NOR3_X1   g250(.A1(new_n669), .A2(new_n672), .A3(new_n675), .ZN(new_n676));
  AOI21_X1  g251(.A(new_n676), .B1(new_n669), .B2(new_n675), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT83), .ZN(new_n680));
  XOR2_X1   g255(.A(new_n678), .B(new_n680), .Z(new_n681));
  XNOR2_X1  g256(.A(G1991), .B(G1996), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1981), .B(G1986), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(G229));
  INV_X1    g261(.A(G16), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n687), .A2(G22), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n688), .B1(G166), .B2(new_n687), .ZN(new_n689));
  INV_X1    g264(.A(G1971), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT32), .B(G1981), .Z(new_n692));
  NOR2_X1   g267(.A1(new_n588), .A2(new_n687), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n693), .B1(G6), .B2(new_n687), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n691), .B1(new_n692), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n694), .A2(new_n692), .ZN(new_n696));
  AND2_X1   g271(.A1(new_n687), .A2(G23), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n697), .B1(G288), .B2(G16), .ZN(new_n698));
  XOR2_X1   g273(.A(KEYINPUT33), .B(G1976), .Z(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n696), .A2(new_n701), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n698), .A2(new_n700), .ZN(new_n703));
  NOR3_X1   g278(.A1(new_n695), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(KEYINPUT34), .ZN(new_n705));
  OR2_X1    g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  XOR2_X1   g281(.A(KEYINPUT84), .B(G29), .Z(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n708), .A2(G25), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n485), .A2(G131), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n480), .A2(G119), .ZN(new_n711));
  OR2_X1    g286(.A1(G95), .A2(G2105), .ZN(new_n712));
  OAI211_X1 g287(.A(new_n712), .B(G2104), .C1(G107), .C2(new_n463), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n710), .A2(new_n711), .A3(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(new_n714), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n709), .B1(new_n715), .B2(new_n708), .ZN(new_n716));
  XOR2_X1   g291(.A(KEYINPUT35), .B(G1991), .Z(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  MUX2_X1   g293(.A(G24), .B(G290), .S(G16), .Z(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(G1986), .Z(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n718), .B1(new_n721), .B2(KEYINPUT85), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(KEYINPUT85), .B2(new_n721), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n704), .A2(new_n705), .ZN(new_n724));
  NAND3_X1  g299(.A1(new_n706), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n725), .B(KEYINPUT36), .Z(new_n726));
  NOR2_X1   g301(.A1(new_n708), .A2(G35), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(G162), .B2(new_n708), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT29), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n729), .A2(G2090), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT95), .ZN(new_n731));
  NAND3_X1  g306(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT88), .ZN(new_n733));
  INV_X1    g308(.A(KEYINPUT26), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n733), .B(new_n734), .ZN(new_n735));
  AOI22_X1  g310(.A1(new_n480), .A2(G129), .B1(G105), .B2(new_n471), .ZN(new_n736));
  INV_X1    g311(.A(G141), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n736), .B1(new_n737), .B2(new_n484), .ZN(new_n738));
  OR3_X1    g313(.A1(new_n735), .A2(new_n738), .A3(KEYINPUT89), .ZN(new_n739));
  OAI21_X1  g314(.A(KEYINPUT89), .B1(new_n735), .B2(new_n738), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(G29), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(new_n743), .B2(G32), .ZN(new_n745));
  XNOR2_X1  g320(.A(KEYINPUT27), .B(G1996), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT90), .ZN(new_n748));
  NOR2_X1   g323(.A1(G4), .A2(G16), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(new_n603), .B2(G16), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n750), .A2(G1348), .ZN(new_n751));
  NAND3_X1  g326(.A1(new_n731), .A2(new_n748), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n687), .A2(G20), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT23), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(new_n610), .B2(new_n687), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(G1956), .ZN(new_n756));
  NAND2_X1  g331(.A1(G168), .A2(G16), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT91), .ZN(new_n758));
  OAI211_X1 g333(.A(new_n757), .B(new_n758), .C1(G16), .C2(G21), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(new_n758), .B2(new_n757), .ZN(new_n760));
  OR2_X1    g335(.A1(new_n760), .A2(G1966), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n708), .A2(G27), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(G164), .B2(new_n708), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(new_n443), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n760), .A2(G1966), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n687), .A2(G19), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(new_n548), .B2(new_n687), .ZN(new_n767));
  INV_X1    g342(.A(G1341), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n767), .B(new_n768), .ZN(new_n769));
  NAND4_X1  g344(.A1(new_n761), .A2(new_n764), .A3(new_n765), .A4(new_n769), .ZN(new_n770));
  NOR2_X1   g345(.A1(G171), .A2(new_n687), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(G5), .B2(new_n687), .ZN(new_n772));
  INV_X1    g347(.A(G1961), .ZN(new_n773));
  INV_X1    g348(.A(KEYINPUT87), .ZN(new_n774));
  XNOR2_X1  g349(.A(KEYINPUT24), .B(G34), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n707), .A2(new_n775), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(KEYINPUT86), .Z(new_n777));
  INV_X1    g352(.A(G160), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n777), .B1(new_n743), .B2(new_n778), .ZN(new_n779));
  INV_X1    g354(.A(G2084), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  AOI22_X1  g356(.A1(new_n772), .A2(new_n773), .B1(new_n774), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n707), .A2(G26), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT28), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n485), .A2(G140), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n480), .A2(G128), .ZN(new_n786));
  OR2_X1    g361(.A1(G104), .A2(G2105), .ZN(new_n787));
  OAI211_X1 g362(.A(new_n787), .B(G2104), .C1(G116), .C2(new_n463), .ZN(new_n788));
  NAND3_X1  g363(.A1(new_n785), .A2(new_n786), .A3(new_n788), .ZN(new_n789));
  INV_X1    g364(.A(new_n789), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n784), .B1(new_n790), .B2(new_n743), .ZN(new_n791));
  INV_X1    g366(.A(G2067), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n782), .A2(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n632), .A2(new_n707), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n795), .A2(KEYINPUT92), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n795), .A2(KEYINPUT92), .ZN(new_n797));
  XNOR2_X1  g372(.A(KEYINPUT31), .B(G11), .ZN(new_n798));
  XOR2_X1   g373(.A(KEYINPUT93), .B(G28), .Z(new_n799));
  NOR2_X1   g374(.A1(new_n799), .A2(KEYINPUT30), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n799), .A2(KEYINPUT30), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n801), .A2(new_n743), .ZN(new_n802));
  OAI211_X1 g377(.A(new_n797), .B(new_n798), .C1(new_n800), .C2(new_n802), .ZN(new_n803));
  AOI211_X1 g378(.A(new_n796), .B(new_n803), .C1(new_n780), .C2(new_n779), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n743), .A2(G33), .ZN(new_n805));
  NAND3_X1  g380(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n806));
  XOR2_X1   g381(.A(new_n806), .B(KEYINPUT25), .Z(new_n807));
  INV_X1    g382(.A(G139), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n807), .B1(new_n808), .B2(new_n484), .ZN(new_n809));
  AOI22_X1  g384(.A1(new_n483), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n810), .A2(new_n463), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n805), .B1(new_n812), .B2(new_n743), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(new_n442), .ZN(new_n814));
  OAI211_X1 g389(.A(new_n804), .B(new_n814), .C1(new_n774), .C2(new_n781), .ZN(new_n815));
  OR4_X1    g390(.A1(new_n756), .A2(new_n770), .A3(new_n794), .A4(new_n815), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n772), .A2(new_n773), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT94), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n818), .B1(new_n729), .B2(G2090), .ZN(new_n819));
  OAI221_X1 g394(.A(new_n819), .B1(G1348), .B2(new_n750), .C1(new_n745), .C2(new_n746), .ZN(new_n820));
  NOR4_X1   g395(.A1(new_n726), .A2(new_n752), .A3(new_n816), .A4(new_n820), .ZN(G311));
  OR4_X1    g396(.A1(new_n726), .A2(new_n752), .A3(new_n816), .A4(new_n820), .ZN(G150));
  NAND2_X1  g397(.A1(new_n526), .A2(G55), .ZN(new_n823));
  INV_X1    g398(.A(G93), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n823), .B1(new_n592), .B2(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT96), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(new_n827));
  AOI22_X1  g402(.A1(new_n506), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n828));
  OR2_X1    g403(.A1(new_n828), .A2(new_n516), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n830), .A2(G860), .ZN(new_n831));
  XOR2_X1   g406(.A(new_n831), .B(KEYINPUT37), .Z(new_n832));
  NAND2_X1  g407(.A1(new_n603), .A2(G559), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT38), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n830), .A2(new_n547), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n827), .A2(new_n548), .A3(new_n829), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  OR2_X1    g412(.A1(new_n834), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n834), .A2(new_n837), .ZN(new_n839));
  AOI21_X1  g414(.A(KEYINPUT39), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n840), .A2(G860), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n838), .A2(new_n839), .A3(KEYINPUT39), .ZN(new_n842));
  AND3_X1   g417(.A1(new_n841), .A2(KEYINPUT97), .A3(new_n842), .ZN(new_n843));
  AOI21_X1  g418(.A(KEYINPUT97), .B1(new_n841), .B2(new_n842), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n832), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT98), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  OAI211_X1 g422(.A(KEYINPUT98), .B(new_n832), .C1(new_n843), .C2(new_n844), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n847), .A2(new_n848), .ZN(G145));
  XNOR2_X1  g424(.A(KEYINPUT101), .B(G37), .ZN(new_n850));
  INV_X1    g425(.A(new_n850), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n741), .A2(new_n789), .ZN(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n790), .B1(new_n739), .B2(new_n740), .ZN(new_n854));
  INV_X1    g429(.A(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT99), .ZN(new_n856));
  AND3_X1   g431(.A1(new_n499), .A2(new_n856), .A3(new_n501), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n856), .B1(new_n499), .B2(new_n501), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n495), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n859), .A2(KEYINPUT100), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT100), .ZN(new_n861));
  OAI211_X1 g436(.A(new_n861), .B(new_n495), .C1(new_n857), .C2(new_n858), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n853), .A2(new_n855), .A3(new_n863), .ZN(new_n864));
  OAI211_X1 g439(.A(new_n860), .B(new_n862), .C1(new_n852), .C2(new_n854), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n866), .B1(new_n811), .B2(new_n809), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n864), .A2(new_n865), .A3(new_n812), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n480), .A2(G130), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n463), .A2(G118), .ZN(new_n871));
  OAI21_X1  g446(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n870), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n873), .B1(G142), .B2(new_n485), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(new_n623), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(new_n715), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n869), .A2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n876), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n867), .A2(new_n878), .A3(new_n868), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n778), .B(new_n632), .ZN(new_n881));
  XOR2_X1   g456(.A(G162), .B(new_n881), .Z(new_n882));
  AOI21_X1  g457(.A(new_n851), .B1(new_n880), .B2(new_n882), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n869), .A2(KEYINPUT102), .A3(new_n876), .ZN(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(KEYINPUT102), .B1(new_n869), .B2(new_n876), .ZN(new_n886));
  INV_X1    g461(.A(new_n882), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n879), .A2(new_n887), .ZN(new_n888));
  NOR4_X1   g463(.A1(new_n885), .A2(new_n886), .A3(new_n888), .A4(KEYINPUT103), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT103), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n886), .A2(new_n888), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n890), .B1(new_n891), .B2(new_n884), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n883), .B1(new_n889), .B2(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n893), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g469(.A1(new_n830), .A2(new_n606), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n837), .B(new_n617), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n603), .A2(new_n610), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n602), .A2(G299), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n896), .A2(new_n899), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n899), .A2(KEYINPUT41), .ZN(new_n901));
  XOR2_X1   g476(.A(KEYINPUT104), .B(KEYINPUT41), .Z(new_n902));
  AOI21_X1  g477(.A(new_n902), .B1(new_n897), .B2(new_n898), .ZN(new_n903));
  OAI21_X1  g478(.A(KEYINPUT105), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n904), .B1(KEYINPUT105), .B2(new_n903), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n900), .B1(new_n905), .B2(new_n896), .ZN(new_n906));
  XNOR2_X1  g481(.A(G288), .B(new_n588), .ZN(new_n907));
  XNOR2_X1  g482(.A(G290), .B(new_n518), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n907), .B(new_n908), .ZN(new_n909));
  XOR2_X1   g484(.A(new_n909), .B(KEYINPUT42), .Z(new_n910));
  NOR2_X1   g485(.A1(new_n910), .A2(KEYINPUT106), .ZN(new_n911));
  OR2_X1    g486(.A1(new_n906), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n906), .A2(new_n911), .ZN(new_n913));
  AOI22_X1  g488(.A1(new_n912), .A2(new_n913), .B1(KEYINPUT106), .B2(new_n910), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n895), .B1(new_n914), .B2(new_n606), .ZN(G295));
  OAI21_X1  g490(.A(new_n895), .B1(new_n914), .B2(new_n606), .ZN(G331));
  NOR3_X1   g491(.A1(new_n522), .A2(new_n531), .A3(KEYINPUT107), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(G286), .A2(KEYINPUT107), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n918), .A2(new_n919), .A3(G171), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT107), .ZN(new_n921));
  NOR2_X1   g496(.A1(G168), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g497(.A(G301), .B1(new_n922), .B2(new_n917), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n920), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n837), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(KEYINPUT108), .ZN(new_n926));
  OR2_X1    g501(.A1(new_n837), .A2(new_n924), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT108), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n837), .A2(new_n924), .A3(new_n928), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n926), .A2(new_n927), .A3(new_n929), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n899), .A2(new_n902), .ZN(new_n931));
  AOI21_X1  g506(.A(KEYINPUT41), .B1(new_n897), .B2(new_n898), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  AND2_X1   g508(.A1(new_n930), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n837), .A2(new_n924), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n935), .A2(new_n899), .ZN(new_n936));
  AND2_X1   g511(.A1(new_n936), .A2(new_n925), .ZN(new_n937));
  OAI211_X1 g512(.A(KEYINPUT109), .B(new_n909), .C1(new_n934), .C2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT109), .ZN(new_n939));
  AOI22_X1  g514(.A1(new_n930), .A2(new_n933), .B1(new_n936), .B2(new_n925), .ZN(new_n940));
  INV_X1    g515(.A(new_n909), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n939), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n938), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n927), .A2(new_n925), .ZN(new_n944));
  AND2_X1   g519(.A1(new_n926), .A2(new_n929), .ZN(new_n945));
  AOI22_X1  g520(.A1(new_n905), .A2(new_n944), .B1(new_n936), .B2(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n851), .B1(new_n946), .B2(new_n941), .ZN(new_n947));
  AND3_X1   g522(.A1(new_n943), .A2(new_n947), .A3(KEYINPUT43), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n945), .A2(new_n936), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n903), .A2(KEYINPUT105), .ZN(new_n950));
  INV_X1    g525(.A(new_n950), .ZN(new_n951));
  AND2_X1   g526(.A1(new_n904), .A2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(new_n944), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n949), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(G37), .B1(new_n954), .B2(new_n909), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n946), .A2(new_n941), .ZN(new_n956));
  AOI21_X1  g531(.A(KEYINPUT43), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  OAI21_X1  g532(.A(KEYINPUT44), .B1(new_n948), .B2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT44), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT43), .ZN(new_n960));
  AND3_X1   g535(.A1(new_n943), .A2(new_n947), .A3(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n960), .B1(new_n955), .B2(new_n956), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n959), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n958), .A2(new_n963), .ZN(G397));
  INV_X1    g539(.A(KEYINPUT126), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT51), .ZN(new_n966));
  INV_X1    g541(.A(G1966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT110), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n968), .B1(G160), .B2(G40), .ZN(new_n969));
  AND2_X1   g544(.A1(new_n469), .A2(new_n472), .ZN(new_n970));
  INV_X1    g545(.A(G125), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n971), .B1(new_n478), .B2(new_n479), .ZN(new_n972));
  INV_X1    g547(.A(new_n467), .ZN(new_n973));
  OAI21_X1  g548(.A(G2105), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  AND4_X1   g549(.A1(new_n968), .A2(new_n970), .A3(new_n974), .A4(G40), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n969), .A2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(G1384), .ZN(new_n977));
  INV_X1    g552(.A(new_n501), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n500), .B1(new_n483), .B2(new_n497), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n483), .A2(G126), .A3(G2105), .ZN(new_n981));
  AOI21_X1  g556(.A(KEYINPUT67), .B1(new_n488), .B2(new_n490), .ZN(new_n982));
  NOR3_X1   g557(.A1(new_n493), .A2(new_n487), .A3(new_n492), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n981), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  OAI211_X1 g559(.A(KEYINPUT45), .B(new_n977), .C1(new_n980), .C2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n976), .A2(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(KEYINPUT45), .B1(new_n859), .B2(new_n977), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n967), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT50), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n859), .A2(new_n989), .A3(new_n977), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n503), .A2(new_n977), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(KEYINPUT50), .ZN(new_n992));
  XOR2_X1   g567(.A(KEYINPUT114), .B(G2084), .Z(new_n993));
  NAND4_X1  g568(.A1(new_n990), .A2(new_n976), .A3(new_n992), .A4(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n988), .A2(new_n994), .ZN(new_n995));
  OAI211_X1 g570(.A(new_n966), .B(G8), .C1(new_n995), .C2(G286), .ZN(new_n996));
  INV_X1    g571(.A(new_n994), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n970), .A2(new_n974), .A3(G40), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(KEYINPUT110), .ZN(new_n999));
  NAND3_X1  g574(.A1(G160), .A2(new_n968), .A3(G40), .ZN(new_n1000));
  AND3_X1   g575(.A1(new_n985), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT45), .ZN(new_n1002));
  OAI21_X1  g577(.A(KEYINPUT99), .B1(new_n978), .B2(new_n979), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n499), .A2(new_n856), .A3(new_n501), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n984), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1002), .B1(new_n1005), .B2(G1384), .ZN(new_n1006));
  AOI21_X1  g581(.A(G1966), .B1(new_n1001), .B2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g582(.A(G8), .B1(new_n997), .B2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(G286), .A2(G8), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1008), .A2(KEYINPUT51), .A3(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT123), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1009), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1011), .B1(new_n995), .B2(new_n1012), .ZN(new_n1013));
  AOI211_X1 g588(.A(KEYINPUT123), .B(new_n1009), .C1(new_n988), .C2(new_n994), .ZN(new_n1014));
  OAI211_X1 g589(.A(new_n996), .B(new_n1010), .C1(new_n1013), .C2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(G8), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n1005), .A2(G1384), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1016), .B1(new_n1017), .B2(new_n976), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n577), .A2(G1976), .A3(new_n579), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(KEYINPUT52), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT49), .ZN(new_n1022));
  NOR3_X1   g597(.A1(new_n582), .A2(new_n587), .A3(G1981), .ZN(new_n1023));
  INV_X1    g598(.A(G1981), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n510), .A2(G86), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1024), .B1(new_n1025), .B2(new_n586), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1022), .B1(new_n1023), .B2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n568), .A2(G86), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1028), .A2(new_n1024), .A3(new_n586), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1026), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1029), .A2(KEYINPUT49), .A3(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1027), .A2(new_n1031), .A3(new_n1018), .ZN(new_n1032));
  INV_X1    g607(.A(G1976), .ZN(new_n1033));
  AOI21_X1  g608(.A(KEYINPUT52), .B1(G288), .B2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1034), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1021), .A2(new_n1032), .A3(new_n1035), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n989), .B1(new_n859), .B2(new_n977), .ZN(new_n1037));
  OAI211_X1 g612(.A(new_n989), .B(new_n977), .C1(new_n980), .C2(new_n984), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1038), .A2(new_n999), .A3(new_n1000), .ZN(new_n1039));
  OAI21_X1  g614(.A(KEYINPUT113), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g615(.A(KEYINPUT50), .B1(new_n1005), .B2(G1384), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT113), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n1041), .A2(new_n1042), .A3(new_n976), .A4(new_n1038), .ZN(new_n1043));
  INV_X1    g618(.A(G2090), .ZN(new_n1044));
  AND3_X1   g619(.A1(new_n1040), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n999), .A2(new_n1000), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT111), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n991), .A2(new_n1047), .A3(new_n1002), .ZN(new_n1048));
  AOI21_X1  g623(.A(G1384), .B1(new_n495), .B2(new_n502), .ZN(new_n1049));
  OAI21_X1  g624(.A(KEYINPUT111), .B1(new_n1049), .B2(KEYINPUT45), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1046), .B1(new_n1048), .B2(new_n1050), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n860), .A2(KEYINPUT45), .A3(new_n977), .A4(new_n862), .ZN(new_n1052));
  AOI21_X1  g627(.A(G1971), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g628(.A(G8), .B1(new_n1045), .B2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n574), .A2(G8), .A3(new_n575), .ZN(new_n1055));
  XNOR2_X1  g630(.A(new_n1055), .B(KEYINPUT55), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1036), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1057));
  XOR2_X1   g632(.A(new_n1055), .B(KEYINPUT55), .Z(new_n1058));
  NAND3_X1  g633(.A1(new_n990), .A2(new_n976), .A3(new_n992), .ZN(new_n1059));
  OAI22_X1  g634(.A1(new_n1053), .A2(KEYINPUT112), .B1(G2090), .B2(new_n1059), .ZN(new_n1060));
  AND2_X1   g635(.A1(new_n1053), .A2(KEYINPUT112), .ZN(new_n1061));
  OAI211_X1 g636(.A(new_n1058), .B(G8), .C1(new_n1060), .C2(new_n1061), .ZN(new_n1062));
  AND3_X1   g637(.A1(new_n1015), .A2(new_n1057), .A3(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1051), .A2(new_n1052), .A3(new_n443), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT53), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1059), .A2(new_n773), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n860), .A2(new_n977), .A3(new_n862), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(new_n1002), .ZN(new_n1069));
  NOR3_X1   g644(.A1(new_n998), .A2(new_n1065), .A3(G2078), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1069), .A2(new_n1052), .A3(new_n1070), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1066), .A2(G301), .A3(new_n1067), .A4(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(KEYINPUT124), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1001), .A2(KEYINPUT53), .A3(new_n1006), .A4(new_n443), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1066), .A2(new_n1067), .A3(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(G171), .ZN(new_n1076));
  AOI22_X1  g651(.A1(new_n1064), .A2(new_n1065), .B1(new_n773), .B2(new_n1059), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT124), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1077), .A2(new_n1078), .A3(G301), .A4(new_n1071), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1073), .A2(new_n1076), .A3(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT54), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1066), .A2(new_n1067), .A3(new_n1071), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT125), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1077), .A2(KEYINPUT125), .A3(new_n1071), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1085), .A2(G171), .A3(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1075), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1081), .B1(new_n1088), .B2(G301), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1063), .A2(new_n1082), .A3(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT122), .ZN(new_n1092));
  INV_X1    g667(.A(G1348), .ZN(new_n1093));
  NOR3_X1   g668(.A1(new_n1046), .A2(G1384), .A3(new_n1005), .ZN(new_n1094));
  AOI22_X1  g669(.A1(new_n1059), .A2(new_n1093), .B1(new_n1094), .B2(new_n792), .ZN(new_n1095));
  OAI211_X1 g670(.A(new_n603), .B(new_n1092), .C1(new_n1095), .C2(KEYINPUT60), .ZN(new_n1096));
  NOR3_X1   g671(.A1(new_n1005), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1097));
  OAI211_X1 g672(.A(new_n999), .B(new_n1000), .C1(new_n1049), .C2(new_n989), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1093), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1017), .A2(new_n976), .A3(new_n792), .ZN(new_n1100));
  AOI21_X1  g675(.A(KEYINPUT60), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  OAI21_X1  g676(.A(KEYINPUT122), .B1(new_n1101), .B2(new_n602), .ZN(new_n1102));
  AND2_X1   g677(.A1(new_n1095), .A2(KEYINPUT60), .ZN(new_n1103));
  AND3_X1   g678(.A1(new_n1096), .A2(new_n1102), .A3(new_n1103), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1103), .B1(new_n1096), .B2(new_n1102), .ZN(new_n1105));
  OR2_X1    g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT57), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n610), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(KEYINPUT117), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT117), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1108), .A2(new_n1109), .A3(new_n1112), .ZN(new_n1113));
  AND2_X1   g688(.A1(new_n1111), .A2(new_n1113), .ZN(new_n1114));
  XNOR2_X1  g689(.A(KEYINPUT56), .B(G2072), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1051), .A2(new_n1052), .A3(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(KEYINPUT116), .ZN(new_n1117));
  INV_X1    g692(.A(G1956), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1118), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT116), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1051), .A2(new_n1052), .A3(new_n1120), .A4(new_n1115), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1117), .A2(new_n1119), .A3(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1114), .A2(new_n1122), .ZN(new_n1123));
  AND2_X1   g698(.A1(new_n1121), .A2(new_n1119), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1124), .A2(new_n1117), .A3(new_n1109), .A4(new_n1108), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1123), .A2(new_n1125), .A3(KEYINPUT61), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1122), .A2(new_n1110), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1125), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT61), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT59), .ZN(new_n1131));
  OAI21_X1  g706(.A(KEYINPUT121), .B1(new_n1131), .B2(KEYINPUT120), .ZN(new_n1132));
  XNOR2_X1  g707(.A(KEYINPUT119), .B(KEYINPUT58), .ZN(new_n1133));
  XNOR2_X1  g708(.A(new_n1133), .B(G1341), .ZN(new_n1134));
  OR2_X1    g709(.A1(new_n1094), .A2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(G1996), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1051), .A2(new_n1052), .A3(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1132), .B1(new_n1138), .B2(new_n548), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1132), .B1(KEYINPUT121), .B2(new_n1131), .ZN(new_n1140));
  AOI211_X1 g715(.A(new_n547), .B(new_n1140), .C1(new_n1135), .C2(new_n1137), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1106), .A2(new_n1126), .A3(new_n1130), .A4(new_n1142), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1095), .A2(new_n602), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1144), .B1(new_n1114), .B2(new_n1122), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1122), .A2(new_n1110), .ZN(new_n1146));
  OAI21_X1  g721(.A(KEYINPUT118), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT118), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1111), .A2(new_n1113), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1149), .B1(new_n1117), .B2(new_n1124), .ZN(new_n1150));
  OAI211_X1 g725(.A(new_n1148), .B(new_n1125), .C1(new_n1150), .C2(new_n1144), .ZN(new_n1151));
  AND2_X1   g726(.A1(new_n1147), .A2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1091), .B1(new_n1143), .B2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n995), .A2(G8), .A3(G168), .ZN(new_n1154));
  XOR2_X1   g729(.A(new_n1154), .B(KEYINPUT115), .Z(new_n1155));
  OAI21_X1  g730(.A(G8), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1156), .A2(new_n1056), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT63), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n1036), .A2(new_n1158), .ZN(new_n1159));
  NAND4_X1  g734(.A1(new_n1155), .A2(new_n1157), .A3(new_n1062), .A4(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1057), .A2(new_n1062), .ZN(new_n1161));
  XNOR2_X1  g736(.A(new_n1154), .B(KEYINPUT115), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1158), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1160), .A2(new_n1163), .ZN(new_n1164));
  NAND4_X1  g739(.A1(new_n1032), .A2(new_n1033), .A3(new_n577), .A4(new_n579), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1165), .A2(new_n1029), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1166), .A2(new_n1018), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1167), .B1(new_n1062), .B2(new_n1036), .ZN(new_n1168));
  INV_X1    g743(.A(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1164), .A2(new_n1169), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n965), .B1(new_n1153), .B2(new_n1170), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1168), .B1(new_n1160), .B2(new_n1163), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1147), .A2(new_n1151), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1142), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1174));
  AOI21_X1  g749(.A(KEYINPUT61), .B1(new_n1125), .B2(new_n1127), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1173), .B1(new_n1176), .B2(new_n1126), .ZN(new_n1177));
  OAI211_X1 g752(.A(KEYINPUT126), .B(new_n1172), .C1(new_n1177), .C2(new_n1091), .ZN(new_n1178));
  INV_X1    g753(.A(new_n1161), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1076), .B1(new_n1015), .B2(KEYINPUT62), .ZN(new_n1180));
  OAI211_X1 g755(.A(new_n1179), .B(new_n1180), .C1(KEYINPUT62), .C2(new_n1015), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1171), .A2(new_n1178), .A3(new_n1181), .ZN(new_n1182));
  NOR2_X1   g757(.A1(new_n1069), .A2(new_n1046), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n742), .A2(new_n1136), .ZN(new_n1184));
  XNOR2_X1  g759(.A(new_n789), .B(new_n792), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n741), .A2(G1996), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n1184), .A2(new_n1185), .A3(new_n1186), .ZN(new_n1187));
  INV_X1    g762(.A(new_n1187), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n715), .A2(new_n717), .ZN(new_n1189));
  OR2_X1    g764(.A1(new_n715), .A2(new_n717), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1188), .A2(new_n1189), .A3(new_n1190), .ZN(new_n1191));
  XNOR2_X1  g766(.A(G290), .B(G1986), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n1183), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1182), .A2(new_n1193), .ZN(new_n1194));
  NOR2_X1   g769(.A1(G290), .A2(G1986), .ZN(new_n1195));
  AOI21_X1  g770(.A(KEYINPUT48), .B1(new_n1183), .B2(new_n1195), .ZN(new_n1196));
  AND3_X1   g771(.A1(new_n1183), .A2(KEYINPUT48), .A3(new_n1195), .ZN(new_n1197));
  AOI211_X1 g772(.A(new_n1196), .B(new_n1197), .C1(new_n1191), .C2(new_n1183), .ZN(new_n1198));
  INV_X1    g773(.A(new_n1185), .ZN(new_n1199));
  OAI21_X1  g774(.A(new_n1183), .B1(new_n741), .B2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1183), .A2(new_n1136), .ZN(new_n1201));
  AND2_X1   g776(.A1(new_n1201), .A2(KEYINPUT46), .ZN(new_n1202));
  NOR2_X1   g777(.A1(new_n1201), .A2(KEYINPUT46), .ZN(new_n1203));
  OAI21_X1  g778(.A(new_n1200), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  XOR2_X1   g779(.A(new_n1204), .B(KEYINPUT47), .Z(new_n1205));
  OAI22_X1  g780(.A1(new_n1187), .A2(new_n1189), .B1(G2067), .B2(new_n789), .ZN(new_n1206));
  AOI211_X1 g781(.A(new_n1198), .B(new_n1205), .C1(new_n1183), .C2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1194), .A2(new_n1207), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g783(.A(G319), .ZN(new_n1210));
  NOR2_X1   g784(.A1(G227), .A2(new_n1210), .ZN(new_n1211));
  XNOR2_X1  g785(.A(new_n1211), .B(KEYINPUT127), .ZN(new_n1212));
  NOR3_X1   g786(.A1(G229), .A2(G401), .A3(new_n1212), .ZN(new_n1213));
  OAI211_X1 g787(.A(new_n893), .B(new_n1213), .C1(new_n961), .C2(new_n962), .ZN(G225));
  INV_X1    g788(.A(G225), .ZN(G308));
endmodule


