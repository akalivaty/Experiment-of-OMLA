

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586;

  INV_X1 U321 ( .A(KEYINPUT94), .ZN(n401) );
  XNOR2_X1 U322 ( .A(n331), .B(n299), .ZN(n300) );
  XNOR2_X1 U323 ( .A(n477), .B(KEYINPUT48), .ZN(n478) );
  XNOR2_X1 U324 ( .A(n408), .B(n407), .ZN(n410) );
  XNOR2_X1 U325 ( .A(n402), .B(n401), .ZN(n408) );
  XNOR2_X1 U326 ( .A(n412), .B(n411), .ZN(n289) );
  AND2_X1 U327 ( .A1(G229GAT), .A2(G233GAT), .ZN(n290) );
  XNOR2_X1 U328 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n361) );
  XNOR2_X1 U329 ( .A(n361), .B(G211GAT), .ZN(n404) );
  XNOR2_X1 U330 ( .A(n419), .B(G99GAT), .ZN(n420) );
  XNOR2_X1 U331 ( .A(n403), .B(n290), .ZN(n299) );
  XNOR2_X1 U332 ( .A(n421), .B(n420), .ZN(n426) );
  XOR2_X1 U333 ( .A(G120GAT), .B(G71GAT), .Z(n418) );
  NOR2_X1 U334 ( .A1(n482), .A2(n513), .ZN(n567) );
  NOR2_X1 U335 ( .A1(n520), .A2(n544), .ZN(n525) );
  XNOR2_X1 U336 ( .A(n479), .B(n478), .ZN(n542) );
  XOR2_X1 U337 ( .A(n430), .B(n429), .Z(n527) );
  NOR2_X1 U338 ( .A1(n527), .A2(n485), .ZN(n565) );
  XOR2_X1 U339 ( .A(n304), .B(n303), .Z(n556) );
  XOR2_X1 U340 ( .A(n289), .B(n416), .Z(n516) );
  XNOR2_X1 U341 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n486) );
  XNOR2_X1 U342 ( .A(G50GAT), .B(KEYINPUT108), .ZN(n451) );
  XNOR2_X1 U343 ( .A(n459), .B(G43GAT), .ZN(n460) );
  XNOR2_X1 U344 ( .A(n487), .B(n486), .ZN(G1351GAT) );
  XNOR2_X1 U345 ( .A(n452), .B(n451), .ZN(G1331GAT) );
  XOR2_X1 U346 ( .A(G113GAT), .B(G141GAT), .Z(n292) );
  XNOR2_X1 U347 ( .A(G197GAT), .B(G22GAT), .ZN(n291) );
  XNOR2_X1 U348 ( .A(n292), .B(n291), .ZN(n296) );
  XOR2_X1 U349 ( .A(KEYINPUT30), .B(KEYINPUT67), .Z(n294) );
  XNOR2_X1 U350 ( .A(KEYINPUT29), .B(KEYINPUT66), .ZN(n293) );
  XNOR2_X1 U351 ( .A(n294), .B(n293), .ZN(n295) );
  XNOR2_X1 U352 ( .A(n296), .B(n295), .ZN(n304) );
  XOR2_X1 U353 ( .A(G29GAT), .B(G43GAT), .Z(n298) );
  XNOR2_X1 U354 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n297) );
  XNOR2_X1 U355 ( .A(n298), .B(n297), .ZN(n331) );
  XOR2_X1 U356 ( .A(G169GAT), .B(G8GAT), .Z(n403) );
  XOR2_X1 U357 ( .A(G15GAT), .B(G1GAT), .Z(n353) );
  XOR2_X1 U358 ( .A(n300), .B(n353), .Z(n302) );
  XNOR2_X1 U359 ( .A(G50GAT), .B(G36GAT), .ZN(n301) );
  XNOR2_X1 U360 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U361 ( .A(KEYINPUT70), .B(KEYINPUT68), .Z(n306) );
  XNOR2_X1 U362 ( .A(KEYINPUT33), .B(KEYINPUT69), .ZN(n305) );
  XNOR2_X1 U363 ( .A(n306), .B(n305), .ZN(n320) );
  XOR2_X1 U364 ( .A(KEYINPUT32), .B(KEYINPUT72), .Z(n308) );
  XOR2_X1 U365 ( .A(G176GAT), .B(G64GAT), .Z(n409) );
  XOR2_X1 U366 ( .A(KEYINPUT13), .B(G57GAT), .Z(n340) );
  XNOR2_X1 U367 ( .A(n409), .B(n340), .ZN(n307) );
  XNOR2_X1 U368 ( .A(n308), .B(n307), .ZN(n313) );
  XNOR2_X1 U369 ( .A(G78GAT), .B(G204GAT), .ZN(n309) );
  XNOR2_X1 U370 ( .A(n309), .B(G148GAT), .ZN(n362) );
  XOR2_X1 U371 ( .A(n362), .B(KEYINPUT31), .Z(n311) );
  NAND2_X1 U372 ( .A1(G230GAT), .A2(G233GAT), .ZN(n310) );
  XNOR2_X1 U373 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U374 ( .A(n313), .B(n312), .Z(n318) );
  XOR2_X1 U375 ( .A(G85GAT), .B(KEYINPUT71), .Z(n315) );
  XNOR2_X1 U376 ( .A(G99GAT), .B(G106GAT), .ZN(n314) );
  XNOR2_X1 U377 ( .A(n315), .B(n314), .ZN(n316) );
  XNOR2_X1 U378 ( .A(G92GAT), .B(n316), .ZN(n336) );
  XOR2_X1 U379 ( .A(n418), .B(n336), .Z(n317) );
  XNOR2_X1 U380 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U381 ( .A(n320), .B(n319), .ZN(n575) );
  NAND2_X1 U382 ( .A1(n556), .A2(n575), .ZN(n494) );
  XNOR2_X1 U383 ( .A(KEYINPUT37), .B(KEYINPUT103), .ZN(n447) );
  XOR2_X1 U384 ( .A(KEYINPUT74), .B(KEYINPUT11), .Z(n322) );
  XNOR2_X1 U385 ( .A(KEYINPUT9), .B(KEYINPUT10), .ZN(n321) );
  XNOR2_X1 U386 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U387 ( .A(n323), .B(KEYINPUT75), .Z(n325) );
  XOR2_X1 U388 ( .A(G50GAT), .B(G162GAT), .Z(n370) );
  XNOR2_X1 U389 ( .A(n370), .B(KEYINPUT76), .ZN(n324) );
  XNOR2_X1 U390 ( .A(n325), .B(n324), .ZN(n335) );
  XOR2_X1 U391 ( .A(KEYINPUT65), .B(KEYINPUT73), .Z(n327) );
  NAND2_X1 U392 ( .A1(G232GAT), .A2(G233GAT), .ZN(n326) );
  XNOR2_X1 U393 ( .A(n327), .B(n326), .ZN(n330) );
  XOR2_X1 U394 ( .A(KEYINPUT77), .B(G218GAT), .Z(n329) );
  XNOR2_X1 U395 ( .A(G36GAT), .B(G190GAT), .ZN(n328) );
  XNOR2_X1 U396 ( .A(n329), .B(n328), .ZN(n400) );
  XOR2_X1 U397 ( .A(n330), .B(n400), .Z(n333) );
  XNOR2_X1 U398 ( .A(n331), .B(G134GAT), .ZN(n332) );
  XNOR2_X1 U399 ( .A(n333), .B(n332), .ZN(n334) );
  XNOR2_X1 U400 ( .A(n335), .B(n334), .ZN(n337) );
  XOR2_X1 U401 ( .A(n337), .B(n336), .Z(n553) );
  INV_X1 U402 ( .A(n553), .ZN(n468) );
  XOR2_X1 U403 ( .A(n468), .B(KEYINPUT78), .Z(n537) );
  XNOR2_X1 U404 ( .A(KEYINPUT36), .B(n537), .ZN(n583) );
  XOR2_X1 U405 ( .A(G78GAT), .B(G211GAT), .Z(n339) );
  XNOR2_X1 U406 ( .A(G183GAT), .B(G127GAT), .ZN(n338) );
  XNOR2_X1 U407 ( .A(n339), .B(n338), .ZN(n341) );
  XOR2_X1 U408 ( .A(n341), .B(n340), .Z(n343) );
  XNOR2_X1 U409 ( .A(G8GAT), .B(G71GAT), .ZN(n342) );
  XNOR2_X1 U410 ( .A(n343), .B(n342), .ZN(n357) );
  XOR2_X1 U411 ( .A(G22GAT), .B(G155GAT), .Z(n369) );
  XOR2_X1 U412 ( .A(KEYINPUT14), .B(n369), .Z(n345) );
  NAND2_X1 U413 ( .A1(G231GAT), .A2(G233GAT), .ZN(n344) );
  XNOR2_X1 U414 ( .A(n345), .B(n344), .ZN(n349) );
  XOR2_X1 U415 ( .A(KEYINPUT79), .B(KEYINPUT15), .Z(n347) );
  XNOR2_X1 U416 ( .A(KEYINPUT83), .B(KEYINPUT12), .ZN(n346) );
  XNOR2_X1 U417 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U418 ( .A(n349), .B(n348), .Z(n355) );
  XOR2_X1 U419 ( .A(KEYINPUT80), .B(KEYINPUT81), .Z(n351) );
  XNOR2_X1 U420 ( .A(G64GAT), .B(KEYINPUT82), .ZN(n350) );
  XNOR2_X1 U421 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U422 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U423 ( .A(n355), .B(n354), .ZN(n356) );
  XNOR2_X1 U424 ( .A(n357), .B(n356), .ZN(n580) );
  XOR2_X1 U425 ( .A(KEYINPUT23), .B(KEYINPUT88), .Z(n359) );
  NAND2_X1 U426 ( .A1(G228GAT), .A2(G233GAT), .ZN(n358) );
  XNOR2_X1 U427 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U428 ( .A(n360), .B(KEYINPUT24), .Z(n364) );
  XNOR2_X1 U429 ( .A(n404), .B(n362), .ZN(n363) );
  XNOR2_X1 U430 ( .A(n364), .B(n363), .ZN(n368) );
  XOR2_X1 U431 ( .A(KEYINPUT22), .B(KEYINPUT89), .Z(n366) );
  XNOR2_X1 U432 ( .A(G218GAT), .B(G106GAT), .ZN(n365) );
  XNOR2_X1 U433 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U434 ( .A(n368), .B(n367), .Z(n372) );
  XNOR2_X1 U435 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U436 ( .A(n372), .B(n371), .ZN(n376) );
  XOR2_X1 U437 ( .A(KEYINPUT3), .B(KEYINPUT87), .Z(n374) );
  XNOR2_X1 U438 ( .A(KEYINPUT2), .B(KEYINPUT86), .ZN(n373) );
  XNOR2_X1 U439 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U440 ( .A(G141GAT), .B(n375), .Z(n383) );
  XOR2_X1 U441 ( .A(n376), .B(n383), .Z(n483) );
  XOR2_X1 U442 ( .A(n483), .B(KEYINPUT28), .Z(n520) );
  XOR2_X1 U443 ( .A(KEYINPUT90), .B(KEYINPUT1), .Z(n378) );
  XNOR2_X1 U444 ( .A(KEYINPUT91), .B(KEYINPUT6), .ZN(n377) );
  XNOR2_X1 U445 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X1 U446 ( .A(KEYINPUT4), .B(n379), .Z(n381) );
  NAND2_X1 U447 ( .A1(G225GAT), .A2(G233GAT), .ZN(n380) );
  XNOR2_X1 U448 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U449 ( .A(n382), .B(KEYINPUT5), .Z(n386) );
  INV_X1 U450 ( .A(n383), .ZN(n384) );
  XOR2_X1 U451 ( .A(n384), .B(KEYINPUT92), .Z(n385) );
  XNOR2_X1 U452 ( .A(n386), .B(n385), .ZN(n390) );
  XOR2_X1 U453 ( .A(G85GAT), .B(G155GAT), .Z(n388) );
  XNOR2_X1 U454 ( .A(G29GAT), .B(G162GAT), .ZN(n387) );
  XNOR2_X1 U455 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U456 ( .A(n390), .B(n389), .Z(n399) );
  XOR2_X1 U457 ( .A(KEYINPUT84), .B(G134GAT), .Z(n392) );
  XNOR2_X1 U458 ( .A(KEYINPUT0), .B(G127GAT), .ZN(n391) );
  XNOR2_X1 U459 ( .A(n392), .B(n391), .ZN(n393) );
  XOR2_X1 U460 ( .A(G113GAT), .B(n393), .Z(n429) );
  INV_X1 U461 ( .A(n429), .ZN(n397) );
  XOR2_X1 U462 ( .A(G57GAT), .B(G148GAT), .Z(n395) );
  XNOR2_X1 U463 ( .A(G1GAT), .B(G120GAT), .ZN(n394) );
  XNOR2_X1 U464 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X1 U465 ( .A(n397), .B(n396), .Z(n398) );
  XOR2_X1 U466 ( .A(n399), .B(n398), .Z(n440) );
  INV_X1 U467 ( .A(n440), .ZN(n513) );
  XNOR2_X1 U468 ( .A(n400), .B(KEYINPUT93), .ZN(n402) );
  XNOR2_X1 U469 ( .A(n404), .B(n403), .ZN(n406) );
  AND2_X1 U470 ( .A1(G226GAT), .A2(G233GAT), .ZN(n405) );
  XNOR2_X1 U471 ( .A(n406), .B(n405), .ZN(n407) );
  XOR2_X1 U472 ( .A(n410), .B(n409), .Z(n412) );
  XNOR2_X1 U473 ( .A(G204GAT), .B(G92GAT), .ZN(n411) );
  XOR2_X1 U474 ( .A(KEYINPUT85), .B(KEYINPUT17), .Z(n414) );
  XNOR2_X1 U475 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n413) );
  XNOR2_X1 U476 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U477 ( .A(KEYINPUT19), .B(n415), .ZN(n428) );
  INV_X1 U478 ( .A(n428), .ZN(n416) );
  XNOR2_X1 U479 ( .A(n516), .B(KEYINPUT27), .ZN(n435) );
  NAND2_X1 U480 ( .A1(n513), .A2(n435), .ZN(n544) );
  INV_X1 U481 ( .A(KEYINPUT95), .ZN(n417) );
  XNOR2_X1 U482 ( .A(n525), .B(n417), .ZN(n431) );
  XOR2_X1 U483 ( .A(G176GAT), .B(n418), .Z(n421) );
  NAND2_X1 U484 ( .A1(G227GAT), .A2(G233GAT), .ZN(n419) );
  XOR2_X1 U485 ( .A(KEYINPUT20), .B(G190GAT), .Z(n423) );
  XNOR2_X1 U486 ( .A(G169GAT), .B(G15GAT), .ZN(n422) );
  XNOR2_X1 U487 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U488 ( .A(G43GAT), .B(n424), .Z(n425) );
  XNOR2_X1 U489 ( .A(n426), .B(n425), .ZN(n427) );
  XOR2_X1 U490 ( .A(n428), .B(n427), .Z(n430) );
  NAND2_X1 U491 ( .A1(n431), .A2(n527), .ZN(n443) );
  XNOR2_X1 U492 ( .A(KEYINPUT97), .B(KEYINPUT26), .ZN(n433) );
  INV_X1 U493 ( .A(n527), .ZN(n518) );
  NOR2_X1 U494 ( .A1(n518), .A2(n483), .ZN(n432) );
  XNOR2_X1 U495 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U496 ( .A(KEYINPUT96), .B(n434), .Z(n568) );
  NAND2_X1 U497 ( .A1(n435), .A2(n568), .ZN(n439) );
  NAND2_X1 U498 ( .A1(n518), .A2(n516), .ZN(n436) );
  NAND2_X1 U499 ( .A1(n483), .A2(n436), .ZN(n437) );
  XOR2_X1 U500 ( .A(KEYINPUT25), .B(n437), .Z(n438) );
  NAND2_X1 U501 ( .A1(n439), .A2(n438), .ZN(n441) );
  NAND2_X1 U502 ( .A1(n441), .A2(n440), .ZN(n442) );
  NAND2_X1 U503 ( .A1(n443), .A2(n442), .ZN(n491) );
  NAND2_X1 U504 ( .A1(n580), .A2(n491), .ZN(n444) );
  XOR2_X1 U505 ( .A(KEYINPUT102), .B(n444), .Z(n445) );
  NAND2_X1 U506 ( .A1(n583), .A2(n445), .ZN(n446) );
  XNOR2_X1 U507 ( .A(n447), .B(n446), .ZN(n512) );
  NOR2_X1 U508 ( .A1(n494), .A2(n512), .ZN(n448) );
  XNOR2_X1 U509 ( .A(n448), .B(KEYINPUT38), .ZN(n458) );
  NAND2_X1 U510 ( .A1(n458), .A2(n516), .ZN(n450) );
  XNOR2_X1 U511 ( .A(G36GAT), .B(KEYINPUT106), .ZN(n449) );
  XNOR2_X1 U512 ( .A(n450), .B(n449), .ZN(G1329GAT) );
  NAND2_X1 U513 ( .A1(n458), .A2(n520), .ZN(n452) );
  NAND2_X1 U514 ( .A1(n458), .A2(n513), .ZN(n457) );
  XOR2_X1 U515 ( .A(KEYINPUT104), .B(KEYINPUT105), .Z(n454) );
  XNOR2_X1 U516 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n453) );
  XNOR2_X1 U517 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U518 ( .A(n455), .B(KEYINPUT101), .ZN(n456) );
  XNOR2_X1 U519 ( .A(n457), .B(n456), .ZN(G1328GAT) );
  NAND2_X1 U520 ( .A1(n458), .A2(n518), .ZN(n461) );
  XOR2_X1 U521 ( .A(KEYINPUT40), .B(KEYINPUT107), .Z(n459) );
  XNOR2_X1 U522 ( .A(n461), .B(n460), .ZN(G1330GAT) );
  XOR2_X1 U523 ( .A(KEYINPUT54), .B(KEYINPUT121), .Z(n481) );
  INV_X1 U524 ( .A(n580), .ZN(n564) );
  INV_X1 U525 ( .A(n556), .ZN(n570) );
  INV_X1 U526 ( .A(KEYINPUT41), .ZN(n462) );
  NAND2_X1 U527 ( .A1(n575), .A2(n462), .ZN(n465) );
  INV_X1 U528 ( .A(n575), .ZN(n463) );
  NAND2_X1 U529 ( .A1(n463), .A2(KEYINPUT41), .ZN(n464) );
  NAND2_X1 U530 ( .A1(n465), .A2(n464), .ZN(n548) );
  NOR2_X1 U531 ( .A1(n570), .A2(n548), .ZN(n466) );
  XNOR2_X1 U532 ( .A(n466), .B(KEYINPUT46), .ZN(n467) );
  NOR2_X1 U533 ( .A1(n564), .A2(n467), .ZN(n469) );
  NAND2_X1 U534 ( .A1(n469), .A2(n468), .ZN(n470) );
  XNOR2_X1 U535 ( .A(KEYINPUT47), .B(n470), .ZN(n476) );
  XOR2_X1 U536 ( .A(KEYINPUT45), .B(KEYINPUT113), .Z(n472) );
  NAND2_X1 U537 ( .A1(n564), .A2(n583), .ZN(n471) );
  XNOR2_X1 U538 ( .A(n472), .B(n471), .ZN(n474) );
  NAND2_X1 U539 ( .A1(n570), .A2(n575), .ZN(n473) );
  NOR2_X1 U540 ( .A1(n474), .A2(n473), .ZN(n475) );
  NOR2_X1 U541 ( .A1(n476), .A2(n475), .ZN(n479) );
  XOR2_X1 U542 ( .A(KEYINPUT64), .B(KEYINPUT114), .Z(n477) );
  NAND2_X1 U543 ( .A1(n542), .A2(n516), .ZN(n480) );
  XNOR2_X1 U544 ( .A(n481), .B(n480), .ZN(n482) );
  NAND2_X1 U545 ( .A1(n483), .A2(n567), .ZN(n484) );
  XOR2_X1 U546 ( .A(KEYINPUT55), .B(n484), .Z(n485) );
  NAND2_X1 U547 ( .A1(n537), .A2(n565), .ZN(n487) );
  XNOR2_X1 U548 ( .A(G1GAT), .B(KEYINPUT99), .ZN(n488) );
  XNOR2_X1 U549 ( .A(n488), .B(KEYINPUT100), .ZN(n489) );
  XOR2_X1 U550 ( .A(KEYINPUT34), .B(n489), .Z(n496) );
  NOR2_X1 U551 ( .A1(n537), .A2(n580), .ZN(n490) );
  XNOR2_X1 U552 ( .A(KEYINPUT16), .B(n490), .ZN(n492) );
  NAND2_X1 U553 ( .A1(n492), .A2(n491), .ZN(n493) );
  XNOR2_X1 U554 ( .A(n493), .B(KEYINPUT98), .ZN(n502) );
  NOR2_X1 U555 ( .A1(n502), .A2(n494), .ZN(n500) );
  NAND2_X1 U556 ( .A1(n500), .A2(n513), .ZN(n495) );
  XNOR2_X1 U557 ( .A(n496), .B(n495), .ZN(G1324GAT) );
  NAND2_X1 U558 ( .A1(n500), .A2(n516), .ZN(n497) );
  XNOR2_X1 U559 ( .A(n497), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U560 ( .A(G15GAT), .B(KEYINPUT35), .Z(n499) );
  NAND2_X1 U561 ( .A1(n500), .A2(n518), .ZN(n498) );
  XNOR2_X1 U562 ( .A(n499), .B(n498), .ZN(G1326GAT) );
  NAND2_X1 U563 ( .A1(n500), .A2(n520), .ZN(n501) );
  XNOR2_X1 U564 ( .A(n501), .B(G22GAT), .ZN(G1327GAT) );
  XNOR2_X1 U565 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n504) );
  XNOR2_X1 U566 ( .A(KEYINPUT109), .B(n548), .ZN(n561) );
  NAND2_X1 U567 ( .A1(n570), .A2(n561), .ZN(n511) );
  NOR2_X1 U568 ( .A1(n502), .A2(n511), .ZN(n508) );
  NAND2_X1 U569 ( .A1(n513), .A2(n508), .ZN(n503) );
  XNOR2_X1 U570 ( .A(n504), .B(n503), .ZN(G1332GAT) );
  NAND2_X1 U571 ( .A1(n508), .A2(n516), .ZN(n505) );
  XNOR2_X1 U572 ( .A(n505), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U573 ( .A1(n508), .A2(n518), .ZN(n506) );
  XNOR2_X1 U574 ( .A(n506), .B(KEYINPUT110), .ZN(n507) );
  XNOR2_X1 U575 ( .A(G71GAT), .B(n507), .ZN(G1334GAT) );
  XOR2_X1 U576 ( .A(G78GAT), .B(KEYINPUT43), .Z(n510) );
  NAND2_X1 U577 ( .A1(n508), .A2(n520), .ZN(n509) );
  XNOR2_X1 U578 ( .A(n510), .B(n509), .ZN(G1335GAT) );
  XOR2_X1 U579 ( .A(G85GAT), .B(KEYINPUT111), .Z(n515) );
  NOR2_X1 U580 ( .A1(n512), .A2(n511), .ZN(n521) );
  NAND2_X1 U581 ( .A1(n521), .A2(n513), .ZN(n514) );
  XNOR2_X1 U582 ( .A(n515), .B(n514), .ZN(G1336GAT) );
  NAND2_X1 U583 ( .A1(n521), .A2(n516), .ZN(n517) );
  XNOR2_X1 U584 ( .A(n517), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U585 ( .A1(n521), .A2(n518), .ZN(n519) );
  XNOR2_X1 U586 ( .A(n519), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U587 ( .A(KEYINPUT112), .B(KEYINPUT44), .Z(n523) );
  NAND2_X1 U588 ( .A1(n521), .A2(n520), .ZN(n522) );
  XNOR2_X1 U589 ( .A(n523), .B(n522), .ZN(n524) );
  XOR2_X1 U590 ( .A(G106GAT), .B(n524), .Z(G1339GAT) );
  NAND2_X1 U591 ( .A1(n542), .A2(n525), .ZN(n526) );
  NOR2_X1 U592 ( .A1(n527), .A2(n526), .ZN(n528) );
  XOR2_X1 U593 ( .A(KEYINPUT115), .B(n528), .Z(n538) );
  NAND2_X1 U594 ( .A1(n556), .A2(n538), .ZN(n529) );
  XNOR2_X1 U595 ( .A(n529), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U596 ( .A(KEYINPUT116), .B(KEYINPUT49), .Z(n531) );
  NAND2_X1 U597 ( .A1(n538), .A2(n561), .ZN(n530) );
  XNOR2_X1 U598 ( .A(n531), .B(n530), .ZN(n532) );
  XNOR2_X1 U599 ( .A(G120GAT), .B(n532), .ZN(G1341GAT) );
  XNOR2_X1 U600 ( .A(G127GAT), .B(KEYINPUT118), .ZN(n536) );
  XOR2_X1 U601 ( .A(KEYINPUT117), .B(KEYINPUT50), .Z(n534) );
  NAND2_X1 U602 ( .A1(n538), .A2(n564), .ZN(n533) );
  XNOR2_X1 U603 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U604 ( .A(n536), .B(n535), .ZN(G1342GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT51), .B(KEYINPUT119), .Z(n540) );
  NAND2_X1 U606 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U607 ( .A(n540), .B(n539), .ZN(n541) );
  XOR2_X1 U608 ( .A(G134GAT), .B(n541), .Z(G1343GAT) );
  NAND2_X1 U609 ( .A1(n542), .A2(n568), .ZN(n543) );
  NOR2_X1 U610 ( .A1(n544), .A2(n543), .ZN(n554) );
  NAND2_X1 U611 ( .A1(n556), .A2(n554), .ZN(n545) );
  XNOR2_X1 U612 ( .A(n545), .B(KEYINPUT120), .ZN(n546) );
  XNOR2_X1 U613 ( .A(G141GAT), .B(n546), .ZN(G1344GAT) );
  INV_X1 U614 ( .A(n554), .ZN(n547) );
  NOR2_X1 U615 ( .A1(n548), .A2(n547), .ZN(n550) );
  XNOR2_X1 U616 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n549) );
  XNOR2_X1 U617 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U618 ( .A(G148GAT), .B(n551), .ZN(G1345GAT) );
  NAND2_X1 U619 ( .A1(n554), .A2(n564), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n552), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U621 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n555), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U623 ( .A1(n556), .A2(n565), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n557), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U625 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n559) );
  XNOR2_X1 U626 ( .A(G176GAT), .B(KEYINPUT122), .ZN(n558) );
  XNOR2_X1 U627 ( .A(n559), .B(n558), .ZN(n560) );
  XOR2_X1 U628 ( .A(KEYINPUT56), .B(n560), .Z(n563) );
  NAND2_X1 U629 ( .A1(n561), .A2(n565), .ZN(n562) );
  XNOR2_X1 U630 ( .A(n563), .B(n562), .ZN(G1349GAT) );
  NAND2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n566), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U633 ( .A1(n567), .A2(n568), .ZN(n569) );
  XOR2_X1 U634 ( .A(KEYINPUT124), .B(n569), .Z(n584) );
  INV_X1 U635 ( .A(n584), .ZN(n581) );
  NOR2_X1 U636 ( .A1(n581), .A2(n570), .ZN(n574) );
  XOR2_X1 U637 ( .A(KEYINPUT60), .B(KEYINPUT125), .Z(n572) );
  XNOR2_X1 U638 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n571) );
  XNOR2_X1 U639 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(G1352GAT) );
  NOR2_X1 U641 ( .A1(n575), .A2(n581), .ZN(n579) );
  XOR2_X1 U642 ( .A(KEYINPUT126), .B(KEYINPUT127), .Z(n577) );
  XNOR2_X1 U643 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n576) );
  XNOR2_X1 U644 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U645 ( .A(n579), .B(n578), .ZN(G1353GAT) );
  NOR2_X1 U646 ( .A1(n581), .A2(n580), .ZN(n582) );
  XOR2_X1 U647 ( .A(G211GAT), .B(n582), .Z(G1354GAT) );
  NAND2_X1 U648 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U649 ( .A(n585), .B(KEYINPUT62), .ZN(n586) );
  XNOR2_X1 U650 ( .A(G218GAT), .B(n586), .ZN(G1355GAT) );
endmodule

