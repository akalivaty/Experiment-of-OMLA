//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 1 1 0 0 1 1 0 0 0 1 0 1 1 1 0 0 0 1 1 1 0 0 1 0 1 1 0 0 0 0 1 0 1 1 1 1 0 1 1 0 1 1 1 1 0 0 1 1 0 0 0 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:02 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n697, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n765, new_n766, new_n767, new_n768, new_n769, new_n771,
    new_n772, new_n773, new_n775, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n806, new_n807, new_n808, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n865, new_n866, new_n867, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n927, new_n928, new_n930, new_n931,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n946, new_n947, new_n948,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n967, new_n968, new_n969, new_n970, new_n971, new_n973,
    new_n974, new_n975, new_n976, new_n978, new_n979;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(G1gat), .ZN(new_n203));
  NAND3_X1  g002(.A1(new_n202), .A2(KEYINPUT16), .A3(new_n203), .ZN(new_n204));
  OR2_X1    g003(.A1(KEYINPUT94), .A2(G8gat), .ZN(new_n205));
  OAI211_X1 g004(.A(new_n204), .B(new_n205), .C1(new_n203), .C2(new_n202), .ZN(new_n206));
  NAND2_X1  g005(.A1(KEYINPUT94), .A2(G8gat), .ZN(new_n207));
  XOR2_X1   g006(.A(new_n206), .B(new_n207), .Z(new_n208));
  INV_X1    g007(.A(KEYINPUT15), .ZN(new_n209));
  OR2_X1    g008(.A1(G43gat), .A2(G50gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(G43gat), .A2(G50gat), .ZN(new_n211));
  AOI21_X1  g010(.A(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(KEYINPUT90), .B(G36gat), .ZN(new_n213));
  INV_X1    g012(.A(G29gat), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(G36gat), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n214), .A2(new_n216), .A3(KEYINPUT14), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT14), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n218), .B1(G29gat), .B2(G36gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n212), .B1(new_n215), .B2(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(KEYINPUT91), .B(G50gat), .ZN(new_n222));
  INV_X1    g021(.A(G43gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  AOI21_X1  g023(.A(KEYINPUT15), .B1(G43gat), .B2(G50gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  XOR2_X1   g025(.A(KEYINPUT90), .B(G36gat), .Z(new_n227));
  INV_X1    g026(.A(KEYINPUT93), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n227), .A2(new_n228), .A3(G29gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n220), .A2(KEYINPUT92), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT92), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n217), .A2(new_n219), .A3(new_n231), .ZN(new_n232));
  NAND4_X1  g031(.A1(new_n226), .A2(new_n229), .A3(new_n230), .A4(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(new_n212), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n234), .B1(new_n215), .B2(new_n228), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n221), .B1(new_n233), .B2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n208), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT17), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n236), .A2(new_n239), .ZN(new_n240));
  AND2_X1   g039(.A1(new_n208), .A2(new_n240), .ZN(new_n241));
  OAI211_X1 g040(.A(KEYINPUT17), .B(new_n221), .C1(new_n233), .C2(new_n235), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n238), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(G229gat), .A2(G233gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT18), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n208), .B(new_n237), .ZN(new_n247));
  XOR2_X1   g046(.A(new_n244), .B(KEYINPUT13), .Z(new_n248));
  AOI22_X1  g047(.A1(new_n245), .A2(new_n246), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT95), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n250), .B1(new_n245), .B2(new_n246), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n243), .A2(KEYINPUT95), .A3(KEYINPUT18), .A4(new_n244), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n249), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(KEYINPUT89), .ZN(new_n254));
  XNOR2_X1  g053(.A(G113gat), .B(G141gat), .ZN(new_n255));
  XNOR2_X1  g054(.A(G169gat), .B(G197gat), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n255), .B(new_n256), .ZN(new_n257));
  XOR2_X1   g056(.A(KEYINPUT88), .B(KEYINPUT11), .Z(new_n258));
  XNOR2_X1  g057(.A(new_n257), .B(new_n258), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n259), .B(KEYINPUT12), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n254), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n253), .A2(KEYINPUT89), .A3(new_n260), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(G197gat), .B(G204gat), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT22), .ZN(new_n266));
  INV_X1    g065(.A(G211gat), .ZN(new_n267));
  INV_X1    g066(.A(G218gat), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n266), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n265), .A2(new_n269), .ZN(new_n270));
  XOR2_X1   g069(.A(G211gat), .B(G218gat), .Z(new_n271));
  OR2_X1    g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n270), .A2(new_n271), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT29), .ZN(new_n275));
  AOI21_X1  g074(.A(KEYINPUT3), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT82), .ZN(new_n277));
  AND2_X1   g076(.A1(G155gat), .A2(G162gat), .ZN(new_n278));
  NOR2_X1   g077(.A1(G155gat), .A2(G162gat), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  XNOR2_X1  g079(.A(G141gat), .B(G148gat), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT2), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n282), .B1(G155gat), .B2(G162gat), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n280), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(G141gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(G148gat), .ZN(new_n286));
  INV_X1    g085(.A(G148gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(G141gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  XNOR2_X1  g088(.A(G155gat), .B(G162gat), .ZN(new_n290));
  INV_X1    g089(.A(G155gat), .ZN(new_n291));
  INV_X1    g090(.A(G162gat), .ZN(new_n292));
  OAI21_X1  g091(.A(KEYINPUT2), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n289), .A2(new_n290), .A3(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n284), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  OR3_X1    g095(.A1(new_n276), .A2(new_n277), .A3(new_n296), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n277), .B1(new_n276), .B2(new_n296), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT76), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n272), .A2(new_n299), .A3(new_n273), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n270), .A2(KEYINPUT76), .A3(new_n271), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT3), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n284), .A2(new_n294), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(new_n275), .ZN(new_n305));
  AOI22_X1  g104(.A1(new_n302), .A2(new_n305), .B1(G228gat), .B2(G233gat), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n297), .A2(new_n298), .A3(new_n306), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n300), .A2(new_n275), .A3(new_n301), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n296), .B1(new_n308), .B2(new_n303), .ZN(new_n309));
  AND2_X1   g108(.A1(new_n302), .A2(new_n305), .ZN(new_n310));
  OAI211_X1 g109(.A(G228gat), .B(G233gat), .C1(new_n309), .C2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n307), .A2(new_n311), .ZN(new_n312));
  XNOR2_X1  g111(.A(KEYINPUT31), .B(G50gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n313), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n307), .A2(new_n311), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(G78gat), .B(G106gat), .ZN(new_n318));
  XNOR2_X1  g117(.A(new_n318), .B(G22gat), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n317), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n314), .A2(new_n319), .A3(new_n316), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(G225gat), .A2(G233gat), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  XNOR2_X1  g124(.A(G113gat), .B(G120gat), .ZN(new_n326));
  INV_X1    g125(.A(G127gat), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n327), .A2(G134gat), .ZN(new_n328));
  INV_X1    g127(.A(G134gat), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n329), .A2(G127gat), .ZN(new_n330));
  OAI22_X1  g129(.A1(new_n326), .A2(KEYINPUT1), .B1(new_n328), .B2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(G120gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(G113gat), .ZN(new_n333));
  INV_X1    g132(.A(G113gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(G120gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  XNOR2_X1  g135(.A(G127gat), .B(G134gat), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT1), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n336), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  NAND4_X1  g138(.A1(new_n331), .A2(new_n284), .A3(new_n294), .A4(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(KEYINPUT4), .ZN(new_n342));
  AND3_X1   g141(.A1(new_n331), .A2(new_n339), .A3(KEYINPUT72), .ZN(new_n343));
  AOI21_X1  g142(.A(KEYINPUT72), .B1(new_n331), .B2(new_n339), .ZN(new_n344));
  NOR3_X1   g143(.A1(new_n343), .A2(new_n344), .A3(new_n295), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n342), .B1(new_n345), .B2(KEYINPUT4), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT78), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n295), .A2(new_n347), .A3(KEYINPUT3), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n331), .A2(new_n339), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n348), .A2(new_n349), .A3(new_n304), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n347), .B1(new_n295), .B2(KEYINPUT3), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n325), .B1(new_n346), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n349), .A2(new_n295), .ZN(new_n354));
  AND2_X1   g153(.A1(new_n354), .A2(new_n340), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(new_n324), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n353), .A2(KEYINPUT39), .A3(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT40), .ZN(new_n359));
  XOR2_X1   g158(.A(G1gat), .B(G29gat), .Z(new_n360));
  XNOR2_X1  g159(.A(G57gat), .B(G85gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n360), .B(new_n361), .ZN(new_n362));
  XNOR2_X1  g161(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n363));
  XNOR2_X1  g162(.A(new_n362), .B(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n365), .B1(new_n353), .B2(KEYINPUT39), .ZN(new_n366));
  OR3_X1    g165(.A1(new_n358), .A2(new_n359), .A3(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT5), .ZN(new_n368));
  OAI211_X1 g167(.A(new_n368), .B(new_n324), .C1(new_n350), .C2(new_n351), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n369), .A2(new_n346), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT4), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n341), .A2(KEYINPUT79), .A3(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT79), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n374), .B1(new_n340), .B2(KEYINPUT4), .ZN(new_n375));
  OAI211_X1 g174(.A(new_n373), .B(new_n375), .C1(new_n345), .C2(new_n372), .ZN(new_n376));
  AOI211_X1 g175(.A(KEYINPUT78), .B(new_n303), .C1(new_n284), .C2(new_n294), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n304), .A2(new_n349), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n351), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n325), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  AND2_X1   g180(.A1(new_n376), .A2(new_n381), .ZN(new_n382));
  OAI21_X1  g181(.A(KEYINPUT5), .B1(new_n355), .B2(new_n324), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n371), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(new_n364), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n359), .B1(new_n358), .B2(new_n366), .ZN(new_n386));
  AND3_X1   g185(.A1(new_n367), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT77), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT30), .ZN(new_n389));
  NAND2_X1  g188(.A1(G226gat), .A2(G233gat), .ZN(new_n390));
  INV_X1    g189(.A(G169gat), .ZN(new_n391));
  INV_X1    g190(.A(G176gat), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n391), .A2(new_n392), .A3(KEYINPUT71), .ZN(new_n393));
  AOI22_X1  g192(.A1(new_n393), .A2(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n394), .B1(KEYINPUT26), .B2(new_n393), .ZN(new_n395));
  NAND2_X1  g194(.A1(G183gat), .A2(G190gat), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT28), .ZN(new_n398));
  XNOR2_X1  g197(.A(KEYINPUT66), .B(G190gat), .ZN(new_n399));
  INV_X1    g198(.A(G183gat), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(KEYINPUT27), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT68), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n400), .A2(KEYINPUT68), .A3(KEYINPUT27), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n399), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  OR2_X1    g204(.A1(KEYINPUT69), .A2(KEYINPUT27), .ZN(new_n406));
  NAND2_X1  g205(.A1(KEYINPUT69), .A2(KEYINPUT27), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n400), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n398), .B1(new_n405), .B2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT70), .ZN(new_n410));
  INV_X1    g209(.A(G190gat), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(KEYINPUT66), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT66), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(G190gat), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n412), .A2(new_n414), .A3(KEYINPUT28), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT27), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(G183gat), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n417), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n410), .B1(new_n415), .B2(new_n418), .ZN(new_n419));
  XNOR2_X1  g218(.A(KEYINPUT27), .B(G183gat), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n399), .A2(new_n420), .A3(KEYINPUT70), .A4(KEYINPUT28), .ZN(new_n421));
  AND2_X1   g220(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n397), .B1(new_n409), .B2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT25), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT24), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n396), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n400), .A2(new_n411), .ZN(new_n428));
  AND3_X1   g227(.A1(new_n426), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n391), .A2(new_n392), .A3(KEYINPUT23), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT23), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n431), .B1(G169gat), .B2(G176gat), .ZN(new_n432));
  NAND2_X1  g231(.A1(G169gat), .A2(G176gat), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n430), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n424), .B1(new_n429), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(KEYINPUT64), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT64), .ZN(new_n437));
  OAI211_X1 g236(.A(new_n437), .B(new_n424), .C1(new_n429), .C2(new_n434), .ZN(new_n438));
  AND2_X1   g237(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n412), .A2(new_n414), .A3(new_n400), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT65), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n426), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n396), .A2(KEYINPUT65), .A3(new_n425), .ZN(new_n443));
  NAND4_X1  g242(.A1(new_n440), .A2(new_n442), .A3(new_n427), .A4(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT67), .ZN(new_n445));
  AND4_X1   g244(.A1(KEYINPUT25), .A2(new_n430), .A3(new_n432), .A4(new_n433), .ZN(new_n446));
  AND3_X1   g245(.A1(new_n444), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n445), .B1(new_n444), .B2(new_n446), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n423), .B1(new_n439), .B2(new_n449), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n390), .B1(new_n450), .B2(KEYINPUT29), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n444), .A2(new_n446), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(KEYINPUT67), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n444), .A2(new_n445), .A3(new_n446), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n453), .A2(new_n436), .A3(new_n438), .A4(new_n454), .ZN(new_n455));
  AND3_X1   g254(.A1(new_n399), .A2(new_n403), .A3(new_n404), .ZN(new_n456));
  INV_X1    g255(.A(new_n408), .ZN(new_n457));
  AOI21_X1  g256(.A(KEYINPUT28), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n419), .A2(new_n421), .ZN(new_n459));
  OAI211_X1 g258(.A(new_n395), .B(new_n396), .C1(new_n458), .C2(new_n459), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n390), .B1(new_n455), .B2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(new_n461), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n302), .B1(new_n451), .B2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n390), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n455), .A2(new_n460), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n464), .B1(new_n465), .B2(new_n275), .ZN(new_n466));
  INV_X1    g265(.A(new_n302), .ZN(new_n467));
  NOR3_X1   g266(.A1(new_n466), .A2(new_n467), .A3(new_n461), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n463), .A2(new_n468), .ZN(new_n469));
  XNOR2_X1  g268(.A(G8gat), .B(G36gat), .ZN(new_n470));
  XNOR2_X1  g269(.A(G64gat), .B(G92gat), .ZN(new_n471));
  XOR2_X1   g270(.A(new_n470), .B(new_n471), .Z(new_n472));
  INV_X1    g271(.A(new_n472), .ZN(new_n473));
  OAI211_X1 g272(.A(new_n388), .B(new_n389), .C1(new_n469), .C2(new_n473), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n467), .B1(new_n466), .B2(new_n461), .ZN(new_n475));
  AOI21_X1  g274(.A(KEYINPUT29), .B1(new_n455), .B2(new_n460), .ZN(new_n476));
  OAI211_X1 g275(.A(new_n462), .B(new_n302), .C1(new_n464), .C2(new_n476), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n473), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  OAI21_X1  g277(.A(KEYINPUT30), .B1(new_n478), .B2(KEYINPUT77), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n469), .A2(new_n473), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n474), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n323), .B1(new_n387), .B2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT87), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n383), .B1(new_n376), .B2(new_n381), .ZN(new_n484));
  OAI211_X1 g283(.A(KEYINPUT6), .B(new_n364), .C1(new_n484), .C2(new_n370), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT81), .ZN(new_n486));
  AND2_X1   g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n485), .A2(new_n486), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n483), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND4_X1  g288(.A1(new_n384), .A2(KEYINPUT81), .A3(KEYINPUT6), .A4(new_n364), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n485), .A2(new_n486), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n490), .A2(KEYINPUT87), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  XNOR2_X1  g292(.A(KEYINPUT85), .B(KEYINPUT37), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n494), .B1(new_n463), .B2(new_n468), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n475), .A2(new_n477), .A3(KEYINPUT37), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n495), .A2(new_n473), .A3(new_n496), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n478), .B1(new_n497), .B2(KEYINPUT38), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT6), .ZN(new_n499));
  OAI211_X1 g298(.A(new_n371), .B(new_n365), .C1(new_n382), .C2(new_n383), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n385), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n493), .A2(new_n498), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n496), .A2(KEYINPUT84), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT84), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n475), .A2(new_n477), .A3(new_n504), .A4(KEYINPUT37), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT38), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n495), .A2(new_n507), .A3(new_n473), .ZN(new_n508));
  OAI21_X1  g307(.A(KEYINPUT86), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(new_n494), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n510), .B1(new_n475), .B2(new_n477), .ZN(new_n511));
  NOR3_X1   g310(.A1(new_n511), .A2(KEYINPUT38), .A3(new_n472), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT86), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n512), .A2(new_n513), .A3(new_n503), .A4(new_n505), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n509), .A2(new_n514), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n482), .B1(new_n502), .B2(new_n515), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n343), .A2(new_n344), .ZN(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  AND3_X1   g317(.A1(new_n455), .A2(new_n518), .A3(new_n460), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n518), .B1(new_n455), .B2(new_n460), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(G227gat), .ZN(new_n522));
  INV_X1    g321(.A(G233gat), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  AOI21_X1  g323(.A(KEYINPUT73), .B1(new_n521), .B2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT73), .ZN(new_n526));
  INV_X1    g325(.A(new_n524), .ZN(new_n527));
  NOR4_X1   g326(.A1(new_n519), .A2(new_n520), .A3(new_n526), .A4(new_n527), .ZN(new_n528));
  OAI21_X1  g327(.A(KEYINPUT32), .B1(new_n525), .B2(new_n528), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n527), .B1(new_n519), .B2(new_n520), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n530), .A2(KEYINPUT34), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT34), .ZN(new_n532));
  OAI211_X1 g331(.A(new_n532), .B(new_n527), .C1(new_n519), .C2(new_n520), .ZN(new_n533));
  AND2_X1   g332(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n529), .A2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT32), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n521), .A2(KEYINPUT73), .A3(new_n524), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n465), .A2(new_n517), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n455), .A2(new_n518), .A3(new_n460), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n538), .A2(new_n524), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(new_n526), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n536), .B1(new_n537), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n531), .A2(new_n533), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  XOR2_X1   g343(.A(G15gat), .B(G43gat), .Z(new_n545));
  XNOR2_X1  g344(.A(new_n545), .B(KEYINPUT74), .ZN(new_n546));
  XNOR2_X1  g345(.A(G71gat), .B(G99gat), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n546), .B(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n537), .A2(new_n541), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT33), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n549), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  AND3_X1   g351(.A1(new_n535), .A2(new_n544), .A3(new_n552), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n552), .B1(new_n535), .B2(new_n544), .ZN(new_n554));
  OAI21_X1  g353(.A(KEYINPUT75), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n552), .A2(KEYINPUT36), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT36), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n555), .A2(new_n559), .ZN(new_n560));
  AND3_X1   g359(.A1(new_n321), .A2(new_n322), .A3(KEYINPUT83), .ZN(new_n561));
  AOI21_X1  g360(.A(KEYINPUT83), .B1(new_n321), .B2(new_n322), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n501), .A2(new_n490), .A3(new_n491), .ZN(new_n564));
  NAND4_X1  g363(.A1(new_n564), .A2(new_n474), .A3(new_n480), .A4(new_n479), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  OAI211_X1 g365(.A(KEYINPUT75), .B(new_n558), .C1(new_n553), .C2(new_n554), .ZN(new_n567));
  NAND4_X1  g366(.A1(new_n516), .A2(new_n560), .A3(new_n566), .A4(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n535), .A2(new_n544), .ZN(new_n569));
  AOI21_X1  g368(.A(KEYINPUT33), .B1(new_n537), .B2(new_n541), .ZN(new_n570));
  OR2_X1    g369(.A1(new_n570), .A2(new_n549), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n323), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n535), .A2(new_n544), .A3(new_n552), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  OAI21_X1  g374(.A(KEYINPUT35), .B1(new_n575), .B2(new_n565), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n553), .A2(new_n554), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n493), .A2(new_n501), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n481), .A2(KEYINPUT35), .ZN(new_n579));
  NAND4_X1  g378(.A1(new_n577), .A2(new_n578), .A3(new_n579), .A4(new_n573), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n576), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n264), .B1(new_n568), .B2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT96), .ZN(new_n583));
  XOR2_X1   g382(.A(G57gat), .B(G64gat), .Z(new_n584));
  NAND2_X1  g383(.A1(G71gat), .A2(G78gat), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT9), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n584), .B1(KEYINPUT97), .B2(new_n587), .ZN(new_n588));
  AND2_X1   g387(.A1(new_n587), .A2(KEYINPUT97), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n583), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(G71gat), .B(G78gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n590), .B(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(G99gat), .A2(G106gat), .ZN(new_n593));
  INV_X1    g392(.A(G85gat), .ZN(new_n594));
  INV_X1    g393(.A(G92gat), .ZN(new_n595));
  AOI22_X1  g394(.A1(KEYINPUT8), .A2(new_n593), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT7), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n597), .B1(new_n594), .B2(new_n595), .ZN(new_n598));
  NAND3_X1  g397(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n596), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(G99gat), .B(G106gat), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  NAND4_X1  g402(.A1(new_n596), .A2(new_n601), .A3(new_n598), .A4(new_n599), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n603), .A2(KEYINPUT100), .A3(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT100), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n600), .A2(new_n606), .A3(new_n602), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n592), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT102), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT10), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n592), .A2(KEYINPUT102), .A3(new_n609), .ZN(new_n614));
  XOR2_X1   g413(.A(new_n590), .B(new_n591), .Z(new_n615));
  AND2_X1   g414(.A1(new_n603), .A2(new_n604), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND4_X1  g416(.A1(new_n612), .A2(new_n613), .A3(new_n614), .A4(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n615), .A2(KEYINPUT10), .A3(new_n608), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(G230gat), .A2(G233gat), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n612), .A2(new_n614), .A3(new_n617), .ZN(new_n623));
  INV_X1    g422(.A(new_n621), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  XOR2_X1   g424(.A(G120gat), .B(G148gat), .Z(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(KEYINPUT103), .ZN(new_n627));
  XNOR2_X1  g426(.A(G176gat), .B(G204gat), .ZN(new_n628));
  XOR2_X1   g427(.A(new_n627), .B(new_n628), .Z(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  AND3_X1   g429(.A1(new_n622), .A2(new_n625), .A3(new_n630), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n630), .B1(new_n622), .B2(new_n625), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT21), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n592), .A2(new_n634), .ZN(new_n635));
  XOR2_X1   g434(.A(G127gat), .B(G155gat), .Z(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n208), .B1(new_n592), .B2(new_n634), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n637), .B(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(G231gat), .A2(G233gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(KEYINPUT98), .ZN(new_n641));
  XOR2_X1   g440(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n642));
  XNOR2_X1  g441(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(G183gat), .B(G211gat), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n639), .B(new_n645), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n608), .B1(new_n236), .B2(new_n239), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n647), .A2(new_n242), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT101), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n647), .A2(KEYINPUT101), .A3(new_n242), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  AND2_X1   g451(.A1(G232gat), .A2(G233gat), .ZN(new_n653));
  AOI22_X1  g452(.A1(new_n236), .A2(new_n608), .B1(KEYINPUT41), .B2(new_n653), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n411), .B1(new_n652), .B2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n654), .ZN(new_n656));
  AOI211_X1 g455(.A(G190gat), .B(new_n656), .C1(new_n650), .C2(new_n651), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n268), .B1(new_n655), .B2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT99), .ZN(new_n659));
  INV_X1    g458(.A(new_n651), .ZN(new_n660));
  AOI21_X1  g459(.A(KEYINPUT101), .B1(new_n647), .B2(new_n242), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n654), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n662), .A2(G190gat), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n652), .A2(new_n411), .A3(new_n654), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n663), .A2(new_n664), .A3(G218gat), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n658), .A2(new_n659), .A3(new_n665), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n653), .A2(KEYINPUT41), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  XOR2_X1   g467(.A(G134gat), .B(G162gat), .Z(new_n669));
  INV_X1    g468(.A(new_n667), .ZN(new_n670));
  NAND4_X1  g469(.A1(new_n658), .A2(new_n659), .A3(new_n665), .A4(new_n670), .ZN(new_n671));
  AND3_X1   g470(.A1(new_n668), .A2(new_n669), .A3(new_n671), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n669), .B1(new_n668), .B2(new_n671), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND4_X1  g473(.A1(new_n582), .A2(new_n633), .A3(new_n646), .A4(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT104), .ZN(new_n676));
  AND2_X1   g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n675), .A2(new_n676), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n679), .A2(new_n564), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n680), .B(new_n203), .ZN(G1324gat));
  INV_X1    g480(.A(new_n481), .ZN(new_n682));
  OAI21_X1  g481(.A(G8gat), .B1(new_n679), .B2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT42), .ZN(new_n684));
  XOR2_X1   g483(.A(KEYINPUT16), .B(G8gat), .Z(new_n685));
  OAI211_X1 g484(.A(new_n481), .B(new_n685), .C1(new_n677), .C2(new_n678), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT105), .ZN(new_n687));
  AND3_X1   g486(.A1(new_n686), .A2(new_n687), .A3(new_n684), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n687), .B1(new_n686), .B2(new_n684), .ZN(new_n689));
  OAI221_X1 g488(.A(new_n683), .B1(new_n684), .B2(new_n686), .C1(new_n688), .C2(new_n689), .ZN(G1325gat));
  NAND2_X1  g489(.A1(new_n560), .A2(new_n567), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(G15gat), .B1(new_n679), .B2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n577), .ZN(new_n694));
  OR2_X1    g493(.A1(new_n694), .A2(G15gat), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n693), .B1(new_n679), .B2(new_n695), .ZN(G1326gat));
  INV_X1    g495(.A(new_n563), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n679), .A2(new_n697), .ZN(new_n698));
  XOR2_X1   g497(.A(KEYINPUT43), .B(G22gat), .Z(new_n699));
  XNOR2_X1  g498(.A(new_n698), .B(new_n699), .ZN(G1327gat));
  NAND2_X1  g499(.A1(new_n622), .A2(new_n625), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(new_n629), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n622), .A2(new_n625), .A3(new_n630), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NOR3_X1   g503(.A1(new_n674), .A2(new_n704), .A3(new_n646), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n582), .A2(new_n705), .ZN(new_n706));
  NOR3_X1   g505(.A1(new_n706), .A2(G29gat), .A3(new_n564), .ZN(new_n707));
  XNOR2_X1  g506(.A(KEYINPUT106), .B(KEYINPUT45), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n707), .B(new_n708), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n704), .B(KEYINPUT107), .ZN(new_n710));
  NOR3_X1   g509(.A1(new_n710), .A2(new_n264), .A3(new_n646), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT44), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n568), .A2(new_n581), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n668), .A2(new_n671), .ZN(new_n714));
  INV_X1    g513(.A(new_n669), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n668), .A2(new_n669), .A3(new_n671), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n712), .B1(new_n713), .B2(new_n718), .ZN(new_n719));
  XOR2_X1   g518(.A(KEYINPUT108), .B(KEYINPUT44), .Z(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  AOI211_X1 g520(.A(new_n674), .B(new_n721), .C1(new_n568), .C2(new_n581), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n711), .B1(new_n719), .B2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT109), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(new_n564), .ZN(new_n726));
  OAI211_X1 g525(.A(KEYINPUT109), .B(new_n711), .C1(new_n719), .C2(new_n722), .ZN(new_n727));
  AND3_X1   g526(.A1(new_n725), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n709), .B1(new_n728), .B2(new_n214), .ZN(G1328gat));
  INV_X1    g528(.A(new_n706), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT46), .ZN(new_n731));
  OR2_X1    g530(.A1(new_n731), .A2(KEYINPUT110), .ZN(new_n732));
  NAND4_X1  g531(.A1(new_n730), .A2(new_n481), .A3(new_n213), .A4(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n731), .A2(KEYINPUT110), .ZN(new_n734));
  XOR2_X1   g533(.A(new_n733), .B(new_n734), .Z(new_n735));
  AND3_X1   g534(.A1(new_n725), .A2(new_n481), .A3(new_n727), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n735), .B1(new_n213), .B2(new_n736), .ZN(G1329gat));
  NOR3_X1   g536(.A1(new_n706), .A2(G43gat), .A3(new_n694), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n725), .A2(new_n691), .A3(new_n727), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n738), .B1(new_n739), .B2(G43gat), .ZN(new_n740));
  INV_X1    g539(.A(new_n723), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n223), .B1(new_n741), .B2(new_n691), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT47), .ZN(new_n743));
  OR2_X1    g542(.A1(new_n738), .A2(new_n743), .ZN(new_n744));
  OAI22_X1  g543(.A1(new_n740), .A2(KEYINPUT47), .B1(new_n742), .B2(new_n744), .ZN(G1330gat));
  INV_X1    g544(.A(new_n222), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n746), .B1(new_n723), .B2(new_n573), .ZN(new_n747));
  AND2_X1   g546(.A1(new_n706), .A2(KEYINPUT112), .ZN(new_n748));
  OAI211_X1 g547(.A(new_n563), .B(new_n222), .C1(new_n706), .C2(KEYINPUT112), .ZN(new_n749));
  OAI211_X1 g548(.A(new_n747), .B(KEYINPUT48), .C1(new_n748), .C2(new_n749), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n749), .A2(new_n748), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n725), .A2(new_n563), .A3(new_n727), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n751), .B1(new_n752), .B2(new_n746), .ZN(new_n753));
  XNOR2_X1  g552(.A(KEYINPUT111), .B(KEYINPUT48), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n750), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(KEYINPUT113), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT113), .ZN(new_n757));
  OAI211_X1 g556(.A(new_n757), .B(new_n750), .C1(new_n753), .C2(new_n754), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n756), .A2(new_n758), .ZN(G1331gat));
  INV_X1    g558(.A(new_n710), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n674), .A2(new_n264), .A3(new_n646), .ZN(new_n761));
  AOI211_X1 g560(.A(new_n760), .B(new_n761), .C1(new_n568), .C2(new_n581), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(new_n726), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n763), .B(G57gat), .ZN(G1332gat));
  XNOR2_X1  g563(.A(new_n481), .B(KEYINPUT114), .ZN(new_n765));
  INV_X1    g564(.A(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n762), .A2(new_n766), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n767), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n768));
  XOR2_X1   g567(.A(KEYINPUT49), .B(G64gat), .Z(new_n769));
  OAI21_X1  g568(.A(new_n768), .B1(new_n767), .B2(new_n769), .ZN(G1333gat));
  NAND2_X1  g569(.A1(new_n762), .A2(new_n691), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n694), .A2(G71gat), .ZN(new_n772));
  AOI22_X1  g571(.A1(new_n771), .A2(G71gat), .B1(new_n762), .B2(new_n772), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n773), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g573(.A1(new_n762), .A2(new_n563), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(G78gat), .ZN(G1335gat));
  OR2_X1    g575(.A1(new_n719), .A2(new_n722), .ZN(new_n777));
  AND3_X1   g576(.A1(new_n253), .A2(KEYINPUT89), .A3(new_n260), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n260), .B1(new_n253), .B2(KEYINPUT89), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n780), .A2(new_n646), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(new_n704), .ZN(new_n782));
  INV_X1    g581(.A(new_n782), .ZN(new_n783));
  AND2_X1   g582(.A1(new_n777), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(new_n726), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(G85gat), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n674), .B1(new_n568), .B2(new_n581), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(new_n781), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT51), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n787), .A2(KEYINPUT51), .A3(new_n781), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n633), .B1(new_n792), .B2(KEYINPUT115), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n793), .B1(KEYINPUT115), .B2(new_n792), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n726), .A2(new_n594), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n786), .B1(new_n794), .B2(new_n795), .ZN(G1336gat));
  AOI21_X1  g595(.A(new_n760), .B1(new_n790), .B2(new_n791), .ZN(new_n797));
  AND3_X1   g596(.A1(new_n797), .A2(new_n595), .A3(new_n766), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n798), .A2(KEYINPUT52), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n784), .A2(new_n766), .ZN(new_n800));
  INV_X1    g599(.A(new_n800), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n799), .B1(new_n595), .B2(new_n801), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n595), .B1(new_n784), .B2(new_n481), .ZN(new_n803));
  OAI21_X1  g602(.A(KEYINPUT52), .B1(new_n803), .B2(new_n798), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n802), .A2(new_n804), .ZN(G1337gat));
  NAND2_X1  g604(.A1(new_n784), .A2(new_n691), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(G99gat), .ZN(new_n807));
  OR2_X1    g606(.A1(new_n694), .A2(G99gat), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n807), .B1(new_n794), .B2(new_n808), .ZN(G1338gat));
  NAND2_X1  g608(.A1(new_n784), .A2(new_n563), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n810), .A2(G106gat), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n573), .A2(G106gat), .ZN(new_n812));
  AND2_X1   g611(.A1(new_n797), .A2(new_n812), .ZN(new_n813));
  OAI21_X1  g612(.A(KEYINPUT53), .B1(new_n811), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n784), .A2(new_n323), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(G106gat), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n813), .A2(KEYINPUT53), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT116), .ZN(new_n818));
  AND3_X1   g617(.A1(new_n816), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n818), .B1(new_n816), .B2(new_n817), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n814), .B1(new_n819), .B2(new_n820), .ZN(G1339gat));
  NAND3_X1  g620(.A1(new_n618), .A2(new_n624), .A3(new_n619), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n622), .A2(KEYINPUT54), .A3(new_n822), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n624), .B1(new_n618), .B2(new_n619), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT54), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n630), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n823), .A2(KEYINPUT55), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(new_n703), .ZN(new_n828));
  AOI21_X1  g627(.A(KEYINPUT55), .B1(new_n823), .B2(new_n826), .ZN(new_n829));
  OAI21_X1  g628(.A(KEYINPUT117), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n823), .A2(new_n826), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT55), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT117), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n833), .A2(new_n834), .A3(new_n703), .A4(new_n827), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n830), .A2(new_n780), .A3(new_n835), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n249), .A2(new_n251), .A3(new_n252), .A4(new_n260), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n243), .A2(new_n244), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n247), .A2(new_n248), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n259), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n837), .A2(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(new_n704), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n836), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(new_n674), .ZN(new_n845));
  NAND4_X1  g644(.A1(new_n718), .A2(new_n842), .A3(new_n830), .A4(new_n835), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n646), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n761), .A2(new_n704), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n766), .A2(new_n564), .ZN(new_n851));
  NAND4_X1  g650(.A1(new_n850), .A2(new_n697), .A3(new_n577), .A4(new_n851), .ZN(new_n852));
  NOR3_X1   g651(.A1(new_n852), .A2(new_n334), .A3(new_n264), .ZN(new_n853));
  OR3_X1    g652(.A1(new_n849), .A2(new_n564), .A3(new_n575), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n854), .A2(new_n766), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(new_n780), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n853), .B1(new_n856), .B2(new_n334), .ZN(G1340gat));
  NOR3_X1   g656(.A1(new_n854), .A2(new_n633), .A3(new_n766), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n710), .A2(G120gat), .ZN(new_n859));
  OAI22_X1  g658(.A1(new_n858), .A2(G120gat), .B1(new_n852), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(KEYINPUT118), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT118), .ZN(new_n862));
  OAI221_X1 g661(.A(new_n862), .B1(new_n852), .B2(new_n859), .C1(new_n858), .C2(G120gat), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n861), .A2(new_n863), .ZN(G1341gat));
  NAND3_X1  g663(.A1(new_n855), .A2(new_n327), .A3(new_n646), .ZN(new_n865));
  INV_X1    g664(.A(new_n646), .ZN(new_n866));
  OAI21_X1  g665(.A(G127gat), .B1(new_n852), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n865), .A2(new_n867), .ZN(G1342gat));
  INV_X1    g667(.A(new_n854), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n674), .A2(new_n481), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n869), .A2(new_n329), .A3(new_n870), .ZN(new_n871));
  OR2_X1    g670(.A1(new_n871), .A2(KEYINPUT56), .ZN(new_n872));
  OAI21_X1  g671(.A(G134gat), .B1(new_n852), .B2(new_n674), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n871), .A2(KEYINPUT56), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(G1343gat));
  OAI21_X1  g674(.A(KEYINPUT121), .B1(new_n849), .B2(new_n564), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT121), .ZN(new_n877));
  OAI211_X1 g676(.A(new_n877), .B(new_n726), .C1(new_n847), .C2(new_n848), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n692), .A2(new_n323), .ZN(new_n880));
  XNOR2_X1  g679(.A(new_n880), .B(KEYINPUT122), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n780), .A2(new_n285), .ZN(new_n882));
  XNOR2_X1  g681(.A(new_n882), .B(KEYINPUT123), .ZN(new_n883));
  NAND4_X1  g682(.A1(new_n879), .A2(new_n881), .A3(new_n765), .A4(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n692), .A2(new_n851), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT57), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n887), .B1(new_n849), .B2(new_n573), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n697), .A2(new_n887), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n833), .A2(new_n703), .A3(new_n827), .ZN(new_n890));
  INV_X1    g689(.A(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(new_n780), .ZN(new_n892));
  OAI21_X1  g691(.A(KEYINPUT119), .B1(new_n633), .B2(new_n841), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT119), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n704), .A2(new_n894), .A3(new_n840), .A4(new_n837), .ZN(new_n895));
  AND2_X1   g694(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(KEYINPUT120), .B1(new_n892), .B2(new_n896), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n264), .A2(new_n890), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n893), .A2(new_n895), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT120), .ZN(new_n900));
  NOR3_X1   g699(.A1(new_n898), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n674), .B1(new_n897), .B2(new_n901), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n646), .B1(new_n902), .B2(new_n846), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n889), .B1(new_n903), .B2(new_n848), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n886), .B1(new_n888), .B2(new_n904), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n285), .B1(new_n905), .B2(new_n780), .ZN(new_n906));
  OAI21_X1  g705(.A(KEYINPUT58), .B1(new_n885), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n888), .A2(new_n904), .ZN(new_n908));
  INV_X1    g707(.A(new_n886), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  OAI21_X1  g709(.A(G141gat), .B1(new_n910), .B2(new_n264), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT58), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n911), .A2(new_n912), .A3(new_n884), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n907), .A2(new_n913), .ZN(G1344gat));
  NAND3_X1  g713(.A1(new_n718), .A2(new_n842), .A3(new_n891), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n646), .B1(new_n902), .B2(new_n915), .ZN(new_n916));
  OAI211_X1 g715(.A(new_n887), .B(new_n563), .C1(new_n916), .C2(new_n848), .ZN(new_n917));
  OAI21_X1  g716(.A(KEYINPUT57), .B1(new_n849), .B2(new_n573), .ZN(new_n918));
  NAND4_X1  g717(.A1(new_n917), .A2(new_n918), .A3(new_n704), .A4(new_n909), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT59), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n920), .A2(new_n287), .ZN(new_n921));
  NOR3_X1   g720(.A1(new_n886), .A2(KEYINPUT59), .A3(new_n633), .ZN(new_n922));
  AOI22_X1  g721(.A1(new_n919), .A2(new_n921), .B1(new_n908), .B2(new_n922), .ZN(new_n923));
  AND3_X1   g722(.A1(new_n879), .A2(new_n765), .A3(new_n881), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n920), .B1(new_n924), .B2(new_n704), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n923), .B1(new_n925), .B2(G148gat), .ZN(G1345gat));
  NAND3_X1  g725(.A1(new_n924), .A2(new_n291), .A3(new_n646), .ZN(new_n927));
  OAI21_X1  g726(.A(G155gat), .B1(new_n910), .B2(new_n866), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(G1346gat));
  OAI21_X1  g728(.A(G162gat), .B1(new_n910), .B2(new_n674), .ZN(new_n930));
  NAND4_X1  g729(.A1(new_n879), .A2(new_n881), .A3(new_n292), .A4(new_n870), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(new_n931), .ZN(G1347gat));
  NOR3_X1   g731(.A1(new_n694), .A2(new_n726), .A3(new_n682), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n850), .A2(new_n697), .A3(new_n933), .ZN(new_n934));
  NOR3_X1   g733(.A1(new_n934), .A2(new_n391), .A3(new_n264), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n849), .A2(new_n726), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n765), .A2(new_n575), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n936), .A2(new_n780), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n935), .B1(new_n391), .B2(new_n938), .ZN(G1348gat));
  OAI21_X1  g738(.A(G176gat), .B1(new_n934), .B2(new_n760), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n936), .A2(new_n937), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n704), .A2(new_n392), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n940), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT124), .ZN(new_n944));
  XNOR2_X1  g743(.A(new_n943), .B(new_n944), .ZN(G1349gat));
  OAI21_X1  g744(.A(G183gat), .B1(new_n934), .B2(new_n866), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n646), .A2(new_n420), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n946), .B1(new_n941), .B2(new_n947), .ZN(new_n948));
  XNOR2_X1  g747(.A(new_n948), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g748(.A(G190gat), .B1(new_n934), .B2(new_n674), .ZN(new_n950));
  XOR2_X1   g749(.A(KEYINPUT126), .B(KEYINPUT61), .Z(new_n951));
  XNOR2_X1  g750(.A(new_n950), .B(new_n951), .ZN(new_n952));
  AND4_X1   g751(.A1(new_n399), .A2(new_n936), .A3(new_n718), .A4(new_n937), .ZN(new_n953));
  XNOR2_X1  g752(.A(new_n953), .B(KEYINPUT125), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n952), .A2(new_n954), .ZN(G1351gat));
  NOR3_X1   g754(.A1(new_n691), .A2(new_n726), .A3(new_n682), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n917), .A2(new_n918), .A3(new_n956), .ZN(new_n957));
  OAI21_X1  g756(.A(G197gat), .B1(new_n957), .B2(new_n264), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT127), .ZN(new_n959));
  NOR2_X1   g758(.A1(new_n880), .A2(new_n765), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n936), .A2(new_n960), .ZN(new_n961));
  INV_X1    g760(.A(new_n961), .ZN(new_n962));
  NOR2_X1   g761(.A1(new_n264), .A2(G197gat), .ZN(new_n963));
  AOI21_X1  g762(.A(new_n959), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NOR4_X1   g763(.A1(new_n961), .A2(KEYINPUT127), .A3(G197gat), .A4(new_n264), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n958), .B1(new_n964), .B2(new_n965), .ZN(G1352gat));
  NOR2_X1   g765(.A1(new_n633), .A2(G204gat), .ZN(new_n967));
  INV_X1    g766(.A(new_n967), .ZN(new_n968));
  OR3_X1    g767(.A1(new_n961), .A2(KEYINPUT62), .A3(new_n968), .ZN(new_n969));
  OAI21_X1  g768(.A(G204gat), .B1(new_n957), .B2(new_n760), .ZN(new_n970));
  OAI21_X1  g769(.A(KEYINPUT62), .B1(new_n961), .B2(new_n968), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n969), .A2(new_n970), .A3(new_n971), .ZN(G1353gat));
  NAND3_X1  g771(.A1(new_n962), .A2(new_n267), .A3(new_n646), .ZN(new_n973));
  NAND4_X1  g772(.A1(new_n917), .A2(new_n918), .A3(new_n646), .A4(new_n956), .ZN(new_n974));
  AND3_X1   g773(.A1(new_n974), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n975));
  AOI21_X1  g774(.A(KEYINPUT63), .B1(new_n974), .B2(G211gat), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n973), .B1(new_n975), .B2(new_n976), .ZN(G1354gat));
  OAI21_X1  g776(.A(G218gat), .B1(new_n957), .B2(new_n674), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n962), .A2(new_n268), .A3(new_n718), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n978), .A2(new_n979), .ZN(G1355gat));
endmodule


