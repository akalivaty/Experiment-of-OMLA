//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 0 0 0 1 0 0 1 1 0 1 0 0 0 1 1 0 0 0 1 0 0 0 1 0 0 1 0 0 1 0 1 1 0 1 1 0 1 1 0 1 0 0 1 0 1 0 0 0 1 1 0 1 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:19 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n543, new_n544, new_n545, new_n546, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n561, new_n563, new_n564, new_n565,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n584, new_n586, new_n587, new_n588, new_n589, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n622, new_n625,
    new_n627, new_n628, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1153, new_n1154,
    new_n1155;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT64), .Z(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(new_n451), .ZN(new_n456));
  INV_X1    g031(.A(new_n452), .ZN(new_n457));
  AOI22_X1  g032(.A1(new_n456), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  INV_X1    g033(.A(G2104), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(KEYINPUT65), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT65), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G2104), .ZN(new_n462));
  AOI21_X1  g037(.A(G2105), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  AND3_X1   g038(.A1(new_n463), .A2(KEYINPUT66), .A3(G101), .ZN(new_n464));
  AOI21_X1  g039(.A(KEYINPUT66), .B1(new_n463), .B2(G101), .ZN(new_n465));
  OR2_X1    g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n460), .A2(new_n462), .A3(KEYINPUT3), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G137), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n459), .A2(KEYINPUT3), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n469), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(G125), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n473), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G2105), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n466), .A2(new_n472), .A3(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G160));
  NAND2_X1  g055(.A1(new_n471), .A2(G136), .ZN(new_n481));
  INV_X1    g056(.A(G2105), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n470), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  OR2_X1    g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(G2104), .C1(G112), .C2(new_n482), .ZN(new_n486));
  XNOR2_X1  g061(.A(new_n486), .B(KEYINPUT67), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n481), .A2(new_n484), .A3(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  OAI21_X1  g064(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  OR2_X1    g066(.A1(new_n482), .A2(G114), .ZN(new_n492));
  AND2_X1   g067(.A1(new_n492), .A2(KEYINPUT68), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n492), .A2(KEYINPUT68), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n491), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n467), .A2(G126), .A3(G2105), .A4(new_n469), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(G138), .ZN(new_n498));
  NOR4_X1   g073(.A1(new_n475), .A2(KEYINPUT4), .A3(new_n498), .A4(G2105), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n498), .A2(G2105), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n467), .A2(new_n469), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT4), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n499), .B1(new_n502), .B2(KEYINPUT69), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT69), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n501), .A2(new_n504), .A3(KEYINPUT4), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n497), .B1(new_n503), .B2(new_n505), .ZN(G164));
  INV_X1    g081(.A(KEYINPUT6), .ZN(new_n507));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(KEYINPUT70), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT70), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G651), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n507), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  NOR2_X1   g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  OAI21_X1  g088(.A(G543), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G50), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT5), .ZN(new_n517));
  INV_X1    g092(.A(G543), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(KEYINPUT5), .A2(G543), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n521), .B1(new_n512), .B2(new_n513), .ZN(new_n522));
  INV_X1    g097(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G88), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n521), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n509), .A2(new_n511), .ZN(new_n526));
  INV_X1    g101(.A(new_n526), .ZN(new_n527));
  OR2_X1    g102(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n516), .A2(new_n524), .A3(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(new_n529), .ZN(G166));
  AND2_X1   g105(.A1(G63), .A2(G651), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n515), .A2(G51), .B1(new_n521), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g107(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n533), .B(KEYINPUT7), .ZN(new_n534));
  INV_X1    g109(.A(G89), .ZN(new_n535));
  OAI211_X1 g110(.A(KEYINPUT71), .B(new_n534), .C1(new_n522), .C2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n532), .A2(new_n536), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n534), .B1(new_n522), .B2(new_n535), .ZN(new_n538));
  INV_X1    g113(.A(KEYINPUT71), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(new_n540), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n537), .A2(new_n541), .ZN(G168));
  NAND2_X1  g117(.A1(new_n523), .A2(G90), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n515), .A2(G52), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n521), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n545));
  OR2_X1    g120(.A1(new_n545), .A2(new_n527), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n543), .A2(new_n544), .A3(new_n546), .ZN(G301));
  INV_X1    g122(.A(G301), .ZN(G171));
  OAI211_X1 g123(.A(G43), .B(G543), .C1(new_n512), .C2(new_n513), .ZN(new_n549));
  OAI211_X1 g124(.A(G81), .B(new_n521), .C1(new_n512), .C2(new_n513), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT72), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n549), .A2(new_n550), .A3(KEYINPUT72), .ZN(new_n554));
  NAND2_X1  g129(.A1(G68), .A2(G543), .ZN(new_n555));
  INV_X1    g130(.A(new_n521), .ZN(new_n556));
  INV_X1    g131(.A(G56), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n555), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n553), .A2(new_n554), .B1(new_n526), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G860), .ZN(G153));
  NAND4_X1  g135(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n561));
  XOR2_X1   g136(.A(new_n561), .B(KEYINPUT73), .Z(G176));
  NAND2_X1  g137(.A1(G1), .A2(G3), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT8), .ZN(new_n564));
  NAND4_X1  g139(.A1(G319), .A2(G483), .A3(G661), .A4(new_n564), .ZN(new_n565));
  XOR2_X1   g140(.A(new_n565), .B(KEYINPUT74), .Z(G188));
  OAI211_X1 g141(.A(G53), .B(G543), .C1(new_n512), .C2(new_n513), .ZN(new_n567));
  NAND2_X1  g142(.A1(KEYINPUT75), .A2(KEYINPUT9), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n567), .B(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(G65), .ZN(new_n570));
  INV_X1    g145(.A(new_n520), .ZN(new_n571));
  NOR2_X1   g146(.A1(KEYINPUT5), .A2(G543), .ZN(new_n572));
  OAI21_X1  g147(.A(KEYINPUT76), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT76), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n519), .A2(new_n574), .A3(new_n520), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n570), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  AND2_X1   g151(.A1(G78), .A2(G543), .ZN(new_n577));
  OAI21_X1  g152(.A(G651), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  OAI211_X1 g153(.A(G91), .B(new_n521), .C1(new_n512), .C2(new_n513), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n569), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(G299));
  INV_X1    g157(.A(G168), .ZN(G286));
  INV_X1    g158(.A(KEYINPUT77), .ZN(new_n584));
  XNOR2_X1  g159(.A(new_n529), .B(new_n584), .ZN(G303));
  NAND2_X1  g160(.A1(new_n515), .A2(G49), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n523), .A2(G87), .ZN(new_n587));
  OAI21_X1  g162(.A(G651), .B1(new_n521), .B2(G74), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  XNOR2_X1  g164(.A(new_n589), .B(KEYINPUT78), .ZN(G288));
  OAI211_X1 g165(.A(G48), .B(G543), .C1(new_n512), .C2(new_n513), .ZN(new_n591));
  INV_X1    g166(.A(G61), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n592), .B1(new_n519), .B2(new_n520), .ZN(new_n593));
  AND2_X1   g168(.A1(G73), .A2(G543), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n526), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(G86), .ZN(new_n596));
  OAI211_X1 g171(.A(new_n591), .B(new_n595), .C1(new_n522), .C2(new_n596), .ZN(G305));
  NAND2_X1  g172(.A1(G72), .A2(G543), .ZN(new_n598));
  INV_X1    g173(.A(G60), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n556), .B2(new_n599), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n515), .A2(G47), .B1(new_n600), .B2(new_n526), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n523), .A2(G85), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n601), .A2(new_n602), .ZN(G290));
  INV_X1    g178(.A(G868), .ZN(new_n604));
  NOR2_X1   g179(.A1(G301), .A2(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(G92), .ZN(new_n606));
  OR3_X1    g181(.A1(new_n522), .A2(KEYINPUT79), .A3(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(KEYINPUT79), .B1(new_n522), .B2(new_n606), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT10), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n515), .A2(G54), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n573), .A2(new_n575), .ZN(new_n613));
  AOI22_X1  g188(.A1(new_n613), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n612), .B1(new_n508), .B2(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(new_n615), .ZN(new_n616));
  NAND3_X1  g191(.A1(new_n607), .A2(KEYINPUT10), .A3(new_n608), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n611), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT80), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n605), .B1(new_n619), .B2(new_n604), .ZN(G284));
  AOI21_X1  g195(.A(new_n605), .B1(new_n619), .B2(new_n604), .ZN(G321));
  NAND2_X1  g196(.A1(G299), .A2(new_n604), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(G168), .B2(new_n604), .ZN(G297));
  OAI21_X1  g198(.A(new_n622), .B1(G168), .B2(new_n604), .ZN(G280));
  INV_X1    g199(.A(G559), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n619), .B1(new_n625), .B2(G860), .ZN(G148));
  NAND2_X1  g201(.A1(new_n619), .A2(new_n625), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n627), .A2(G868), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n628), .B1(G868), .B2(new_n559), .ZN(G323));
  XNOR2_X1  g204(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g205(.A(new_n475), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n631), .A2(new_n463), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT12), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT13), .ZN(new_n634));
  INV_X1    g209(.A(G2100), .ZN(new_n635));
  AOI21_X1  g210(.A(new_n634), .B1(KEYINPUT81), .B2(new_n635), .ZN(new_n636));
  NOR2_X1   g211(.A1(new_n635), .A2(KEYINPUT81), .ZN(new_n637));
  MUX2_X1   g212(.A(new_n636), .B(new_n634), .S(new_n637), .Z(new_n638));
  NAND2_X1  g213(.A1(new_n471), .A2(G135), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n483), .A2(G123), .ZN(new_n640));
  NOR2_X1   g215(.A1(new_n482), .A2(G111), .ZN(new_n641));
  OAI21_X1  g216(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n642));
  OAI211_X1 g217(.A(new_n639), .B(new_n640), .C1(new_n641), .C2(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT82), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n644), .B(G2096), .Z(new_n645));
  NAND2_X1  g220(.A1(new_n638), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT83), .ZN(G156));
  XNOR2_X1  g222(.A(G2427), .B(G2438), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(G2430), .ZN(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT15), .B(G2435), .ZN(new_n650));
  OR2_X1    g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n649), .A2(new_n650), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n651), .A2(KEYINPUT14), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G1341), .B(G1348), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2443), .B(G2446), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n653), .B(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G2451), .B(G2454), .Z(new_n658));
  XNOR2_X1  g233(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n661), .A2(G14), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n657), .A2(new_n660), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n662), .A2(new_n663), .ZN(G401));
  XOR2_X1   g239(.A(KEYINPUT85), .B(KEYINPUT18), .Z(new_n665));
  XOR2_X1   g240(.A(G2084), .B(G2090), .Z(new_n666));
  XNOR2_X1  g241(.A(G2067), .B(G2678), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  AND2_X1   g243(.A1(new_n668), .A2(KEYINPUT17), .ZN(new_n669));
  OR2_X1    g244(.A1(new_n666), .A2(new_n667), .ZN(new_n670));
  AOI21_X1  g245(.A(new_n665), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(G2072), .B(G2078), .Z(new_n672));
  AOI21_X1  g247(.A(new_n672), .B1(new_n668), .B2(new_n665), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n671), .B(new_n673), .Z(new_n674));
  XNOR2_X1  g249(.A(G2096), .B(G2100), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(G227));
  XOR2_X1   g251(.A(G1971), .B(G1976), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT19), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1956), .B(G2474), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1961), .B(G1966), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  AND2_X1   g256(.A1(new_n679), .A2(new_n680), .ZN(new_n682));
  NOR3_X1   g257(.A1(new_n678), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n678), .A2(new_n681), .ZN(new_n684));
  XOR2_X1   g259(.A(new_n684), .B(KEYINPUT20), .Z(new_n685));
  AOI211_X1 g260(.A(new_n683), .B(new_n685), .C1(new_n678), .C2(new_n682), .ZN(new_n686));
  XOR2_X1   g261(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1991), .B(G1996), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1981), .B(G1986), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(G229));
  INV_X1    g267(.A(G16), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n693), .A2(G23), .ZN(new_n694));
  INV_X1    g269(.A(new_n589), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n694), .B1(new_n695), .B2(new_n693), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT33), .B(G1976), .ZN(new_n697));
  XOR2_X1   g272(.A(new_n696), .B(new_n697), .Z(new_n698));
  NAND2_X1  g273(.A1(new_n693), .A2(G22), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(G166), .B2(new_n693), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(G1971), .ZN(new_n701));
  MUX2_X1   g276(.A(G6), .B(G305), .S(G16), .Z(new_n702));
  XOR2_X1   g277(.A(KEYINPUT32), .B(G1981), .Z(new_n703));
  XOR2_X1   g278(.A(new_n702), .B(new_n703), .Z(new_n704));
  NOR3_X1   g279(.A1(new_n698), .A2(new_n701), .A3(new_n704), .ZN(new_n705));
  XOR2_X1   g280(.A(KEYINPUT87), .B(KEYINPUT34), .Z(new_n706));
  OR2_X1    g281(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  MUX2_X1   g282(.A(G24), .B(G290), .S(G16), .Z(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT86), .ZN(new_n709));
  INV_X1    g284(.A(G1986), .ZN(new_n710));
  OR2_X1    g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n471), .A2(G131), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n483), .A2(G119), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n482), .A2(G107), .ZN(new_n714));
  OAI21_X1  g289(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n715));
  OAI211_X1 g290(.A(new_n712), .B(new_n713), .C1(new_n714), .C2(new_n715), .ZN(new_n716));
  MUX2_X1   g291(.A(G25), .B(new_n716), .S(G29), .Z(new_n717));
  XOR2_X1   g292(.A(KEYINPUT35), .B(G1991), .Z(new_n718));
  INV_X1    g293(.A(new_n718), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n717), .B(new_n719), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(KEYINPUT88), .B2(KEYINPUT36), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n709), .A2(new_n710), .ZN(new_n722));
  AND3_X1   g297(.A1(new_n711), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n705), .A2(new_n706), .ZN(new_n724));
  NAND3_X1  g299(.A1(new_n707), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  NOR2_X1   g300(.A1(KEYINPUT88), .A2(KEYINPUT36), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n725), .B(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n471), .A2(G139), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n482), .A2(G103), .A3(G2104), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n729), .B(KEYINPUT25), .Z(new_n730));
  AOI22_X1  g305(.A1(new_n631), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n731));
  OAI211_X1 g306(.A(new_n728), .B(new_n730), .C1(new_n482), .C2(new_n731), .ZN(new_n732));
  MUX2_X1   g307(.A(G33), .B(new_n732), .S(G29), .Z(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(G2072), .ZN(new_n734));
  INV_X1    g309(.A(G29), .ZN(new_n735));
  NOR2_X1   g310(.A1(G162), .A2(new_n735), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(new_n735), .B2(G35), .ZN(new_n737));
  XOR2_X1   g312(.A(KEYINPUT29), .B(G2090), .Z(new_n738));
  NAND2_X1  g313(.A1(new_n735), .A2(G26), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(KEYINPUT28), .Z(new_n740));
  NAND2_X1  g315(.A1(new_n471), .A2(G140), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n483), .A2(G128), .ZN(new_n742));
  INV_X1    g317(.A(G104), .ZN(new_n743));
  AND3_X1   g318(.A1(new_n743), .A2(new_n482), .A3(KEYINPUT90), .ZN(new_n744));
  AOI21_X1  g319(.A(KEYINPUT90), .B1(new_n743), .B2(new_n482), .ZN(new_n745));
  OAI221_X1 g320(.A(G2104), .B1(G116), .B2(new_n482), .C1(new_n744), .C2(new_n745), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n741), .A2(new_n742), .A3(new_n746), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n740), .B1(new_n747), .B2(G29), .ZN(new_n748));
  XOR2_X1   g323(.A(KEYINPUT91), .B(G2067), .Z(new_n749));
  OAI22_X1  g324(.A1(new_n737), .A2(new_n738), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  AOI211_X1 g325(.A(new_n734), .B(new_n750), .C1(new_n737), .C2(new_n738), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n471), .A2(G141), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n752), .B(KEYINPUT92), .Z(new_n753));
  NAND3_X1  g328(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT26), .ZN(new_n755));
  AND2_X1   g330(.A1(new_n463), .A2(G105), .ZN(new_n756));
  AOI211_X1 g331(.A(new_n755), .B(new_n756), .C1(new_n483), .C2(G129), .ZN(new_n757));
  AND2_X1   g332(.A1(new_n753), .A2(new_n757), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n758), .A2(new_n735), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(new_n735), .B2(G32), .ZN(new_n760));
  XNOR2_X1  g335(.A(KEYINPUT27), .B(G1996), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT93), .ZN(new_n762));
  INV_X1    g337(.A(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n760), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n748), .A2(new_n749), .ZN(new_n765));
  INV_X1    g340(.A(G2084), .ZN(new_n766));
  INV_X1    g341(.A(G34), .ZN(new_n767));
  AOI21_X1  g342(.A(G29), .B1(new_n767), .B2(KEYINPUT24), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(KEYINPUT24), .B2(new_n767), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(new_n479), .B2(new_n735), .ZN(new_n770));
  NOR2_X1   g345(.A1(G171), .A2(new_n693), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(G5), .B2(new_n693), .ZN(new_n772));
  INV_X1    g347(.A(G1961), .ZN(new_n773));
  OAI221_X1 g348(.A(new_n765), .B1(new_n766), .B2(new_n770), .C1(new_n772), .C2(new_n773), .ZN(new_n774));
  INV_X1    g349(.A(G1341), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n559), .A2(G16), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(G16), .B2(G19), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n774), .B1(new_n775), .B2(new_n777), .ZN(new_n778));
  NAND3_X1  g353(.A1(new_n751), .A2(new_n764), .A3(new_n778), .ZN(new_n779));
  NOR2_X1   g354(.A1(G168), .A2(new_n693), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(new_n693), .B2(G21), .ZN(new_n781));
  INV_X1    g356(.A(G1966), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT96), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n693), .A2(G20), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(KEYINPUT23), .Z(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(G299), .B2(G16), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(G1956), .ZN(new_n788));
  OAI221_X1 g363(.A(new_n788), .B1(new_n775), .B2(new_n777), .C1(new_n781), .C2(new_n782), .ZN(new_n789));
  OR3_X1    g364(.A1(new_n779), .A2(new_n784), .A3(new_n789), .ZN(new_n790));
  XNOR2_X1  g365(.A(KEYINPUT31), .B(G11), .ZN(new_n791));
  XOR2_X1   g366(.A(KEYINPUT94), .B(G28), .Z(new_n792));
  NOR2_X1   g367(.A1(new_n792), .A2(KEYINPUT30), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n792), .A2(KEYINPUT30), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n794), .A2(new_n735), .ZN(new_n795));
  OAI221_X1 g370(.A(new_n791), .B1(new_n793), .B2(new_n795), .C1(new_n644), .C2(new_n735), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(KEYINPUT95), .Z(new_n797));
  AOI22_X1  g372(.A1(new_n772), .A2(new_n773), .B1(new_n766), .B2(new_n770), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(new_n760), .B2(new_n763), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n797), .B1(KEYINPUT97), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n735), .A2(G27), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(G164), .B2(new_n735), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT98), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(G2078), .ZN(new_n804));
  OAI211_X1 g379(.A(new_n800), .B(new_n804), .C1(KEYINPUT97), .C2(new_n799), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n693), .A2(G4), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(new_n619), .B2(new_n693), .ZN(new_n807));
  XOR2_X1   g382(.A(KEYINPUT89), .B(G1348), .Z(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NOR4_X1   g384(.A1(new_n727), .A2(new_n790), .A3(new_n805), .A4(new_n809), .ZN(G311));
  INV_X1    g385(.A(G311), .ZN(G150));
  NAND2_X1  g386(.A1(new_n619), .A2(G559), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT38), .ZN(new_n813));
  OAI211_X1 g388(.A(G55), .B(G543), .C1(new_n512), .C2(new_n513), .ZN(new_n814));
  AOI22_X1  g389(.A1(new_n521), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n815));
  INV_X1    g390(.A(G93), .ZN(new_n816));
  OAI221_X1 g391(.A(new_n814), .B1(new_n815), .B2(new_n527), .C1(new_n522), .C2(new_n816), .ZN(new_n817));
  OAI21_X1  g392(.A(KEYINPUT100), .B1(new_n559), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n558), .A2(new_n526), .ZN(new_n819));
  INV_X1    g394(.A(new_n554), .ZN(new_n820));
  AOI21_X1  g395(.A(KEYINPUT72), .B1(new_n549), .B2(new_n550), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n819), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT100), .ZN(new_n823));
  INV_X1    g398(.A(new_n817), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n822), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  AND2_X1   g400(.A1(new_n818), .A2(new_n825), .ZN(new_n826));
  OAI211_X1 g401(.A(new_n817), .B(new_n819), .C1(new_n820), .C2(new_n821), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT99), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n826), .A2(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n813), .B(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT39), .ZN(new_n832));
  AOI21_X1  g407(.A(G860), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n833), .B1(new_n832), .B2(new_n831), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n817), .A2(G860), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT101), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT37), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n834), .A2(new_n837), .ZN(G145));
  XNOR2_X1  g413(.A(new_n758), .B(G164), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(new_n716), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n747), .B(KEYINPUT102), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(new_n732), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n483), .A2(G130), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n482), .A2(G118), .ZN(new_n844));
  OAI21_X1  g419(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n843), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n846), .B1(G142), .B2(new_n471), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n847), .B(new_n633), .Z(new_n848));
  XNOR2_X1  g423(.A(new_n842), .B(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n840), .B(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n644), .B(new_n488), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(new_n479), .ZN(new_n852));
  AOI21_X1  g427(.A(G37), .B1(new_n850), .B2(new_n852), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n853), .B1(new_n852), .B2(new_n850), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g430(.A1(new_n817), .A2(new_n604), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n627), .B(new_n830), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n618), .A2(G299), .ZN(new_n858));
  NAND4_X1  g433(.A1(new_n611), .A2(new_n581), .A3(new_n617), .A4(new_n616), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  AND3_X1   g436(.A1(new_n858), .A2(KEYINPUT41), .A3(new_n859), .ZN(new_n862));
  AOI21_X1  g437(.A(KEYINPUT41), .B1(new_n858), .B2(new_n859), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n861), .B1(new_n857), .B2(new_n864), .ZN(new_n865));
  XOR2_X1   g440(.A(G290), .B(G305), .Z(new_n866));
  XOR2_X1   g441(.A(new_n529), .B(new_n589), .Z(new_n867));
  OR2_X1    g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n866), .A2(new_n867), .ZN(new_n869));
  AOI21_X1  g444(.A(KEYINPUT42), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  AOI21_X1  g445(.A(KEYINPUT103), .B1(new_n868), .B2(new_n869), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n868), .A2(KEYINPUT103), .A3(new_n869), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n870), .B1(new_n874), .B2(KEYINPUT42), .ZN(new_n875));
  XOR2_X1   g450(.A(new_n865), .B(new_n875), .Z(new_n876));
  OAI21_X1  g451(.A(new_n856), .B1(new_n876), .B2(new_n604), .ZN(G295));
  OAI21_X1  g452(.A(new_n856), .B1(new_n876), .B2(new_n604), .ZN(G331));
  NAND4_X1  g453(.A1(G171), .A2(new_n540), .A3(new_n536), .A4(new_n532), .ZN(new_n879));
  OAI21_X1  g454(.A(G301), .B1(new_n537), .B2(new_n541), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n882), .B1(new_n826), .B2(new_n829), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT104), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n827), .B(KEYINPUT99), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n818), .A2(new_n825), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n885), .A2(new_n886), .A3(new_n881), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n883), .A2(new_n884), .A3(new_n887), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n830), .A2(KEYINPUT104), .A3(new_n881), .ZN(new_n889));
  AND3_X1   g464(.A1(new_n888), .A2(new_n889), .A3(new_n864), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n883), .A2(KEYINPUT105), .A3(new_n887), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT105), .ZN(new_n892));
  OAI211_X1 g467(.A(new_n882), .B(new_n892), .C1(new_n826), .C2(new_n829), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n860), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n890), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n873), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n896), .A2(new_n871), .ZN(new_n897));
  AOI21_X1  g472(.A(G37), .B1(new_n895), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n874), .B1(new_n890), .B2(new_n894), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n900), .A2(KEYINPUT43), .ZN(new_n901));
  AND3_X1   g476(.A1(new_n891), .A2(new_n864), .A3(new_n893), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n860), .B1(new_n888), .B2(new_n889), .ZN(new_n903));
  OAI211_X1 g478(.A(KEYINPUT106), .B(new_n874), .C1(new_n902), .C2(new_n903), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n874), .B1(new_n902), .B2(new_n903), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT106), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n898), .A2(new_n904), .A3(new_n907), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n901), .B1(KEYINPUT43), .B2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT44), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n910), .B1(new_n908), .B2(KEYINPUT43), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT43), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n898), .A2(KEYINPUT107), .A3(new_n913), .A4(new_n899), .ZN(new_n914));
  INV_X1    g489(.A(new_n894), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n888), .A2(new_n864), .A3(new_n889), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n915), .A2(new_n897), .A3(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(G37), .ZN(new_n918));
  NAND4_X1  g493(.A1(new_n917), .A2(new_n899), .A3(new_n913), .A4(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT107), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n914), .A2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT108), .ZN(new_n923));
  AND3_X1   g498(.A1(new_n912), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n923), .B1(new_n912), .B2(new_n922), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n911), .B1(new_n924), .B2(new_n925), .ZN(G397));
  NAND2_X1  g501(.A1(new_n502), .A2(KEYINPUT69), .ZN(new_n927));
  INV_X1    g502(.A(new_n499), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n927), .A2(new_n505), .A3(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(new_n497), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  XNOR2_X1  g506(.A(KEYINPUT109), .B(G1384), .ZN(new_n932));
  AOI21_X1  g507(.A(KEYINPUT45), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND4_X1  g508(.A1(new_n466), .A2(G40), .A3(new_n472), .A4(new_n478), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(new_n936), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n758), .B(G1996), .ZN(new_n938));
  XOR2_X1   g513(.A(new_n747), .B(G2067), .Z(new_n939));
  AND2_X1   g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  XNOR2_X1  g516(.A(new_n716), .B(new_n719), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n937), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n601), .A2(new_n710), .A3(new_n602), .ZN(new_n944));
  NAND2_X1  g519(.A1(G290), .A2(G1986), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n936), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  XNOR2_X1  g521(.A(new_n946), .B(KEYINPUT110), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n943), .A2(new_n947), .ZN(new_n948));
  XOR2_X1   g523(.A(new_n948), .B(KEYINPUT111), .Z(new_n949));
  INV_X1    g524(.A(KEYINPUT112), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n950), .B1(G164), .B2(G1384), .ZN(new_n951));
  INV_X1    g526(.A(G1384), .ZN(new_n952));
  AND3_X1   g527(.A1(new_n501), .A2(new_n504), .A3(KEYINPUT4), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n504), .B1(new_n501), .B2(KEYINPUT4), .ZN(new_n954));
  NOR3_X1   g529(.A1(new_n953), .A2(new_n954), .A3(new_n499), .ZN(new_n955));
  OAI211_X1 g530(.A(KEYINPUT112), .B(new_n952), .C1(new_n955), .C2(new_n497), .ZN(new_n956));
  AOI21_X1  g531(.A(KEYINPUT45), .B1(new_n951), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n931), .A2(new_n952), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT45), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n935), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT53), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n961), .A2(G2078), .ZN(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  OR3_X1    g538(.A1(new_n957), .A2(new_n960), .A3(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n934), .B1(new_n958), .B2(KEYINPUT50), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n951), .A2(new_n956), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n965), .B1(new_n966), .B2(KEYINPUT50), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(new_n773), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n931), .A2(KEYINPUT45), .A3(new_n932), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n959), .B1(G164), .B2(G1384), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n969), .A2(new_n970), .A3(new_n935), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n961), .B1(new_n971), .B2(G2078), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n964), .A2(new_n968), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(G171), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n933), .A2(new_n963), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n975), .A2(new_n935), .A3(new_n969), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n968), .A2(G301), .A3(new_n972), .A4(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(KEYINPUT54), .B1(new_n974), .B2(new_n977), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n968), .A2(new_n972), .A3(new_n976), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(G171), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT125), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n979), .A2(KEYINPUT125), .A3(G171), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT54), .ZN(new_n985));
  INV_X1    g560(.A(new_n973), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n985), .B1(new_n986), .B2(G301), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n978), .B1(new_n984), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(G303), .A2(G8), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT55), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND3_X1  g566(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(new_n993), .ZN(new_n994));
  AOI21_X1  g569(.A(KEYINPUT112), .B1(new_n931), .B2(new_n952), .ZN(new_n995));
  NOR3_X1   g570(.A1(G164), .A2(new_n950), .A3(G1384), .ZN(new_n996));
  OAI21_X1  g571(.A(KEYINPUT50), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT50), .ZN(new_n998));
  OAI211_X1 g573(.A(new_n998), .B(new_n952), .C1(new_n955), .C2(new_n497), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT116), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n931), .A2(KEYINPUT116), .A3(new_n998), .A4(new_n952), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n997), .A2(new_n1003), .A3(new_n935), .ZN(new_n1004));
  OR2_X1    g579(.A1(new_n1004), .A2(KEYINPUT117), .ZN(new_n1005));
  AOI21_X1  g580(.A(G2090), .B1(new_n1004), .B2(KEYINPUT117), .ZN(new_n1006));
  INV_X1    g581(.A(G1971), .ZN(new_n1007));
  AOI22_X1  g582(.A1(new_n1005), .A2(new_n1006), .B1(new_n1007), .B2(new_n971), .ZN(new_n1008));
  INV_X1    g583(.A(G8), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n994), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n951), .A2(new_n956), .A3(new_n935), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(G8), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1012), .ZN(new_n1013));
  AOI21_X1  g588(.A(KEYINPUT114), .B1(new_n695), .B2(G1976), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT52), .ZN(new_n1016));
  INV_X1    g591(.A(G1976), .ZN(new_n1017));
  NAND2_X1  g592(.A1(G288), .A2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1016), .B1(new_n1012), .B2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1015), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT115), .ZN(new_n1021));
  OR2_X1    g596(.A1(G305), .A2(G1981), .ZN(new_n1022));
  NAND2_X1  g597(.A1(G305), .A2(G1981), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT49), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1022), .A2(KEYINPUT49), .A3(new_n1023), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1021), .B1(new_n1012), .B2(new_n1028), .ZN(new_n1029));
  AND2_X1   g604(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1030), .A2(new_n1011), .A3(KEYINPUT115), .A4(G8), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n1013), .A2(new_n1016), .A3(new_n1014), .A4(new_n1018), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1020), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n971), .A2(new_n1007), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1035), .B1(new_n967), .B2(G2090), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(G8), .ZN(new_n1037));
  OAI21_X1  g612(.A(KEYINPUT113), .B1(new_n1037), .B2(new_n994), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT113), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n1036), .A2(new_n993), .A3(new_n1039), .A4(G8), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1034), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n782), .B1(new_n957), .B2(new_n960), .ZN(new_n1042));
  OAI211_X1 g617(.A(new_n965), .B(new_n766), .C1(new_n966), .C2(KEYINPUT50), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g619(.A(G8), .B1(new_n1044), .B2(G286), .ZN(new_n1045));
  AOI21_X1  g620(.A(G168), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1046));
  OAI21_X1  g621(.A(KEYINPUT51), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT51), .ZN(new_n1048));
  OAI211_X1 g623(.A(new_n1048), .B(G8), .C1(new_n1044), .C2(G286), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1047), .A2(new_n1049), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n988), .A2(new_n1010), .A3(new_n1041), .A4(new_n1050), .ZN(new_n1051));
  OAI21_X1  g626(.A(KEYINPUT119), .B1(new_n569), .B2(new_n580), .ZN(new_n1052));
  INV_X1    g627(.A(new_n568), .ZN(new_n1053));
  XNOR2_X1  g628(.A(new_n567), .B(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT118), .ZN(new_n1055));
  AOI21_X1  g630(.A(KEYINPUT57), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT119), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1054), .A2(new_n1057), .A3(new_n578), .A4(new_n579), .ZN(new_n1058));
  AND3_X1   g633(.A1(new_n1052), .A2(new_n1056), .A3(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1056), .B1(new_n1052), .B2(new_n1058), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n934), .B1(new_n966), .B2(KEYINPUT50), .ZN(new_n1062));
  AOI21_X1  g637(.A(G1956), .B1(new_n1062), .B2(new_n1003), .ZN(new_n1063));
  XNOR2_X1  g638(.A(KEYINPUT120), .B(KEYINPUT56), .ZN(new_n1064));
  XNOR2_X1  g639(.A(new_n1064), .B(G2072), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n969), .A2(new_n970), .A3(new_n935), .A4(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1066), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1061), .B1(new_n1063), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(G1956), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1004), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1061), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1070), .A2(new_n1066), .A3(new_n1071), .ZN(new_n1072));
  AND3_X1   g647(.A1(new_n1068), .A2(new_n1072), .A3(KEYINPUT61), .ZN(new_n1073));
  AOI21_X1  g648(.A(KEYINPUT61), .B1(new_n1068), .B2(new_n1072), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT123), .ZN(new_n1076));
  XOR2_X1   g651(.A(KEYINPUT58), .B(G1341), .Z(new_n1077));
  NAND2_X1  g652(.A1(new_n1011), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(G1996), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n969), .A2(new_n970), .A3(new_n935), .A4(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1078), .A2(KEYINPUT121), .A3(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(KEYINPUT121), .B1(new_n1078), .B2(new_n1080), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n559), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT122), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  OAI211_X1 g661(.A(KEYINPUT122), .B(new_n559), .C1(new_n1082), .C2(new_n1083), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1086), .A2(KEYINPUT59), .A3(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT59), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1084), .A2(new_n1085), .A3(new_n1089), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1075), .A2(new_n1076), .A3(new_n1088), .A4(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT61), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1071), .B1(new_n1070), .B2(new_n1066), .ZN(new_n1093));
  AOI211_X1 g668(.A(new_n1067), .B(new_n1061), .C1(new_n1004), .C2(new_n1069), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1092), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1068), .A2(new_n1072), .A3(KEYINPUT61), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1095), .A2(new_n1090), .A3(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1087), .A2(KEYINPUT59), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1078), .A2(new_n1080), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT121), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(new_n1081), .ZN(new_n1102));
  AOI21_X1  g677(.A(KEYINPUT122), .B1(new_n1102), .B2(new_n559), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1098), .A2(new_n1103), .ZN(new_n1104));
  OAI21_X1  g679(.A(KEYINPUT123), .B1(new_n1097), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(G1348), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n967), .A2(new_n1106), .ZN(new_n1107));
  OR2_X1    g682(.A1(new_n1011), .A2(G2067), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1107), .A2(KEYINPUT60), .A3(new_n1108), .ZN(new_n1109));
  AND3_X1   g684(.A1(new_n1109), .A2(KEYINPUT124), .A3(new_n618), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n618), .B1(new_n1109), .B2(KEYINPUT124), .ZN(new_n1111));
  OAI22_X1  g686(.A1(new_n1110), .A2(new_n1111), .B1(KEYINPUT124), .B2(new_n1109), .ZN(new_n1112));
  AND2_X1   g687(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1112), .B1(KEYINPUT60), .B2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1091), .A2(new_n1105), .A3(new_n1114), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1068), .B1(new_n1113), .B2(new_n618), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(new_n1072), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1051), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1118));
  AOI211_X1 g693(.A(G1976), .B(G288), .C1(new_n1029), .C2(new_n1031), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1022), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1013), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1038), .A2(new_n1040), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1121), .B1(new_n1122), .B2(new_n1034), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT62), .ZN(new_n1124));
  AND3_X1   g699(.A1(new_n1047), .A2(new_n1124), .A3(new_n1049), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1124), .B1(new_n1047), .B2(new_n1049), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(new_n974), .ZN(new_n1128));
  AND3_X1   g703(.A1(new_n1041), .A2(new_n1010), .A3(new_n1128), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1123), .B1(new_n1127), .B2(new_n1129), .ZN(new_n1130));
  AOI211_X1 g705(.A(new_n1009), .B(G286), .C1(new_n1042), .C2(new_n1043), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1037), .A2(new_n994), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1041), .A2(KEYINPUT63), .A3(new_n1131), .A4(new_n1132), .ZN(new_n1133));
  AND3_X1   g708(.A1(new_n1041), .A2(new_n1010), .A3(new_n1131), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1133), .B1(new_n1134), .B2(KEYINPUT63), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1130), .A2(new_n1135), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n949), .B1(new_n1118), .B2(new_n1136), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n716), .A2(new_n719), .ZN(new_n1138));
  XNOR2_X1  g713(.A(new_n1138), .B(KEYINPUT126), .ZN(new_n1139));
  OAI22_X1  g714(.A1(new_n941), .A2(new_n1139), .B1(G2067), .B2(new_n747), .ZN(new_n1140));
  AND2_X1   g715(.A1(new_n1140), .A2(new_n937), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n937), .A2(new_n1079), .ZN(new_n1142));
  XNOR2_X1  g717(.A(new_n1142), .B(KEYINPUT46), .ZN(new_n1143));
  AND2_X1   g718(.A1(new_n758), .A2(new_n939), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1143), .B1(new_n936), .B2(new_n1144), .ZN(new_n1145));
  XOR2_X1   g720(.A(new_n1145), .B(KEYINPUT47), .Z(new_n1146));
  NOR2_X1   g721(.A1(new_n936), .A2(new_n944), .ZN(new_n1147));
  XOR2_X1   g722(.A(new_n1147), .B(KEYINPUT48), .Z(new_n1148));
  XNOR2_X1  g723(.A(new_n943), .B(KEYINPUT127), .ZN(new_n1149));
  AOI211_X1 g724(.A(new_n1141), .B(new_n1146), .C1(new_n1148), .C2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1137), .A2(new_n1150), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g726(.A(G227), .ZN(new_n1153));
  NAND2_X1  g727(.A1(new_n1153), .A2(G319), .ZN(new_n1154));
  NOR3_X1   g728(.A1(G229), .A2(G401), .A3(new_n1154), .ZN(new_n1155));
  NAND3_X1  g729(.A1(new_n909), .A2(new_n1155), .A3(new_n854), .ZN(G225));
  INV_X1    g730(.A(G225), .ZN(G308));
endmodule


