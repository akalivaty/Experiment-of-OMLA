//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 1 1 1 0 1 1 1 0 1 0 0 1 1 1 0 0 1 1 0 0 0 0 0 1 1 0 0 0 1 1 0 0 1 0 0 1 0 1 0 1 0 0 1 0 0 0 0 0 1 0 1 0 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:55 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n450, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n555, new_n556, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n580, new_n581,
    new_n584, new_n585, new_n586, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n626, new_n627, new_n630, new_n632, new_n633,
    new_n634, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1228, new_n1229, new_n1230;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT65), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT66), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  XOR2_X1   g014(.A(KEYINPUT67), .B(G69), .Z(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT68), .Z(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G221), .A3(G219), .A4(G218), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  NOR4_X1   g029(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n460));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(G2105), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G137), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT70), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n466), .B1(new_n461), .B2(G2105), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n468), .A2(KEYINPUT70), .A3(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G101), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n465), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n462), .A2(new_n463), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n474), .B1(new_n475), .B2(G125), .ZN(new_n476));
  OAI21_X1  g051(.A(KEYINPUT69), .B1(new_n476), .B2(new_n468), .ZN(new_n477));
  AND2_X1   g052(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n478));
  NOR2_X1   g053(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n479));
  OAI21_X1  g054(.A(G125), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n468), .B1(new_n480), .B2(new_n473), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT69), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n472), .B1(new_n477), .B2(new_n483), .ZN(G160));
  NAND2_X1  g059(.A1(new_n464), .A2(G136), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n468), .B1(new_n462), .B2(new_n463), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G124), .ZN(new_n487));
  OR2_X1    g062(.A1(G100), .A2(G2105), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n488), .B(G2104), .C1(G112), .C2(new_n468), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n485), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  OAI21_X1  g066(.A(G2104), .B1(new_n468), .B2(G114), .ZN(new_n492));
  NOR2_X1   g067(.A1(G102), .A2(G2105), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(G126), .A2(G2105), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n495), .B1(new_n462), .B2(new_n463), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n464), .A2(KEYINPUT4), .A3(G138), .ZN(new_n498));
  OAI211_X1 g073(.A(G138), .B(new_n468), .C1(new_n478), .C2(new_n479), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n497), .A2(new_n498), .A3(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(G164));
  INV_X1    g078(.A(G651), .ZN(new_n504));
  NAND2_X1  g079(.A1(KEYINPUT71), .A2(KEYINPUT5), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G543), .ZN(new_n506));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n507), .A2(KEYINPUT71), .A3(KEYINPUT5), .ZN(new_n508));
  AND2_X1   g083(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G62), .ZN(new_n510));
  NAND2_X1  g085(.A1(G75), .A2(G543), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n504), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n504), .A2(KEYINPUT6), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT6), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G651), .ZN(new_n515));
  AND2_X1   g090(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G543), .ZN(new_n517));
  INV_X1    g092(.A(G50), .ZN(new_n518));
  NAND4_X1  g093(.A1(new_n506), .A2(new_n508), .A3(new_n513), .A4(new_n515), .ZN(new_n519));
  INV_X1    g094(.A(G88), .ZN(new_n520));
  OAI22_X1  g095(.A1(new_n517), .A2(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n512), .A2(new_n521), .ZN(G166));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  XNOR2_X1  g098(.A(new_n523), .B(KEYINPUT7), .ZN(new_n524));
  NAND4_X1  g099(.A1(new_n513), .A2(new_n515), .A3(G51), .A4(G543), .ZN(new_n525));
  INV_X1    g100(.A(G89), .ZN(new_n526));
  OAI211_X1 g101(.A(new_n524), .B(new_n525), .C1(new_n519), .C2(new_n526), .ZN(new_n527));
  AND2_X1   g102(.A1(G63), .A2(G651), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n506), .A2(new_n508), .A3(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT72), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n509), .A2(KEYINPUT72), .A3(new_n528), .ZN(new_n532));
  AOI21_X1  g107(.A(new_n527), .B1(new_n531), .B2(new_n532), .ZN(G168));
  INV_X1    g108(.A(G52), .ZN(new_n534));
  INV_X1    g109(.A(G90), .ZN(new_n535));
  OAI22_X1  g110(.A1(new_n517), .A2(new_n534), .B1(new_n519), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n506), .A2(new_n508), .A3(G64), .ZN(new_n537));
  NAND2_X1  g112(.A1(G77), .A2(G543), .ZN(new_n538));
  AOI21_X1  g113(.A(new_n504), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n536), .A2(new_n539), .ZN(G171));
  NAND2_X1  g115(.A1(G68), .A2(G543), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n506), .A2(new_n508), .ZN(new_n542));
  INV_X1    g117(.A(G56), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT73), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n504), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n546), .B1(new_n545), .B2(new_n544), .ZN(new_n547));
  AND2_X1   g122(.A1(new_n516), .A2(G543), .ZN(new_n548));
  AND4_X1   g123(.A1(new_n506), .A2(new_n508), .A3(new_n513), .A4(new_n515), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n548), .A2(G43), .B1(G81), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n547), .A2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  NAND4_X1  g128(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND4_X1  g131(.A1(G319), .A2(G483), .A3(G661), .A4(new_n556), .ZN(G188));
  INV_X1    g132(.A(KEYINPUT74), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n549), .A2(new_n558), .A3(G91), .ZN(new_n559));
  INV_X1    g134(.A(G91), .ZN(new_n560));
  OAI21_X1  g135(.A(KEYINPUT74), .B1(new_n519), .B2(new_n560), .ZN(new_n561));
  NAND4_X1  g136(.A1(new_n513), .A2(new_n515), .A3(G53), .A4(G543), .ZN(new_n562));
  OR2_X1    g137(.A1(new_n562), .A2(KEYINPUT9), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n562), .A2(KEYINPUT9), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n559), .A2(new_n561), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  AND3_X1   g140(.A1(new_n506), .A2(new_n508), .A3(KEYINPUT76), .ZN(new_n566));
  AOI21_X1  g141(.A(KEYINPUT76), .B1(new_n506), .B2(new_n508), .ZN(new_n567));
  INV_X1    g142(.A(G65), .ZN(new_n568));
  NOR3_X1   g143(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(G78), .A2(G543), .ZN(new_n570));
  XOR2_X1   g145(.A(new_n570), .B(KEYINPUT75), .Z(new_n571));
  OAI21_X1  g146(.A(G651), .B1(new_n569), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n565), .A2(new_n572), .ZN(G299));
  AOI22_X1  g148(.A1(new_n548), .A2(G52), .B1(G90), .B2(new_n549), .ZN(new_n574));
  INV_X1    g149(.A(new_n539), .ZN(new_n575));
  AOI21_X1  g150(.A(KEYINPUT77), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT77), .ZN(new_n577));
  NOR3_X1   g152(.A1(new_n536), .A2(new_n577), .A3(new_n539), .ZN(new_n578));
  NOR2_X1   g153(.A1(new_n576), .A2(new_n578), .ZN(G301));
  NAND2_X1  g154(.A1(new_n532), .A2(new_n531), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n549), .A2(G89), .ZN(new_n581));
  NAND4_X1  g156(.A1(new_n580), .A2(new_n581), .A3(new_n524), .A4(new_n525), .ZN(G286));
  INV_X1    g157(.A(G166), .ZN(G303));
  NAND2_X1  g158(.A1(new_n548), .A2(G49), .ZN(new_n584));
  OAI21_X1  g159(.A(G651), .B1(new_n509), .B2(G74), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n549), .A2(G87), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(G288));
  NAND2_X1  g162(.A1(G73), .A2(G543), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT78), .ZN(new_n589));
  XNOR2_X1  g164(.A(new_n588), .B(new_n589), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n506), .A2(new_n508), .A3(G61), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n504), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND4_X1  g167(.A1(new_n513), .A2(new_n515), .A3(G48), .A4(G543), .ZN(new_n593));
  INV_X1    g168(.A(G86), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n519), .B2(new_n594), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(G305));
  NAND2_X1  g172(.A1(new_n509), .A2(G60), .ZN(new_n598));
  NAND2_X1  g173(.A1(G72), .A2(G543), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n504), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(G47), .ZN(new_n601));
  INV_X1    g176(.A(G85), .ZN(new_n602));
  OAI22_X1  g177(.A1(new_n517), .A2(new_n601), .B1(new_n519), .B2(new_n602), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  OR2_X1    g179(.A1(new_n604), .A2(KEYINPUT79), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n604), .A2(KEYINPUT79), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(new_n606), .ZN(G290));
  INV_X1    g182(.A(G868), .ZN(new_n608));
  NOR2_X1   g183(.A1(G301), .A2(new_n608), .ZN(new_n609));
  NOR2_X1   g184(.A1(new_n566), .A2(new_n567), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n610), .A2(G66), .ZN(new_n611));
  NAND2_X1  g186(.A1(G79), .A2(G543), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n504), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  XOR2_X1   g188(.A(KEYINPUT80), .B(KEYINPUT10), .Z(new_n614));
  INV_X1    g189(.A(new_n614), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n549), .A2(new_n615), .A3(G92), .ZN(new_n616));
  INV_X1    g191(.A(G92), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n614), .B1(new_n519), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n548), .A2(G54), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NOR2_X1   g196(.A1(new_n613), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT81), .ZN(new_n623));
  AOI21_X1  g198(.A(new_n609), .B1(new_n623), .B2(new_n608), .ZN(G284));
  AOI21_X1  g199(.A(new_n609), .B1(new_n623), .B2(new_n608), .ZN(G321));
  NAND2_X1  g200(.A1(G286), .A2(G868), .ZN(new_n626));
  INV_X1    g201(.A(G299), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n626), .B1(new_n627), .B2(G868), .ZN(G297));
  OAI21_X1  g203(.A(new_n626), .B1(new_n627), .B2(G868), .ZN(G280));
  INV_X1    g204(.A(G559), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n623), .B1(new_n630), .B2(G860), .ZN(G148));
  AOI21_X1  g206(.A(new_n608), .B1(new_n623), .B2(new_n630), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n632), .A2(KEYINPUT82), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n632), .A2(KEYINPUT82), .ZN(new_n634));
  OAI211_X1 g209(.A(new_n633), .B(new_n634), .C1(G868), .C2(new_n552), .ZN(G323));
  XNOR2_X1  g210(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g211(.A1(new_n470), .A2(new_n475), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(KEYINPUT12), .Z(new_n638));
  XOR2_X1   g213(.A(new_n638), .B(KEYINPUT13), .Z(new_n639));
  INV_X1    g214(.A(G2100), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n639), .A2(new_n640), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n464), .A2(G135), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n486), .A2(G123), .ZN(new_n644));
  NOR2_X1   g219(.A1(G99), .A2(G2105), .ZN(new_n645));
  OAI21_X1  g220(.A(G2104), .B1(new_n468), .B2(G111), .ZN(new_n646));
  OAI211_X1 g221(.A(new_n643), .B(new_n644), .C1(new_n645), .C2(new_n646), .ZN(new_n647));
  INV_X1    g222(.A(G2096), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n641), .A2(new_n642), .A3(new_n649), .ZN(G156));
  XNOR2_X1  g225(.A(G2427), .B(G2438), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2430), .ZN(new_n652));
  XNOR2_X1  g227(.A(KEYINPUT15), .B(G2435), .ZN(new_n653));
  OR2_X1    g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n652), .A2(new_n653), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n654), .A2(KEYINPUT14), .A3(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT85), .ZN(new_n657));
  XOR2_X1   g232(.A(G1341), .B(G1348), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n660));
  XOR2_X1   g235(.A(new_n659), .B(new_n660), .Z(new_n661));
  XNOR2_X1  g236(.A(G2451), .B(G2454), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT84), .ZN(new_n663));
  XOR2_X1   g238(.A(G2443), .B(G2446), .Z(new_n664));
  XOR2_X1   g239(.A(new_n663), .B(new_n664), .Z(new_n665));
  NAND2_X1  g240(.A1(new_n661), .A2(new_n665), .ZN(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n661), .A2(new_n665), .ZN(new_n668));
  INV_X1    g243(.A(G14), .ZN(new_n669));
  NOR3_X1   g244(.A1(new_n667), .A2(new_n668), .A3(new_n669), .ZN(G401));
  XNOR2_X1  g245(.A(G2072), .B(G2078), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT17), .ZN(new_n672));
  XOR2_X1   g247(.A(G2084), .B(G2090), .Z(new_n673));
  XNOR2_X1  g248(.A(G2067), .B(G2678), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n672), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n673), .A2(new_n674), .ZN(new_n676));
  OR3_X1    g251(.A1(new_n673), .A2(new_n671), .A3(new_n674), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n675), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n673), .A2(new_n671), .A3(new_n674), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n679), .B(KEYINPUT18), .Z(new_n680));
  NAND2_X1  g255(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(new_n648), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(G2100), .ZN(G227));
  XNOR2_X1  g258(.A(G1971), .B(G1976), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT19), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  XOR2_X1   g261(.A(G1956), .B(G2474), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT86), .ZN(new_n688));
  XOR2_X1   g263(.A(G1961), .B(G1966), .Z(new_n689));
  NAND3_X1  g264(.A1(new_n686), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT87), .B(KEYINPUT20), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n688), .A2(new_n689), .ZN(new_n692));
  AOI22_X1  g267(.A1(new_n690), .A2(new_n691), .B1(new_n692), .B2(new_n686), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n688), .A2(new_n689), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n694), .A2(new_n685), .ZN(new_n695));
  OAI221_X1 g270(.A(new_n693), .B1(new_n690), .B2(new_n691), .C1(new_n692), .C2(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(G1986), .ZN(new_n697));
  XOR2_X1   g272(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n698));
  NOR2_X1   g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(G1986), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n696), .B(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(new_n698), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n699), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(G1991), .B(G1996), .ZN(new_n705));
  INV_X1    g280(.A(G1981), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n704), .B(new_n708), .ZN(G229));
  AND2_X1   g284(.A1(new_n605), .A2(new_n606), .ZN(new_n710));
  INV_X1    g285(.A(G16), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n711), .A2(KEYINPUT89), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n711), .A2(KEYINPUT89), .ZN(new_n713));
  AND2_X1   g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n710), .A2(new_n714), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n715), .B1(G24), .B2(new_n714), .ZN(new_n716));
  AND2_X1   g291(.A1(new_n716), .A2(new_n700), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n716), .A2(new_n700), .ZN(new_n718));
  OR2_X1    g293(.A1(G95), .A2(G2105), .ZN(new_n719));
  OAI211_X1 g294(.A(new_n719), .B(G2104), .C1(G107), .C2(new_n468), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n720), .B(KEYINPUT88), .Z(new_n721));
  AOI22_X1  g296(.A1(G119), .A2(new_n486), .B1(new_n464), .B2(G131), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  MUX2_X1   g298(.A(G25), .B(new_n723), .S(G29), .Z(new_n724));
  XOR2_X1   g299(.A(KEYINPUT35), .B(G1991), .Z(new_n725));
  XOR2_X1   g300(.A(new_n724), .B(new_n725), .Z(new_n726));
  NOR3_X1   g301(.A1(new_n717), .A2(new_n718), .A3(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(new_n714), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n728), .A2(G22), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(G166), .B2(new_n728), .ZN(new_n730));
  INV_X1    g305(.A(G1971), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  NOR2_X1   g307(.A1(G16), .A2(G23), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT90), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(G288), .B2(new_n711), .ZN(new_n735));
  XOR2_X1   g310(.A(KEYINPUT33), .B(G1976), .Z(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  NOR2_X1   g312(.A1(G6), .A2(G16), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(new_n596), .B2(G16), .ZN(new_n739));
  XOR2_X1   g314(.A(KEYINPUT32), .B(G1981), .Z(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n732), .A2(new_n737), .A3(new_n741), .ZN(new_n742));
  OR2_X1    g317(.A1(new_n742), .A2(KEYINPUT34), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n742), .A2(KEYINPUT34), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n727), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT36), .ZN(new_n746));
  AOI22_X1  g321(.A1(G129), .A2(new_n486), .B1(new_n470), .B2(G105), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n464), .A2(G141), .ZN(new_n748));
  NAND3_X1  g323(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT26), .Z(new_n750));
  NAND3_X1  g325(.A1(new_n747), .A2(new_n748), .A3(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(KEYINPUT94), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  MUX2_X1   g328(.A(G32), .B(new_n753), .S(G29), .Z(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT27), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(G1996), .ZN(new_n756));
  XNOR2_X1  g331(.A(KEYINPUT91), .B(G1348), .ZN(new_n757));
  NOR2_X1   g332(.A1(G4), .A2(G16), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(new_n623), .B2(G16), .ZN(new_n759));
  INV_X1    g334(.A(new_n759), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n756), .B1(new_n757), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n714), .A2(G20), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(KEYINPUT97), .Z(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT23), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(G16), .B2(G299), .ZN(new_n765));
  INV_X1    g340(.A(G1956), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n728), .A2(G19), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(new_n552), .B2(new_n728), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(G1341), .ZN(new_n770));
  NOR2_X1   g345(.A1(new_n767), .A2(new_n770), .ZN(new_n771));
  XOR2_X1   g346(.A(KEYINPUT31), .B(G11), .Z(new_n772));
  INV_X1    g347(.A(G28), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n773), .A2(KEYINPUT30), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT95), .ZN(new_n775));
  AOI21_X1  g350(.A(G29), .B1(new_n773), .B2(KEYINPUT30), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n772), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  INV_X1    g352(.A(G29), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n777), .B1(new_n647), .B2(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n778), .A2(G33), .ZN(new_n780));
  NAND3_X1  g355(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n781));
  XOR2_X1   g356(.A(new_n781), .B(KEYINPUT25), .Z(new_n782));
  NAND2_X1  g357(.A1(new_n464), .A2(G139), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  AOI22_X1  g359(.A1(new_n475), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n785), .A2(new_n468), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n780), .B1(new_n787), .B2(new_n778), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n779), .B1(new_n788), .B2(G2072), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(G2072), .B2(new_n788), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n711), .A2(G21), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(G168), .B2(new_n711), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(G1966), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n711), .A2(G5), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(G171), .B2(new_n711), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(G1961), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n778), .A2(G27), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(G164), .B2(new_n778), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(G2078), .ZN(new_n799));
  NOR4_X1   g374(.A1(new_n790), .A2(new_n793), .A3(new_n796), .A4(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n778), .A2(G26), .ZN(new_n801));
  XOR2_X1   g376(.A(new_n801), .B(KEYINPUT93), .Z(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT28), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n486), .A2(G128), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT92), .ZN(new_n805));
  OR2_X1    g380(.A1(G104), .A2(G2105), .ZN(new_n806));
  INV_X1    g381(.A(G116), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n461), .B1(new_n807), .B2(G2105), .ZN(new_n808));
  AOI22_X1  g383(.A1(new_n464), .A2(G140), .B1(new_n806), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n805), .A2(new_n809), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n803), .B1(new_n810), .B2(G29), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(G2067), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT24), .ZN(new_n813));
  INV_X1    g388(.A(G34), .ZN(new_n814));
  AOI21_X1  g389(.A(G29), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(new_n813), .B2(new_n814), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(G160), .B2(new_n778), .ZN(new_n817));
  INV_X1    g392(.A(G2084), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  NAND4_X1  g394(.A1(new_n771), .A2(new_n800), .A3(new_n812), .A4(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n778), .A2(G35), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(G162), .B2(new_n778), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT96), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT29), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(G2090), .ZN(new_n825));
  INV_X1    g400(.A(new_n757), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n825), .B1(new_n826), .B2(new_n759), .ZN(new_n827));
  NOR3_X1   g402(.A1(new_n761), .A2(new_n820), .A3(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n746), .A2(new_n828), .ZN(G150));
  INV_X1    g404(.A(G150), .ZN(G311));
  NAND2_X1  g405(.A1(new_n509), .A2(G67), .ZN(new_n831));
  NAND2_X1  g406(.A1(G80), .A2(G543), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n504), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(G55), .ZN(new_n834));
  INV_X1    g409(.A(G93), .ZN(new_n835));
  OAI22_X1  g410(.A1(new_n517), .A2(new_n834), .B1(new_n519), .B2(new_n835), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n833), .A2(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(G860), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT37), .ZN(new_n840));
  INV_X1    g415(.A(new_n837), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n551), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n547), .A2(new_n837), .A3(new_n550), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT38), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n623), .A2(G559), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n845), .B(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(KEYINPUT39), .ZN(new_n849));
  XOR2_X1   g424(.A(new_n849), .B(KEYINPUT98), .Z(new_n850));
  OAI21_X1  g425(.A(new_n838), .B1(new_n848), .B2(KEYINPUT39), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n840), .B1(new_n850), .B2(new_n851), .ZN(G145));
  XNOR2_X1  g427(.A(G160), .B(new_n490), .ZN(new_n853));
  XOR2_X1   g428(.A(new_n853), .B(new_n647), .Z(new_n854));
  INV_X1    g429(.A(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n723), .B(new_n638), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n464), .A2(G142), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n486), .A2(G130), .ZN(new_n858));
  NOR2_X1   g433(.A1(G106), .A2(G2105), .ZN(new_n859));
  OAI21_X1  g434(.A(G2104), .B1(new_n468), .B2(G118), .ZN(new_n860));
  OAI211_X1 g435(.A(new_n857), .B(new_n858), .C1(new_n859), .C2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n856), .B(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT101), .ZN(new_n863));
  INV_X1    g438(.A(new_n787), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT99), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n865), .B1(new_n494), .B2(new_n496), .ZN(new_n866));
  INV_X1    g441(.A(G114), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n867), .A2(G2105), .ZN(new_n868));
  OAI211_X1 g443(.A(new_n868), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n869));
  INV_X1    g444(.A(new_n495), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n870), .B1(new_n478), .B2(new_n479), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n869), .A2(new_n871), .A3(KEYINPUT99), .ZN(new_n872));
  NAND4_X1  g447(.A1(new_n866), .A2(new_n501), .A3(new_n498), .A4(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  OR2_X1    g449(.A1(new_n753), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n753), .A2(new_n874), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  XOR2_X1   g452(.A(new_n810), .B(KEYINPUT100), .Z(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n878), .A2(new_n875), .A3(new_n876), .ZN(new_n881));
  AOI211_X1 g456(.A(new_n863), .B(new_n864), .C1(new_n880), .C2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n864), .A2(new_n863), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n880), .A2(new_n884), .A3(new_n881), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n864), .A2(new_n863), .ZN(new_n886));
  OR2_X1    g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n862), .B1(new_n883), .B2(new_n887), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n885), .A2(new_n886), .ZN(new_n889));
  INV_X1    g464(.A(new_n862), .ZN(new_n890));
  NOR3_X1   g465(.A1(new_n889), .A2(new_n882), .A3(new_n890), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n855), .B1(new_n888), .B2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(G37), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n883), .A2(new_n887), .A3(new_n862), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n890), .B1(new_n889), .B2(new_n882), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n894), .A2(new_n854), .A3(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n892), .A2(new_n893), .A3(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n897), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g473(.A1(new_n710), .A2(G305), .ZN(new_n899));
  XNOR2_X1  g474(.A(G166), .B(G288), .ZN(new_n900));
  NOR2_X1   g475(.A1(G290), .A2(new_n596), .ZN(new_n901));
  OR3_X1    g476(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n900), .B1(new_n899), .B2(new_n901), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  XOR2_X1   g479(.A(new_n904), .B(KEYINPUT42), .Z(new_n905));
  NAND2_X1  g480(.A1(new_n623), .A2(new_n630), .ZN(new_n906));
  INV_X1    g481(.A(new_n844), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n906), .B(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(new_n622), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT102), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n909), .A2(new_n627), .A3(new_n910), .ZN(new_n911));
  OAI21_X1  g486(.A(KEYINPUT102), .B1(new_n622), .B2(G299), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n622), .A2(G299), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT41), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n909), .A2(new_n627), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n915), .B1(new_n622), .B2(G299), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n916), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n908), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n917), .A2(new_n913), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n921), .B1(new_n923), .B2(new_n908), .ZN(new_n924));
  AND2_X1   g499(.A1(new_n905), .A2(new_n924), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n905), .A2(new_n924), .ZN(new_n926));
  OAI21_X1  g501(.A(G868), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n927), .B1(G868), .B2(new_n837), .ZN(G295));
  OAI21_X1  g503(.A(new_n927), .B1(G868), .B2(new_n837), .ZN(G331));
  INV_X1    g504(.A(KEYINPUT43), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT103), .ZN(new_n931));
  OAI21_X1  g506(.A(G168), .B1(new_n576), .B2(new_n578), .ZN(new_n932));
  OAI21_X1  g507(.A(G286), .B1(new_n539), .B2(new_n536), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n931), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n548), .A2(G52), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n549), .A2(G90), .ZN(new_n936));
  NAND4_X1  g511(.A1(new_n935), .A2(new_n575), .A3(KEYINPUT77), .A4(new_n936), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n577), .B1(new_n536), .B2(new_n539), .ZN(new_n938));
  AOI21_X1  g513(.A(G286), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NOR2_X1   g514(.A1(G168), .A2(G171), .ZN(new_n940));
  NOR3_X1   g515(.A1(new_n939), .A2(new_n940), .A3(KEYINPUT103), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n907), .B1(new_n934), .B2(new_n941), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n932), .A2(new_n931), .A3(new_n933), .ZN(new_n943));
  OAI21_X1  g518(.A(KEYINPUT103), .B1(new_n939), .B2(new_n940), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n943), .A2(new_n944), .A3(new_n844), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n942), .A2(KEYINPUT104), .A3(new_n945), .ZN(new_n946));
  OR2_X1    g521(.A1(new_n945), .A2(KEYINPUT104), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n920), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n942), .A2(new_n922), .A3(new_n945), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n948), .A2(new_n904), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(new_n893), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n946), .A2(new_n947), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(new_n922), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n911), .A2(new_n912), .A3(new_n918), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n954), .B1(new_n923), .B2(KEYINPUT41), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n942), .A2(new_n945), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n904), .B1(new_n953), .B2(new_n957), .ZN(new_n958));
  OAI21_X1  g533(.A(KEYINPUT105), .B1(new_n951), .B2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(new_n904), .ZN(new_n960));
  INV_X1    g535(.A(new_n957), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n923), .B1(new_n946), .B2(new_n947), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n960), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT105), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n963), .A2(new_n964), .A3(new_n950), .A4(new_n893), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n930), .B1(new_n959), .B2(new_n965), .ZN(new_n966));
  AND2_X1   g541(.A1(new_n950), .A2(new_n893), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n948), .A2(new_n949), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(new_n960), .ZN(new_n969));
  AOI21_X1  g544(.A(KEYINPUT43), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  OAI21_X1  g545(.A(KEYINPUT44), .B1(new_n966), .B2(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n967), .A2(new_n930), .A3(new_n963), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n951), .B1(new_n960), .B2(new_n968), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n972), .B1(new_n973), .B2(new_n930), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT44), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n971), .A2(new_n976), .ZN(G397));
  INV_X1    g552(.A(G1384), .ZN(new_n978));
  AOI21_X1  g553(.A(KEYINPUT45), .B1(new_n873), .B2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(new_n979), .ZN(new_n980));
  AOI22_X1  g555(.A1(G137), .A2(new_n464), .B1(new_n470), .B2(G101), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n480), .A2(new_n473), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n482), .B1(new_n982), .B2(G2105), .ZN(new_n983));
  AOI211_X1 g558(.A(KEYINPUT69), .B(new_n468), .C1(new_n480), .C2(new_n473), .ZN(new_n984));
  OAI211_X1 g559(.A(G40), .B(new_n981), .C1(new_n983), .C2(new_n984), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n980), .A2(new_n985), .ZN(new_n986));
  XNOR2_X1  g561(.A(new_n753), .B(G1996), .ZN(new_n987));
  XNOR2_X1  g562(.A(new_n810), .B(G2067), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  XNOR2_X1  g564(.A(new_n723), .B(new_n725), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n710), .A2(new_n700), .ZN(new_n992));
  NAND2_X1  g567(.A1(G290), .A2(G1986), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n986), .B1(new_n991), .B2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT53), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT45), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n997), .A2(G1384), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n502), .A2(new_n998), .ZN(new_n999));
  NAND3_X1  g574(.A1(G160), .A2(G40), .A3(new_n999), .ZN(new_n1000));
  OR4_X1    g575(.A1(new_n996), .A2(new_n1000), .A3(G2078), .A4(new_n979), .ZN(new_n1001));
  INV_X1    g576(.A(new_n985), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n502), .A2(new_n978), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(new_n997), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT106), .ZN(new_n1005));
  AND3_X1   g580(.A1(new_n873), .A2(new_n1005), .A3(new_n998), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1005), .B1(new_n873), .B2(new_n998), .ZN(new_n1007));
  OAI211_X1 g582(.A(new_n1002), .B(new_n1004), .C1(new_n1006), .C2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n996), .B1(new_n1008), .B2(G2078), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n873), .A2(new_n978), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT50), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n985), .B1(KEYINPUT50), .B2(new_n1003), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(G1961), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1001), .A2(new_n1009), .A3(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(G301), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n996), .A2(G2078), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n981), .A2(G40), .A3(new_n1021), .ZN(new_n1022));
  NOR3_X1   g597(.A1(new_n979), .A2(new_n481), .A3(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1007), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n873), .A2(new_n1005), .A3(new_n998), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1023), .A2(new_n1026), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n1009), .A2(new_n1017), .A3(G301), .A4(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(KEYINPUT54), .B1(new_n1020), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(G1966), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1030), .B1(new_n1000), .B2(new_n979), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(KEYINPUT115), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1013), .A2(new_n1014), .A3(new_n818), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT115), .ZN(new_n1034));
  OAI211_X1 g609(.A(new_n1034), .B(new_n1030), .C1(new_n1000), .C2(new_n979), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n1032), .A2(new_n1033), .A3(G168), .A4(new_n1035), .ZN(new_n1036));
  AOI21_X1  g611(.A(KEYINPUT51), .B1(new_n1036), .B2(G8), .ZN(new_n1037));
  NAND2_X1  g612(.A1(KEYINPUT51), .A2(G8), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1032), .A2(new_n1033), .A3(new_n1035), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(G168), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1032), .A2(new_n1033), .A3(G286), .A4(new_n1035), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1038), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  NOR3_X1   g617(.A1(new_n1029), .A2(new_n1037), .A3(new_n1042), .ZN(new_n1043));
  OAI211_X1 g618(.A(KEYINPUT55), .B(G8), .C1(new_n512), .C2(new_n521), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT107), .ZN(new_n1045));
  XNOR2_X1  g620(.A(new_n1044), .B(new_n1045), .ZN(new_n1046));
  OAI21_X1  g621(.A(G8), .B1(new_n512), .B2(new_n521), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT108), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT55), .ZN(new_n1049));
  AND3_X1   g624(.A1(new_n1047), .A2(new_n1048), .A3(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1048), .B1(new_n1047), .B2(new_n1049), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n502), .A2(new_n1012), .A3(new_n978), .ZN(new_n1054));
  OAI211_X1 g629(.A(new_n1002), .B(new_n1054), .C1(new_n1011), .C2(new_n1012), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT114), .ZN(new_n1056));
  AOI21_X1  g631(.A(G2090), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1012), .B1(new_n873), .B2(new_n978), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1054), .ZN(new_n1059));
  NOR3_X1   g634(.A1(new_n1058), .A2(new_n1059), .A3(new_n985), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(KEYINPUT114), .ZN(new_n1061));
  AOI22_X1  g636(.A1(new_n1057), .A2(new_n1061), .B1(new_n731), .B2(new_n1008), .ZN(new_n1062));
  INV_X1    g637(.A(G8), .ZN(new_n1063));
  OAI211_X1 g638(.A(new_n1046), .B(new_n1053), .C1(new_n1062), .C2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(G1976), .ZN(new_n1065));
  NOR2_X1   g640(.A1(G288), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(KEYINPUT52), .B1(G288), .B2(new_n1065), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT110), .ZN(new_n1069));
  NAND4_X1  g644(.A1(G160), .A2(G40), .A3(new_n978), .A4(new_n873), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1069), .B1(new_n1070), .B2(G8), .ZN(new_n1071));
  OAI211_X1 g646(.A(new_n1069), .B(G8), .C1(new_n1010), .C2(new_n985), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1072), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n1067), .B(new_n1068), .C1(new_n1071), .C2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n590), .A2(new_n591), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(G651), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n549), .A2(G86), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1076), .A2(new_n706), .A3(new_n1077), .A4(new_n593), .ZN(new_n1078));
  NAND2_X1  g653(.A1(KEYINPUT111), .A2(KEYINPUT49), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1079), .ZN(new_n1080));
  OAI21_X1  g655(.A(G1981), .B1(new_n592), .B2(new_n595), .ZN(new_n1081));
  AND3_X1   g656(.A1(new_n1078), .A2(new_n1080), .A3(new_n1081), .ZN(new_n1082));
  OAI211_X1 g657(.A(new_n1078), .B(new_n1081), .C1(KEYINPUT111), .C2(KEYINPUT49), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1082), .B1(new_n1079), .B2(new_n1083), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1084), .B1(new_n1073), .B2(new_n1071), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1074), .A2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g661(.A(G8), .B1(new_n1010), .B2(new_n985), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(KEYINPUT110), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1066), .B1(new_n1088), .B2(new_n1072), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT52), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1086), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1008), .A2(new_n731), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1093), .B1(G2090), .B2(new_n1015), .ZN(new_n1094));
  XNOR2_X1  g669(.A(new_n1044), .B(KEYINPUT107), .ZN(new_n1095));
  OAI21_X1  g670(.A(KEYINPUT109), .B1(new_n1052), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT109), .ZN(new_n1097));
  OAI211_X1 g672(.A(new_n1046), .B(new_n1097), .C1(new_n1051), .C2(new_n1050), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1094), .A2(new_n1096), .A3(new_n1098), .A4(G8), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1064), .A2(new_n1092), .A3(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1009), .A2(new_n1017), .A3(new_n1027), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(G171), .ZN(new_n1103));
  OAI211_X1 g678(.A(new_n1103), .B(KEYINPUT54), .C1(new_n1019), .C2(new_n1018), .ZN(new_n1104));
  AND2_X1   g679(.A1(new_n1104), .A2(KEYINPUT125), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1104), .A2(KEYINPUT125), .ZN(new_n1106));
  OAI211_X1 g681(.A(new_n1043), .B(new_n1101), .C1(new_n1105), .C2(new_n1106), .ZN(new_n1107));
  XNOR2_X1  g682(.A(KEYINPUT121), .B(KEYINPUT61), .ZN(new_n1108));
  XNOR2_X1  g683(.A(KEYINPUT56), .B(G2072), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1109), .ZN(new_n1110));
  OAI22_X1  g685(.A1(new_n1008), .A2(new_n1110), .B1(new_n1060), .B2(G1956), .ZN(new_n1111));
  AOI21_X1  g686(.A(KEYINPUT57), .B1(G299), .B2(KEYINPUT117), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT117), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT57), .ZN(new_n1114));
  AOI211_X1 g689(.A(new_n1113), .B(new_n1114), .C1(new_n565), .C2(new_n572), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1112), .A2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1116), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1111), .A2(new_n1117), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1026), .A2(new_n1002), .A3(new_n1004), .A4(new_n1109), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1055), .A2(new_n766), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1116), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1108), .B1(new_n1118), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT59), .ZN(new_n1123));
  XOR2_X1   g698(.A(KEYINPUT119), .B(G1996), .Z(new_n1124));
  INV_X1    g699(.A(new_n1124), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n985), .A2(new_n1125), .ZN(new_n1126));
  OAI211_X1 g701(.A(new_n1126), .B(new_n1004), .C1(new_n1007), .C2(new_n1006), .ZN(new_n1127));
  XOR2_X1   g702(.A(KEYINPUT58), .B(G1341), .Z(new_n1128));
  NAND2_X1  g703(.A1(new_n1070), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT120), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1127), .A2(KEYINPUT120), .A3(new_n1129), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1123), .B1(new_n1134), .B2(new_n552), .ZN(new_n1135));
  AND3_X1   g710(.A1(new_n1127), .A2(KEYINPUT120), .A3(new_n1129), .ZN(new_n1136));
  AOI21_X1  g711(.A(KEYINPUT120), .B1(new_n1127), .B2(new_n1129), .ZN(new_n1137));
  OAI211_X1 g712(.A(new_n1123), .B(new_n552), .C1(new_n1136), .C2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1138), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1122), .B1(new_n1135), .B2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT122), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1141), .B1(new_n1111), .B2(new_n1117), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1119), .A2(new_n1116), .A3(new_n1120), .A4(KEYINPUT122), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1142), .A2(KEYINPUT61), .A3(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT118), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1111), .A2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1119), .A2(new_n1120), .A3(KEYINPUT118), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1116), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1144), .A2(new_n1148), .ZN(new_n1149));
  OAI21_X1  g724(.A(KEYINPUT123), .B1(new_n1140), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1151), .A2(new_n1117), .ZN(new_n1152));
  AND2_X1   g727(.A1(new_n1143), .A2(KEYINPUT61), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1152), .A2(new_n1142), .A3(new_n1153), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n552), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1155), .A2(KEYINPUT59), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1156), .A2(new_n1138), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT123), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1154), .A2(new_n1157), .A3(new_n1158), .A4(new_n1122), .ZN(new_n1159));
  AND2_X1   g734(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1160));
  OAI22_X1  g735(.A1(new_n1160), .A2(G1348), .B1(G2067), .B2(new_n1070), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT60), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT124), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1163), .A2(new_n1164), .A3(new_n623), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1166));
  XNOR2_X1  g741(.A(new_n623), .B(new_n1164), .ZN(new_n1167));
  OAI211_X1 g742(.A(new_n1165), .B(new_n1166), .C1(new_n1163), .C2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1150), .A2(new_n1159), .A3(new_n1168), .ZN(new_n1169));
  AND2_X1   g744(.A1(new_n1161), .A2(new_n623), .ZN(new_n1170));
  OAI22_X1  g745(.A1(new_n1148), .A2(new_n1170), .B1(new_n1117), .B2(new_n1111), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1107), .B1(new_n1169), .B2(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(new_n1099), .ZN(new_n1173));
  NOR3_X1   g748(.A1(new_n1086), .A2(new_n1091), .A3(KEYINPUT112), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT112), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1088), .A2(new_n1072), .ZN(new_n1176));
  AOI22_X1  g751(.A1(new_n1089), .A2(new_n1068), .B1(new_n1176), .B2(new_n1084), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1067), .B1(new_n1071), .B2(new_n1073), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1178), .A2(KEYINPUT52), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1175), .B1(new_n1177), .B2(new_n1179), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1173), .B1(new_n1174), .B2(new_n1180), .ZN(new_n1181));
  XOR2_X1   g756(.A(new_n1176), .B(KEYINPUT113), .Z(new_n1182));
  AOI211_X1 g757(.A(G1976), .B(G288), .C1(new_n1176), .C2(new_n1084), .ZN(new_n1183));
  INV_X1    g758(.A(new_n1078), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n1182), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1181), .A2(new_n1185), .ZN(new_n1186));
  INV_X1    g761(.A(KEYINPUT62), .ZN(new_n1187));
  NOR3_X1   g762(.A1(new_n1042), .A2(new_n1187), .A3(new_n1037), .ZN(new_n1188));
  INV_X1    g763(.A(new_n1020), .ZN(new_n1189));
  NAND4_X1  g764(.A1(new_n1064), .A2(new_n1189), .A3(new_n1092), .A4(new_n1099), .ZN(new_n1190));
  NOR2_X1   g765(.A1(new_n1188), .A2(new_n1190), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1187), .B1(new_n1042), .B2(new_n1037), .ZN(new_n1192));
  AOI21_X1  g767(.A(new_n1186), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  INV_X1    g768(.A(KEYINPUT63), .ZN(new_n1194));
  NAND3_X1  g769(.A1(new_n1039), .A2(G8), .A3(G168), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n1194), .B1(new_n1100), .B2(new_n1195), .ZN(new_n1196));
  NOR3_X1   g771(.A1(new_n1173), .A2(new_n1194), .A3(new_n1195), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1053), .A2(new_n1046), .ZN(new_n1198));
  AOI21_X1  g773(.A(new_n1198), .B1(new_n1094), .B2(G8), .ZN(new_n1199));
  OAI21_X1  g774(.A(KEYINPUT112), .B1(new_n1086), .B2(new_n1091), .ZN(new_n1200));
  NAND3_X1  g775(.A1(new_n1177), .A2(new_n1175), .A3(new_n1179), .ZN(new_n1201));
  AOI21_X1  g776(.A(new_n1199), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  OAI21_X1  g777(.A(new_n1197), .B1(new_n1202), .B2(KEYINPUT116), .ZN(new_n1203));
  INV_X1    g778(.A(KEYINPUT116), .ZN(new_n1204));
  AOI211_X1 g779(.A(new_n1204), .B(new_n1199), .C1(new_n1200), .C2(new_n1201), .ZN(new_n1205));
  OAI21_X1  g780(.A(new_n1196), .B1(new_n1203), .B2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1193), .A2(new_n1206), .ZN(new_n1207));
  OAI21_X1  g782(.A(new_n995), .B1(new_n1172), .B2(new_n1207), .ZN(new_n1208));
  INV_X1    g783(.A(new_n986), .ZN(new_n1209));
  NAND4_X1  g784(.A1(new_n989), .A2(new_n725), .A3(new_n721), .A4(new_n722), .ZN(new_n1210));
  OR2_X1    g785(.A1(new_n810), .A2(G2067), .ZN(new_n1211));
  AOI21_X1  g786(.A(new_n1209), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g787(.A1(new_n991), .A2(new_n986), .ZN(new_n1213));
  NOR2_X1   g788(.A1(new_n992), .A2(new_n1209), .ZN(new_n1214));
  XNOR2_X1  g789(.A(KEYINPUT127), .B(KEYINPUT48), .ZN(new_n1215));
  XNOR2_X1  g790(.A(new_n1214), .B(new_n1215), .ZN(new_n1216));
  AOI21_X1  g791(.A(new_n1212), .B1(new_n1213), .B2(new_n1216), .ZN(new_n1217));
  INV_X1    g792(.A(KEYINPUT46), .ZN(new_n1218));
  OR3_X1    g793(.A1(new_n1209), .A2(new_n1218), .A3(G1996), .ZN(new_n1219));
  OAI21_X1  g794(.A(new_n986), .B1(new_n988), .B2(new_n753), .ZN(new_n1220));
  OAI21_X1  g795(.A(new_n1218), .B1(new_n1209), .B2(G1996), .ZN(new_n1221));
  NAND3_X1  g796(.A1(new_n1219), .A2(new_n1220), .A3(new_n1221), .ZN(new_n1222));
  XOR2_X1   g797(.A(new_n1222), .B(KEYINPUT47), .Z(new_n1223));
  OAI21_X1  g798(.A(new_n1217), .B1(new_n1223), .B2(KEYINPUT126), .ZN(new_n1224));
  AOI21_X1  g799(.A(new_n1224), .B1(KEYINPUT126), .B2(new_n1223), .ZN(new_n1225));
  NAND2_X1  g800(.A1(new_n1208), .A2(new_n1225), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g801(.A(G401), .ZN(new_n1228));
  INV_X1    g802(.A(G319), .ZN(new_n1229));
  NOR3_X1   g803(.A1(G229), .A2(new_n1229), .A3(G227), .ZN(new_n1230));
  AND4_X1   g804(.A1(new_n1228), .A2(new_n974), .A3(new_n1230), .A4(new_n897), .ZN(G308));
  NAND4_X1  g805(.A1(new_n974), .A2(new_n1228), .A3(new_n1230), .A4(new_n897), .ZN(G225));
endmodule


