//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 1 1 0 0 0 1 0 0 1 0 0 1 0 1 1 0 1 0 0 0 0 0 1 1 0 0 0 0 1 1 0 0 1 0 1 0 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 1 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:53 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n451, new_n452, new_n453, new_n457, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n546, new_n548, new_n549, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n564, new_n565, new_n566, new_n567,
    new_n570, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n607, new_n608, new_n609, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n826, new_n827, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1161, new_n1162, new_n1163, new_n1164;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT64), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XNOR2_X1  g012(.A(KEYINPUT65), .B(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT66), .Z(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  OR4_X1    g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  AOI22_X1  g030(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n453), .ZN(G319));
  INV_X1    g031(.A(G2104), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n457), .A2(KEYINPUT3), .ZN(new_n458));
  INV_X1    g033(.A(KEYINPUT3), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G2104), .ZN(new_n460));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  AND3_X1   g036(.A1(new_n458), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G137), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT67), .ZN(new_n464));
  NOR3_X1   g039(.A1(new_n464), .A2(new_n457), .A3(G2105), .ZN(new_n465));
  AOI21_X1  g040(.A(KEYINPUT67), .B1(new_n461), .B2(G2104), .ZN(new_n466));
  OAI21_X1  g041(.A(G101), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n463), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n458), .A2(new_n460), .A3(G125), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n461), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n468), .A2(new_n471), .ZN(G160));
  NAND2_X1  g047(.A1(new_n462), .A2(G136), .ZN(new_n473));
  NOR2_X1   g048(.A1(G100), .A2(G2105), .ZN(new_n474));
  OAI21_X1  g049(.A(G2104), .B1(new_n461), .B2(G112), .ZN(new_n475));
  AND2_X1   g050(.A1(new_n458), .A2(new_n460), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G2105), .ZN(new_n477));
  INV_X1    g052(.A(G124), .ZN(new_n478));
  OAI221_X1 g053(.A(new_n473), .B1(new_n474), .B2(new_n475), .C1(new_n477), .C2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G162));
  INV_X1    g055(.A(KEYINPUT4), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(KEYINPUT69), .ZN(new_n482));
  OR2_X1    g057(.A1(new_n481), .A2(KEYINPUT69), .ZN(new_n483));
  NAND4_X1  g058(.A1(new_n462), .A2(G138), .A3(new_n482), .A4(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(G114), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n457), .B1(new_n485), .B2(G2105), .ZN(new_n486));
  NOR2_X1   g061(.A1(G102), .A2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n486), .A2(KEYINPUT68), .A3(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT68), .ZN(new_n490));
  OAI21_X1  g065(.A(G2104), .B1(new_n461), .B2(G114), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n490), .B1(new_n491), .B2(new_n487), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n476), .A2(G126), .A3(G2105), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n458), .A2(new_n460), .A3(G138), .A4(new_n461), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n495), .A2(KEYINPUT69), .A3(new_n481), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n484), .A2(new_n493), .A3(new_n494), .A4(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(G164));
  NAND2_X1  g073(.A1(KEYINPUT70), .A2(KEYINPUT5), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(G543), .ZN(new_n500));
  INV_X1    g075(.A(G543), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n501), .A2(KEYINPUT70), .A3(KEYINPUT5), .ZN(new_n502));
  AND2_X1   g077(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  XNOR2_X1  g078(.A(KEYINPUT6), .B(G651), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  XNOR2_X1  g080(.A(KEYINPUT71), .B(G88), .ZN(new_n506));
  INV_X1    g081(.A(G50), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n504), .A2(G543), .ZN(new_n508));
  OAI22_X1  g083(.A1(new_n505), .A2(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n503), .A2(G62), .ZN(new_n511));
  NAND2_X1  g086(.A1(G75), .A2(G543), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n509), .A2(new_n513), .ZN(G166));
  NAND3_X1  g089(.A1(new_n503), .A2(G63), .A3(G651), .ZN(new_n515));
  NAND3_X1  g090(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n516));
  XNOR2_X1  g091(.A(new_n516), .B(KEYINPUT7), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n504), .A2(G51), .A3(G543), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n515), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  AND3_X1   g094(.A1(new_n503), .A2(G89), .A3(new_n504), .ZN(new_n520));
  OAI21_X1  g095(.A(KEYINPUT72), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  AND2_X1   g096(.A1(new_n517), .A2(new_n518), .ZN(new_n522));
  AND3_X1   g097(.A1(new_n504), .A2(new_n500), .A3(new_n502), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G89), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT72), .ZN(new_n525));
  NAND4_X1  g100(.A1(new_n522), .A2(new_n524), .A3(new_n525), .A4(new_n515), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n521), .A2(new_n526), .ZN(G168));
  NAND2_X1  g102(.A1(new_n523), .A2(G90), .ZN(new_n528));
  INV_X1    g103(.A(new_n508), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(G52), .ZN(new_n530));
  NAND2_X1  g105(.A1(G77), .A2(G543), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n500), .A2(new_n502), .ZN(new_n532));
  INV_X1    g107(.A(G64), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  AND3_X1   g109(.A1(new_n534), .A2(KEYINPUT73), .A3(G651), .ZN(new_n535));
  AOI21_X1  g110(.A(KEYINPUT73), .B1(new_n534), .B2(G651), .ZN(new_n536));
  OAI211_X1 g111(.A(new_n528), .B(new_n530), .C1(new_n535), .C2(new_n536), .ZN(G301));
  INV_X1    g112(.A(G301), .ZN(G171));
  NAND2_X1  g113(.A1(new_n503), .A2(G56), .ZN(new_n539));
  NAND2_X1  g114(.A1(G68), .A2(G543), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G651), .ZN(new_n542));
  AOI22_X1  g117(.A1(G81), .A2(new_n523), .B1(new_n529), .B2(G43), .ZN(new_n543));
  AND2_X1   g118(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G860), .ZN(G153));
  AND3_X1   g120(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G36), .ZN(G176));
  NAND2_X1  g122(.A1(G1), .A2(G3), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT8), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n546), .A2(new_n549), .ZN(G188));
  NAND2_X1  g125(.A1(G78), .A2(G543), .ZN(new_n551));
  INV_X1    g126(.A(G65), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n551), .B1(new_n532), .B2(new_n552), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT74), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G651), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n529), .A2(G53), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT9), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n523), .A2(G91), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n555), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT75), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND4_X1  g136(.A1(new_n555), .A2(new_n557), .A3(KEYINPUT75), .A4(new_n558), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n561), .A2(new_n562), .ZN(G299));
  AOI21_X1  g138(.A(KEYINPUT76), .B1(new_n521), .B2(new_n526), .ZN(new_n564));
  INV_X1    g139(.A(new_n564), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n521), .A2(KEYINPUT76), .A3(new_n526), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(new_n567), .ZN(G286));
  INV_X1    g143(.A(G166), .ZN(G303));
  INV_X1    g144(.A(G74), .ZN(new_n570));
  AOI21_X1  g145(.A(new_n510), .B1(new_n532), .B2(new_n570), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n571), .B1(G49), .B2(new_n529), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n523), .A2(G87), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n572), .A2(new_n573), .ZN(G288));
  NAND3_X1  g149(.A1(new_n500), .A2(new_n502), .A3(G61), .ZN(new_n575));
  NAND2_X1  g150(.A1(G73), .A2(G543), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  AOI21_X1  g152(.A(KEYINPUT77), .B1(new_n577), .B2(G651), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT77), .ZN(new_n579));
  AOI211_X1 g154(.A(new_n579), .B(new_n510), .C1(new_n575), .C2(new_n576), .ZN(new_n580));
  NAND4_X1  g155(.A1(new_n504), .A2(G86), .A3(new_n500), .A4(new_n502), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n504), .A2(G48), .A3(G543), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NOR3_X1   g158(.A1(new_n578), .A2(new_n580), .A3(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(new_n584), .ZN(G305));
  NAND2_X1  g160(.A1(G72), .A2(G543), .ZN(new_n586));
  INV_X1    g161(.A(G60), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n532), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n588), .A2(G651), .ZN(new_n589));
  INV_X1    g164(.A(G85), .ZN(new_n590));
  INV_X1    g165(.A(G47), .ZN(new_n591));
  OAI22_X1  g166(.A1(new_n505), .A2(new_n590), .B1(new_n591), .B2(new_n508), .ZN(new_n592));
  AND2_X1   g167(.A1(new_n592), .A2(KEYINPUT78), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n592), .A2(KEYINPUT78), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n589), .B1(new_n593), .B2(new_n594), .ZN(G290));
  NAND2_X1  g170(.A1(G301), .A2(G868), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n523), .A2(G92), .ZN(new_n597));
  XOR2_X1   g172(.A(new_n597), .B(KEYINPUT10), .Z(new_n598));
  NAND2_X1  g173(.A1(new_n529), .A2(G54), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n503), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n600));
  OR2_X1    g175(.A1(new_n600), .A2(new_n510), .ZN(new_n601));
  AND3_X1   g176(.A1(new_n598), .A2(new_n599), .A3(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n596), .B1(new_n602), .B2(G868), .ZN(G284));
  OAI21_X1  g178(.A(new_n596), .B1(new_n602), .B2(G868), .ZN(G321));
  MUX2_X1   g179(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g180(.A(G299), .B(G286), .S(G868), .Z(G280));
  NAND3_X1  g181(.A1(new_n598), .A2(new_n599), .A3(new_n601), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n607), .A2(G559), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n608), .B1(G860), .B2(new_n602), .ZN(new_n609));
  XOR2_X1   g184(.A(new_n609), .B(KEYINPUT79), .Z(G148));
  INV_X1    g185(.A(G868), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n613), .B1(G868), .B2(new_n544), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(KEYINPUT80), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(KEYINPUT80), .B2(new_n612), .ZN(G323));
  XNOR2_X1  g191(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OR2_X1    g192(.A1(new_n465), .A2(new_n466), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n618), .A2(new_n476), .ZN(new_n619));
  XNOR2_X1  g194(.A(KEYINPUT81), .B(KEYINPUT12), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n619), .B(new_n620), .ZN(new_n621));
  XOR2_X1   g196(.A(KEYINPUT13), .B(G2100), .Z(new_n622));
  XNOR2_X1  g197(.A(new_n621), .B(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n462), .A2(G135), .ZN(new_n624));
  NOR2_X1   g199(.A1(G99), .A2(G2105), .ZN(new_n625));
  OAI21_X1  g200(.A(G2104), .B1(new_n461), .B2(G111), .ZN(new_n626));
  INV_X1    g201(.A(G123), .ZN(new_n627));
  OAI221_X1 g202(.A(new_n624), .B1(new_n625), .B2(new_n626), .C1(new_n477), .C2(new_n627), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n628), .B(G2096), .Z(new_n629));
  NAND2_X1  g204(.A1(new_n623), .A2(new_n629), .ZN(G156));
  XNOR2_X1  g205(.A(G2451), .B(G2454), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT82), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT16), .ZN(new_n633));
  XOR2_X1   g208(.A(G2443), .B(G2446), .Z(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(G1341), .B(G1348), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(KEYINPUT15), .B(G2435), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2438), .ZN(new_n639));
  XOR2_X1   g214(.A(G2427), .B(G2430), .Z(new_n640));
  NOR2_X1   g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n639), .A2(new_n640), .ZN(new_n642));
  INV_X1    g217(.A(KEYINPUT83), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n642), .B1(new_n643), .B2(KEYINPUT14), .ZN(new_n644));
  AOI211_X1 g219(.A(new_n641), .B(new_n644), .C1(new_n643), .C2(KEYINPUT14), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n637), .B(new_n645), .ZN(new_n646));
  INV_X1    g221(.A(G14), .ZN(new_n647));
  NOR2_X1   g222(.A1(new_n646), .A2(new_n647), .ZN(G401));
  XNOR2_X1  g223(.A(G2067), .B(G2678), .ZN(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2084), .B(G2090), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n650), .A2(new_n651), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n652), .A2(new_n653), .A3(KEYINPUT17), .ZN(new_n654));
  INV_X1    g229(.A(KEYINPUT18), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n652), .A2(KEYINPUT18), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2072), .B(G2078), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n656), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  OAI21_X1  g234(.A(new_n659), .B1(new_n658), .B2(new_n656), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(G2100), .ZN(new_n661));
  XOR2_X1   g236(.A(KEYINPUT84), .B(G2096), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(G227));
  XNOR2_X1  g238(.A(G1971), .B(G1976), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT19), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(G1961), .B(G1966), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT85), .ZN(new_n668));
  XOR2_X1   g243(.A(G1956), .B(G2474), .Z(new_n669));
  NAND2_X1  g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(KEYINPUT20), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n668), .A2(new_n669), .ZN(new_n673));
  OAI21_X1  g248(.A(new_n666), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n671), .B1(new_n670), .B2(new_n665), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n673), .A2(new_n666), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n676), .A2(new_n670), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n674), .A2(new_n675), .A3(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT21), .ZN(new_n679));
  INV_X1    g254(.A(G1986), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1991), .B(G1996), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT88), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(G1981), .ZN(new_n684));
  XOR2_X1   g259(.A(KEYINPUT86), .B(KEYINPUT87), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT22), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n684), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n681), .B(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(G229));
  INV_X1    g264(.A(G29), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n690), .A2(G35), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n691), .B1(G162), .B2(new_n690), .ZN(new_n692));
  XOR2_X1   g267(.A(new_n692), .B(KEYINPUT29), .Z(new_n693));
  INV_X1    g268(.A(G2090), .ZN(new_n694));
  OR2_X1    g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT95), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n693), .A2(new_n694), .ZN(new_n697));
  INV_X1    g272(.A(G16), .ZN(new_n698));
  AND2_X1   g273(.A1(new_n698), .A2(G4), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n699), .B1(new_n607), .B2(G16), .ZN(new_n700));
  INV_X1    g275(.A(G1348), .ZN(new_n701));
  OR2_X1    g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(G164), .A2(G29), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n703), .B1(G27), .B2(G29), .ZN(new_n704));
  INV_X1    g279(.A(G2078), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n700), .A2(new_n701), .ZN(new_n707));
  NAND4_X1  g282(.A1(new_n697), .A2(new_n702), .A3(new_n706), .A4(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n690), .A2(G26), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT91), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT28), .ZN(new_n711));
  INV_X1    g286(.A(new_n477), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(G128), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n462), .A2(G140), .ZN(new_n714));
  OR2_X1    g289(.A1(G104), .A2(G2105), .ZN(new_n715));
  OAI211_X1 g290(.A(new_n715), .B(G2104), .C1(G116), .C2(new_n461), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n713), .A2(new_n714), .A3(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(new_n717), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n711), .B1(new_n718), .B2(new_n690), .ZN(new_n719));
  INV_X1    g294(.A(G2067), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(KEYINPUT24), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n690), .B1(new_n722), .B2(G34), .ZN(new_n723));
  INV_X1    g298(.A(KEYINPUT93), .ZN(new_n724));
  OR2_X1    g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n722), .A2(G34), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n723), .A2(new_n724), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n725), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(G160), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n728), .B1(new_n729), .B2(new_n690), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(G2084), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n698), .A2(G19), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(new_n544), .B2(new_n698), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n733), .A2(G1341), .ZN(new_n734));
  OR2_X1    g309(.A1(new_n733), .A2(G1341), .ZN(new_n735));
  NAND4_X1  g310(.A1(new_n721), .A2(new_n731), .A3(new_n734), .A4(new_n735), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n704), .A2(new_n705), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n712), .A2(G129), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n618), .A2(G105), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n462), .A2(G141), .ZN(new_n740));
  NAND3_X1  g315(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n741));
  XOR2_X1   g316(.A(new_n741), .B(KEYINPUT26), .Z(new_n742));
  NAND4_X1  g317(.A1(new_n738), .A2(new_n739), .A3(new_n740), .A4(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n744), .A2(G29), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(G29), .B2(G32), .ZN(new_n746));
  XNOR2_X1  g321(.A(KEYINPUT27), .B(G1996), .ZN(new_n747));
  OR2_X1    g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n746), .A2(new_n747), .ZN(new_n749));
  XNOR2_X1  g324(.A(KEYINPUT94), .B(G28), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT30), .ZN(new_n751));
  MUX2_X1   g326(.A(new_n751), .B(new_n628), .S(G29), .Z(new_n752));
  NAND3_X1  g327(.A1(new_n748), .A2(new_n749), .A3(new_n752), .ZN(new_n753));
  NOR4_X1   g328(.A1(new_n708), .A2(new_n736), .A3(new_n737), .A4(new_n753), .ZN(new_n754));
  XNOR2_X1  g329(.A(KEYINPUT31), .B(G11), .ZN(new_n755));
  NOR2_X1   g330(.A1(G16), .A2(G21), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(G168), .B2(G16), .ZN(new_n757));
  INV_X1    g332(.A(G1966), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n757), .B(new_n758), .ZN(new_n759));
  AND3_X1   g334(.A1(new_n754), .A2(new_n755), .A3(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(G299), .ZN(new_n761));
  OAI21_X1  g336(.A(KEYINPUT23), .B1(new_n761), .B2(new_n698), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n698), .A2(G20), .ZN(new_n763));
  MUX2_X1   g338(.A(KEYINPUT23), .B(new_n762), .S(new_n763), .Z(new_n764));
  NOR2_X1   g339(.A1(new_n764), .A2(G1956), .ZN(new_n765));
  INV_X1    g340(.A(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n764), .A2(G1956), .ZN(new_n767));
  NAND2_X1  g342(.A1(G171), .A2(G16), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G5), .B2(G16), .ZN(new_n769));
  INV_X1    g344(.A(G1961), .ZN(new_n770));
  AND2_X1   g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT25), .Z(new_n773));
  NAND2_X1  g348(.A1(new_n462), .A2(G139), .ZN(new_n774));
  AOI22_X1  g349(.A1(new_n476), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n775));
  OAI211_X1 g350(.A(new_n773), .B(new_n774), .C1(new_n775), .C2(new_n461), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT92), .ZN(new_n777));
  AND2_X1   g352(.A1(new_n777), .A2(G29), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(new_n690), .B2(G33), .ZN(new_n779));
  INV_X1    g354(.A(G2072), .ZN(new_n780));
  OAI22_X1  g355(.A1(new_n769), .A2(new_n770), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  AOI211_X1 g356(.A(new_n771), .B(new_n781), .C1(new_n780), .C2(new_n779), .ZN(new_n782));
  NAND4_X1  g357(.A1(new_n760), .A2(new_n766), .A3(new_n767), .A4(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n698), .A2(G23), .ZN(new_n784));
  AND2_X1   g359(.A1(new_n572), .A2(new_n573), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n784), .B1(new_n785), .B2(new_n698), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT33), .ZN(new_n787));
  INV_X1    g362(.A(G1976), .ZN(new_n788));
  OR2_X1    g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n787), .A2(new_n788), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n698), .A2(G22), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(G166), .B2(new_n698), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n792), .A2(G1971), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n789), .A2(new_n790), .A3(new_n793), .ZN(new_n794));
  XOR2_X1   g369(.A(KEYINPUT32), .B(G1981), .Z(new_n795));
  NAND2_X1  g370(.A1(new_n698), .A2(G6), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(new_n584), .B2(new_n698), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT90), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n794), .B1(new_n795), .B2(new_n798), .ZN(new_n799));
  OR2_X1    g374(.A1(new_n792), .A2(G1971), .ZN(new_n800));
  OR2_X1    g375(.A1(new_n798), .A2(new_n795), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n799), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  OR2_X1    g377(.A1(new_n802), .A2(KEYINPUT34), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n802), .A2(KEYINPUT34), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n698), .A2(G24), .ZN(new_n805));
  INV_X1    g380(.A(G290), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n805), .B1(new_n806), .B2(new_n698), .ZN(new_n807));
  INV_X1    g382(.A(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n808), .A2(new_n680), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n712), .A2(G119), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT89), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n811), .B1(G131), .B2(new_n462), .ZN(new_n812));
  OR2_X1    g387(.A1(G95), .A2(G2105), .ZN(new_n813));
  OAI211_X1 g388(.A(new_n813), .B(G2104), .C1(G107), .C2(new_n461), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  MUX2_X1   g390(.A(G25), .B(new_n815), .S(G29), .Z(new_n816));
  XOR2_X1   g391(.A(KEYINPUT35), .B(G1991), .Z(new_n817));
  XOR2_X1   g392(.A(new_n816), .B(new_n817), .Z(new_n818));
  AOI21_X1  g393(.A(new_n818), .B1(G1986), .B2(new_n807), .ZN(new_n819));
  NAND4_X1  g394(.A1(new_n803), .A2(new_n804), .A3(new_n809), .A4(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n820), .A2(KEYINPUT36), .ZN(new_n821));
  AND2_X1   g396(.A1(new_n804), .A2(new_n819), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT36), .ZN(new_n823));
  NAND4_X1  g398(.A1(new_n822), .A2(new_n823), .A3(new_n803), .A4(new_n809), .ZN(new_n824));
  AOI211_X1 g399(.A(new_n696), .B(new_n783), .C1(new_n821), .C2(new_n824), .ZN(G311));
  AOI21_X1  g400(.A(new_n783), .B1(new_n821), .B2(new_n824), .ZN(new_n826));
  INV_X1    g401(.A(new_n696), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n826), .A2(new_n827), .ZN(G150));
  INV_X1    g403(.A(G93), .ZN(new_n829));
  INV_X1    g404(.A(G55), .ZN(new_n830));
  OAI22_X1  g405(.A1(new_n505), .A2(new_n829), .B1(new_n830), .B2(new_n508), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n503), .A2(G67), .ZN(new_n832));
  NAND2_X1  g407(.A1(G80), .A2(G543), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n510), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  OAI21_X1  g409(.A(G860), .B1(new_n831), .B2(new_n834), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n835), .B(KEYINPUT37), .Z(new_n836));
  NAND2_X1  g411(.A1(new_n602), .A2(G559), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT39), .ZN(new_n838));
  XNOR2_X1  g413(.A(KEYINPUT96), .B(KEYINPUT38), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n838), .B(new_n839), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n831), .A2(new_n834), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n544), .B(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n840), .B(new_n842), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n836), .B1(new_n843), .B2(G860), .ZN(G145));
  XNOR2_X1  g419(.A(G160), .B(new_n628), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(G162), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n777), .B(new_n743), .ZN(new_n847));
  XNOR2_X1  g422(.A(G164), .B(new_n717), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n847), .B(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n462), .A2(G142), .ZN(new_n850));
  NOR2_X1   g425(.A1(G106), .A2(G2105), .ZN(new_n851));
  OAI21_X1  g426(.A(G2104), .B1(new_n461), .B2(G118), .ZN(new_n852));
  INV_X1    g427(.A(G130), .ZN(new_n853));
  OAI221_X1 g428(.A(new_n850), .B1(new_n851), .B2(new_n852), .C1(new_n477), .C2(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n621), .B(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n815), .B(new_n855), .ZN(new_n856));
  OR2_X1    g431(.A1(new_n849), .A2(new_n856), .ZN(new_n857));
  XOR2_X1   g432(.A(new_n857), .B(KEYINPUT98), .Z(new_n858));
  NAND2_X1  g433(.A1(new_n849), .A2(new_n856), .ZN(new_n859));
  XOR2_X1   g434(.A(new_n859), .B(KEYINPUT97), .Z(new_n860));
  OAI21_X1  g435(.A(new_n846), .B1(new_n858), .B2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(G37), .ZN(new_n862));
  INV_X1    g437(.A(new_n846), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n857), .A2(new_n859), .A3(new_n863), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n861), .A2(new_n862), .A3(new_n864), .ZN(new_n865));
  XOR2_X1   g440(.A(KEYINPUT99), .B(KEYINPUT40), .Z(new_n866));
  XNOR2_X1  g441(.A(new_n865), .B(new_n866), .ZN(G395));
  NAND3_X1  g442(.A1(new_n602), .A2(new_n561), .A3(new_n562), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n602), .B1(new_n561), .B2(new_n562), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n608), .B(new_n842), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT41), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n874), .B1(new_n869), .B2(new_n870), .ZN(new_n875));
  NAND2_X1  g450(.A1(G299), .A2(new_n607), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n876), .A2(KEYINPUT41), .A3(new_n868), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n873), .B1(new_n878), .B2(new_n872), .ZN(new_n879));
  NAND2_X1  g454(.A1(G303), .A2(new_n785), .ZN(new_n880));
  NAND2_X1  g455(.A1(G166), .A2(G288), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(new_n584), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n880), .A2(G305), .A3(new_n881), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n885), .A2(G290), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n883), .A2(new_n806), .A3(new_n884), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(KEYINPUT42), .ZN(new_n889));
  OR2_X1    g464(.A1(new_n879), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n879), .A2(new_n889), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n890), .A2(G868), .A3(new_n891), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n841), .A2(G868), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n892), .B1(KEYINPUT100), .B2(new_n893), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n894), .B1(KEYINPUT100), .B2(new_n892), .ZN(G295));
  OAI21_X1  g470(.A(new_n894), .B1(KEYINPUT100), .B2(new_n892), .ZN(G331));
  INV_X1    g471(.A(KEYINPUT44), .ZN(new_n897));
  AND3_X1   g472(.A1(new_n883), .A2(new_n806), .A3(new_n884), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n806), .B1(new_n883), .B2(new_n884), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT102), .ZN(new_n900));
  NOR3_X1   g475(.A1(new_n898), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(KEYINPUT102), .B1(new_n886), .B2(new_n887), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  XOR2_X1   g478(.A(new_n544), .B(new_n841), .Z(new_n904));
  AND3_X1   g479(.A1(new_n521), .A2(KEYINPUT76), .A3(new_n526), .ZN(new_n905));
  NOR3_X1   g480(.A1(new_n905), .A2(new_n564), .A3(G301), .ZN(new_n906));
  NAND2_X1  g481(.A1(G168), .A2(G301), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n904), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n565), .A2(G171), .A3(new_n566), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n910), .A2(new_n842), .A3(new_n907), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  AND3_X1   g487(.A1(new_n875), .A2(new_n912), .A3(new_n877), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n876), .A2(new_n868), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n909), .A2(KEYINPUT101), .A3(new_n911), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT101), .ZN(new_n916));
  OAI211_X1 g491(.A(new_n904), .B(new_n916), .C1(new_n906), .C2(new_n908), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n914), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n903), .B1(new_n913), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n915), .A2(new_n917), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(new_n871), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n875), .A2(new_n912), .A3(new_n877), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n921), .A2(new_n888), .A3(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT43), .ZN(new_n924));
  NAND4_X1  g499(.A1(new_n919), .A2(new_n923), .A3(new_n924), .A4(new_n862), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT103), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n897), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n871), .A2(new_n911), .A3(new_n909), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n928), .B1(new_n878), .B2(new_n920), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(new_n903), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n930), .A2(new_n862), .A3(new_n923), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n931), .A2(KEYINPUT43), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n913), .A2(new_n918), .ZN(new_n933));
  AOI21_X1  g508(.A(G37), .B1(new_n933), .B2(new_n888), .ZN(new_n934));
  NAND4_X1  g509(.A1(new_n934), .A2(KEYINPUT103), .A3(new_n924), .A4(new_n919), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n927), .A2(new_n932), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n924), .B1(new_n934), .B2(new_n919), .ZN(new_n937));
  AND4_X1   g512(.A1(new_n924), .A2(new_n930), .A3(new_n862), .A4(new_n923), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n897), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n936), .A2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT104), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n936), .A2(new_n939), .A3(KEYINPUT104), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(G397));
  INV_X1    g519(.A(new_n583), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(KEYINPUT113), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n577), .A2(KEYINPUT77), .A3(G651), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n577), .A2(G651), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(new_n579), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT113), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n583), .A2(new_n950), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n946), .A2(new_n947), .A3(new_n949), .A4(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(G1981), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT112), .ZN(new_n954));
  INV_X1    g529(.A(G1981), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n954), .B1(new_n584), .B2(new_n955), .ZN(new_n956));
  NAND4_X1  g531(.A1(new_n949), .A2(new_n955), .A3(new_n947), .A4(new_n945), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n957), .A2(KEYINPUT112), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n953), .B1(new_n956), .B2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT49), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  XNOR2_X1  g536(.A(new_n957), .B(KEYINPUT112), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n962), .A2(KEYINPUT49), .A3(new_n953), .ZN(new_n963));
  XOR2_X1   g538(.A(KEYINPUT105), .B(G40), .Z(new_n964));
  NOR3_X1   g539(.A1(new_n468), .A2(new_n471), .A3(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(G1384), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n965), .A2(new_n966), .A3(new_n497), .ZN(new_n967));
  INV_X1    g542(.A(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(G8), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n961), .A2(new_n963), .A3(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n572), .A2(G1976), .A3(new_n573), .ZN(new_n972));
  AND3_X1   g547(.A1(new_n967), .A2(G8), .A3(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT111), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT52), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n785), .A2(G1976), .ZN(new_n976));
  INV_X1    g551(.A(new_n976), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n973), .A2(new_n974), .A3(new_n975), .A4(new_n977), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n967), .A2(new_n975), .A3(G8), .A4(new_n972), .ZN(new_n979));
  OAI21_X1  g554(.A(KEYINPUT111), .B1(new_n979), .B2(new_n976), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n973), .A2(KEYINPUT110), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n967), .A2(G8), .A3(new_n972), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT110), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n982), .A2(KEYINPUT52), .A3(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n971), .A2(new_n981), .A3(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT50), .ZN(new_n988));
  AND3_X1   g563(.A1(new_n497), .A2(new_n988), .A3(new_n966), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n988), .B1(new_n497), .B2(new_n966), .ZN(new_n990));
  OR3_X1    g565(.A1(new_n468), .A2(new_n471), .A3(new_n964), .ZN(new_n991));
  NOR3_X1   g566(.A1(new_n989), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(new_n694), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n497), .A2(new_n966), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT45), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n497), .A2(KEYINPUT45), .A3(new_n966), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n996), .A2(new_n965), .A3(new_n997), .ZN(new_n998));
  XNOR2_X1  g573(.A(KEYINPUT108), .B(G1971), .ZN(new_n999));
  INV_X1    g574(.A(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n969), .B1(new_n993), .B2(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g577(.A(KEYINPUT109), .B(KEYINPUT55), .ZN(new_n1003));
  NAND3_X1  g578(.A1(G303), .A2(G8), .A3(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(KEYINPUT109), .A2(KEYINPUT55), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1005), .B1(G166), .B2(new_n969), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n1002), .A2(new_n1007), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n987), .A2(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g584(.A(KEYINPUT116), .B(G2084), .ZN(new_n1010));
  AOI22_X1  g585(.A1(new_n992), .A2(new_n1010), .B1(new_n998), .B2(new_n758), .ZN(new_n1011));
  NOR3_X1   g586(.A1(new_n1011), .A2(G286), .A3(new_n969), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1009), .A2(new_n1012), .ZN(new_n1013));
  AND2_X1   g588(.A1(new_n961), .A2(new_n963), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n785), .A2(new_n788), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n962), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  AOI22_X1  g591(.A1(new_n1013), .A2(KEYINPUT63), .B1(new_n970), .B2(new_n1016), .ZN(new_n1017));
  AND2_X1   g592(.A1(new_n1002), .A2(new_n1007), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1018), .A2(new_n981), .A3(new_n971), .A4(new_n986), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT115), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n987), .A2(new_n1020), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n971), .A2(new_n981), .A3(KEYINPUT115), .A4(new_n986), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n990), .A2(new_n991), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT114), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g601(.A(KEYINPUT114), .B1(new_n990), .B2(new_n991), .ZN(new_n1027));
  AOI211_X1 g602(.A(G2090), .B(new_n989), .C1(new_n1026), .C2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1001), .ZN(new_n1029));
  OAI21_X1  g604(.A(G8), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1007), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1018), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT63), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n1023), .A2(new_n1032), .A3(new_n1033), .A4(new_n1012), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1017), .A2(new_n1019), .A3(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT53), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1036), .B1(new_n998), .B2(G2078), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n497), .A2(new_n988), .A3(new_n966), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1024), .A2(new_n1038), .ZN(new_n1039));
  XOR2_X1   g614(.A(KEYINPUT123), .B(G1961), .Z(new_n1040));
  INV_X1    g615(.A(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n996), .A2(new_n997), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1036), .A2(G2078), .ZN(new_n1044));
  NAND3_X1  g619(.A1(G160), .A2(G40), .A3(new_n1044), .ZN(new_n1045));
  OAI211_X1 g620(.A(new_n1037), .B(new_n1042), .C1(new_n1043), .C2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(G171), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT124), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1044), .ZN(new_n1049));
  OAI211_X1 g624(.A(new_n1042), .B(new_n1048), .C1(new_n998), .C2(new_n1049), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n992), .A2(new_n1040), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n998), .A2(new_n1049), .ZN(new_n1052));
  OAI21_X1  g627(.A(KEYINPUT124), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1050), .A2(new_n1053), .A3(new_n1037), .ZN(new_n1054));
  OAI211_X1 g629(.A(KEYINPUT54), .B(new_n1047), .C1(new_n1054), .C2(G171), .ZN(new_n1055));
  AND3_X1   g630(.A1(new_n1023), .A2(new_n1032), .A3(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT54), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1054), .A2(G171), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1058), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1046), .A2(G171), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1057), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  OAI21_X1  g636(.A(KEYINPUT121), .B1(new_n1011), .B2(new_n969), .ZN(new_n1062));
  NOR2_X1   g637(.A1(G168), .A2(new_n969), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1063), .A2(KEYINPUT51), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n994), .A2(KEYINPUT50), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1065), .A2(new_n965), .A3(new_n1038), .A4(new_n1010), .ZN(new_n1066));
  AND3_X1   g641(.A1(new_n996), .A2(new_n965), .A3(new_n997), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1066), .B1(new_n1067), .B2(G1966), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT121), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1068), .A2(new_n1069), .A3(G8), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1062), .A2(new_n1064), .A3(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(KEYINPUT122), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n969), .B1(new_n1011), .B2(G168), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(KEYINPUT51), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT122), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1062), .A2(new_n1070), .A3(new_n1075), .A4(new_n1064), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1072), .A2(new_n1074), .A3(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1068), .A2(new_n1063), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  AND3_X1   g654(.A1(new_n1056), .A2(new_n1061), .A3(new_n1079), .ZN(new_n1080));
  XNOR2_X1  g655(.A(KEYINPUT58), .B(G1341), .ZN(new_n1081));
  OAI22_X1  g656(.A1(new_n998), .A2(G1996), .B1(new_n968), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT118), .ZN(new_n1083));
  AND3_X1   g658(.A1(new_n1082), .A2(new_n1083), .A3(new_n544), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1084), .A2(KEYINPUT59), .ZN(new_n1085));
  XOR2_X1   g660(.A(new_n559), .B(KEYINPUT57), .Z(new_n1086));
  INV_X1    g661(.A(new_n1086), .ZN(new_n1087));
  XNOR2_X1  g662(.A(KEYINPUT56), .B(G2072), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1067), .A2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n989), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1089), .B1(new_n1090), .B2(G1956), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1087), .A2(new_n1091), .ZN(new_n1092));
  OAI211_X1 g667(.A(new_n1086), .B(new_n1089), .C1(new_n1090), .C2(G1956), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT61), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1085), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  OAI22_X1  g671(.A1(new_n992), .A2(G1348), .B1(G2067), .B2(new_n967), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT60), .ZN(new_n1098));
  OAI211_X1 g673(.A(KEYINPUT119), .B(new_n607), .C1(new_n1097), .C2(new_n1098), .ZN(new_n1099));
  AOI22_X1  g674(.A1(new_n1039), .A2(new_n701), .B1(new_n720), .B2(new_n968), .ZN(new_n1100));
  OR2_X1    g675(.A1(new_n607), .A2(KEYINPUT119), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n607), .A2(KEYINPUT119), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1100), .A2(new_n1101), .A3(KEYINPUT60), .A4(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1099), .A2(new_n1103), .A3(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(KEYINPUT120), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT120), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1099), .A2(new_n1103), .A3(new_n1107), .A4(new_n1104), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1106), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1084), .A2(KEYINPUT59), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1092), .A2(new_n1093), .A3(KEYINPUT61), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1096), .A2(new_n1109), .A3(new_n1110), .A4(new_n1111), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1092), .B1(new_n607), .B2(new_n1100), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(new_n1093), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT117), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1113), .A2(KEYINPUT117), .A3(new_n1093), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1112), .A2(new_n1116), .A3(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1035), .B1(new_n1080), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1079), .A2(KEYINPUT62), .ZN(new_n1120));
  AND2_X1   g695(.A1(new_n1023), .A2(new_n1032), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT62), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1077), .A2(new_n1122), .A3(new_n1078), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1120), .A2(new_n1121), .A3(new_n1059), .A4(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(KEYINPUT125), .ZN(new_n1125));
  AND2_X1   g700(.A1(new_n1123), .A2(new_n1059), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT125), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1126), .A2(new_n1127), .A3(new_n1121), .A4(new_n1120), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1119), .A2(new_n1125), .A3(new_n1128), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n996), .A2(new_n991), .ZN(new_n1130));
  XNOR2_X1  g705(.A(new_n1130), .B(KEYINPUT106), .ZN(new_n1131));
  INV_X1    g706(.A(G1996), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n744), .A2(new_n1132), .ZN(new_n1133));
  XNOR2_X1  g708(.A(new_n717), .B(G2067), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1131), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1135), .B1(new_n743), .B2(new_n1136), .ZN(new_n1137));
  XNOR2_X1  g712(.A(new_n815), .B(new_n817), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT107), .ZN(new_n1139));
  OR2_X1    g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1140), .A2(new_n1131), .A3(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1142), .ZN(new_n1143));
  XNOR2_X1  g718(.A(G290), .B(G1986), .ZN(new_n1144));
  AOI211_X1 g719(.A(new_n1137), .B(new_n1143), .C1(new_n1130), .C2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1129), .A2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1131), .B1(new_n743), .B2(new_n1134), .ZN(new_n1147));
  NOR2_X1   g722(.A1(KEYINPUT126), .A2(KEYINPUT46), .ZN(new_n1148));
  AND2_X1   g723(.A1(KEYINPUT126), .A2(KEYINPUT46), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1136), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  OAI211_X1 g725(.A(new_n1147), .B(new_n1150), .C1(new_n1136), .C2(new_n1148), .ZN(new_n1151));
  XOR2_X1   g726(.A(new_n1151), .B(KEYINPUT47), .Z(new_n1152));
  NAND3_X1  g727(.A1(new_n806), .A2(new_n680), .A3(new_n1130), .ZN(new_n1153));
  XOR2_X1   g728(.A(new_n1153), .B(KEYINPUT48), .Z(new_n1154));
  NOR3_X1   g729(.A1(new_n1143), .A2(new_n1137), .A3(new_n1154), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n812), .A2(new_n817), .A3(new_n814), .ZN(new_n1156));
  OAI22_X1  g731(.A1(new_n1137), .A2(new_n1156), .B1(G2067), .B2(new_n717), .ZN(new_n1157));
  AOI211_X1 g732(.A(new_n1152), .B(new_n1155), .C1(new_n1131), .C2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1146), .A2(new_n1158), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g734(.A1(G401), .A2(G227), .ZN(new_n1161));
  NAND3_X1  g735(.A1(new_n688), .A2(G319), .A3(new_n1161), .ZN(new_n1162));
  XOR2_X1   g736(.A(new_n1162), .B(KEYINPUT127), .Z(new_n1163));
  OR2_X1    g737(.A1(new_n937), .A2(new_n938), .ZN(new_n1164));
  AND3_X1   g738(.A1(new_n1163), .A2(new_n865), .A3(new_n1164), .ZN(G308));
  NAND3_X1  g739(.A1(new_n1163), .A2(new_n865), .A3(new_n1164), .ZN(G225));
endmodule


