//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 1 0 1 1 1 0 0 1 1 1 1 1 0 1 1 1 1 1 1 1 1 1 1 0 0 1 1 1 0 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 1 1 1 0 0 1 1 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:44 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n699,
    new_n700, new_n701, new_n702, new_n704, new_n705, new_n706, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n763, new_n764, new_n765, new_n766,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n797,
    new_n798, new_n799, new_n800, new_n802, new_n803, new_n804, new_n806,
    new_n807, new_n808, new_n810, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n837, new_n838,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n888, new_n889, new_n891,
    new_n892, new_n893, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n960, new_n961, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n980, new_n981, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1022, new_n1023, new_n1024, new_n1025;
  XOR2_X1   g000(.A(KEYINPUT95), .B(KEYINPUT13), .Z(new_n202));
  NAND2_X1  g001(.A1(G229gat), .A2(G233gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT15), .ZN(new_n205));
  XNOR2_X1  g004(.A(G43gat), .B(G50gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT91), .ZN(new_n207));
  AOI21_X1  g006(.A(new_n205), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n208), .B1(new_n207), .B2(new_n206), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT94), .ZN(new_n210));
  OR2_X1    g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n209), .A2(new_n210), .ZN(new_n212));
  NAND2_X1  g011(.A1(G29gat), .A2(G36gat), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT92), .ZN(new_n214));
  XNOR2_X1  g013(.A(new_n213), .B(new_n214), .ZN(new_n215));
  OR3_X1    g014(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n216));
  OAI21_X1  g015(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n206), .A2(KEYINPUT15), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n211), .A2(new_n212), .A3(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(new_n219), .ZN(new_n223));
  OAI21_X1  g022(.A(KEYINPUT93), .B1(new_n209), .B2(new_n223), .ZN(new_n224));
  OR3_X1    g023(.A1(new_n209), .A2(new_n223), .A3(KEYINPUT93), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n222), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(G15gat), .B(G22gat), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT16), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n227), .B1(new_n228), .B2(G1gat), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n229), .B1(G1gat), .B2(new_n227), .ZN(new_n230));
  INV_X1    g029(.A(G8gat), .ZN(new_n231));
  XNOR2_X1  g030(.A(new_n230), .B(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  AND2_X1   g032(.A1(new_n226), .A2(new_n233), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n226), .A2(new_n233), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n204), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(KEYINPUT96), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT96), .ZN(new_n238));
  OAI211_X1 g037(.A(new_n238), .B(new_n204), .C1(new_n234), .C2(new_n235), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT17), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n226), .A2(new_n240), .ZN(new_n241));
  NAND4_X1  g040(.A1(new_n222), .A2(new_n224), .A3(KEYINPUT17), .A4(new_n225), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n241), .A2(new_n232), .A3(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n226), .A2(new_n233), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n243), .A2(new_n203), .A3(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT18), .ZN(new_n246));
  AOI22_X1  g045(.A1(new_n237), .A2(new_n239), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  AND2_X1   g046(.A1(new_n243), .A2(new_n244), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n248), .A2(KEYINPUT18), .A3(new_n203), .ZN(new_n249));
  XNOR2_X1  g048(.A(G113gat), .B(G141gat), .ZN(new_n250));
  XNOR2_X1  g049(.A(KEYINPUT90), .B(KEYINPUT11), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XOR2_X1   g051(.A(G169gat), .B(G197gat), .Z(new_n253));
  XNOR2_X1  g052(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n254), .B(KEYINPUT12), .ZN(new_n255));
  AND3_X1   g054(.A1(new_n247), .A2(new_n249), .A3(new_n255), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n255), .B1(new_n247), .B2(new_n249), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT97), .ZN(new_n258));
  NOR3_X1   g057(.A1(new_n256), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n247), .A2(new_n249), .ZN(new_n260));
  INV_X1    g059(.A(new_n255), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n247), .A2(new_n249), .A3(new_n255), .ZN(new_n263));
  AOI21_X1  g062(.A(KEYINPUT97), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n259), .A2(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(G78gat), .B(G106gat), .ZN(new_n266));
  XNOR2_X1  g065(.A(KEYINPUT31), .B(G50gat), .ZN(new_n267));
  XOR2_X1   g066(.A(new_n266), .B(new_n267), .Z(new_n268));
  NAND2_X1  g067(.A1(G228gat), .A2(G233gat), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n269), .B(KEYINPUT78), .ZN(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT29), .ZN(new_n272));
  NAND2_X1  g071(.A1(G211gat), .A2(G218gat), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT22), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT71), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  OR2_X1    g076(.A1(G197gat), .A2(G204gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(G197gat), .A2(G204gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  AOI21_X1  g079(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(KEYINPUT71), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n277), .A2(new_n280), .A3(new_n282), .ZN(new_n283));
  XNOR2_X1  g082(.A(G211gat), .B(G218gat), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  AOI22_X1  g085(.A1(new_n278), .A2(new_n279), .B1(new_n281), .B2(KEYINPUT71), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n284), .B1(new_n287), .B2(new_n277), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n272), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  XOR2_X1   g088(.A(KEYINPUT73), .B(KEYINPUT3), .Z(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  AND2_X1   g090(.A1(G155gat), .A2(G162gat), .ZN(new_n292));
  NOR2_X1   g091(.A1(G155gat), .A2(G162gat), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(G141gat), .B(G148gat), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT2), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n296), .B1(G155gat), .B2(G162gat), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n294), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(G141gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(G148gat), .ZN(new_n300));
  INV_X1    g099(.A(G148gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(G141gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  XNOR2_X1  g102(.A(G155gat), .B(G162gat), .ZN(new_n304));
  INV_X1    g103(.A(G155gat), .ZN(new_n305));
  INV_X1    g104(.A(G162gat), .ZN(new_n306));
  OAI21_X1  g105(.A(KEYINPUT2), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n303), .A2(new_n304), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n298), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n291), .A2(new_n309), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n286), .A2(new_n288), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n298), .A2(new_n308), .A3(new_n290), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(new_n272), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n271), .B1(new_n310), .B2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT81), .ZN(new_n316));
  INV_X1    g115(.A(new_n269), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT80), .ZN(new_n318));
  AND3_X1   g117(.A1(new_n311), .A2(new_n313), .A3(new_n318), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n318), .B1(new_n311), .B2(new_n313), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n317), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  AND2_X1   g120(.A1(new_n298), .A2(new_n308), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT79), .ZN(new_n323));
  AOI21_X1  g122(.A(KEYINPUT3), .B1(new_n289), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n283), .A2(new_n285), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n287), .A2(new_n284), .A3(new_n277), .ZN(new_n326));
  AOI21_X1  g125(.A(KEYINPUT29), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(KEYINPUT79), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n322), .B1(new_n324), .B2(new_n328), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n316), .B1(new_n321), .B2(new_n329), .ZN(new_n330));
  AND2_X1   g129(.A1(new_n312), .A2(new_n272), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n325), .A2(new_n326), .ZN(new_n332));
  OAI21_X1  g131(.A(KEYINPUT80), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n311), .A2(new_n313), .A3(new_n318), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n269), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT3), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n336), .B1(new_n327), .B2(KEYINPUT79), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n289), .A2(new_n323), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n309), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n335), .A2(new_n339), .A3(KEYINPUT81), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n315), .B1(new_n330), .B2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT82), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n342), .A2(G22gat), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n268), .B1(new_n341), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n342), .A2(G22gat), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  AOI211_X1 g146(.A(new_n315), .B(new_n347), .C1(new_n330), .C2(new_n340), .ZN(new_n348));
  OR2_X1    g147(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n315), .ZN(new_n350));
  NAND2_X1  g149(.A1(KEYINPUT83), .A2(G22gat), .ZN(new_n351));
  AND3_X1   g150(.A1(new_n335), .A2(new_n339), .A3(KEYINPUT81), .ZN(new_n352));
  AOI21_X1  g151(.A(KEYINPUT81), .B1(new_n335), .B2(new_n339), .ZN(new_n353));
  OAI211_X1 g152(.A(new_n350), .B(new_n351), .C1(new_n352), .C2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n268), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n330), .A2(new_n340), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n351), .B1(new_n357), .B2(new_n350), .ZN(new_n358));
  NOR3_X1   g157(.A1(new_n356), .A2(new_n358), .A3(KEYINPUT84), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT84), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n268), .B1(new_n341), .B2(new_n351), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n350), .B1(new_n352), .B2(new_n353), .ZN(new_n362));
  INV_X1    g161(.A(new_n351), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n360), .B1(new_n361), .B2(new_n364), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n349), .B1(new_n359), .B2(new_n365), .ZN(new_n366));
  XNOR2_X1  g165(.A(KEYINPUT27), .B(G183gat), .ZN(new_n367));
  INV_X1    g166(.A(G190gat), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n367), .A2(KEYINPUT28), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(KEYINPUT67), .A2(G183gat), .ZN(new_n370));
  AOI21_X1  g169(.A(G190gat), .B1(new_n370), .B2(KEYINPUT27), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT27), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n372), .A2(KEYINPUT67), .A3(G183gat), .ZN(new_n373));
  AND2_X1   g172(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n369), .B1(new_n374), .B2(KEYINPUT28), .ZN(new_n375));
  NAND2_X1  g174(.A1(G183gat), .A2(G190gat), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(G169gat), .A2(G176gat), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(KEYINPUT64), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT64), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n380), .A2(G169gat), .A3(G176gat), .ZN(new_n381));
  INV_X1    g180(.A(G169gat), .ZN(new_n382));
  INV_X1    g181(.A(G176gat), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  AOI22_X1  g183(.A1(new_n379), .A2(new_n381), .B1(new_n384), .B2(KEYINPUT26), .ZN(new_n385));
  NOR2_X1   g184(.A1(G169gat), .A2(G176gat), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT66), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT26), .ZN(new_n389));
  OAI21_X1  g188(.A(KEYINPUT66), .B1(G169gat), .B2(G176gat), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n388), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n377), .B1(new_n385), .B2(new_n391), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n375), .B1(new_n392), .B2(KEYINPUT68), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT68), .ZN(new_n394));
  AOI211_X1 g193(.A(new_n394), .B(new_n377), .C1(new_n385), .C2(new_n391), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n381), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT65), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n379), .A2(new_n381), .A3(KEYINPUT65), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n388), .A2(KEYINPUT23), .A3(new_n390), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n398), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT25), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT23), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n402), .B1(new_n384), .B2(new_n403), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n376), .A2(KEYINPUT24), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT24), .ZN(new_n407));
  XNOR2_X1  g206(.A(G183gat), .B(G190gat), .ZN(new_n408));
  OAI211_X1 g207(.A(new_n404), .B(new_n406), .C1(new_n407), .C2(new_n408), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n401), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n384), .A2(new_n403), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n386), .A2(KEYINPUT23), .ZN(new_n412));
  AND3_X1   g211(.A1(new_n396), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  XOR2_X1   g212(.A(G183gat), .B(G190gat), .Z(new_n414));
  AOI21_X1  g213(.A(new_n405), .B1(new_n414), .B2(KEYINPUT24), .ZN(new_n415));
  AOI21_X1  g214(.A(KEYINPUT25), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  OAI22_X1  g215(.A1(new_n393), .A2(new_n395), .B1(new_n410), .B2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(G134gat), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(G127gat), .ZN(new_n419));
  INV_X1    g218(.A(G127gat), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(G134gat), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  XNOR2_X1  g221(.A(G113gat), .B(G120gat), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n422), .B1(new_n423), .B2(KEYINPUT1), .ZN(new_n424));
  INV_X1    g223(.A(G120gat), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(G113gat), .ZN(new_n426));
  INV_X1    g225(.A(G113gat), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(G120gat), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  XNOR2_X1  g228(.A(G127gat), .B(G134gat), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT1), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n429), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  AND3_X1   g231(.A1(new_n424), .A2(new_n432), .A3(KEYINPUT69), .ZN(new_n433));
  AOI21_X1  g232(.A(KEYINPUT69), .B1(new_n424), .B2(new_n432), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n417), .A2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(G227gat), .ZN(new_n438));
  INV_X1    g237(.A(G233gat), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n406), .B1(new_n408), .B2(new_n407), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n396), .A2(new_n411), .A3(new_n412), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n402), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n443), .B1(new_n409), .B2(new_n401), .ZN(new_n444));
  OAI211_X1 g243(.A(new_n444), .B(new_n435), .C1(new_n395), .C2(new_n393), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n437), .A2(new_n440), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(KEYINPUT32), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(KEYINPUT70), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT70), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n446), .A2(new_n449), .A3(KEYINPUT32), .ZN(new_n450));
  XNOR2_X1  g249(.A(G15gat), .B(G43gat), .ZN(new_n451));
  XNOR2_X1  g250(.A(G71gat), .B(G99gat), .ZN(new_n452));
  XNOR2_X1  g251(.A(new_n451), .B(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT33), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n453), .B1(new_n446), .B2(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n448), .A2(new_n450), .A3(new_n455), .ZN(new_n456));
  OAI211_X1 g255(.A(new_n446), .B(KEYINPUT32), .C1(new_n454), .C2(new_n453), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n440), .B1(new_n437), .B2(new_n445), .ZN(new_n459));
  XNOR2_X1  g258(.A(new_n459), .B(KEYINPUT34), .ZN(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n458), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n456), .A2(new_n460), .A3(new_n457), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n366), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  XNOR2_X1  g263(.A(G1gat), .B(G29gat), .ZN(new_n465));
  XNOR2_X1  g264(.A(new_n465), .B(KEYINPUT0), .ZN(new_n466));
  XNOR2_X1  g265(.A(G57gat), .B(G85gat), .ZN(new_n467));
  XOR2_X1   g266(.A(new_n466), .B(new_n467), .Z(new_n468));
  INV_X1    g267(.A(new_n468), .ZN(new_n469));
  XNOR2_X1  g268(.A(KEYINPUT75), .B(KEYINPUT5), .ZN(new_n470));
  INV_X1    g269(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n424), .A2(new_n432), .ZN(new_n472));
  AND2_X1   g271(.A1(new_n309), .A2(new_n472), .ZN(new_n473));
  AND2_X1   g272(.A1(new_n424), .A2(new_n432), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n322), .A2(new_n474), .A3(KEYINPUT74), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT74), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n476), .B1(new_n309), .B2(new_n472), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n473), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(G225gat), .A2(G233gat), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n471), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  AND2_X1   g279(.A1(new_n312), .A2(new_n472), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT72), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n482), .B1(new_n309), .B2(KEYINPUT3), .ZN(new_n483));
  AOI211_X1 g282(.A(KEYINPUT72), .B(new_n336), .C1(new_n298), .C2(new_n308), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n481), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(new_n479), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  AOI21_X1  g287(.A(KEYINPUT4), .B1(new_n475), .B2(new_n477), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT4), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT69), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n472), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n424), .A2(new_n432), .A3(KEYINPUT69), .ZN(new_n493));
  AOI211_X1 g292(.A(new_n490), .B(new_n309), .C1(new_n492), .C2(new_n493), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n489), .A2(new_n494), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n480), .B1(new_n488), .B2(new_n495), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n309), .B1(new_n492), .B2(new_n493), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT76), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n497), .A2(new_n498), .A3(new_n490), .ZN(new_n499));
  OAI211_X1 g298(.A(new_n490), .B(new_n322), .C1(new_n433), .C2(new_n434), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(KEYINPUT76), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n490), .B1(new_n475), .B2(new_n477), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n499), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n485), .A2(new_n479), .A3(new_n470), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  OAI211_X1 g304(.A(KEYINPUT6), .B(new_n469), .C1(new_n496), .C2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT77), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n500), .A2(KEYINPUT76), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n498), .B1(new_n497), .B2(new_n490), .ZN(new_n510));
  AOI21_X1  g309(.A(KEYINPUT74), .B1(new_n322), .B2(new_n474), .ZN(new_n511));
  NOR3_X1   g310(.A1(new_n309), .A2(new_n472), .A3(new_n476), .ZN(new_n512));
  OAI21_X1  g311(.A(KEYINPUT4), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n509), .B1(new_n510), .B2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(new_n504), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  OAI22_X1  g315(.A1(new_n511), .A2(new_n512), .B1(new_n322), .B2(new_n474), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n470), .B1(new_n517), .B2(new_n487), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n490), .B1(new_n511), .B2(new_n512), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n497), .A2(KEYINPUT4), .ZN(new_n520));
  NAND4_X1  g319(.A1(new_n519), .A2(new_n520), .A3(new_n479), .A4(new_n485), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n518), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n468), .B1(new_n516), .B2(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n523), .A2(KEYINPUT77), .A3(KEYINPUT6), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n523), .A2(KEYINPUT6), .ZN(new_n527));
  AOI22_X1  g326(.A1(new_n514), .A2(new_n515), .B1(new_n518), .B2(new_n521), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(new_n468), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n526), .A2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(G226gat), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n532), .A2(new_n439), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n533), .B1(new_n417), .B2(new_n272), .ZN(new_n534));
  INV_X1    g333(.A(new_n533), .ZN(new_n535));
  AND2_X1   g334(.A1(new_n385), .A2(new_n391), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n394), .B1(new_n536), .B2(new_n377), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n392), .A2(KEYINPUT68), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n537), .A2(new_n538), .A3(new_n375), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n535), .B1(new_n539), .B2(new_n444), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n311), .B1(new_n534), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n417), .A2(new_n533), .ZN(new_n542));
  AOI21_X1  g341(.A(KEYINPUT29), .B1(new_n539), .B2(new_n444), .ZN(new_n543));
  OAI211_X1 g342(.A(new_n542), .B(new_n332), .C1(new_n543), .C2(new_n533), .ZN(new_n544));
  XNOR2_X1  g343(.A(G8gat), .B(G36gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(G64gat), .B(G92gat), .ZN(new_n546));
  XOR2_X1   g345(.A(new_n545), .B(new_n546), .Z(new_n547));
  AND3_X1   g346(.A1(new_n541), .A2(new_n544), .A3(new_n547), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n547), .B1(new_n541), .B2(new_n544), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT30), .ZN(new_n550));
  NOR3_X1   g349(.A1(new_n548), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n541), .ZN(new_n552));
  INV_X1    g351(.A(new_n544), .ZN(new_n553));
  INV_X1    g352(.A(new_n547), .ZN(new_n554));
  NOR4_X1   g353(.A1(new_n552), .A2(new_n553), .A3(KEYINPUT30), .A4(new_n554), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n551), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n531), .A2(new_n557), .ZN(new_n558));
  OAI21_X1  g357(.A(KEYINPUT35), .B1(new_n464), .B2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT89), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n345), .A2(new_n348), .ZN(new_n561));
  OAI21_X1  g360(.A(KEYINPUT84), .B1(new_n356), .B2(new_n358), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n361), .A2(new_n360), .A3(new_n364), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n561), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT6), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n565), .B1(new_n528), .B2(new_n468), .ZN(new_n566));
  NOR3_X1   g365(.A1(new_n496), .A2(new_n505), .A3(new_n469), .ZN(new_n567));
  OAI21_X1  g366(.A(KEYINPUT86), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT86), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n527), .A2(new_n569), .A3(new_n529), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n525), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(KEYINPUT88), .B(KEYINPUT35), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n573), .B1(new_n551), .B2(new_n555), .ZN(new_n574));
  NOR3_X1   g373(.A1(new_n564), .A2(new_n571), .A3(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT87), .ZN(new_n576));
  AND3_X1   g375(.A1(new_n456), .A2(new_n460), .A3(new_n457), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n460), .B1(new_n456), .B2(new_n457), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n576), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n462), .A2(KEYINPUT87), .A3(new_n463), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n560), .B1(new_n575), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n570), .A2(new_n568), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n574), .B1(new_n583), .B2(new_n526), .ZN(new_n584));
  AND4_X1   g383(.A1(new_n560), .A2(new_n581), .A3(new_n584), .A4(new_n366), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n559), .B1(new_n582), .B2(new_n585), .ZN(new_n586));
  OAI21_X1  g385(.A(KEYINPUT37), .B1(new_n552), .B2(new_n553), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT37), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n541), .A2(new_n544), .A3(new_n588), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n587), .A2(new_n554), .A3(new_n589), .ZN(new_n590));
  OR2_X1    g389(.A1(new_n590), .A2(KEYINPUT38), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n548), .B1(new_n590), .B2(KEYINPUT38), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n571), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n487), .B1(new_n503), .B2(new_n486), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT39), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n595), .B1(new_n478), .B2(new_n479), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  OAI211_X1 g396(.A(new_n595), .B(new_n487), .C1(new_n503), .C2(new_n486), .ZN(new_n598));
  NAND4_X1  g397(.A1(new_n597), .A2(KEYINPUT40), .A3(new_n468), .A4(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(KEYINPUT85), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n597), .A2(new_n468), .A3(new_n598), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT40), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n523), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n600), .A2(new_n556), .A3(new_n603), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n593), .A2(new_n604), .A3(new_n366), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n558), .A2(new_n564), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n462), .A2(new_n463), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT36), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n605), .A2(new_n606), .A3(new_n609), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n265), .B1(new_n586), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(G85gat), .A2(G92gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(KEYINPUT7), .ZN(new_n613));
  INV_X1    g412(.A(G99gat), .ZN(new_n614));
  INV_X1    g413(.A(G106gat), .ZN(new_n615));
  OAI21_X1  g414(.A(KEYINPUT8), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(KEYINPUT101), .B(G85gat), .ZN(new_n617));
  OAI211_X1 g416(.A(new_n613), .B(new_n616), .C1(G92gat), .C2(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(G99gat), .B(G106gat), .ZN(new_n619));
  XOR2_X1   g418(.A(new_n618), .B(new_n619), .Z(new_n620));
  NAND3_X1  g419(.A1(new_n241), .A2(new_n242), .A3(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n618), .B(new_n619), .ZN(new_n622));
  AND2_X1   g421(.A1(G232gat), .A2(G233gat), .ZN(new_n623));
  AOI22_X1  g422(.A1(new_n226), .A2(new_n622), .B1(KEYINPUT41), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n621), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(G190gat), .B(G218gat), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n621), .A2(new_n624), .A3(new_n626), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n623), .A2(KEYINPUT41), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(KEYINPUT99), .ZN(new_n631));
  XNOR2_X1  g430(.A(G134gat), .B(G162gat), .ZN(new_n632));
  XOR2_X1   g431(.A(new_n631), .B(new_n632), .Z(new_n633));
  XOR2_X1   g432(.A(new_n633), .B(KEYINPUT100), .Z(new_n634));
  NAND3_X1  g433(.A1(new_n628), .A2(new_n629), .A3(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(KEYINPUT102), .ZN(new_n636));
  INV_X1    g435(.A(new_n633), .ZN(new_n637));
  INV_X1    g436(.A(new_n629), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n626), .B1(new_n621), .B2(new_n624), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n637), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n640), .A2(KEYINPUT103), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT103), .ZN(new_n642));
  OAI211_X1 g441(.A(new_n642), .B(new_n637), .C1(new_n638), .C2(new_n639), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  AND2_X1   g443(.A1(new_n636), .A2(new_n644), .ZN(new_n645));
  XOR2_X1   g444(.A(G57gat), .B(G64gat), .Z(new_n646));
  INV_X1    g445(.A(KEYINPUT9), .ZN(new_n647));
  INV_X1    g446(.A(G71gat), .ZN(new_n648));
  INV_X1    g447(.A(G78gat), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n647), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n646), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(G71gat), .B(G78gat), .ZN(new_n652));
  XOR2_X1   g451(.A(new_n651), .B(new_n652), .Z(new_n653));
  INV_X1    g452(.A(KEYINPUT21), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(G231gat), .A2(G233gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(new_n420), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n232), .B1(new_n654), .B2(new_n653), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n658), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g459(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(KEYINPUT98), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(G155gat), .ZN(new_n663));
  XOR2_X1   g462(.A(G183gat), .B(G211gat), .Z(new_n664));
  XNOR2_X1  g463(.A(new_n663), .B(new_n664), .ZN(new_n665));
  OR2_X1    g464(.A1(new_n660), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n660), .A2(new_n665), .ZN(new_n667));
  AND2_X1   g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT104), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n645), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n636), .A2(new_n644), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n666), .A2(new_n667), .ZN(new_n672));
  OAI21_X1  g471(.A(KEYINPUT104), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(G230gat), .A2(G233gat), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n651), .B(new_n652), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n622), .A2(KEYINPUT10), .A3(new_n676), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n677), .A2(KEYINPUT105), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n620), .A2(new_n653), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT10), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n622), .A2(new_n676), .ZN(new_n682));
  AND3_X1   g481(.A1(new_n680), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n677), .A2(KEYINPUT105), .ZN(new_n684));
  OAI211_X1 g483(.A(new_n675), .B(new_n679), .C1(new_n683), .C2(new_n684), .ZN(new_n685));
  AND2_X1   g484(.A1(new_n680), .A2(new_n682), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n685), .B1(new_n675), .B2(new_n686), .ZN(new_n687));
  XNOR2_X1  g486(.A(G120gat), .B(G148gat), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(KEYINPUT106), .ZN(new_n689));
  XOR2_X1   g488(.A(G176gat), .B(G204gat), .Z(new_n690));
  XNOR2_X1  g489(.A(new_n689), .B(new_n690), .ZN(new_n691));
  OR2_X1    g490(.A1(new_n687), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n687), .A2(new_n691), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n674), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n611), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n696), .A2(new_n531), .ZN(new_n697));
  XOR2_X1   g496(.A(new_n697), .B(G1gat), .Z(G1324gat));
  NOR2_X1   g497(.A1(new_n696), .A2(new_n557), .ZN(new_n699));
  XOR2_X1   g498(.A(KEYINPUT16), .B(G8gat), .Z(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n701), .B1(new_n231), .B2(new_n699), .ZN(new_n702));
  MUX2_X1   g501(.A(new_n701), .B(new_n702), .S(KEYINPUT42), .Z(G1325gat));
  OAI21_X1  g502(.A(G15gat), .B1(new_n696), .B2(new_n609), .ZN(new_n704));
  AND2_X1   g503(.A1(new_n579), .A2(new_n580), .ZN(new_n705));
  OR2_X1    g504(.A1(new_n705), .A2(G15gat), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n704), .B1(new_n696), .B2(new_n706), .ZN(G1326gat));
  NOR2_X1   g506(.A1(new_n696), .A2(new_n366), .ZN(new_n708));
  XOR2_X1   g507(.A(KEYINPUT43), .B(G22gat), .Z(new_n709));
  XNOR2_X1  g508(.A(new_n708), .B(new_n709), .ZN(G1327gat));
  INV_X1    g509(.A(G29gat), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT109), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT35), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n564), .A2(new_n607), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n556), .B1(new_n526), .B2(new_n530), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n713), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NOR3_X1   g515(.A1(new_n566), .A2(new_n567), .A3(KEYINPUT86), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n569), .B1(new_n527), .B2(new_n529), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n526), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(new_n574), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n366), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  OAI21_X1  g520(.A(KEYINPUT89), .B1(new_n721), .B2(new_n705), .ZN(new_n722));
  NAND4_X1  g521(.A1(new_n581), .A2(new_n584), .A3(new_n560), .A4(new_n366), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n716), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  AND3_X1   g523(.A1(new_n605), .A2(new_n606), .A3(new_n609), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n671), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n606), .A2(KEYINPUT107), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT107), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n558), .A2(new_n564), .A3(new_n728), .ZN(new_n729));
  NAND4_X1  g528(.A1(new_n727), .A2(new_n609), .A3(new_n605), .A4(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n586), .A2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT108), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n636), .A2(new_n644), .A3(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(new_n733), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n732), .B1(new_n636), .B2(new_n644), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT44), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(new_n738), .ZN(new_n739));
  AOI22_X1  g538(.A1(KEYINPUT44), .A2(new_n726), .B1(new_n731), .B2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(new_n694), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n672), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n262), .A2(new_n263), .ZN(new_n743));
  INV_X1    g542(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(new_n745), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n712), .B1(new_n740), .B2(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(new_n531), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n586), .A2(new_n610), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n737), .B1(new_n749), .B2(new_n671), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n738), .B1(new_n586), .B2(new_n730), .ZN(new_n751));
  OAI211_X1 g550(.A(KEYINPUT109), .B(new_n745), .C1(new_n750), .C2(new_n751), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n747), .A2(new_n748), .A3(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT110), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n711), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n755), .B1(new_n754), .B2(new_n753), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n742), .A2(new_n645), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n611), .A2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(new_n758), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n759), .A2(new_n711), .A3(new_n748), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(KEYINPUT45), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n756), .A2(new_n761), .ZN(G1328gat));
  NAND3_X1  g561(.A1(new_n747), .A2(new_n556), .A3(new_n752), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(G36gat), .ZN(new_n764));
  NOR3_X1   g563(.A1(new_n758), .A2(G36gat), .A3(new_n557), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(KEYINPUT46), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n764), .A2(new_n766), .ZN(G1329gat));
  NOR3_X1   g566(.A1(new_n758), .A2(G43gat), .A3(new_n705), .ZN(new_n768));
  INV_X1    g567(.A(new_n768), .ZN(new_n769));
  NOR3_X1   g568(.A1(new_n740), .A2(new_n609), .A3(new_n746), .ZN(new_n770));
  INV_X1    g569(.A(G43gat), .ZN(new_n771));
  OAI211_X1 g570(.A(new_n769), .B(KEYINPUT47), .C1(new_n770), .C2(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(new_n609), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n747), .A2(new_n773), .A3(new_n752), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(G43gat), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(new_n769), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT47), .ZN(new_n777));
  AOI21_X1  g576(.A(KEYINPUT111), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n768), .B1(new_n774), .B2(G43gat), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT111), .ZN(new_n780));
  NOR3_X1   g579(.A1(new_n779), .A2(new_n780), .A3(KEYINPUT47), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n772), .B1(new_n778), .B2(new_n781), .ZN(G1330gat));
  INV_X1    g581(.A(KEYINPUT112), .ZN(new_n783));
  OR2_X1    g582(.A1(new_n783), .A2(KEYINPUT48), .ZN(new_n784));
  OR2_X1    g583(.A1(new_n366), .A2(G50gat), .ZN(new_n785));
  NOR3_X1   g584(.A1(new_n740), .A2(new_n366), .A3(new_n746), .ZN(new_n786));
  NAND2_X1  g585(.A1(KEYINPUT48), .A2(G50gat), .ZN(new_n787));
  OAI221_X1 g586(.A(new_n784), .B1(new_n758), .B2(new_n785), .C1(new_n786), .C2(new_n787), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n758), .A2(new_n783), .A3(new_n785), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n747), .A2(new_n564), .A3(new_n752), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n789), .B1(new_n790), .B2(G50gat), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n788), .B1(new_n791), .B2(KEYINPUT48), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT113), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  OAI211_X1 g593(.A(new_n788), .B(KEYINPUT113), .C1(new_n791), .C2(KEYINPUT48), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(G1331gat));
  INV_X1    g595(.A(new_n674), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n731), .A2(new_n744), .A3(new_n797), .A4(new_n694), .ZN(new_n798));
  INV_X1    g597(.A(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(new_n748), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n800), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g600(.A1(new_n799), .A2(new_n556), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n802), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n803));
  XOR2_X1   g602(.A(KEYINPUT49), .B(G64gat), .Z(new_n804));
  OAI21_X1  g603(.A(new_n803), .B1(new_n802), .B2(new_n804), .ZN(G1333gat));
  OAI21_X1  g604(.A(G71gat), .B1(new_n798), .B2(new_n609), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n581), .A2(new_n648), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n806), .B1(new_n798), .B2(new_n807), .ZN(new_n808));
  XOR2_X1   g607(.A(new_n808), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g608(.A1(new_n799), .A2(new_n564), .ZN(new_n810));
  XNOR2_X1  g609(.A(new_n810), .B(G78gat), .ZN(G1335gat));
  INV_X1    g610(.A(new_n740), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n668), .A2(new_n743), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n812), .A2(new_n694), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(KEYINPUT114), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT114), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n812), .A2(new_n816), .A3(new_n694), .A4(new_n813), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n617), .B1(new_n818), .B2(new_n531), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n731), .A2(new_n671), .A3(new_n813), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT51), .ZN(new_n821));
  OR2_X1    g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(new_n822), .ZN(new_n823));
  AND2_X1   g622(.A1(new_n820), .A2(new_n821), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n694), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  OR2_X1    g624(.A1(new_n531), .A2(new_n617), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n819), .B1(new_n825), .B2(new_n826), .ZN(G1336gat));
  OAI21_X1  g626(.A(G92gat), .B1(new_n814), .B2(new_n557), .ZN(new_n828));
  XOR2_X1   g627(.A(KEYINPUT115), .B(KEYINPUT52), .Z(new_n829));
  OR2_X1    g628(.A1(new_n557), .A2(G92gat), .ZN(new_n830));
  OAI211_X1 g629(.A(new_n828), .B(new_n829), .C1(new_n825), .C2(new_n830), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n825), .A2(new_n830), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n815), .A2(new_n556), .A3(new_n817), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n832), .B1(G92gat), .B2(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT52), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n831), .B1(new_n834), .B2(new_n835), .ZN(G1337gat));
  OAI21_X1  g635(.A(G99gat), .B1(new_n818), .B2(new_n609), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n581), .A2(new_n614), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n837), .B1(new_n825), .B2(new_n838), .ZN(G1338gat));
  OAI21_X1  g638(.A(G106gat), .B1(new_n814), .B2(new_n366), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT53), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n564), .A2(new_n615), .ZN(new_n842));
  OAI211_X1 g641(.A(new_n840), .B(new_n841), .C1(new_n825), .C2(new_n842), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n825), .A2(new_n842), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n815), .A2(new_n564), .A3(new_n817), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n844), .B1(G106gat), .B2(new_n845), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n843), .B1(new_n846), .B2(new_n841), .ZN(G1339gat));
  INV_X1    g646(.A(new_n735), .ZN(new_n848));
  INV_X1    g647(.A(new_n684), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n680), .A2(new_n681), .A3(new_n682), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n678), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT54), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n851), .A2(new_n852), .A3(new_n675), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n685), .A2(KEYINPUT54), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n851), .A2(new_n675), .ZN(new_n855));
  OAI211_X1 g654(.A(new_n691), .B(new_n853), .C1(new_n854), .C2(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT55), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n692), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(KEYINPUT116), .ZN(new_n859));
  AND2_X1   g658(.A1(new_n853), .A2(new_n691), .ZN(new_n860));
  OAI211_X1 g659(.A(new_n860), .B(KEYINPUT55), .C1(new_n855), .C2(new_n854), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT116), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n861), .A2(new_n862), .A3(new_n692), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n856), .A2(new_n857), .ZN(new_n864));
  NAND4_X1  g663(.A1(new_n743), .A2(new_n859), .A3(new_n863), .A4(new_n864), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n248), .A2(new_n203), .ZN(new_n866));
  NOR3_X1   g665(.A1(new_n234), .A2(new_n235), .A3(new_n204), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n254), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  AND2_X1   g667(.A1(new_n263), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(new_n694), .ZN(new_n870));
  AOI22_X1  g669(.A1(new_n848), .A2(new_n733), .B1(new_n865), .B2(new_n870), .ZN(new_n871));
  NAND4_X1  g670(.A1(new_n859), .A2(new_n869), .A3(new_n863), .A4(new_n864), .ZN(new_n872));
  NOR3_X1   g671(.A1(new_n872), .A2(new_n734), .A3(new_n735), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n672), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n670), .A2(new_n673), .A3(new_n744), .A4(new_n741), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n531), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n464), .A2(new_n556), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(new_n878), .ZN(new_n879));
  AOI21_X1  g678(.A(G113gat), .B1(new_n879), .B2(new_n743), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n874), .A2(new_n875), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n705), .A2(new_n564), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n748), .A2(new_n557), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n265), .A2(new_n427), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n880), .B1(new_n885), .B2(new_n886), .ZN(G1340gat));
  AOI21_X1  g686(.A(G120gat), .B1(new_n879), .B2(new_n694), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n741), .A2(new_n425), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n888), .B1(new_n885), .B2(new_n889), .ZN(G1341gat));
  INV_X1    g689(.A(new_n885), .ZN(new_n891));
  OAI21_X1  g690(.A(G127gat), .B1(new_n891), .B2(new_n672), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n879), .A2(new_n420), .A3(new_n668), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(G1342gat));
  NOR3_X1   g693(.A1(new_n878), .A2(G134gat), .A3(new_n645), .ZN(new_n895));
  INV_X1    g694(.A(new_n895), .ZN(new_n896));
  OR2_X1    g695(.A1(new_n896), .A2(KEYINPUT56), .ZN(new_n897));
  OAI21_X1  g696(.A(G134gat), .B1(new_n891), .B2(new_n645), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n896), .A2(KEYINPUT56), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n897), .A2(new_n898), .A3(new_n899), .ZN(G1343gat));
  NOR2_X1   g699(.A1(new_n773), .A2(new_n884), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT57), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n366), .A2(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(new_n903), .ZN(new_n904));
  INV_X1    g703(.A(new_n875), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n861), .A2(new_n864), .A3(new_n692), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n258), .B1(new_n256), .B2(new_n257), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n262), .A2(KEYINPUT97), .A3(new_n263), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n906), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  INV_X1    g708(.A(new_n870), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n645), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  AND3_X1   g710(.A1(new_n859), .A2(new_n863), .A3(new_n864), .ZN(new_n912));
  NAND4_X1  g711(.A1(new_n912), .A2(new_n848), .A3(new_n733), .A4(new_n869), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n668), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT117), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n905), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  INV_X1    g715(.A(new_n906), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n917), .B1(new_n259), .B2(new_n264), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n671), .B1(new_n918), .B2(new_n870), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n672), .B1(new_n919), .B2(new_n873), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(KEYINPUT117), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n904), .B1(new_n916), .B2(new_n921), .ZN(new_n922));
  AOI21_X1  g721(.A(KEYINPUT57), .B1(new_n881), .B2(new_n564), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n901), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  OAI21_X1  g723(.A(G141gat), .B1(new_n924), .B2(new_n265), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT58), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n299), .B1(new_n259), .B2(new_n264), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n773), .A2(new_n366), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n876), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n929), .A2(KEYINPUT119), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT119), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n876), .A2(new_n931), .A3(new_n928), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n930), .A2(new_n557), .A3(new_n932), .ZN(new_n933));
  OAI211_X1 g732(.A(new_n925), .B(new_n926), .C1(new_n927), .C2(new_n933), .ZN(new_n934));
  OAI211_X1 g733(.A(new_n743), .B(new_n901), .C1(new_n922), .C2(new_n923), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT118), .ZN(new_n936));
  AND3_X1   g735(.A1(new_n935), .A2(new_n936), .A3(G141gat), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n936), .B1(new_n935), .B2(G141gat), .ZN(new_n938));
  NOR3_X1   g737(.A1(new_n929), .A2(new_n556), .A3(new_n927), .ZN(new_n939));
  NOR3_X1   g738(.A1(new_n937), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n934), .B1(new_n940), .B2(new_n926), .ZN(G1344gat));
  NAND2_X1  g740(.A1(new_n695), .A2(new_n265), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n872), .A2(new_n645), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n672), .B1(new_n919), .B2(new_n943), .ZN(new_n944));
  AND2_X1   g743(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  OAI211_X1 g744(.A(KEYINPUT120), .B(new_n902), .C1(new_n945), .C2(new_n366), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT120), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n366), .B1(new_n942), .B2(new_n944), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n947), .B1(new_n948), .B2(KEYINPUT57), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n881), .A2(new_n903), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n946), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n951), .A2(new_n694), .A3(new_n901), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n952), .A2(KEYINPUT59), .A3(G148gat), .ZN(new_n953));
  OAI21_X1  g752(.A(KEYINPUT59), .B1(new_n933), .B2(new_n741), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n954), .A2(new_n301), .ZN(new_n955));
  OR3_X1    g754(.A1(new_n924), .A2(KEYINPUT59), .A3(new_n741), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n953), .A2(new_n955), .A3(new_n956), .ZN(G1345gat));
  OR2_X1    g756(.A1(new_n933), .A2(new_n672), .ZN(new_n958));
  INV_X1    g757(.A(new_n924), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n668), .A2(G155gat), .ZN(new_n960));
  XNOR2_X1  g759(.A(new_n960), .B(KEYINPUT121), .ZN(new_n961));
  AOI22_X1  g760(.A1(new_n958), .A2(new_n305), .B1(new_n959), .B2(new_n961), .ZN(G1346gat));
  NAND3_X1  g761(.A1(new_n959), .A2(G162gat), .A3(new_n736), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n306), .B1(new_n933), .B2(new_n645), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT122), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n963), .A2(new_n964), .A3(KEYINPUT122), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n967), .A2(new_n968), .ZN(G1347gat));
  INV_X1    g768(.A(new_n883), .ZN(new_n970));
  NOR2_X1   g769(.A1(new_n748), .A2(new_n557), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NOR3_X1   g771(.A1(new_n972), .A2(new_n382), .A3(new_n265), .ZN(new_n973));
  AOI21_X1  g772(.A(new_n748), .B1(new_n874), .B2(new_n875), .ZN(new_n974));
  XNOR2_X1  g773(.A(new_n974), .B(KEYINPUT123), .ZN(new_n975));
  NOR2_X1   g774(.A1(new_n464), .A2(new_n557), .ZN(new_n976));
  AND2_X1   g775(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n977), .A2(new_n743), .ZN(new_n978));
  AOI21_X1  g777(.A(new_n973), .B1(new_n978), .B2(new_n382), .ZN(G1348gat));
  NAND3_X1  g778(.A1(new_n977), .A2(new_n383), .A3(new_n694), .ZN(new_n980));
  OAI21_X1  g779(.A(G176gat), .B1(new_n972), .B2(new_n741), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n980), .A2(new_n981), .ZN(G1349gat));
  NAND4_X1  g781(.A1(new_n975), .A2(new_n367), .A3(new_n668), .A4(new_n976), .ZN(new_n983));
  INV_X1    g782(.A(KEYINPUT124), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n984), .A2(KEYINPUT60), .ZN(new_n985));
  OAI21_X1  g784(.A(G183gat), .B1(new_n972), .B2(new_n672), .ZN(new_n986));
  NAND3_X1  g785(.A1(new_n983), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  OR2_X1    g786(.A1(new_n984), .A2(KEYINPUT60), .ZN(new_n988));
  XNOR2_X1  g787(.A(new_n987), .B(new_n988), .ZN(G1350gat));
  NAND3_X1  g788(.A1(new_n977), .A2(new_n368), .A3(new_n736), .ZN(new_n990));
  INV_X1    g789(.A(KEYINPUT125), .ZN(new_n991));
  NAND3_X1  g790(.A1(new_n970), .A2(new_n671), .A3(new_n971), .ZN(new_n992));
  INV_X1    g791(.A(KEYINPUT61), .ZN(new_n993));
  AND4_X1   g792(.A1(new_n991), .A2(new_n992), .A3(new_n993), .A4(G190gat), .ZN(new_n994));
  AOI21_X1  g793(.A(new_n368), .B1(KEYINPUT125), .B2(KEYINPUT61), .ZN(new_n995));
  AOI22_X1  g794(.A1(new_n992), .A2(new_n995), .B1(new_n991), .B2(new_n993), .ZN(new_n996));
  OAI21_X1  g795(.A(new_n990), .B1(new_n994), .B2(new_n996), .ZN(G1351gat));
  NOR3_X1   g796(.A1(new_n773), .A2(new_n557), .A3(new_n366), .ZN(new_n998));
  AND2_X1   g797(.A1(new_n975), .A2(new_n998), .ZN(new_n999));
  AOI21_X1  g798(.A(G197gat), .B1(new_n999), .B2(new_n743), .ZN(new_n1000));
  AND2_X1   g799(.A1(new_n609), .A2(new_n971), .ZN(new_n1001));
  AND2_X1   g800(.A1(new_n951), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g801(.A(G197gat), .ZN(new_n1003));
  NOR2_X1   g802(.A1(new_n265), .A2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g803(.A(new_n1000), .B1(new_n1002), .B2(new_n1004), .ZN(G1352gat));
  NAND3_X1  g804(.A1(new_n951), .A2(new_n694), .A3(new_n1001), .ZN(new_n1006));
  INV_X1    g805(.A(KEYINPUT127), .ZN(new_n1007));
  NAND2_X1  g806(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND4_X1  g807(.A1(new_n951), .A2(KEYINPUT127), .A3(new_n694), .A4(new_n1001), .ZN(new_n1009));
  NAND3_X1  g808(.A1(new_n1008), .A2(G204gat), .A3(new_n1009), .ZN(new_n1010));
  NOR2_X1   g809(.A1(new_n741), .A2(G204gat), .ZN(new_n1011));
  NAND3_X1  g810(.A1(new_n975), .A2(new_n998), .A3(new_n1011), .ZN(new_n1012));
  XOR2_X1   g811(.A(KEYINPUT126), .B(KEYINPUT62), .Z(new_n1013));
  XNOR2_X1  g812(.A(new_n1012), .B(new_n1013), .ZN(new_n1014));
  NAND2_X1  g813(.A1(new_n1010), .A2(new_n1014), .ZN(G1353gat));
  INV_X1    g814(.A(G211gat), .ZN(new_n1016));
  NAND3_X1  g815(.A1(new_n999), .A2(new_n1016), .A3(new_n668), .ZN(new_n1017));
  NAND3_X1  g816(.A1(new_n951), .A2(new_n668), .A3(new_n1001), .ZN(new_n1018));
  AND3_X1   g817(.A1(new_n1018), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1019));
  AOI21_X1  g818(.A(KEYINPUT63), .B1(new_n1018), .B2(G211gat), .ZN(new_n1020));
  OAI21_X1  g819(.A(new_n1017), .B1(new_n1019), .B2(new_n1020), .ZN(G1354gat));
  NAND2_X1  g820(.A1(new_n1002), .A2(new_n671), .ZN(new_n1022));
  NAND2_X1  g821(.A1(new_n1022), .A2(G218gat), .ZN(new_n1023));
  INV_X1    g822(.A(G218gat), .ZN(new_n1024));
  NAND3_X1  g823(.A1(new_n999), .A2(new_n1024), .A3(new_n736), .ZN(new_n1025));
  NAND2_X1  g824(.A1(new_n1023), .A2(new_n1025), .ZN(G1355gat));
endmodule


