//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 1 0 0 1 1 0 0 0 1 1 0 1 0 1 1 0 0 1 1 1 0 1 1 0 1 1 0 1 0 0 0 1 1 1 0 0 0 0 0 0 0 1 0 1 1 0 0 0 0 1 0 0 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:53 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n788, new_n790,
    new_n791, new_n792, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n810, new_n811, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n825, new_n826, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1004, new_n1005, new_n1006, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1061, new_n1062, new_n1063, new_n1064, new_n1065, new_n1066,
    new_n1067, new_n1068, new_n1069, new_n1070, new_n1071, new_n1072,
    new_n1073, new_n1074, new_n1075, new_n1076, new_n1077, new_n1078,
    new_n1079, new_n1080, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1091,
    new_n1092, new_n1093, new_n1094, new_n1095, new_n1096, new_n1097,
    new_n1098, new_n1099, new_n1100, new_n1101, new_n1102, new_n1103,
    new_n1104, new_n1105;
  XNOR2_X1  g000(.A(G110), .B(G140), .ZN(new_n187));
  XNOR2_X1  g001(.A(new_n187), .B(KEYINPUT80), .ZN(new_n188));
  INV_X1    g002(.A(G227), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n189), .A2(G953), .ZN(new_n190));
  XOR2_X1   g004(.A(new_n188), .B(new_n190), .Z(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT11), .ZN(new_n193));
  INV_X1    g007(.A(G134), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n193), .B1(new_n194), .B2(G137), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(G137), .ZN(new_n196));
  INV_X1    g010(.A(G137), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n197), .A2(KEYINPUT11), .A3(G134), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n195), .A2(new_n196), .A3(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G131), .ZN(new_n200));
  INV_X1    g014(.A(G131), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n195), .A2(new_n198), .A3(new_n201), .A4(new_n196), .ZN(new_n202));
  AND2_X1   g016(.A1(new_n200), .A2(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(KEYINPUT0), .A2(G128), .ZN(new_n204));
  NOR2_X1   g018(.A1(KEYINPUT0), .A2(G128), .ZN(new_n205));
  INV_X1    g019(.A(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G143), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n207), .A2(G146), .ZN(new_n208));
  INV_X1    g022(.A(G146), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n209), .A2(G143), .ZN(new_n210));
  OAI211_X1 g024(.A(new_n204), .B(new_n206), .C1(new_n208), .C2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n209), .A2(G143), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n207), .A2(G146), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n212), .A2(new_n213), .A3(KEYINPUT0), .A4(G128), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n211), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G101), .ZN(new_n216));
  INV_X1    g030(.A(G107), .ZN(new_n217));
  OAI21_X1  g031(.A(KEYINPUT81), .B1(new_n217), .B2(G104), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT81), .ZN(new_n219));
  INV_X1    g033(.A(G104), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n219), .A2(new_n220), .A3(G107), .ZN(new_n221));
  AND2_X1   g035(.A1(new_n218), .A2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n223), .B1(new_n220), .B2(G107), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n217), .A2(KEYINPUT3), .A3(G104), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n216), .B1(new_n222), .B2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT4), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n215), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  AND2_X1   g043(.A1(new_n224), .A2(new_n225), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n218), .A2(new_n221), .ZN(new_n231));
  OAI21_X1  g045(.A(G101), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  NAND4_X1  g046(.A1(new_n226), .A2(new_n216), .A3(new_n218), .A4(new_n221), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n232), .A2(KEYINPUT4), .A3(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT10), .ZN(new_n235));
  INV_X1    g049(.A(G128), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n236), .A2(KEYINPUT1), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n237), .A2(new_n212), .A3(new_n213), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n236), .B1(new_n212), .B2(KEYINPUT1), .ZN(new_n239));
  XNOR2_X1  g053(.A(G143), .B(G146), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n238), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n220), .A2(G107), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n217), .A2(G104), .ZN(new_n243));
  OAI21_X1  g057(.A(G101), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n241), .A2(new_n233), .A3(new_n244), .ZN(new_n245));
  AOI22_X1  g059(.A1(new_n229), .A2(new_n234), .B1(new_n235), .B2(new_n245), .ZN(new_n246));
  AND2_X1   g060(.A1(new_n233), .A2(new_n244), .ZN(new_n247));
  INV_X1    g061(.A(new_n240), .ZN(new_n248));
  OAI211_X1 g062(.A(KEYINPUT65), .B(KEYINPUT1), .C1(new_n207), .C2(G146), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G128), .ZN(new_n250));
  AOI21_X1  g064(.A(KEYINPUT65), .B1(new_n212), .B2(KEYINPUT1), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n248), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(new_n238), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n247), .A2(KEYINPUT10), .A3(new_n253), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n203), .B1(new_n246), .B2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(new_n215), .ZN(new_n256));
  OAI211_X1 g070(.A(new_n228), .B(G101), .C1(new_n230), .C2(new_n231), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n233), .A2(KEYINPUT4), .ZN(new_n258));
  OAI211_X1 g072(.A(new_n256), .B(new_n257), .C1(new_n258), .C2(new_n227), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n245), .A2(new_n235), .ZN(new_n260));
  AND4_X1   g074(.A1(new_n203), .A2(new_n254), .A3(new_n259), .A4(new_n260), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n192), .B1(new_n255), .B2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT83), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n261), .A2(new_n192), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n233), .A2(new_n244), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n266), .A2(new_n238), .A3(new_n252), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n267), .A2(KEYINPUT82), .A3(new_n245), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n200), .A2(new_n202), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n270), .B1(new_n267), .B2(KEYINPUT82), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT12), .ZN(new_n272));
  NOR3_X1   g086(.A1(new_n269), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n247), .A2(new_n253), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT82), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n203), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  AOI21_X1  g090(.A(KEYINPUT12), .B1(new_n276), .B2(new_n268), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n265), .B1(new_n273), .B2(new_n277), .ZN(new_n278));
  OAI211_X1 g092(.A(KEYINPUT83), .B(new_n192), .C1(new_n255), .C2(new_n261), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n264), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(G469), .ZN(new_n281));
  INV_X1    g095(.A(G902), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n280), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n255), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n265), .A2(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n272), .B1(new_n269), .B2(new_n271), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n276), .A2(KEYINPUT12), .A3(new_n268), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n261), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  OAI211_X1 g102(.A(new_n285), .B(G469), .C1(new_n288), .C2(new_n191), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n281), .A2(new_n282), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n283), .A2(new_n289), .A3(new_n291), .ZN(new_n292));
  XNOR2_X1  g106(.A(KEYINPUT9), .B(G234), .ZN(new_n293));
  OAI21_X1  g107(.A(G221), .B1(new_n293), .B2(G902), .ZN(new_n294));
  AND2_X1   g108(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  OAI21_X1  g109(.A(G214), .B1(G237), .B2(G902), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  OAI21_X1  g111(.A(G210), .B1(G237), .B2(G902), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(G119), .ZN(new_n300));
  OAI21_X1  g114(.A(KEYINPUT69), .B1(new_n300), .B2(G116), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT69), .ZN(new_n302));
  INV_X1    g116(.A(G116), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n302), .A2(new_n303), .A3(G119), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n301), .A2(new_n304), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n303), .A2(G119), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT2), .ZN(new_n309));
  INV_X1    g123(.A(G113), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n309), .A2(new_n310), .A3(KEYINPUT67), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT67), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n312), .B1(KEYINPUT2), .B2(G113), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(KEYINPUT2), .A2(G113), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(KEYINPUT68), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT68), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n317), .A2(KEYINPUT2), .A3(G113), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n314), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n308), .A2(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n306), .B1(new_n301), .B2(new_n304), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n322), .A2(new_n314), .A3(new_n319), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n234), .A2(new_n324), .A3(new_n257), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT84), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n305), .A2(KEYINPUT5), .A3(new_n307), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT5), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n310), .B1(new_n306), .B2(new_n328), .ZN(new_n329));
  AOI22_X1  g143(.A1(new_n313), .A2(new_n311), .B1(new_n316), .B2(new_n318), .ZN(new_n330));
  AOI22_X1  g144(.A1(new_n327), .A2(new_n329), .B1(new_n330), .B2(new_n322), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n247), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n325), .A2(new_n326), .A3(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n326), .B1(new_n325), .B2(new_n332), .ZN(new_n335));
  XNOR2_X1  g149(.A(G110), .B(G122), .ZN(new_n336));
  NOR4_X1   g150(.A1(new_n334), .A2(new_n335), .A3(KEYINPUT6), .A4(new_n336), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n308), .A2(new_n320), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n330), .A2(new_n322), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n257), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n258), .A2(new_n227), .ZN(new_n341));
  OAI211_X1 g155(.A(new_n332), .B(new_n336), .C1(new_n340), .C2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(KEYINPUT6), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n325), .A2(new_n332), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n336), .B1(new_n344), .B2(KEYINPUT84), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n343), .B1(new_n345), .B2(new_n333), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n215), .A2(G125), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n347), .B1(new_n253), .B2(G125), .ZN(new_n348));
  INV_X1    g162(.A(G224), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n349), .A2(G953), .ZN(new_n350));
  XNOR2_X1  g164(.A(new_n350), .B(KEYINPUT85), .ZN(new_n351));
  XNOR2_X1  g165(.A(new_n348), .B(new_n351), .ZN(new_n352));
  NOR3_X1   g166(.A1(new_n337), .A2(new_n346), .A3(new_n352), .ZN(new_n353));
  AND3_X1   g167(.A1(new_n233), .A2(KEYINPUT86), .A3(new_n244), .ZN(new_n354));
  AOI211_X1 g168(.A(new_n328), .B(new_n306), .C1(new_n304), .C2(new_n301), .ZN(new_n355));
  INV_X1    g169(.A(new_n329), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n323), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n354), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n233), .A2(KEYINPUT86), .A3(new_n244), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n331), .A2(new_n359), .ZN(new_n360));
  XNOR2_X1  g174(.A(new_n336), .B(KEYINPUT8), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n358), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  OAI21_X1  g176(.A(KEYINPUT7), .B1(new_n349), .B2(G953), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n348), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(new_n363), .ZN(new_n365));
  OAI211_X1 g179(.A(new_n347), .B(new_n365), .C1(new_n253), .C2(G125), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n342), .A2(new_n362), .A3(new_n364), .A4(new_n366), .ZN(new_n367));
  AND3_X1   g181(.A1(new_n367), .A2(KEYINPUT87), .A3(new_n282), .ZN(new_n368));
  AOI21_X1  g182(.A(KEYINPUT87), .B1(new_n367), .B2(new_n282), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n299), .B1(new_n353), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n367), .A2(new_n282), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT87), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n367), .A2(KEYINPUT87), .A3(new_n282), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT6), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n345), .A2(new_n377), .A3(new_n333), .ZN(new_n378));
  INV_X1    g192(.A(new_n352), .ZN(new_n379));
  NOR3_X1   g193(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n380));
  OAI211_X1 g194(.A(new_n378), .B(new_n379), .C1(new_n380), .C2(new_n343), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n376), .A2(new_n298), .A3(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n297), .B1(new_n371), .B2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(G237), .ZN(new_n384));
  INV_X1    g198(.A(G953), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n384), .A2(new_n385), .A3(G214), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(new_n207), .ZN(new_n387));
  NOR2_X1   g201(.A1(G237), .A2(G953), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n388), .A2(G143), .A3(G214), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g204(.A(KEYINPUT90), .B1(new_n390), .B2(G131), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT90), .ZN(new_n392));
  AOI211_X1 g206(.A(new_n392), .B(new_n201), .C1(new_n387), .C2(new_n389), .ZN(new_n393));
  OAI21_X1  g207(.A(KEYINPUT17), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  AND4_X1   g208(.A1(G143), .A2(new_n384), .A3(new_n385), .A4(G214), .ZN(new_n395));
  AOI21_X1  g209(.A(G143), .B1(new_n388), .B2(G214), .ZN(new_n396));
  OAI21_X1  g210(.A(G131), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(new_n392), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT17), .ZN(new_n399));
  OAI211_X1 g213(.A(KEYINPUT90), .B(G131), .C1(new_n395), .C2(new_n396), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n387), .A2(new_n201), .A3(new_n389), .ZN(new_n401));
  NAND4_X1  g215(.A1(new_n398), .A2(new_n399), .A3(new_n400), .A4(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT78), .ZN(new_n403));
  INV_X1    g217(.A(G140), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(G125), .ZN(new_n405));
  INV_X1    g219(.A(G125), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(G140), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n405), .A2(new_n407), .A3(KEYINPUT16), .ZN(new_n408));
  OR3_X1    g222(.A1(new_n406), .A2(KEYINPUT16), .A3(G140), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n403), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NOR3_X1   g224(.A1(new_n406), .A2(KEYINPUT16), .A3(G140), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n411), .A2(KEYINPUT78), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n209), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n409), .A2(new_n403), .ZN(new_n414));
  XNOR2_X1  g228(.A(G125), .B(G140), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n411), .B1(new_n415), .B2(KEYINPUT16), .ZN(new_n416));
  OAI211_X1 g230(.A(G146), .B(new_n414), .C1(new_n416), .C2(new_n403), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n394), .A2(new_n402), .A3(new_n413), .A4(new_n417), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n390), .A2(KEYINPUT88), .A3(KEYINPUT18), .A4(G131), .ZN(new_n419));
  NAND3_X1  g233(.A1(KEYINPUT88), .A2(KEYINPUT18), .A3(G131), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n387), .A2(new_n389), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n405), .A2(new_n407), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(G146), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n415), .A2(new_n209), .ZN(new_n424));
  AND3_X1   g238(.A1(new_n423), .A2(new_n424), .A3(KEYINPUT89), .ZN(new_n425));
  AOI21_X1  g239(.A(KEYINPUT89), .B1(new_n423), .B2(new_n424), .ZN(new_n426));
  OAI211_X1 g240(.A(new_n419), .B(new_n421), .C1(new_n425), .C2(new_n426), .ZN(new_n427));
  XOR2_X1   g241(.A(KEYINPUT92), .B(G104), .Z(new_n428));
  XNOR2_X1  g242(.A(G113), .B(G122), .ZN(new_n429));
  XNOR2_X1  g243(.A(new_n428), .B(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n418), .A2(new_n427), .A3(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n431), .B1(new_n418), .B2(new_n427), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n282), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(G475), .ZN(new_n436));
  AND3_X1   g250(.A1(new_n398), .A2(new_n400), .A3(new_n401), .ZN(new_n437));
  AND3_X1   g251(.A1(new_n405), .A2(new_n407), .A3(KEYINPUT19), .ZN(new_n438));
  AOI21_X1  g252(.A(KEYINPUT19), .B1(new_n405), .B2(new_n407), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n209), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT91), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  OAI211_X1 g256(.A(KEYINPUT91), .B(new_n209), .C1(new_n438), .C2(new_n439), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n442), .A2(new_n417), .A3(new_n443), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n427), .B1(new_n437), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(new_n430), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(new_n432), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT20), .ZN(new_n448));
  NOR2_X1   g262(.A1(G475), .A2(G902), .ZN(new_n449));
  NAND4_X1  g263(.A1(new_n447), .A2(KEYINPUT93), .A3(new_n448), .A4(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(new_n449), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n451), .B1(new_n446), .B2(new_n432), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n450), .B1(new_n448), .B2(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(KEYINPUT93), .B1(new_n452), .B2(new_n448), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n436), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  AND2_X1   g269(.A1(new_n385), .A2(G952), .ZN(new_n456));
  NAND2_X1  g270(.A1(G234), .A2(G237), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  XNOR2_X1  g273(.A(KEYINPUT21), .B(G898), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n457), .A2(G902), .A3(G953), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n459), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(G478), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT15), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n464), .B1(KEYINPUT95), .B2(new_n465), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n466), .B1(KEYINPUT95), .B2(new_n465), .ZN(new_n467));
  INV_X1    g281(.A(G217), .ZN(new_n468));
  NOR3_X1   g282(.A1(new_n293), .A2(new_n468), .A3(G953), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n303), .A2(KEYINPUT14), .A3(G122), .ZN(new_n471));
  INV_X1    g285(.A(G122), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(G116), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n303), .A2(G122), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  OAI211_X1 g289(.A(G107), .B(new_n471), .C1(new_n475), .C2(KEYINPUT14), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n473), .A2(new_n474), .A3(new_n217), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n207), .A2(G128), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n236), .A2(G143), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n478), .A2(new_n479), .A3(new_n194), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n194), .B1(new_n478), .B2(new_n479), .ZN(new_n482));
  OAI211_X1 g296(.A(new_n476), .B(new_n477), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT13), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n484), .B1(new_n236), .B2(G143), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n207), .A2(KEYINPUT13), .A3(G128), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n485), .A2(new_n486), .A3(new_n479), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(G134), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n217), .B1(new_n473), .B2(new_n474), .ZN(new_n489));
  INV_X1    g303(.A(new_n477), .ZN(new_n490));
  OAI211_X1 g304(.A(new_n488), .B(new_n480), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT94), .ZN(new_n492));
  AND3_X1   g306(.A1(new_n483), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n492), .B1(new_n483), .B2(new_n491), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n470), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n483), .A2(new_n491), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(KEYINPUT94), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n483), .A2(new_n491), .A3(new_n492), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n497), .A2(new_n469), .A3(new_n498), .ZN(new_n499));
  AOI21_X1  g313(.A(G902), .B1(new_n495), .B2(new_n499), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n500), .A2(KEYINPUT96), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT96), .ZN(new_n502));
  AOI211_X1 g316(.A(new_n502), .B(G902), .C1(new_n495), .C2(new_n499), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n467), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  OR2_X1    g318(.A1(new_n503), .A2(new_n467), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NOR3_X1   g320(.A1(new_n455), .A2(new_n463), .A3(new_n506), .ZN(new_n507));
  AND3_X1   g321(.A1(new_n295), .A2(new_n383), .A3(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(G234), .ZN(new_n509));
  OAI21_X1  g323(.A(G217), .B1(new_n509), .B2(G902), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n510), .B(KEYINPUT76), .ZN(new_n511));
  XNOR2_X1  g325(.A(KEYINPUT22), .B(G137), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n385), .A2(G221), .A3(G234), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n512), .B(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n413), .A2(new_n417), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT23), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n516), .B1(new_n300), .B2(G128), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n300), .A2(G128), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n236), .A2(KEYINPUT23), .A3(G119), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(G110), .ZN(new_n521));
  XNOR2_X1  g335(.A(KEYINPUT24), .B(G110), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT77), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n523), .B1(new_n300), .B2(G128), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n236), .A2(KEYINPUT77), .A3(G119), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n524), .A2(new_n525), .A3(new_n518), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n521), .B1(new_n522), .B2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n526), .A2(new_n522), .ZN(new_n529));
  INV_X1    g343(.A(G110), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n517), .A2(new_n519), .A3(new_n530), .A4(new_n518), .ZN(new_n531));
  AOI22_X1  g345(.A1(new_n529), .A2(new_n531), .B1(new_n209), .B2(new_n415), .ZN(new_n532));
  AOI22_X1  g346(.A1(new_n515), .A2(new_n528), .B1(new_n417), .B2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT79), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n514), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  AND2_X1   g349(.A1(new_n532), .A2(new_n417), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n527), .B1(new_n413), .B2(new_n417), .ZN(new_n537));
  OAI21_X1  g351(.A(KEYINPUT79), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n515), .A2(new_n528), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n532), .A2(new_n417), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n539), .A2(new_n534), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n538), .A2(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n535), .B1(new_n542), .B2(new_n514), .ZN(new_n543));
  AOI21_X1  g357(.A(KEYINPUT25), .B1(new_n543), .B2(new_n282), .ZN(new_n544));
  INV_X1    g358(.A(new_n514), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n545), .B1(new_n538), .B2(new_n541), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT25), .ZN(new_n547));
  NOR4_X1   g361(.A1(new_n546), .A2(new_n535), .A3(new_n547), .A4(G902), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n511), .B1(new_n544), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n510), .A2(new_n282), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n543), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n388), .A2(G210), .ZN(new_n554));
  XNOR2_X1  g368(.A(new_n554), .B(KEYINPUT27), .ZN(new_n555));
  XNOR2_X1  g369(.A(KEYINPUT26), .B(G101), .ZN(new_n556));
  XNOR2_X1  g370(.A(new_n555), .B(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT28), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n338), .A2(new_n339), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT64), .ZN(new_n561));
  INV_X1    g375(.A(new_n204), .ZN(new_n562));
  NOR3_X1   g376(.A1(new_n240), .A2(new_n562), .A3(new_n205), .ZN(new_n563));
  INV_X1    g377(.A(new_n214), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n561), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n211), .A2(KEYINPUT64), .A3(new_n214), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n565), .A2(new_n270), .A3(new_n566), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n197), .A2(G134), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n194), .A2(G137), .ZN(new_n569));
  OAI21_X1  g383(.A(G131), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n202), .A2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n253), .A2(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n560), .B1(new_n567), .B2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT71), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n571), .B1(new_n252), .B2(new_n238), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n576), .B1(new_n270), .B2(new_n256), .ZN(new_n577));
  AOI22_X1  g391(.A1(new_n574), .A2(new_n575), .B1(new_n577), .B2(new_n560), .ZN(new_n578));
  AOI22_X1  g392(.A1(new_n215), .A2(new_n561), .B1(new_n200), .B2(new_n202), .ZN(new_n579));
  AOI22_X1  g393(.A1(new_n579), .A2(new_n566), .B1(new_n253), .B2(new_n572), .ZN(new_n580));
  OAI21_X1  g394(.A(KEYINPUT71), .B1(new_n580), .B2(new_n560), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n559), .B1(new_n578), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n256), .A2(new_n270), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n573), .A2(new_n560), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(new_n559), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n558), .B1(new_n582), .B2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT66), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n588), .B1(new_n580), .B2(KEYINPUT30), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n567), .A2(new_n573), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT30), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n590), .A2(KEYINPUT66), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT70), .ZN(new_n594));
  OAI21_X1  g408(.A(KEYINPUT30), .B1(new_n203), .B2(new_n215), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n594), .B1(new_n595), .B2(new_n576), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n591), .B1(new_n256), .B2(new_n270), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n597), .A2(new_n573), .A3(KEYINPUT70), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n560), .B1(new_n596), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n593), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n584), .A2(new_n557), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  AOI21_X1  g416(.A(KEYINPUT31), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT31), .ZN(new_n604));
  AOI211_X1 g418(.A(new_n604), .B(new_n601), .C1(new_n593), .C2(new_n599), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n587), .B1(new_n603), .B2(new_n605), .ZN(new_n606));
  NOR2_X1   g420(.A1(G472), .A2(G902), .ZN(new_n607));
  AND3_X1   g421(.A1(new_n606), .A2(KEYINPUT32), .A3(new_n607), .ZN(new_n608));
  XNOR2_X1  g422(.A(KEYINPUT72), .B(KEYINPUT32), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n609), .B1(new_n606), .B2(new_n607), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT29), .ZN(new_n612));
  INV_X1    g426(.A(new_n584), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n613), .B1(new_n593), .B2(new_n599), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n612), .B1(new_n614), .B2(new_n557), .ZN(new_n615));
  NOR3_X1   g429(.A1(new_n582), .A2(new_n586), .A3(new_n558), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n282), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n573), .A2(new_n583), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(new_n324), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n619), .A2(KEYINPUT73), .A3(new_n584), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT73), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n618), .A2(new_n621), .A3(new_n324), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n620), .A2(KEYINPUT28), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n585), .A2(KEYINPUT74), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT74), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n584), .A2(new_n625), .A3(new_n559), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n558), .A2(new_n612), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n623), .A2(new_n624), .A3(new_n626), .A4(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(KEYINPUT75), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n624), .A2(new_n626), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT75), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n631), .A2(new_n632), .A3(new_n623), .A4(new_n627), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n629), .A2(new_n633), .ZN(new_n634));
  OAI21_X1  g448(.A(G472), .B1(new_n617), .B2(new_n634), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n553), .B1(new_n611), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n508), .A2(new_n636), .ZN(new_n637));
  XOR2_X1   g451(.A(KEYINPUT97), .B(G101), .Z(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(G3));
  INV_X1    g453(.A(KEYINPUT98), .ZN(new_n640));
  INV_X1    g454(.A(new_n553), .ZN(new_n641));
  AOI21_X1  g455(.A(KEYINPUT66), .B1(new_n590), .B2(new_n591), .ZN(new_n642));
  AOI211_X1 g456(.A(new_n588), .B(KEYINPUT30), .C1(new_n567), .C2(new_n573), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n598), .ZN(new_n645));
  AOI21_X1  g459(.A(KEYINPUT70), .B1(new_n597), .B2(new_n573), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n324), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n602), .B1(new_n644), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(new_n604), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n600), .A2(KEYINPUT31), .A3(new_n602), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n590), .A2(new_n575), .A3(new_n324), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n581), .A2(new_n584), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(KEYINPUT28), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n653), .A2(new_n585), .ZN(new_n654));
  AOI22_X1  g468(.A1(new_n649), .A2(new_n650), .B1(new_n654), .B2(new_n558), .ZN(new_n655));
  OAI21_X1  g469(.A(G472), .B1(new_n655), .B2(G902), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n606), .A2(new_n607), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n641), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n292), .A2(new_n294), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n640), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(G472), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n661), .B1(new_n606), .B2(new_n282), .ZN(new_n662));
  INV_X1    g476(.A(new_n607), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n655), .A2(new_n663), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n295), .A2(new_n665), .A3(KEYINPUT98), .A4(new_n641), .ZN(new_n666));
  AND2_X1   g480(.A1(new_n660), .A2(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(new_n463), .ZN(new_n668));
  AND3_X1   g482(.A1(new_n376), .A2(new_n298), .A3(new_n381), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n298), .B1(new_n376), .B2(new_n381), .ZN(new_n670));
  OAI211_X1 g484(.A(new_n296), .B(new_n668), .C1(new_n669), .C2(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n455), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n464), .A2(G902), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n495), .A2(new_n499), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT99), .ZN(new_n676));
  AOI21_X1  g490(.A(KEYINPUT33), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT33), .ZN(new_n678));
  AOI211_X1 g492(.A(KEYINPUT99), .B(new_n678), .C1(new_n495), .C2(new_n499), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n674), .B1(new_n677), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n675), .A2(new_n282), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(new_n464), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n673), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n672), .A2(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n667), .A2(new_n687), .ZN(new_n688));
  XOR2_X1   g502(.A(KEYINPUT34), .B(G104), .Z(new_n689));
  XNOR2_X1  g503(.A(new_n688), .B(new_n689), .ZN(G6));
  NOR2_X1   g504(.A1(new_n503), .A2(new_n467), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n681), .A2(new_n502), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n500), .A2(KEYINPUT96), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n691), .B1(new_n694), .B2(new_n467), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n447), .A2(new_n448), .A3(new_n449), .ZN(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n452), .A2(new_n448), .ZN(new_n698));
  OAI21_X1  g512(.A(new_n436), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n695), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n672), .A2(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n667), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(KEYINPUT100), .ZN(new_n704));
  XOR2_X1   g518(.A(KEYINPUT35), .B(G107), .Z(new_n705));
  XNOR2_X1  g519(.A(new_n704), .B(new_n705), .ZN(G9));
  NAND2_X1  g520(.A1(new_n539), .A2(new_n540), .ZN(new_n707));
  OR2_X1    g521(.A1(new_n545), .A2(KEYINPUT36), .ZN(new_n708));
  OR2_X1    g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n707), .A2(new_n708), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n709), .A2(new_n551), .A3(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT101), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n709), .A2(KEYINPUT101), .A3(new_n551), .A4(new_n710), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NOR3_X1   g529(.A1(new_n536), .A2(new_n537), .A3(KEYINPUT79), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n534), .B1(new_n539), .B2(new_n540), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n514), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(new_n535), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n718), .A2(new_n282), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(new_n547), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n543), .A2(KEYINPUT25), .A3(new_n282), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n715), .B1(new_n723), .B2(new_n511), .ZN(new_n724));
  NOR3_X1   g538(.A1(new_n662), .A2(new_n664), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n508), .A2(new_n725), .ZN(new_n726));
  XOR2_X1   g540(.A(KEYINPUT37), .B(G110), .Z(new_n727));
  XNOR2_X1  g541(.A(new_n726), .B(new_n727), .ZN(G12));
  INV_X1    g542(.A(new_n609), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n729), .B1(new_n655), .B2(new_n663), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n606), .A2(KEYINPUT32), .A3(new_n607), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n635), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n447), .A2(new_n449), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n733), .A2(KEYINPUT20), .ZN(new_n734));
  AOI22_X1  g548(.A1(new_n734), .A2(new_n696), .B1(G475), .B2(new_n435), .ZN(new_n735));
  XOR2_X1   g549(.A(new_n458), .B(KEYINPUT103), .Z(new_n736));
  INV_X1    g550(.A(G900), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n457), .A2(new_n737), .A3(G902), .A4(G953), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(KEYINPUT102), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n736), .A2(new_n739), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n506), .A2(new_n735), .A3(new_n740), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n741), .A2(new_n724), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n732), .A2(new_n295), .A3(new_n383), .A4(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G128), .ZN(G30));
  NAND2_X1  g558(.A1(new_n371), .A2(new_n382), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(KEYINPUT38), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n600), .A2(new_n584), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(new_n557), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n620), .A2(new_n622), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(new_n558), .ZN(new_n750));
  AOI21_X1  g564(.A(KEYINPUT104), .B1(new_n748), .B2(new_n750), .ZN(new_n751));
  OAI211_X1 g565(.A(KEYINPUT104), .B(new_n750), .C1(new_n614), .C2(new_n558), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(new_n282), .ZN(new_n753));
  OAI21_X1  g567(.A(G472), .B1(new_n751), .B2(new_n753), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n754), .A2(new_n730), .A3(new_n731), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n455), .A2(new_n506), .ZN(new_n756));
  INV_X1    g570(.A(new_n715), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n549), .A2(new_n757), .ZN(new_n758));
  NOR3_X1   g572(.A1(new_n756), .A2(new_n758), .A3(new_n297), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n746), .A2(new_n755), .A3(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n740), .B(KEYINPUT39), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n295), .A2(KEYINPUT105), .A3(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n292), .A2(new_n294), .A3(new_n761), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT105), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n762), .A2(new_n765), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n760), .B1(KEYINPUT40), .B2(new_n766), .ZN(new_n767));
  OR2_X1    g581(.A1(new_n766), .A2(KEYINPUT40), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G143), .ZN(G45));
  OAI21_X1  g584(.A(new_n296), .B1(new_n669), .B2(new_n670), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n659), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n455), .A2(new_n683), .A3(new_n740), .ZN(new_n773));
  INV_X1    g587(.A(new_n773), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n772), .A2(new_n732), .A3(new_n758), .A4(new_n774), .ZN(new_n775));
  XOR2_X1   g589(.A(KEYINPUT106), .B(G146), .Z(new_n776));
  XNOR2_X1  g590(.A(new_n775), .B(new_n776), .ZN(G48));
  NAND2_X1  g591(.A1(new_n280), .A2(new_n282), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(G469), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n779), .A2(new_n294), .A3(new_n283), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT107), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n779), .A2(KEYINPUT107), .A3(new_n294), .A4(new_n283), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n732), .A2(new_n782), .A3(new_n641), .A4(new_n783), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n784), .A2(new_n686), .ZN(new_n785));
  XOR2_X1   g599(.A(KEYINPUT41), .B(G113), .Z(new_n786));
  XNOR2_X1  g600(.A(new_n785), .B(new_n786), .ZN(G15));
  NOR2_X1   g601(.A1(new_n784), .A2(new_n701), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(new_n303), .ZN(G18));
  NOR2_X1   g603(.A1(new_n780), .A2(new_n771), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n790), .A2(new_n732), .A3(new_n507), .A4(new_n758), .ZN(new_n791));
  XOR2_X1   g605(.A(KEYINPUT108), .B(G119), .Z(new_n792));
  XNOR2_X1  g606(.A(new_n791), .B(new_n792), .ZN(G21));
  NOR3_X1   g607(.A1(new_n771), .A2(new_n756), .A3(KEYINPUT109), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT109), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT93), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n696), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n797), .A2(new_n450), .A3(new_n734), .ZN(new_n798));
  AOI22_X1  g612(.A1(new_n798), .A2(new_n436), .B1(new_n504), .B2(new_n505), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n795), .B1(new_n383), .B2(new_n799), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n794), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n649), .A2(new_n650), .ZN(new_n802));
  INV_X1    g616(.A(new_n623), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n558), .B1(new_n803), .B2(new_n630), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n663), .B1(new_n802), .B2(new_n804), .ZN(new_n805));
  NOR3_X1   g619(.A1(new_n662), .A2(new_n553), .A3(new_n805), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n806), .A2(new_n782), .A3(new_n668), .A4(new_n783), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n801), .A2(new_n807), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(new_n472), .ZN(G24));
  NOR3_X1   g623(.A1(new_n662), .A2(new_n724), .A3(new_n805), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n790), .A2(new_n810), .A3(new_n774), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n811), .B(G125), .ZN(G27));
  INV_X1    g626(.A(KEYINPUT32), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n657), .A2(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n814), .A2(new_n635), .A3(new_n731), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(new_n641), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n669), .A2(new_n670), .A3(new_n297), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n295), .A2(new_n774), .A3(new_n817), .ZN(new_n818));
  OAI21_X1  g632(.A(KEYINPUT42), .B1(new_n816), .B2(new_n818), .ZN(new_n819));
  AND3_X1   g633(.A1(new_n817), .A2(new_n294), .A3(new_n292), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n773), .A2(KEYINPUT42), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n636), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n819), .A2(new_n822), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n823), .B(new_n201), .ZN(G33));
  INV_X1    g638(.A(new_n741), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n820), .A2(new_n732), .A3(new_n641), .A4(new_n825), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n826), .B(G134), .ZN(G36));
  NAND3_X1  g641(.A1(new_n683), .A2(new_n798), .A3(new_n436), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n828), .A2(KEYINPUT110), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT111), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT43), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n832), .B1(new_n828), .B2(KEYINPUT111), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n665), .A2(new_n724), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n829), .A2(new_n830), .A3(new_n832), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n834), .A2(new_n835), .A3(KEYINPUT44), .A4(new_n836), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n285), .B1(new_n288), .B2(new_n191), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT45), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  OAI211_X1 g654(.A(new_n285), .B(KEYINPUT45), .C1(new_n288), .C2(new_n191), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n840), .A2(G469), .A3(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT46), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n842), .A2(new_n843), .A3(new_n283), .A4(new_n291), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(new_n294), .ZN(new_n845));
  INV_X1    g659(.A(new_n761), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n843), .B1(new_n842), .B2(new_n291), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n845), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n848), .A2(new_n817), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n834), .A2(new_n835), .A3(new_n836), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT112), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT44), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n850), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(new_n853), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n851), .B1(new_n850), .B2(new_n852), .ZN(new_n855));
  OAI211_X1 g669(.A(new_n837), .B(new_n849), .C1(new_n854), .C2(new_n855), .ZN(new_n856));
  XNOR2_X1  g670(.A(new_n856), .B(G137), .ZN(G39));
  INV_X1    g671(.A(KEYINPUT47), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n858), .B1(new_n845), .B2(new_n847), .ZN(new_n859));
  INV_X1    g673(.A(new_n847), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n860), .A2(KEYINPUT47), .A3(new_n294), .A4(new_n844), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n817), .A2(new_n553), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n732), .A2(new_n863), .A3(new_n773), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n865), .B(G140), .ZN(G42));
  NAND3_X1  g680(.A1(new_n641), .A2(new_n294), .A3(new_n296), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n746), .A2(new_n755), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n779), .A2(new_n283), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n828), .B1(new_n869), .B2(KEYINPUT49), .ZN(new_n870));
  OAI211_X1 g684(.A(new_n868), .B(new_n870), .C1(KEYINPUT49), .C2(new_n869), .ZN(new_n871));
  INV_X1    g685(.A(new_n736), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n834), .A2(new_n872), .A3(new_n836), .ZN(new_n873));
  INV_X1    g687(.A(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n874), .A2(new_n806), .ZN(new_n875));
  OR3_X1    g689(.A1(new_n746), .A2(new_n296), .A3(new_n780), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  XNOR2_X1  g691(.A(new_n877), .B(KEYINPUT50), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT51), .ZN(new_n879));
  OAI211_X1 g693(.A(new_n859), .B(new_n861), .C1(new_n294), .C2(new_n869), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n880), .A2(new_n817), .ZN(new_n881));
  INV_X1    g695(.A(new_n875), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n879), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(new_n755), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n780), .A2(new_n297), .A3(new_n745), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n884), .A2(new_n885), .A3(new_n641), .A4(new_n459), .ZN(new_n886));
  OR3_X1    g700(.A1(new_n886), .A2(new_n455), .A3(new_n683), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n874), .A2(new_n810), .A3(new_n885), .ZN(new_n888));
  AOI21_X1  g702(.A(KEYINPUT118), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n887), .A2(new_n888), .A3(KEYINPUT118), .ZN(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  OAI211_X1 g705(.A(new_n878), .B(new_n883), .C1(new_n889), .C2(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT50), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n877), .B(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n881), .A2(new_n882), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n895), .A2(new_n888), .A3(new_n887), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n879), .B1(new_n894), .B2(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(new_n816), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n874), .A2(new_n898), .A3(new_n885), .ZN(new_n899));
  XOR2_X1   g713(.A(new_n899), .B(KEYINPUT48), .Z(new_n900));
  INV_X1    g714(.A(new_n685), .ZN(new_n901));
  INV_X1    g715(.A(new_n790), .ZN(new_n902));
  OAI221_X1 g716(.A(new_n456), .B1(new_n901), .B2(new_n886), .C1(new_n875), .C2(new_n902), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n900), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n892), .A2(new_n897), .A3(new_n904), .ZN(new_n905));
  AND2_X1   g719(.A1(new_n819), .A2(new_n822), .ZN(new_n906));
  INV_X1    g720(.A(new_n807), .ZN(new_n907));
  OAI21_X1  g721(.A(KEYINPUT109), .B1(new_n771), .B2(new_n756), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n383), .A2(new_n795), .A3(new_n799), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  AND4_X1   g724(.A1(new_n732), .A2(new_n782), .A3(new_n641), .A4(new_n783), .ZN(new_n911));
  AOI22_X1  g725(.A1(new_n907), .A2(new_n910), .B1(new_n911), .B2(new_n702), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT53), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n811), .A2(new_n743), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n913), .B1(new_n914), .B2(KEYINPUT52), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n791), .B1(new_n784), .B2(new_n686), .ZN(new_n916));
  INV_X1    g730(.A(new_n916), .ZN(new_n917));
  AND4_X1   g731(.A1(new_n906), .A2(new_n912), .A3(new_n915), .A4(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n732), .A2(new_n758), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n295), .A2(new_n383), .A3(new_n774), .ZN(new_n920));
  OAI211_X1 g734(.A(new_n811), .B(new_n743), .C1(new_n919), .C2(new_n920), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n755), .A2(new_n295), .A3(new_n724), .A4(new_n740), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n801), .A2(new_n922), .ZN(new_n923));
  OAI21_X1  g737(.A(KEYINPUT52), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n700), .A2(new_n758), .A3(new_n740), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n925), .B1(new_n611), .B2(new_n635), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n804), .B1(new_n603), .B2(new_n605), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(new_n607), .ZN(new_n928));
  AOI21_X1  g742(.A(G902), .B1(new_n802), .B2(new_n587), .ZN(new_n929));
  OAI211_X1 g743(.A(new_n928), .B(new_n758), .C1(new_n929), .C2(new_n661), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n930), .A2(new_n773), .ZN(new_n931));
  AOI22_X1  g745(.A1(new_n926), .A2(new_n772), .B1(new_n931), .B2(new_n790), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT52), .ZN(new_n933));
  INV_X1    g747(.A(new_n740), .ZN(new_n934));
  NOR3_X1   g748(.A1(new_n659), .A2(new_n758), .A3(new_n934), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n910), .A2(new_n755), .A3(new_n935), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n932), .A2(new_n933), .A3(new_n775), .A4(new_n936), .ZN(new_n937));
  AND2_X1   g751(.A1(new_n924), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n508), .B1(new_n636), .B2(new_n725), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT113), .ZN(new_n940));
  AND3_X1   g754(.A1(new_n455), .A2(new_n940), .A3(new_n683), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n940), .B1(new_n455), .B2(new_n683), .ZN(new_n942));
  NOR3_X1   g756(.A1(new_n941), .A2(new_n671), .A3(new_n942), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n660), .A2(new_n666), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n673), .A2(new_n506), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n945), .A2(new_n671), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n660), .A2(new_n666), .A3(new_n946), .ZN(new_n947));
  AND3_X1   g761(.A1(new_n939), .A2(new_n944), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n931), .A2(new_n820), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n695), .A2(KEYINPUT114), .A3(new_n735), .A4(new_n740), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT114), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n504), .A2(new_n505), .A3(new_n740), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n951), .B1(new_n952), .B2(new_n699), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n817), .A2(new_n950), .A3(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT115), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n817), .A2(new_n953), .A3(KEYINPUT115), .A4(new_n950), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n732), .A2(new_n295), .A3(new_n758), .ZN(new_n959));
  OAI211_X1 g773(.A(new_n826), .B(new_n949), .C1(new_n958), .C2(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(new_n960), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n948), .A2(new_n961), .A3(KEYINPUT116), .ZN(new_n962));
  INV_X1    g776(.A(KEYINPUT116), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n939), .A2(new_n944), .A3(new_n947), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n963), .B1(new_n964), .B2(new_n960), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n918), .A2(new_n938), .A3(new_n962), .A4(new_n965), .ZN(new_n966));
  OAI22_X1  g780(.A1(new_n801), .A2(new_n807), .B1(new_n784), .B2(new_n701), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n967), .A2(new_n916), .ZN(new_n968));
  NAND4_X1  g782(.A1(new_n968), .A2(new_n924), .A3(new_n906), .A4(new_n937), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n948), .A2(new_n961), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n913), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT54), .ZN(new_n972));
  AND3_X1   g786(.A1(new_n966), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n964), .A2(new_n960), .ZN(new_n974));
  NOR3_X1   g788(.A1(new_n823), .A2(new_n967), .A3(new_n916), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n913), .B1(new_n932), .B2(new_n933), .ZN(new_n976));
  NAND4_X1  g790(.A1(new_n938), .A2(new_n974), .A3(new_n975), .A4(new_n976), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n972), .B1(new_n971), .B2(new_n977), .ZN(new_n978));
  OAI21_X1  g792(.A(KEYINPUT117), .B1(new_n973), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n971), .A2(new_n977), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n980), .A2(KEYINPUT54), .ZN(new_n981));
  INV_X1    g795(.A(KEYINPUT117), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n966), .A2(new_n971), .A3(new_n972), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n981), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n905), .B1(new_n979), .B2(new_n984), .ZN(new_n985));
  NOR2_X1   g799(.A1(G952), .A2(G953), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n871), .B1(new_n985), .B2(new_n986), .ZN(G75));
  NOR2_X1   g801(.A1(new_n385), .A2(G952), .ZN(new_n988));
  INV_X1    g802(.A(new_n988), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n282), .B1(new_n966), .B2(new_n971), .ZN(new_n990));
  AOI21_X1  g804(.A(KEYINPUT56), .B1(new_n990), .B2(G210), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n378), .B1(new_n380), .B2(new_n343), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n992), .B(new_n379), .ZN(new_n993));
  XOR2_X1   g807(.A(KEYINPUT119), .B(KEYINPUT55), .Z(new_n994));
  XNOR2_X1  g808(.A(new_n993), .B(new_n994), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n989), .B1(new_n991), .B2(new_n995), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n996), .B1(new_n991), .B2(new_n995), .ZN(G51));
  XNOR2_X1  g811(.A(new_n290), .B(KEYINPUT57), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n972), .B1(new_n966), .B2(new_n971), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n998), .B1(new_n973), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n1000), .A2(new_n280), .ZN(new_n1001));
  NAND4_X1  g815(.A1(new_n990), .A2(G469), .A3(new_n841), .A4(new_n840), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n988), .B1(new_n1001), .B2(new_n1002), .ZN(G54));
  AND2_X1   g817(.A1(KEYINPUT58), .A2(G475), .ZN(new_n1004));
  AND3_X1   g818(.A1(new_n990), .A2(new_n447), .A3(new_n1004), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n447), .B1(new_n990), .B2(new_n1004), .ZN(new_n1006));
  NOR3_X1   g820(.A1(new_n1005), .A2(new_n1006), .A3(new_n988), .ZN(G60));
  OR2_X1    g821(.A1(new_n677), .A2(new_n679), .ZN(new_n1008));
  INV_X1    g822(.A(new_n1008), .ZN(new_n1009));
  NAND2_X1  g823(.A1(G478), .A2(G902), .ZN(new_n1010));
  XOR2_X1   g824(.A(new_n1010), .B(KEYINPUT59), .Z(new_n1011));
  NOR2_X1   g825(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g826(.A(new_n1012), .B1(new_n973), .B2(new_n999), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1013), .A2(new_n989), .ZN(new_n1014));
  INV_X1    g828(.A(new_n1011), .ZN(new_n1015));
  NAND3_X1  g829(.A1(new_n979), .A2(new_n984), .A3(new_n1015), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n1014), .B1(new_n1016), .B2(new_n1009), .ZN(G63));
  NAND2_X1  g831(.A1(new_n966), .A2(new_n971), .ZN(new_n1018));
  NAND2_X1  g832(.A1(G217), .A2(G902), .ZN(new_n1019));
  XNOR2_X1  g833(.A(new_n1019), .B(KEYINPUT60), .ZN(new_n1020));
  INV_X1    g834(.A(new_n1020), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1018), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g836(.A(new_n543), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n988), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n709), .A2(new_n710), .ZN(new_n1025));
  OAI211_X1 g839(.A(new_n1024), .B(KEYINPUT61), .C1(new_n1025), .C2(new_n1022), .ZN(new_n1026));
  INV_X1    g840(.A(KEYINPUT61), .ZN(new_n1027));
  NOR2_X1   g841(.A1(new_n1022), .A2(new_n1025), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n1020), .B1(new_n966), .B2(new_n971), .ZN(new_n1029));
  OAI21_X1  g843(.A(new_n989), .B1(new_n1029), .B2(new_n543), .ZN(new_n1030));
  OAI21_X1  g844(.A(new_n1027), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n1026), .A2(new_n1031), .ZN(G66));
  OAI21_X1  g846(.A(G953), .B1(new_n460), .B2(new_n349), .ZN(new_n1033));
  NAND2_X1  g847(.A1(new_n948), .A2(new_n968), .ZN(new_n1034));
  INV_X1    g848(.A(new_n1034), .ZN(new_n1035));
  OAI21_X1  g849(.A(new_n1033), .B1(new_n1035), .B2(G953), .ZN(new_n1036));
  OAI21_X1  g850(.A(new_n992), .B1(G898), .B2(new_n385), .ZN(new_n1037));
  XNOR2_X1  g851(.A(new_n1036), .B(new_n1037), .ZN(G69));
  OAI21_X1  g852(.A(G953), .B1(new_n189), .B2(new_n737), .ZN(new_n1039));
  XOR2_X1   g853(.A(new_n1039), .B(KEYINPUT125), .Z(new_n1040));
  INV_X1    g854(.A(new_n1040), .ZN(new_n1041));
  OAI21_X1  g855(.A(new_n593), .B1(new_n646), .B2(new_n645), .ZN(new_n1042));
  NOR2_X1   g856(.A1(new_n438), .A2(new_n439), .ZN(new_n1043));
  XOR2_X1   g857(.A(new_n1042), .B(new_n1043), .Z(new_n1044));
  INV_X1    g858(.A(new_n1044), .ZN(new_n1045));
  INV_X1    g859(.A(KEYINPUT120), .ZN(new_n1046));
  NAND3_X1  g860(.A1(new_n932), .A2(new_n1046), .A3(new_n775), .ZN(new_n1047));
  NAND2_X1  g861(.A1(new_n921), .A2(KEYINPUT120), .ZN(new_n1048));
  NAND2_X1  g862(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g863(.A1(new_n1049), .A2(new_n769), .ZN(new_n1050));
  NAND3_X1  g864(.A1(new_n1050), .A2(KEYINPUT121), .A3(KEYINPUT62), .ZN(new_n1051));
  INV_X1    g865(.A(KEYINPUT121), .ZN(new_n1052));
  AOI22_X1  g866(.A1(new_n1047), .A2(new_n1048), .B1(new_n767), .B2(new_n768), .ZN(new_n1053));
  INV_X1    g867(.A(KEYINPUT62), .ZN(new_n1054));
  OAI21_X1  g868(.A(new_n1052), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g869(.A1(new_n1051), .A2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g870(.A1(new_n1049), .A2(new_n1054), .A3(new_n769), .ZN(new_n1057));
  NAND3_X1  g871(.A1(new_n732), .A2(new_n641), .A3(new_n817), .ZN(new_n1058));
  NOR2_X1   g872(.A1(new_n766), .A2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g873(.A(new_n945), .B1(new_n941), .B2(new_n942), .ZN(new_n1060));
  INV_X1    g874(.A(KEYINPUT122), .ZN(new_n1061));
  NAND2_X1  g875(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  OAI211_X1 g876(.A(KEYINPUT122), .B(new_n945), .C1(new_n941), .C2(new_n942), .ZN(new_n1063));
  NAND2_X1  g877(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g878(.A1(new_n1059), .A2(KEYINPUT123), .A3(new_n1064), .ZN(new_n1065));
  NAND2_X1  g879(.A1(new_n1065), .A2(new_n865), .ZN(new_n1066));
  AOI21_X1  g880(.A(KEYINPUT123), .B1(new_n1059), .B2(new_n1064), .ZN(new_n1067));
  NOR2_X1   g881(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND4_X1  g882(.A1(new_n1056), .A2(new_n856), .A3(new_n1057), .A4(new_n1068), .ZN(new_n1069));
  AOI21_X1  g883(.A(new_n1045), .B1(new_n1069), .B2(new_n385), .ZN(new_n1070));
  NAND3_X1  g884(.A1(new_n819), .A2(new_n822), .A3(new_n826), .ZN(new_n1071));
  NAND2_X1  g885(.A1(new_n1071), .A2(KEYINPUT124), .ZN(new_n1072));
  INV_X1    g886(.A(KEYINPUT124), .ZN(new_n1073));
  NAND4_X1  g887(.A1(new_n819), .A2(new_n822), .A3(new_n1073), .A4(new_n826), .ZN(new_n1074));
  NOR2_X1   g888(.A1(new_n801), .A2(new_n816), .ZN(new_n1075));
  AOI22_X1  g889(.A1(new_n1075), .A2(new_n848), .B1(new_n862), .B2(new_n864), .ZN(new_n1076));
  NAND4_X1  g890(.A1(new_n1049), .A2(new_n1072), .A3(new_n1074), .A4(new_n1076), .ZN(new_n1077));
  NAND2_X1  g891(.A1(new_n849), .A2(new_n837), .ZN(new_n1078));
  INV_X1    g892(.A(new_n855), .ZN(new_n1079));
  AOI21_X1  g893(.A(new_n1078), .B1(new_n1079), .B2(new_n853), .ZN(new_n1080));
  OAI21_X1  g894(.A(new_n385), .B1(new_n1077), .B2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g895(.A1(new_n737), .A2(G953), .ZN(new_n1082));
  AND2_X1   g896(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NOR2_X1   g897(.A1(new_n1083), .A2(new_n1044), .ZN(new_n1084));
  OAI21_X1  g898(.A(new_n1041), .B1(new_n1070), .B2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g899(.A1(new_n1068), .A2(new_n856), .A3(new_n1057), .ZN(new_n1086));
  AOI21_X1  g900(.A(new_n1086), .B1(new_n1055), .B2(new_n1051), .ZN(new_n1087));
  OAI21_X1  g901(.A(new_n1044), .B1(new_n1087), .B2(G953), .ZN(new_n1088));
  OAI211_X1 g902(.A(new_n1088), .B(new_n1040), .C1(new_n1044), .C2(new_n1083), .ZN(new_n1089));
  NAND2_X1  g903(.A1(new_n1085), .A2(new_n1089), .ZN(G72));
  NOR2_X1   g904(.A1(new_n747), .A2(new_n557), .ZN(new_n1091));
  NOR3_X1   g905(.A1(new_n1077), .A2(new_n1080), .A3(new_n1034), .ZN(new_n1092));
  XOR2_X1   g906(.A(KEYINPUT126), .B(KEYINPUT63), .Z(new_n1093));
  NOR2_X1   g907(.A1(new_n661), .A2(new_n282), .ZN(new_n1094));
  XNOR2_X1  g908(.A(new_n1093), .B(new_n1094), .ZN(new_n1095));
  OAI21_X1  g909(.A(new_n1091), .B1(new_n1092), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g910(.A(KEYINPUT127), .ZN(new_n1097));
  AND3_X1   g911(.A1(new_n1096), .A2(new_n1097), .A3(new_n989), .ZN(new_n1098));
  AOI21_X1  g912(.A(new_n1097), .B1(new_n1096), .B2(new_n989), .ZN(new_n1099));
  NOR2_X1   g913(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g914(.A(new_n748), .ZN(new_n1101));
  NOR3_X1   g915(.A1(new_n1101), .A2(new_n1091), .A3(new_n1095), .ZN(new_n1102));
  NAND2_X1  g916(.A1(new_n980), .A2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g917(.A(new_n1095), .B1(new_n1087), .B2(new_n1035), .ZN(new_n1104));
  OAI21_X1  g918(.A(new_n1103), .B1(new_n1104), .B2(new_n748), .ZN(new_n1105));
  NOR2_X1   g919(.A1(new_n1100), .A2(new_n1105), .ZN(G57));
endmodule


