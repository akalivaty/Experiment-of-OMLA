//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 0 0 0 1 0 0 1 1 0 1 1 0 0 0 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 1 1 0 1 1 1 0 1 0 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:19 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n492, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n511,
    new_n512, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n543,
    new_n544, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n563, new_n564, new_n565, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n607, new_n610, new_n611,
    new_n613, new_n614, new_n616, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1177;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT65), .B(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT66), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT67), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT68), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT69), .Z(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G219), .A2(G221), .A3(G220), .A4(G218), .ZN(new_n451));
  XNOR2_X1  g026(.A(KEYINPUT70), .B(KEYINPUT2), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n453), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n453), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT71), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  OAI21_X1  g039(.A(G125), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n462), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  OAI211_X1 g042(.A(G137), .B(new_n462), .C1(new_n463), .C2(new_n464), .ZN(new_n468));
  AND2_X1   g043(.A1(new_n462), .A2(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G101), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n467), .A2(new_n471), .ZN(G160));
  XNOR2_X1  g047(.A(KEYINPUT3), .B(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G2105), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G124), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n462), .A2(G112), .ZN(new_n477));
  OAI21_X1  g052(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  AND2_X1   g054(.A1(new_n473), .A2(new_n462), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n479), .B1(G136), .B2(new_n480), .ZN(new_n481));
  XOR2_X1   g056(.A(new_n481), .B(KEYINPUT72), .Z(G162));
  OAI211_X1 g057(.A(G138), .B(new_n462), .C1(new_n463), .C2(new_n464), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT4), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND4_X1  g060(.A1(new_n473), .A2(KEYINPUT4), .A3(G138), .A4(new_n462), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n473), .A2(G126), .A3(G2105), .ZN(new_n487));
  OR2_X1    g062(.A1(G102), .A2(G2105), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n488), .B(G2104), .C1(G114), .C2(new_n462), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n485), .A2(new_n486), .A3(new_n487), .A4(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G164));
  INV_X1    g066(.A(G543), .ZN(new_n492));
  NAND2_X1  g067(.A1(KEYINPUT73), .A2(G651), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT6), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g070(.A1(KEYINPUT73), .A2(KEYINPUT6), .A3(G651), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n492), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(G50), .ZN(new_n498));
  INV_X1    g073(.A(G88), .ZN(new_n499));
  AND3_X1   g074(.A1(KEYINPUT73), .A2(KEYINPUT6), .A3(G651), .ZN(new_n500));
  AOI21_X1  g075(.A(KEYINPUT6), .B1(KEYINPUT73), .B2(G651), .ZN(new_n501));
  AND2_X1   g076(.A1(KEYINPUT5), .A2(G543), .ZN(new_n502));
  NOR2_X1   g077(.A1(KEYINPUT5), .A2(G543), .ZN(new_n503));
  OAI22_X1  g078(.A1(new_n500), .A2(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n498), .B1(new_n499), .B2(new_n504), .ZN(new_n505));
  XNOR2_X1  g080(.A(KEYINPUT5), .B(G543), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n506), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n507));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n505), .A2(new_n509), .ZN(G166));
  NAND3_X1  g085(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n511));
  XNOR2_X1  g086(.A(new_n511), .B(KEYINPUT7), .ZN(new_n512));
  INV_X1    g087(.A(G89), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n512), .B1(new_n513), .B2(new_n504), .ZN(new_n514));
  OAI211_X1 g089(.A(G51), .B(G543), .C1(new_n500), .C2(new_n501), .ZN(new_n515));
  OAI211_X1 g090(.A(G63), .B(G651), .C1(new_n502), .C2(new_n503), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT74), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n515), .A2(KEYINPUT74), .A3(new_n516), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n514), .B1(new_n519), .B2(new_n520), .ZN(G168));
  INV_X1    g096(.A(G90), .ZN(new_n522));
  OAI21_X1  g097(.A(G543), .B1(new_n500), .B2(new_n501), .ZN(new_n523));
  INV_X1    g098(.A(G52), .ZN(new_n524));
  OAI22_X1  g099(.A1(new_n504), .A2(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  OAI21_X1  g100(.A(G64), .B1(new_n502), .B2(new_n503), .ZN(new_n526));
  NAND2_X1  g101(.A1(G77), .A2(G543), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g103(.A(new_n508), .B1(new_n528), .B2(KEYINPUT75), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT75), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n526), .A2(new_n530), .A3(new_n527), .ZN(new_n531));
  AOI21_X1  g106(.A(new_n525), .B1(new_n529), .B2(new_n531), .ZN(G171));
  NAND2_X1  g107(.A1(new_n495), .A2(new_n496), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n533), .A2(G43), .A3(G543), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n533), .A2(G81), .A3(new_n506), .ZN(new_n535));
  INV_X1    g110(.A(G68), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n536), .A2(new_n492), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n537), .B1(new_n506), .B2(G56), .ZN(new_n538));
  OAI211_X1 g113(.A(new_n534), .B(new_n535), .C1(new_n538), .C2(new_n508), .ZN(new_n539));
  INV_X1    g114(.A(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G860), .ZN(G153));
  NAND4_X1  g116(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g117(.A1(G1), .A2(G3), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT8), .ZN(new_n544));
  NAND4_X1  g119(.A1(G319), .A2(G483), .A3(G661), .A4(new_n544), .ZN(G188));
  NAND2_X1  g120(.A1(G78), .A2(G543), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n502), .A2(new_n503), .ZN(new_n547));
  INV_X1    g122(.A(G65), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  OR2_X1    g124(.A1(KEYINPUT5), .A2(G543), .ZN(new_n550));
  NAND2_X1  g125(.A1(KEYINPUT5), .A2(G543), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n495), .A2(new_n496), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n549), .A2(G651), .B1(new_n552), .B2(G91), .ZN(new_n553));
  INV_X1    g128(.A(G53), .ZN(new_n554));
  OAI21_X1  g129(.A(KEYINPUT9), .B1(new_n523), .B2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT9), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n497), .A2(new_n556), .A3(G53), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n553), .A2(new_n558), .ZN(G299));
  INV_X1    g134(.A(G171), .ZN(G301));
  INV_X1    g135(.A(G168), .ZN(G286));
  OAI221_X1 g136(.A(new_n498), .B1(new_n499), .B2(new_n504), .C1(new_n507), .C2(new_n508), .ZN(G303));
  NAND2_X1  g137(.A1(new_n552), .A2(G87), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n497), .A2(G49), .ZN(new_n564));
  OAI21_X1  g139(.A(G651), .B1(new_n506), .B2(G74), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(G288));
  INV_X1    g141(.A(KEYINPUT76), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n552), .A2(new_n567), .A3(G86), .ZN(new_n568));
  INV_X1    g143(.A(G86), .ZN(new_n569));
  OAI21_X1  g144(.A(KEYINPUT76), .B1(new_n504), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(G73), .A2(G543), .ZN(new_n572));
  INV_X1    g147(.A(G61), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n572), .B1(new_n547), .B2(new_n573), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n574), .A2(G651), .B1(G48), .B2(new_n497), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n571), .A2(new_n575), .ZN(G305));
  NAND2_X1  g151(.A1(G72), .A2(G543), .ZN(new_n577));
  INV_X1    g152(.A(G60), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n547), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n579), .A2(G651), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n497), .A2(G47), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n552), .A2(G85), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(G290));
  INV_X1    g158(.A(G66), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n584), .B1(new_n550), .B2(new_n551), .ZN(new_n585));
  NAND2_X1  g160(.A1(G79), .A2(G543), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(new_n587));
  OAI21_X1  g162(.A(KEYINPUT78), .B1(new_n585), .B2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT78), .ZN(new_n589));
  OAI211_X1 g164(.A(new_n589), .B(new_n586), .C1(new_n547), .C2(new_n584), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n588), .A2(G651), .A3(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT10), .ZN(new_n592));
  INV_X1    g167(.A(G92), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n504), .B2(new_n593), .ZN(new_n594));
  NAND4_X1  g169(.A1(new_n533), .A2(KEYINPUT10), .A3(new_n506), .A4(G92), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(G54), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT77), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n597), .B1(new_n523), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n497), .A2(KEYINPUT77), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n591), .A2(new_n596), .A3(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(G868), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n604), .B1(new_n603), .B2(G171), .ZN(G284));
  OAI21_X1  g180(.A(new_n604), .B1(new_n603), .B2(G171), .ZN(G321));
  NAND2_X1  g181(.A1(G299), .A2(new_n603), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n607), .B1(new_n603), .B2(G168), .ZN(G297));
  OAI21_X1  g183(.A(new_n607), .B1(new_n603), .B2(G168), .ZN(G280));
  AND3_X1   g184(.A1(new_n591), .A2(new_n596), .A3(new_n601), .ZN(new_n610));
  INV_X1    g185(.A(G559), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n611), .B2(G860), .ZN(G148));
  NAND2_X1  g187(.A1(new_n610), .A2(new_n611), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n613), .A2(G868), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n614), .B1(G868), .B2(new_n540), .ZN(G323));
  XOR2_X1   g190(.A(KEYINPUT79), .B(KEYINPUT11), .Z(new_n616));
  XNOR2_X1  g191(.A(G323), .B(new_n616), .ZN(G282));
  NAND2_X1  g192(.A1(new_n473), .A2(new_n469), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT12), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT13), .ZN(new_n620));
  INV_X1    g195(.A(G2100), .ZN(new_n621));
  OR2_X1    g196(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n620), .A2(new_n621), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n475), .A2(G123), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n480), .A2(G135), .ZN(new_n625));
  NOR2_X1   g200(.A1(new_n462), .A2(G111), .ZN(new_n626));
  OAI21_X1  g201(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n627));
  OAI211_X1 g202(.A(new_n624), .B(new_n625), .C1(new_n626), .C2(new_n627), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n628), .B(G2096), .Z(new_n629));
  NAND3_X1  g204(.A1(new_n622), .A2(new_n623), .A3(new_n629), .ZN(G156));
  XNOR2_X1  g205(.A(G2427), .B(G2438), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2430), .ZN(new_n632));
  XNOR2_X1  g207(.A(KEYINPUT15), .B(G2435), .ZN(new_n633));
  OR2_X1    g208(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n632), .A2(new_n633), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n634), .A2(KEYINPUT14), .A3(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT80), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2451), .B(G2454), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT16), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2443), .B(G2446), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n637), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(G1341), .B(G1348), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n642), .A2(new_n643), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n644), .A2(new_n645), .A3(G14), .ZN(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(G401));
  XOR2_X1   g222(.A(G2072), .B(G2078), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT17), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2067), .B(G2678), .ZN(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(new_n651));
  NOR2_X1   g226(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(G2084), .B(G2090), .Z(new_n653));
  AOI21_X1  g228(.A(new_n653), .B1(new_n651), .B2(new_n648), .ZN(new_n654));
  AOI21_X1  g229(.A(new_n652), .B1(KEYINPUT81), .B2(new_n654), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n655), .B1(KEYINPUT81), .B2(new_n654), .ZN(new_n656));
  INV_X1    g231(.A(new_n648), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n657), .A2(new_n653), .A3(new_n650), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(KEYINPUT18), .Z(new_n659));
  NAND3_X1  g234(.A1(new_n649), .A2(new_n653), .A3(new_n651), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n656), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(G2096), .B(G2100), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(G227));
  XOR2_X1   g238(.A(G1971), .B(G1976), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT19), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1956), .B(G2474), .ZN(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G1961), .B(G1966), .Z(new_n668));
  AND2_X1   g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n665), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT20), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n667), .A2(new_n668), .ZN(new_n672));
  NOR3_X1   g247(.A1(new_n665), .A2(new_n669), .A3(new_n672), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n673), .B1(new_n665), .B2(new_n672), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n676), .B(KEYINPUT82), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n675), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1981), .B(G1986), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT83), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n678), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1991), .B(G1996), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(G229));
  INV_X1    g258(.A(G16), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n684), .A2(G23), .ZN(new_n685));
  INV_X1    g260(.A(G288), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n685), .B1(new_n686), .B2(new_n684), .ZN(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT33), .B(G1976), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n684), .A2(G22), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n690), .B1(G166), .B2(new_n684), .ZN(new_n691));
  INV_X1    g266(.A(G1971), .ZN(new_n692));
  AND2_X1   g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n691), .A2(new_n692), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n689), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  MUX2_X1   g270(.A(G6), .B(G305), .S(G16), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT85), .ZN(new_n697));
  XOR2_X1   g272(.A(KEYINPUT32), .B(G1981), .Z(new_n698));
  AOI21_X1  g273(.A(new_n695), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(new_n697), .B2(new_n698), .ZN(new_n700));
  OR2_X1    g275(.A1(new_n700), .A2(KEYINPUT34), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n700), .A2(KEYINPUT34), .ZN(new_n702));
  AND2_X1   g277(.A1(new_n684), .A2(G24), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n703), .B1(G290), .B2(G16), .ZN(new_n704));
  INV_X1    g279(.A(G1986), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  AOI22_X1  g281(.A1(new_n475), .A2(G119), .B1(new_n480), .B2(G131), .ZN(new_n707));
  NOR2_X1   g282(.A1(G95), .A2(G2105), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT84), .ZN(new_n709));
  OAI21_X1  g284(.A(G2104), .B1(new_n462), .B2(G107), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n707), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  MUX2_X1   g286(.A(G25), .B(new_n711), .S(G29), .Z(new_n712));
  XOR2_X1   g287(.A(KEYINPUT35), .B(G1991), .Z(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n712), .B(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(new_n704), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n715), .B1(G1986), .B2(new_n716), .ZN(new_n717));
  NAND4_X1  g292(.A1(new_n701), .A2(new_n702), .A3(new_n706), .A4(new_n717), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT36), .ZN(new_n719));
  INV_X1    g294(.A(G29), .ZN(new_n720));
  AND2_X1   g295(.A1(new_n720), .A2(G33), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n480), .A2(G139), .ZN(new_n722));
  XOR2_X1   g297(.A(new_n722), .B(KEYINPUT89), .Z(new_n723));
  NAND3_X1  g298(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT88), .ZN(new_n725));
  XNOR2_X1  g300(.A(KEYINPUT87), .B(KEYINPUT25), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n725), .B(new_n726), .ZN(new_n727));
  AOI22_X1  g302(.A1(new_n473), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n728));
  OAI211_X1 g303(.A(new_n723), .B(new_n727), .C1(new_n462), .C2(new_n728), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n721), .B1(new_n729), .B2(G29), .ZN(new_n730));
  INV_X1    g305(.A(G2072), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n720), .A2(G32), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n475), .A2(G129), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n480), .A2(G141), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n469), .A2(G105), .ZN(new_n736));
  NAND3_X1  g311(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT26), .Z(new_n738));
  NAND4_X1  g313(.A1(new_n734), .A2(new_n735), .A3(new_n736), .A4(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(new_n739), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n733), .B1(new_n740), .B2(new_n720), .ZN(new_n741));
  XNOR2_X1  g316(.A(KEYINPUT27), .B(G1996), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n741), .B(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(KEYINPUT24), .ZN(new_n744));
  INV_X1    g319(.A(G34), .ZN(new_n745));
  AOI21_X1  g320(.A(G29), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(new_n744), .B2(new_n745), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(G160), .B2(new_n720), .ZN(new_n748));
  OAI211_X1 g323(.A(new_n732), .B(new_n743), .C1(G2084), .C2(new_n748), .ZN(new_n749));
  NOR2_X1   g324(.A1(G171), .A2(new_n684), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(G5), .B2(new_n684), .ZN(new_n751));
  INV_X1    g326(.A(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n684), .A2(G20), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT23), .ZN(new_n754));
  AND2_X1   g329(.A1(new_n553), .A2(new_n558), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n754), .B1(new_n755), .B2(new_n684), .ZN(new_n756));
  INV_X1    g331(.A(new_n756), .ZN(new_n757));
  XOR2_X1   g332(.A(KEYINPUT93), .B(G1956), .Z(new_n758));
  AOI22_X1  g333(.A1(new_n752), .A2(G1961), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(new_n757), .B2(new_n758), .ZN(new_n760));
  OAI22_X1  g335(.A1(new_n730), .A2(new_n731), .B1(G1961), .B2(new_n752), .ZN(new_n761));
  NOR3_X1   g336(.A1(new_n749), .A2(new_n760), .A3(new_n761), .ZN(new_n762));
  NOR2_X1   g337(.A1(G164), .A2(new_n720), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(G27), .B2(new_n720), .ZN(new_n764));
  INV_X1    g339(.A(G2078), .ZN(new_n765));
  OR2_X1    g340(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n475), .A2(G128), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n480), .A2(G140), .ZN(new_n768));
  OR2_X1    g343(.A1(G104), .A2(G2105), .ZN(new_n769));
  OAI211_X1 g344(.A(new_n769), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n770));
  NAND3_X1  g345(.A1(new_n767), .A2(new_n768), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n771), .A2(G29), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n720), .A2(G26), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT28), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  INV_X1    g350(.A(G2067), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  XOR2_X1   g352(.A(KEYINPUT31), .B(G11), .Z(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT90), .ZN(new_n779));
  INV_X1    g354(.A(KEYINPUT30), .ZN(new_n780));
  AND2_X1   g355(.A1(new_n780), .A2(G28), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n720), .B1(new_n780), .B2(G28), .ZN(new_n782));
  OAI221_X1 g357(.A(new_n779), .B1(new_n781), .B2(new_n782), .C1(new_n628), .C2(new_n720), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(G2084), .B2(new_n748), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n764), .A2(new_n765), .ZN(new_n785));
  NAND4_X1  g360(.A1(new_n766), .A2(new_n777), .A3(new_n784), .A4(new_n785), .ZN(new_n786));
  NOR2_X1   g361(.A1(G29), .A2(G35), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(G162), .B2(G29), .ZN(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT92), .B(KEYINPUT29), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(G2090), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n788), .B(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n684), .A2(G21), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(G168), .B2(new_n684), .ZN(new_n793));
  AOI211_X1 g368(.A(new_n786), .B(new_n791), .C1(G1966), .C2(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(G16), .A2(G19), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(new_n540), .B2(G16), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT86), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(G1341), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n684), .A2(G4), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(new_n610), .B2(new_n684), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(G1348), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n798), .A2(new_n801), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n793), .A2(G1966), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT91), .ZN(new_n804));
  AND4_X1   g379(.A1(new_n762), .A2(new_n794), .A3(new_n802), .A4(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n719), .A2(new_n805), .ZN(G150));
  INV_X1    g381(.A(G150), .ZN(G311));
  NAND2_X1  g382(.A1(new_n610), .A2(G559), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT38), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n533), .A2(G93), .A3(new_n506), .ZN(new_n810));
  OAI211_X1 g385(.A(G55), .B(G543), .C1(new_n500), .C2(new_n501), .ZN(new_n811));
  NAND2_X1  g386(.A1(G80), .A2(G543), .ZN(new_n812));
  INV_X1    g387(.A(new_n812), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n813), .B1(new_n506), .B2(G67), .ZN(new_n814));
  OAI211_X1 g389(.A(new_n810), .B(new_n811), .C1(new_n814), .C2(new_n508), .ZN(new_n815));
  AND2_X1   g390(.A1(new_n539), .A2(new_n815), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n539), .A2(new_n815), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n809), .B(new_n818), .ZN(new_n819));
  AND2_X1   g394(.A1(new_n819), .A2(KEYINPUT39), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n819), .A2(KEYINPUT39), .ZN(new_n821));
  NOR3_X1   g396(.A1(new_n820), .A2(new_n821), .A3(G860), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n815), .A2(G860), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT37), .ZN(new_n824));
  OR2_X1    g399(.A1(new_n822), .A2(new_n824), .ZN(G145));
  XNOR2_X1  g400(.A(new_n771), .B(new_n490), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n729), .B(new_n826), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(new_n740), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n711), .B(new_n619), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n475), .A2(G130), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n480), .A2(G142), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT94), .ZN(new_n832));
  NOR3_X1   g407(.A1(new_n832), .A2(new_n462), .A3(G118), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n832), .B1(new_n462), .B2(G118), .ZN(new_n834));
  OR2_X1    g409(.A1(G106), .A2(G2105), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n834), .A2(G2104), .A3(new_n835), .ZN(new_n836));
  OAI211_X1 g411(.A(new_n830), .B(new_n831), .C1(new_n833), .C2(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n829), .B(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT95), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  OR2_X1    g415(.A1(new_n828), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n828), .A2(new_n840), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n628), .B(G160), .Z(new_n843));
  XNOR2_X1  g418(.A(G162), .B(new_n843), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n841), .A2(new_n842), .A3(new_n844), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n844), .B1(new_n828), .B2(new_n838), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n846), .B1(new_n828), .B2(new_n838), .ZN(new_n847));
  INV_X1    g422(.A(G37), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n845), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(KEYINPUT40), .ZN(G395));
  AND3_X1   g425(.A1(new_n755), .A2(new_n602), .A3(KEYINPUT97), .ZN(new_n851));
  AOI21_X1  g426(.A(KEYINPUT97), .B1(new_n755), .B2(new_n602), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n610), .A2(KEYINPUT96), .A3(G299), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT96), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n855), .B1(new_n755), .B2(new_n602), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n853), .A2(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(KEYINPUT98), .ZN(new_n859));
  XOR2_X1   g434(.A(new_n613), .B(new_n818), .Z(new_n860));
  INV_X1    g435(.A(KEYINPUT41), .ZN(new_n861));
  AOI21_X1  g436(.A(KEYINPUT96), .B1(new_n610), .B2(G299), .ZN(new_n862));
  AOI22_X1  g437(.A1(new_n594), .A2(new_n595), .B1(new_n599), .B2(new_n600), .ZN(new_n863));
  AND4_X1   g438(.A1(KEYINPUT96), .A2(G299), .A3(new_n863), .A4(new_n591), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT97), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n866), .B1(new_n610), .B2(G299), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n755), .A2(new_n602), .A3(KEYINPUT97), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n861), .B1(new_n865), .B2(new_n869), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n853), .A2(KEYINPUT41), .A3(new_n857), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n860), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT99), .ZN(new_n873));
  AOI22_X1  g448(.A1(new_n859), .A2(new_n860), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n872), .A2(new_n873), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(G305), .B(G303), .ZN(new_n878));
  INV_X1    g453(.A(G74), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n508), .B1(new_n547), .B2(new_n879), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n880), .B1(G87), .B2(new_n552), .ZN(new_n881));
  AOI22_X1  g456(.A1(new_n579), .A2(G651), .B1(new_n552), .B2(G85), .ZN(new_n882));
  NAND4_X1  g457(.A1(new_n881), .A2(new_n882), .A3(new_n564), .A4(new_n581), .ZN(new_n883));
  NAND2_X1  g458(.A1(G290), .A2(G288), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT100), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g462(.A(KEYINPUT100), .B1(new_n883), .B2(new_n884), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n878), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(new_n888), .ZN(new_n890));
  XNOR2_X1  g465(.A(G305), .B(G166), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n889), .A2(new_n892), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n893), .A2(KEYINPUT42), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(KEYINPUT101), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT101), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n889), .A2(new_n896), .A3(new_n892), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n894), .B1(new_n898), .B2(KEYINPUT42), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  OAI21_X1  g475(.A(KEYINPUT103), .B1(new_n877), .B2(new_n900), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n877), .A2(KEYINPUT102), .A3(new_n900), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT102), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n874), .B1(new_n873), .B2(new_n872), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n903), .B1(new_n904), .B2(new_n899), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT103), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n904), .A2(new_n906), .A3(new_n899), .ZN(new_n907));
  NAND4_X1  g482(.A1(new_n901), .A2(new_n902), .A3(new_n905), .A4(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(G868), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n815), .A2(new_n603), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(G295));
  NAND2_X1  g486(.A1(new_n909), .A2(new_n910), .ZN(G331));
  INV_X1    g487(.A(KEYINPUT44), .ZN(new_n913));
  AND3_X1   g488(.A1(new_n889), .A2(new_n896), .A3(new_n892), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n896), .B1(new_n889), .B2(new_n892), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(G64), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n917), .B1(new_n550), .B2(new_n551), .ZN(new_n918));
  INV_X1    g493(.A(new_n527), .ZN(new_n919));
  OAI21_X1  g494(.A(KEYINPUT75), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n920), .A2(G651), .A3(new_n531), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT104), .ZN(new_n922));
  AOI22_X1  g497(.A1(new_n552), .A2(G90), .B1(new_n497), .B2(G52), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n921), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(G168), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(KEYINPUT105), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT105), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n924), .A2(G168), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(G56), .ZN(new_n930));
  OAI22_X1  g505(.A1(new_n547), .A2(new_n930), .B1(new_n536), .B2(new_n492), .ZN(new_n931));
  AOI22_X1  g506(.A1(new_n931), .A2(G651), .B1(new_n552), .B2(G81), .ZN(new_n932));
  INV_X1    g507(.A(G67), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n812), .B1(new_n547), .B2(new_n933), .ZN(new_n934));
  AOI22_X1  g509(.A1(new_n934), .A2(G651), .B1(new_n552), .B2(G93), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n932), .A2(new_n935), .A3(new_n534), .A4(new_n811), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n539), .A2(new_n815), .ZN(new_n937));
  OAI211_X1 g512(.A(new_n936), .B(new_n937), .C1(new_n922), .C2(G171), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n922), .B1(new_n921), .B2(new_n923), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n939), .B1(new_n816), .B2(new_n817), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n929), .A2(new_n941), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n926), .A2(new_n938), .A3(new_n940), .A4(new_n928), .ZN(new_n943));
  AND2_X1   g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n870), .A2(new_n871), .ZN(new_n945));
  AND2_X1   g520(.A1(new_n945), .A2(KEYINPUT107), .ZN(new_n946));
  INV_X1    g521(.A(new_n871), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n944), .B1(new_n947), .B2(KEYINPUT107), .ZN(new_n948));
  OAI221_X1 g523(.A(new_n916), .B1(new_n859), .B2(new_n944), .C1(new_n946), .C2(new_n948), .ZN(new_n949));
  AOI22_X1  g524(.A1(new_n942), .A2(new_n943), .B1(new_n857), .B2(new_n853), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n950), .B1(new_n945), .B2(new_n944), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(new_n898), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n949), .A2(new_n848), .A3(new_n952), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n913), .B1(new_n953), .B2(KEYINPUT43), .ZN(new_n954));
  OAI211_X1 g529(.A(KEYINPUT106), .B(new_n848), .C1(new_n951), .C2(new_n898), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(new_n952), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n942), .A2(new_n943), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n957), .B1(new_n870), .B2(new_n871), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n916), .B1(new_n958), .B2(new_n950), .ZN(new_n959));
  AOI21_X1  g534(.A(KEYINPUT106), .B1(new_n959), .B2(new_n848), .ZN(new_n960));
  OR2_X1    g535(.A1(new_n956), .A2(new_n960), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n954), .B1(new_n961), .B2(KEYINPUT43), .ZN(new_n962));
  OAI21_X1  g537(.A(KEYINPUT43), .B1(new_n956), .B2(new_n960), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT43), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n949), .A2(new_n964), .A3(new_n848), .A4(new_n952), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(KEYINPUT108), .B1(new_n966), .B2(new_n913), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT108), .ZN(new_n968));
  AOI211_X1 g543(.A(new_n968), .B(KEYINPUT44), .C1(new_n963), .C2(new_n965), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n962), .B1(new_n967), .B2(new_n969), .ZN(G397));
  INV_X1    g545(.A(G8), .ZN(new_n971));
  NOR2_X1   g546(.A1(G168), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT50), .ZN(new_n974));
  INV_X1    g549(.A(G1384), .ZN(new_n975));
  AND3_X1   g550(.A1(new_n490), .A2(new_n974), .A3(new_n975), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n974), .B1(new_n490), .B2(new_n975), .ZN(new_n977));
  NAND2_X1  g552(.A1(G160), .A2(G40), .ZN(new_n978));
  NOR3_X1   g553(.A1(new_n976), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(G2084), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n490), .A2(new_n975), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT45), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(new_n978), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n490), .A2(KEYINPUT45), .A3(new_n975), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n983), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(G1966), .ZN(new_n987));
  AOI22_X1  g562(.A1(new_n979), .A2(new_n980), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  OAI211_X1 g563(.A(KEYINPUT51), .B(new_n973), .C1(new_n988), .C2(new_n971), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT51), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n986), .A2(new_n987), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n981), .A2(KEYINPUT50), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n490), .A2(new_n974), .A3(new_n975), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n992), .A2(new_n984), .A3(new_n980), .A4(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n991), .A2(new_n994), .ZN(new_n995));
  OAI211_X1 g570(.A(new_n990), .B(G8), .C1(new_n995), .C2(G286), .ZN(new_n996));
  AOI21_X1  g571(.A(KEYINPUT122), .B1(new_n995), .B2(new_n972), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT122), .ZN(new_n998));
  AOI211_X1 g573(.A(new_n998), .B(new_n973), .C1(new_n991), .C2(new_n994), .ZN(new_n999));
  OAI211_X1 g574(.A(new_n989), .B(new_n996), .C1(new_n997), .C2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(KEYINPUT123), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n998), .B1(new_n988), .B2(new_n973), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n995), .A2(KEYINPUT122), .A3(new_n972), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT123), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n1004), .A2(new_n1005), .A3(new_n989), .A4(new_n996), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1001), .A2(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g582(.A(KEYINPUT111), .B(G1971), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n986), .A2(new_n1009), .ZN(new_n1010));
  OR3_X1    g585(.A1(new_n977), .A2(KEYINPUT116), .A3(new_n978), .ZN(new_n1011));
  OAI21_X1  g586(.A(KEYINPUT116), .B1(new_n977), .B2(new_n978), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1011), .A2(new_n993), .A3(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1010), .B1(new_n1013), .B2(G2090), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(G8), .ZN(new_n1015));
  NAND3_X1  g590(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT112), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND4_X1  g593(.A1(G303), .A2(KEYINPUT112), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1019));
  NOR2_X1   g594(.A1(G166), .A2(new_n971), .ZN(new_n1020));
  OAI211_X1 g595(.A(new_n1018), .B(new_n1019), .C1(KEYINPUT55), .C2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1015), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(G2090), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n992), .A2(new_n984), .A3(new_n1024), .A4(new_n993), .ZN(new_n1025));
  AND3_X1   g600(.A1(new_n490), .A2(KEYINPUT45), .A3(new_n975), .ZN(new_n1026));
  AOI21_X1  g601(.A(KEYINPUT45), .B1(new_n490), .B2(new_n975), .ZN(new_n1027));
  NOR3_X1   g602(.A1(new_n1026), .A2(new_n1027), .A3(new_n978), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1025), .B1(new_n1028), .B2(new_n1008), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1029), .A2(G8), .A3(new_n1021), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(KEYINPUT113), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n971), .B1(new_n1010), .B2(new_n1025), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT113), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1032), .A2(new_n1033), .A3(new_n1021), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1031), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT114), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n490), .A2(G160), .A3(G40), .A4(new_n975), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1036), .B1(new_n1037), .B2(G8), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1037), .A2(new_n1036), .A3(G8), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n497), .A2(G48), .ZN(new_n1042));
  AOI22_X1  g617(.A1(new_n506), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1042), .B1(new_n1043), .B2(new_n508), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n504), .A2(new_n569), .ZN(new_n1045));
  OAI21_X1  g620(.A(G1981), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1046), .B1(G305), .B2(G1981), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(KEYINPUT115), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(KEYINPUT49), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT49), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1047), .A2(KEYINPUT115), .A3(new_n1050), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1041), .A2(new_n1049), .A3(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n686), .A2(G1976), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1040), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1053), .B1(new_n1054), .B2(new_n1038), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(KEYINPUT52), .ZN(new_n1056));
  INV_X1    g631(.A(G1976), .ZN(new_n1057));
  AOI21_X1  g632(.A(KEYINPUT52), .B1(G288), .B2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1041), .A2(new_n1053), .A3(new_n1058), .ZN(new_n1059));
  AND3_X1   g634(.A1(new_n1052), .A2(new_n1056), .A3(new_n1059), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n983), .A2(new_n984), .A3(new_n765), .A4(new_n985), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT53), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n992), .A2(new_n984), .A3(new_n993), .ZN(new_n1064));
  INV_X1    g639(.A(G1961), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1062), .A2(G2078), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(G40), .ZN(new_n1068));
  AOI21_X1  g643(.A(KEYINPUT124), .B1(new_n465), .B2(new_n466), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1069), .A2(new_n462), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n465), .A2(KEYINPUT124), .A3(new_n466), .ZN(new_n1071));
  AOI211_X1 g646(.A(new_n471), .B(new_n1068), .C1(new_n1070), .C2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1072), .A2(new_n983), .A3(new_n985), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1063), .A2(new_n1066), .A3(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(G171), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1028), .A2(new_n1067), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1076), .A2(new_n1063), .A3(G301), .A4(new_n1066), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1075), .A2(KEYINPUT54), .A3(new_n1077), .ZN(new_n1078));
  AND4_X1   g653(.A1(new_n1023), .A2(new_n1035), .A3(new_n1060), .A4(new_n1078), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1063), .A2(new_n1066), .A3(G301), .A4(new_n1073), .ZN(new_n1080));
  OR2_X1    g655(.A1(new_n1080), .A2(KEYINPUT125), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(KEYINPUT125), .ZN(new_n1082));
  AND2_X1   g657(.A1(new_n1063), .A2(new_n1066), .ZN(new_n1083));
  AND2_X1   g658(.A1(new_n1083), .A2(new_n1076), .ZN(new_n1084));
  OAI211_X1 g659(.A(new_n1081), .B(new_n1082), .C1(new_n1084), .C2(G301), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT54), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1007), .A2(new_n1079), .A3(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT126), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(G1956), .ZN(new_n1091));
  XNOR2_X1  g666(.A(KEYINPUT118), .B(KEYINPUT56), .ZN(new_n1092));
  XNOR2_X1  g667(.A(new_n1092), .B(new_n731), .ZN(new_n1093));
  AOI22_X1  g668(.A1(new_n1013), .A2(new_n1091), .B1(new_n1028), .B2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT117), .ZN(new_n1095));
  AOI21_X1  g670(.A(KEYINPUT57), .B1(new_n558), .B2(new_n1095), .ZN(new_n1096));
  XNOR2_X1  g671(.A(new_n1096), .B(G299), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1094), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(KEYINPUT119), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT119), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1094), .A2(new_n1100), .A3(new_n1097), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1102));
  OR2_X1    g677(.A1(new_n1037), .A2(KEYINPUT120), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1037), .A2(KEYINPUT120), .ZN(new_n1104));
  AOI21_X1  g679(.A(G2067), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n979), .A2(G1348), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1107), .A2(new_n602), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1094), .A2(new_n1097), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1102), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1109), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1111), .A2(KEYINPUT61), .A3(new_n1098), .ZN(new_n1112));
  NOR3_X1   g687(.A1(new_n1105), .A2(new_n1106), .A3(new_n610), .ZN(new_n1113));
  OAI21_X1  g688(.A(KEYINPUT60), .B1(new_n1108), .B2(new_n1113), .ZN(new_n1114));
  XOR2_X1   g689(.A(KEYINPUT58), .B(G1341), .Z(new_n1115));
  NAND3_X1  g690(.A1(new_n1103), .A2(new_n1104), .A3(new_n1115), .ZN(new_n1116));
  XOR2_X1   g691(.A(KEYINPUT121), .B(G1996), .Z(new_n1117));
  NAND2_X1  g692(.A1(new_n1028), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1119));
  AND3_X1   g694(.A1(new_n1119), .A2(KEYINPUT59), .A3(new_n540), .ZN(new_n1120));
  NOR4_X1   g695(.A1(new_n1105), .A2(new_n1106), .A3(KEYINPUT60), .A4(new_n602), .ZN(new_n1121));
  AOI21_X1  g696(.A(KEYINPUT59), .B1(new_n1119), .B2(new_n540), .ZN(new_n1122));
  NOR3_X1   g697(.A1(new_n1120), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1112), .A2(new_n1114), .A3(new_n1123), .ZN(new_n1124));
  AOI21_X1  g699(.A(KEYINPUT61), .B1(new_n1102), .B2(new_n1111), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1110), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1007), .A2(new_n1079), .A3(new_n1087), .A4(KEYINPUT126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1090), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1060), .ZN(new_n1129));
  NOR3_X1   g704(.A1(new_n988), .A2(new_n971), .A3(G286), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1130), .B1(new_n1021), .B2(new_n1032), .ZN(new_n1131));
  OAI21_X1  g706(.A(KEYINPUT63), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1132));
  AND3_X1   g707(.A1(new_n1052), .A2(new_n1057), .A3(new_n686), .ZN(new_n1133));
  NOR2_X1   g708(.A1(G305), .A2(G1981), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1041), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  NOR4_X1   g710(.A1(new_n988), .A2(KEYINPUT63), .A3(new_n971), .A4(G286), .ZN(new_n1136));
  AOI22_X1  g711(.A1(new_n1023), .A2(new_n1136), .B1(new_n1031), .B2(new_n1034), .ZN(new_n1137));
  OAI211_X1 g712(.A(new_n1132), .B(new_n1135), .C1(new_n1137), .C2(new_n1129), .ZN(new_n1138));
  OR2_X1    g713(.A1(new_n1007), .A2(KEYINPUT62), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1084), .A2(G301), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1140), .A2(new_n1023), .A3(new_n1060), .A4(new_n1035), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1141), .B1(new_n1007), .B2(KEYINPUT62), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1138), .B1(new_n1139), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1128), .A2(new_n1143), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n983), .A2(new_n978), .ZN(new_n1145));
  INV_X1    g720(.A(G1996), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n1147), .A2(new_n739), .ZN(new_n1148));
  XOR2_X1   g723(.A(new_n1148), .B(KEYINPUT109), .Z(new_n1149));
  XNOR2_X1  g724(.A(new_n771), .B(new_n776), .ZN(new_n1150));
  XNOR2_X1  g725(.A(new_n1150), .B(KEYINPUT110), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1151), .A2(new_n740), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1151), .A2(new_n1146), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1152), .A2(new_n1153), .A3(new_n1145), .ZN(new_n1154));
  INV_X1    g729(.A(new_n1145), .ZN(new_n1155));
  XNOR2_X1  g730(.A(new_n711), .B(new_n713), .ZN(new_n1156));
  OAI211_X1 g731(.A(new_n1149), .B(new_n1154), .C1(new_n1155), .C2(new_n1156), .ZN(new_n1157));
  XNOR2_X1  g732(.A(G290), .B(G1986), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1157), .B1(new_n1145), .B2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1144), .A2(new_n1159), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n711), .A2(new_n714), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1149), .A2(new_n1154), .A3(new_n1161), .ZN(new_n1162));
  OR2_X1    g737(.A1(new_n771), .A2(G2067), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1155), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  AND2_X1   g739(.A1(new_n1164), .A2(KEYINPUT127), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1152), .A2(new_n1145), .ZN(new_n1166));
  XNOR2_X1  g741(.A(new_n1147), .B(KEYINPUT46), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  XNOR2_X1  g743(.A(new_n1168), .B(KEYINPUT47), .ZN(new_n1169));
  NOR3_X1   g744(.A1(new_n1155), .A2(G1986), .A3(G290), .ZN(new_n1170));
  XNOR2_X1  g745(.A(new_n1170), .B(KEYINPUT48), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1169), .B1(new_n1157), .B2(new_n1171), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1164), .A2(KEYINPUT127), .ZN(new_n1173));
  NOR3_X1   g748(.A1(new_n1165), .A2(new_n1172), .A3(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1160), .A2(new_n1174), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g750(.A1(G229), .A2(new_n460), .A3(G401), .A4(G227), .ZN(new_n1177));
  NAND3_X1  g751(.A1(new_n1177), .A2(new_n849), .A3(new_n966), .ZN(G225));
  INV_X1    g752(.A(G225), .ZN(G308));
endmodule


