

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U550 ( .A(n734), .ZN(n713) );
  NAND2_X1 U551 ( .A1(G8), .A2(n707), .ZN(n769) );
  NOR2_X2 U552 ( .A1(n531), .A2(n530), .ZN(n532) );
  NOR2_X2 U553 ( .A1(n537), .A2(n536), .ZN(n538) );
  NOR2_X1 U554 ( .A1(n745), .A2(n693), .ZN(n694) );
  OR2_X1 U555 ( .A1(n751), .A2(n750), .ZN(n518) );
  OR2_X1 U556 ( .A1(n707), .A2(n942), .ZN(n708) );
  NOR2_X1 U557 ( .A1(n700), .A2(n699), .ZN(n701) );
  INV_X1 U558 ( .A(n961), .ZN(n753) );
  AND2_X1 U559 ( .A1(n754), .A2(n753), .ZN(n755) );
  INV_X1 U560 ( .A(KEYINPUT103), .ZN(n757) );
  XNOR2_X1 U561 ( .A(n758), .B(n757), .ZN(n759) );
  NOR2_X1 U562 ( .A1(G2104), .A2(G2105), .ZN(n523) );
  OR2_X1 U563 ( .A1(n768), .A2(n767), .ZN(n812) );
  NOR2_X2 U564 ( .A1(G2105), .A2(n519), .ZN(n887) );
  NOR2_X1 U565 ( .A1(G651), .A2(n650), .ZN(n661) );
  NOR2_X1 U566 ( .A1(n527), .A2(n526), .ZN(G160) );
  AND2_X2 U567 ( .A1(G2104), .A2(G2105), .ZN(n892) );
  NAND2_X1 U568 ( .A1(n892), .A2(G113), .ZN(n522) );
  INV_X1 U569 ( .A(G2104), .ZN(n519) );
  NAND2_X1 U570 ( .A1(G101), .A2(n887), .ZN(n520) );
  XOR2_X1 U571 ( .A(KEYINPUT23), .B(n520), .Z(n521) );
  NAND2_X1 U572 ( .A1(n522), .A2(n521), .ZN(n527) );
  AND2_X4 U573 ( .A1(n519), .A2(G2105), .ZN(n891) );
  NAND2_X1 U574 ( .A1(G125), .A2(n891), .ZN(n525) );
  XOR2_X2 U575 ( .A(KEYINPUT17), .B(n523), .Z(n886) );
  NAND2_X1 U576 ( .A1(G137), .A2(n886), .ZN(n524) );
  NAND2_X1 U577 ( .A1(n525), .A2(n524), .ZN(n526) );
  NAND2_X1 U578 ( .A1(n892), .A2(G114), .ZN(n528) );
  XNOR2_X1 U579 ( .A(KEYINPUT87), .B(n528), .ZN(n531) );
  NAND2_X1 U580 ( .A1(n891), .A2(G126), .ZN(n529) );
  XOR2_X1 U581 ( .A(n529), .B(KEYINPUT86), .Z(n530) );
  XNOR2_X1 U582 ( .A(n532), .B(KEYINPUT88), .ZN(n534) );
  NAND2_X1 U583 ( .A1(G102), .A2(n887), .ZN(n533) );
  NAND2_X1 U584 ( .A1(n534), .A2(n533), .ZN(n537) );
  NAND2_X1 U585 ( .A1(G138), .A2(n886), .ZN(n535) );
  XNOR2_X1 U586 ( .A(KEYINPUT89), .B(n535), .ZN(n536) );
  XNOR2_X1 U587 ( .A(n538), .B(KEYINPUT90), .ZN(n690) );
  BUF_X1 U588 ( .A(n690), .Z(G164) );
  NOR2_X1 U589 ( .A1(G651), .A2(G543), .ZN(n653) );
  NAND2_X1 U590 ( .A1(G85), .A2(n653), .ZN(n540) );
  XOR2_X1 U591 ( .A(KEYINPUT0), .B(G543), .Z(n650) );
  INV_X1 U592 ( .A(G651), .ZN(n541) );
  NOR2_X1 U593 ( .A1(n650), .A2(n541), .ZN(n657) );
  NAND2_X1 U594 ( .A1(G72), .A2(n657), .ZN(n539) );
  NAND2_X1 U595 ( .A1(n540), .A2(n539), .ZN(n546) );
  NOR2_X1 U596 ( .A1(G543), .A2(n541), .ZN(n542) );
  XOR2_X1 U597 ( .A(KEYINPUT1), .B(n542), .Z(n654) );
  NAND2_X1 U598 ( .A1(G60), .A2(n654), .ZN(n544) );
  NAND2_X1 U599 ( .A1(G47), .A2(n661), .ZN(n543) );
  NAND2_X1 U600 ( .A1(n544), .A2(n543), .ZN(n545) );
  OR2_X1 U601 ( .A1(n546), .A2(n545), .ZN(G290) );
  XOR2_X1 U602 ( .A(G2443), .B(G2446), .Z(n548) );
  XNOR2_X1 U603 ( .A(G2427), .B(G2451), .ZN(n547) );
  XNOR2_X1 U604 ( .A(n548), .B(n547), .ZN(n554) );
  XOR2_X1 U605 ( .A(G2430), .B(G2454), .Z(n550) );
  XNOR2_X1 U606 ( .A(G1341), .B(G1348), .ZN(n549) );
  XNOR2_X1 U607 ( .A(n550), .B(n549), .ZN(n552) );
  XOR2_X1 U608 ( .A(G2435), .B(G2438), .Z(n551) );
  XNOR2_X1 U609 ( .A(n552), .B(n551), .ZN(n553) );
  XOR2_X1 U610 ( .A(n554), .B(n553), .Z(n555) );
  AND2_X1 U611 ( .A1(G14), .A2(n555), .ZN(G401) );
  AND2_X1 U612 ( .A1(G452), .A2(G94), .ZN(G173) );
  XOR2_X1 U613 ( .A(KEYINPUT76), .B(KEYINPUT18), .Z(n557) );
  NAND2_X1 U614 ( .A1(G123), .A2(n891), .ZN(n556) );
  XNOR2_X1 U615 ( .A(n557), .B(n556), .ZN(n562) );
  NAND2_X1 U616 ( .A1(G111), .A2(n892), .ZN(n559) );
  NAND2_X1 U617 ( .A1(G99), .A2(n887), .ZN(n558) );
  NAND2_X1 U618 ( .A1(n559), .A2(n558), .ZN(n560) );
  XOR2_X1 U619 ( .A(KEYINPUT77), .B(n560), .Z(n561) );
  NOR2_X1 U620 ( .A1(n562), .A2(n561), .ZN(n564) );
  NAND2_X1 U621 ( .A1(n886), .A2(G135), .ZN(n563) );
  NAND2_X1 U622 ( .A1(n564), .A2(n563), .ZN(n918) );
  XNOR2_X1 U623 ( .A(G2096), .B(n918), .ZN(n565) );
  OR2_X1 U624 ( .A1(G2100), .A2(n565), .ZN(G156) );
  INV_X1 U625 ( .A(G57), .ZN(G237) );
  INV_X1 U626 ( .A(G132), .ZN(G219) );
  INV_X1 U627 ( .A(G82), .ZN(G220) );
  NAND2_X1 U628 ( .A1(G64), .A2(n654), .ZN(n567) );
  NAND2_X1 U629 ( .A1(G52), .A2(n661), .ZN(n566) );
  NAND2_X1 U630 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U631 ( .A(KEYINPUT64), .B(n568), .ZN(n575) );
  NAND2_X1 U632 ( .A1(n653), .A2(G90), .ZN(n569) );
  XNOR2_X1 U633 ( .A(KEYINPUT65), .B(n569), .ZN(n572) );
  NAND2_X1 U634 ( .A1(n657), .A2(G77), .ZN(n570) );
  XOR2_X1 U635 ( .A(KEYINPUT66), .B(n570), .Z(n571) );
  NOR2_X1 U636 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U637 ( .A(n573), .B(KEYINPUT9), .ZN(n574) );
  NOR2_X1 U638 ( .A1(n575), .A2(n574), .ZN(G171) );
  NAND2_X1 U639 ( .A1(G88), .A2(n653), .ZN(n577) );
  NAND2_X1 U640 ( .A1(G75), .A2(n657), .ZN(n576) );
  NAND2_X1 U641 ( .A1(n577), .A2(n576), .ZN(n581) );
  NAND2_X1 U642 ( .A1(G62), .A2(n654), .ZN(n579) );
  NAND2_X1 U643 ( .A1(G50), .A2(n661), .ZN(n578) );
  NAND2_X1 U644 ( .A1(n579), .A2(n578), .ZN(n580) );
  NOR2_X1 U645 ( .A1(n581), .A2(n580), .ZN(G166) );
  XNOR2_X1 U646 ( .A(KEYINPUT74), .B(KEYINPUT7), .ZN(n593) );
  NAND2_X1 U647 ( .A1(n653), .A2(G89), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n582), .B(KEYINPUT4), .ZN(n584) );
  NAND2_X1 U649 ( .A1(G76), .A2(n657), .ZN(n583) );
  NAND2_X1 U650 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U651 ( .A(n585), .B(KEYINPUT5), .ZN(n591) );
  XNOR2_X1 U652 ( .A(KEYINPUT73), .B(KEYINPUT6), .ZN(n589) );
  NAND2_X1 U653 ( .A1(G63), .A2(n654), .ZN(n587) );
  NAND2_X1 U654 ( .A1(G51), .A2(n661), .ZN(n586) );
  NAND2_X1 U655 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U656 ( .A(n589), .B(n588), .ZN(n590) );
  NAND2_X1 U657 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U658 ( .A(n593), .B(n592), .ZN(G168) );
  XOR2_X1 U659 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  XOR2_X1 U660 ( .A(KEYINPUT67), .B(KEYINPUT10), .Z(n595) );
  NAND2_X1 U661 ( .A1(G7), .A2(G661), .ZN(n594) );
  XNOR2_X1 U662 ( .A(n595), .B(n594), .ZN(G223) );
  XOR2_X1 U663 ( .A(G223), .B(KEYINPUT68), .Z(n828) );
  NAND2_X1 U664 ( .A1(n828), .A2(G567), .ZN(n596) );
  XNOR2_X1 U665 ( .A(n596), .B(KEYINPUT69), .ZN(n597) );
  XNOR2_X1 U666 ( .A(KEYINPUT11), .B(n597), .ZN(G234) );
  NAND2_X1 U667 ( .A1(n654), .A2(G56), .ZN(n598) );
  XOR2_X1 U668 ( .A(KEYINPUT14), .B(n598), .Z(n604) );
  NAND2_X1 U669 ( .A1(n653), .A2(G81), .ZN(n599) );
  XNOR2_X1 U670 ( .A(n599), .B(KEYINPUT12), .ZN(n601) );
  NAND2_X1 U671 ( .A1(G68), .A2(n657), .ZN(n600) );
  NAND2_X1 U672 ( .A1(n601), .A2(n600), .ZN(n602) );
  XOR2_X1 U673 ( .A(KEYINPUT13), .B(n602), .Z(n603) );
  NOR2_X1 U674 ( .A1(n604), .A2(n603), .ZN(n605) );
  XNOR2_X1 U675 ( .A(n605), .B(KEYINPUT70), .ZN(n607) );
  NAND2_X1 U676 ( .A1(G43), .A2(n661), .ZN(n606) );
  NAND2_X1 U677 ( .A1(n607), .A2(n606), .ZN(n980) );
  INV_X1 U678 ( .A(G860), .ZN(n628) );
  OR2_X1 U679 ( .A1(n980), .A2(n628), .ZN(n608) );
  XOR2_X1 U680 ( .A(KEYINPUT71), .B(n608), .Z(G153) );
  INV_X1 U681 ( .A(G171), .ZN(G301) );
  NAND2_X1 U682 ( .A1(G868), .A2(G301), .ZN(n618) );
  NAND2_X1 U683 ( .A1(G54), .A2(n661), .ZN(n615) );
  NAND2_X1 U684 ( .A1(G92), .A2(n653), .ZN(n610) );
  NAND2_X1 U685 ( .A1(G66), .A2(n654), .ZN(n609) );
  NAND2_X1 U686 ( .A1(n610), .A2(n609), .ZN(n613) );
  NAND2_X1 U687 ( .A1(n657), .A2(G79), .ZN(n611) );
  XOR2_X1 U688 ( .A(KEYINPUT72), .B(n611), .Z(n612) );
  NOR2_X1 U689 ( .A1(n613), .A2(n612), .ZN(n614) );
  NAND2_X1 U690 ( .A1(n615), .A2(n614), .ZN(n616) );
  XNOR2_X1 U691 ( .A(n616), .B(KEYINPUT15), .ZN(n970) );
  OR2_X1 U692 ( .A1(n970), .A2(G868), .ZN(n617) );
  NAND2_X1 U693 ( .A1(n618), .A2(n617), .ZN(G284) );
  NAND2_X1 U694 ( .A1(G65), .A2(n654), .ZN(n620) );
  NAND2_X1 U695 ( .A1(G53), .A2(n661), .ZN(n619) );
  NAND2_X1 U696 ( .A1(n620), .A2(n619), .ZN(n624) );
  NAND2_X1 U697 ( .A1(G91), .A2(n653), .ZN(n622) );
  NAND2_X1 U698 ( .A1(G78), .A2(n657), .ZN(n621) );
  NAND2_X1 U699 ( .A1(n622), .A2(n621), .ZN(n623) );
  NOR2_X1 U700 ( .A1(n624), .A2(n623), .ZN(n973) );
  INV_X1 U701 ( .A(n973), .ZN(G299) );
  INV_X1 U702 ( .A(G868), .ZN(n673) );
  NOR2_X1 U703 ( .A1(G286), .A2(n673), .ZN(n625) );
  XOR2_X1 U704 ( .A(KEYINPUT75), .B(n625), .Z(n627) );
  NOR2_X1 U705 ( .A1(G868), .A2(G299), .ZN(n626) );
  NOR2_X1 U706 ( .A1(n627), .A2(n626), .ZN(G297) );
  NAND2_X1 U707 ( .A1(n628), .A2(G559), .ZN(n629) );
  NAND2_X1 U708 ( .A1(n629), .A2(n970), .ZN(n630) );
  XNOR2_X1 U709 ( .A(n630), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U710 ( .A1(G868), .A2(n980), .ZN(n633) );
  NAND2_X1 U711 ( .A1(n970), .A2(G868), .ZN(n631) );
  NOR2_X1 U712 ( .A1(G559), .A2(n631), .ZN(n632) );
  NOR2_X1 U713 ( .A1(n633), .A2(n632), .ZN(G282) );
  NAND2_X1 U714 ( .A1(n657), .A2(G80), .ZN(n634) );
  XNOR2_X1 U715 ( .A(n634), .B(KEYINPUT80), .ZN(n636) );
  NAND2_X1 U716 ( .A1(G93), .A2(n653), .ZN(n635) );
  NAND2_X1 U717 ( .A1(n636), .A2(n635), .ZN(n637) );
  XNOR2_X1 U718 ( .A(n637), .B(KEYINPUT81), .ZN(n639) );
  NAND2_X1 U719 ( .A1(G55), .A2(n661), .ZN(n638) );
  NAND2_X1 U720 ( .A1(n639), .A2(n638), .ZN(n642) );
  NAND2_X1 U721 ( .A1(n654), .A2(G67), .ZN(n640) );
  XOR2_X1 U722 ( .A(KEYINPUT82), .B(n640), .Z(n641) );
  OR2_X1 U723 ( .A1(n642), .A2(n641), .ZN(n672) );
  NAND2_X1 U724 ( .A1(G559), .A2(n970), .ZN(n643) );
  XOR2_X1 U725 ( .A(n980), .B(n643), .Z(n670) );
  XOR2_X1 U726 ( .A(n670), .B(KEYINPUT78), .Z(n644) );
  NOR2_X1 U727 ( .A1(G860), .A2(n644), .ZN(n645) );
  XOR2_X1 U728 ( .A(KEYINPUT79), .B(n645), .Z(n646) );
  XOR2_X1 U729 ( .A(n672), .B(n646), .Z(G145) );
  NAND2_X1 U730 ( .A1(G49), .A2(n661), .ZN(n648) );
  NAND2_X1 U731 ( .A1(G74), .A2(G651), .ZN(n647) );
  NAND2_X1 U732 ( .A1(n648), .A2(n647), .ZN(n649) );
  NOR2_X1 U733 ( .A1(n654), .A2(n649), .ZN(n652) );
  NAND2_X1 U734 ( .A1(n650), .A2(G87), .ZN(n651) );
  NAND2_X1 U735 ( .A1(n652), .A2(n651), .ZN(G288) );
  NAND2_X1 U736 ( .A1(G86), .A2(n653), .ZN(n656) );
  NAND2_X1 U737 ( .A1(G61), .A2(n654), .ZN(n655) );
  NAND2_X1 U738 ( .A1(n656), .A2(n655), .ZN(n660) );
  NAND2_X1 U739 ( .A1(n657), .A2(G73), .ZN(n658) );
  XOR2_X1 U740 ( .A(KEYINPUT2), .B(n658), .Z(n659) );
  NOR2_X1 U741 ( .A1(n660), .A2(n659), .ZN(n663) );
  NAND2_X1 U742 ( .A1(n661), .A2(G48), .ZN(n662) );
  NAND2_X1 U743 ( .A1(n663), .A2(n662), .ZN(G305) );
  XNOR2_X1 U744 ( .A(G166), .B(G288), .ZN(n669) );
  XNOR2_X1 U745 ( .A(KEYINPUT83), .B(KEYINPUT19), .ZN(n665) );
  XOR2_X1 U746 ( .A(G290), .B(n672), .Z(n664) );
  XNOR2_X1 U747 ( .A(n665), .B(n664), .ZN(n666) );
  XNOR2_X1 U748 ( .A(n973), .B(n666), .ZN(n667) );
  XNOR2_X1 U749 ( .A(n667), .B(G305), .ZN(n668) );
  XNOR2_X1 U750 ( .A(n669), .B(n668), .ZN(n836) );
  XNOR2_X1 U751 ( .A(n836), .B(n670), .ZN(n671) );
  NAND2_X1 U752 ( .A1(n671), .A2(G868), .ZN(n675) );
  NAND2_X1 U753 ( .A1(n673), .A2(n672), .ZN(n674) );
  NAND2_X1 U754 ( .A1(n675), .A2(n674), .ZN(G295) );
  NAND2_X1 U755 ( .A1(G2078), .A2(G2084), .ZN(n677) );
  XOR2_X1 U756 ( .A(KEYINPUT84), .B(KEYINPUT20), .Z(n676) );
  XNOR2_X1 U757 ( .A(n677), .B(n676), .ZN(n678) );
  NAND2_X1 U758 ( .A1(G2090), .A2(n678), .ZN(n679) );
  XNOR2_X1 U759 ( .A(KEYINPUT21), .B(n679), .ZN(n680) );
  NAND2_X1 U760 ( .A1(n680), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U761 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U762 ( .A1(G220), .A2(G219), .ZN(n681) );
  XOR2_X1 U763 ( .A(KEYINPUT22), .B(n681), .Z(n682) );
  NOR2_X1 U764 ( .A1(G218), .A2(n682), .ZN(n683) );
  NAND2_X1 U765 ( .A1(G96), .A2(n683), .ZN(n834) );
  NAND2_X1 U766 ( .A1(n834), .A2(G2106), .ZN(n687) );
  NAND2_X1 U767 ( .A1(G69), .A2(G120), .ZN(n684) );
  NOR2_X1 U768 ( .A1(G237), .A2(n684), .ZN(n685) );
  NAND2_X1 U769 ( .A1(G108), .A2(n685), .ZN(n835) );
  NAND2_X1 U770 ( .A1(n835), .A2(G567), .ZN(n686) );
  NAND2_X1 U771 ( .A1(n687), .A2(n686), .ZN(n909) );
  NAND2_X1 U772 ( .A1(G483), .A2(G661), .ZN(n688) );
  NOR2_X1 U773 ( .A1(n909), .A2(n688), .ZN(n831) );
  NAND2_X1 U774 ( .A1(G36), .A2(n831), .ZN(n689) );
  XOR2_X1 U775 ( .A(KEYINPUT85), .B(n689), .Z(G176) );
  INV_X1 U776 ( .A(G166), .ZN(G303) );
  NOR2_X2 U777 ( .A1(n690), .A2(G1384), .ZN(n793) );
  NAND2_X1 U778 ( .A1(G160), .A2(G40), .ZN(n792) );
  INV_X1 U779 ( .A(n792), .ZN(n691) );
  NAND2_X2 U780 ( .A1(n793), .A2(n691), .ZN(n707) );
  BUF_X2 U781 ( .A(n707), .Z(n734) );
  NOR2_X1 U782 ( .A1(G2084), .A2(n734), .ZN(n745) );
  NOR2_X1 U783 ( .A1(n769), .A2(G1966), .ZN(n692) );
  XNOR2_X1 U784 ( .A(n692), .B(KEYINPUT97), .ZN(n743) );
  NAND2_X1 U785 ( .A1(n743), .A2(G8), .ZN(n693) );
  XOR2_X1 U786 ( .A(n694), .B(KEYINPUT30), .Z(n695) );
  NOR2_X1 U787 ( .A1(G168), .A2(n695), .ZN(n700) );
  XOR2_X1 U788 ( .A(G2078), .B(KEYINPUT25), .Z(n945) );
  NOR2_X1 U789 ( .A1(n945), .A2(n734), .ZN(n696) );
  XNOR2_X1 U790 ( .A(n696), .B(KEYINPUT98), .ZN(n698) );
  NOR2_X1 U791 ( .A1(n713), .A2(G1961), .ZN(n697) );
  NOR2_X1 U792 ( .A1(n698), .A2(n697), .ZN(n727) );
  AND2_X1 U793 ( .A1(G301), .A2(n727), .ZN(n699) );
  XNOR2_X1 U794 ( .A(n701), .B(KEYINPUT31), .ZN(n731) );
  NAND2_X1 U795 ( .A1(n713), .A2(G2072), .ZN(n702) );
  XNOR2_X1 U796 ( .A(n702), .B(KEYINPUT27), .ZN(n704) );
  INV_X1 U797 ( .A(G1956), .ZN(n990) );
  NOR2_X1 U798 ( .A1(n990), .A2(n713), .ZN(n703) );
  NOR2_X1 U799 ( .A1(n704), .A2(n703), .ZN(n721) );
  NOR2_X1 U800 ( .A1(n973), .A2(n721), .ZN(n706) );
  XNOR2_X1 U801 ( .A(KEYINPUT99), .B(KEYINPUT28), .ZN(n705) );
  XNOR2_X1 U802 ( .A(n706), .B(n705), .ZN(n725) );
  INV_X1 U803 ( .A(G1996), .ZN(n942) );
  XNOR2_X1 U804 ( .A(n708), .B(KEYINPUT26), .ZN(n710) );
  NAND2_X1 U805 ( .A1(n734), .A2(G1341), .ZN(n709) );
  NAND2_X1 U806 ( .A1(n710), .A2(n709), .ZN(n711) );
  NOR2_X1 U807 ( .A1(n980), .A2(n711), .ZN(n718) );
  NAND2_X1 U808 ( .A1(n970), .A2(n718), .ZN(n717) );
  NAND2_X1 U809 ( .A1(n734), .A2(G1348), .ZN(n712) );
  XNOR2_X1 U810 ( .A(n712), .B(KEYINPUT100), .ZN(n715) );
  NAND2_X1 U811 ( .A1(n713), .A2(G2067), .ZN(n714) );
  NAND2_X1 U812 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U813 ( .A1(n717), .A2(n716), .ZN(n720) );
  OR2_X1 U814 ( .A1(n970), .A2(n718), .ZN(n719) );
  NAND2_X1 U815 ( .A1(n720), .A2(n719), .ZN(n723) );
  NAND2_X1 U816 ( .A1(n973), .A2(n721), .ZN(n722) );
  NAND2_X1 U817 ( .A1(n723), .A2(n722), .ZN(n724) );
  NAND2_X1 U818 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U819 ( .A(n726), .B(KEYINPUT29), .ZN(n729) );
  NOR2_X1 U820 ( .A1(G301), .A2(n727), .ZN(n728) );
  NOR2_X1 U821 ( .A1(n729), .A2(n728), .ZN(n730) );
  NOR2_X1 U822 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U823 ( .A(n732), .B(KEYINPUT101), .ZN(n744) );
  AND2_X1 U824 ( .A1(G286), .A2(G8), .ZN(n733) );
  NAND2_X1 U825 ( .A1(n744), .A2(n733), .ZN(n741) );
  INV_X1 U826 ( .A(G8), .ZN(n739) );
  NOR2_X1 U827 ( .A1(G1971), .A2(n769), .ZN(n736) );
  NOR2_X1 U828 ( .A1(G2090), .A2(n734), .ZN(n735) );
  NOR2_X1 U829 ( .A1(n736), .A2(n735), .ZN(n737) );
  NAND2_X1 U830 ( .A1(n737), .A2(G303), .ZN(n738) );
  OR2_X1 U831 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U832 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U833 ( .A(KEYINPUT32), .B(n742), .ZN(n751) );
  INV_X1 U834 ( .A(n743), .ZN(n749) );
  BUF_X1 U835 ( .A(n744), .Z(n747) );
  NAND2_X1 U836 ( .A1(G8), .A2(n745), .ZN(n746) );
  NAND2_X1 U837 ( .A1(n747), .A2(n746), .ZN(n748) );
  NOR2_X1 U838 ( .A1(n749), .A2(n748), .ZN(n750) );
  NOR2_X1 U839 ( .A1(G1971), .A2(G303), .ZN(n752) );
  XOR2_X1 U840 ( .A(n752), .B(KEYINPUT102), .Z(n754) );
  NOR2_X1 U841 ( .A1(G1976), .A2(G288), .ZN(n961) );
  NAND2_X1 U842 ( .A1(n518), .A2(n755), .ZN(n756) );
  NAND2_X1 U843 ( .A1(G1976), .A2(G288), .ZN(n962) );
  NAND2_X1 U844 ( .A1(n756), .A2(n962), .ZN(n758) );
  NOR2_X1 U845 ( .A1(n769), .A2(n759), .ZN(n768) );
  NOR2_X1 U846 ( .A1(G2090), .A2(G303), .ZN(n760) );
  NAND2_X1 U847 ( .A1(G8), .A2(n760), .ZN(n761) );
  NAND2_X1 U848 ( .A1(n518), .A2(n761), .ZN(n762) );
  NAND2_X1 U849 ( .A1(n762), .A2(n769), .ZN(n766) );
  NOR2_X1 U850 ( .A1(G1981), .A2(G305), .ZN(n763) );
  XOR2_X1 U851 ( .A(n763), .B(KEYINPUT24), .Z(n764) );
  OR2_X1 U852 ( .A1(n769), .A2(n764), .ZN(n765) );
  NAND2_X1 U853 ( .A1(n766), .A2(n765), .ZN(n774) );
  OR2_X2 U854 ( .A1(KEYINPUT33), .A2(n774), .ZN(n767) );
  NAND2_X1 U855 ( .A1(n961), .A2(KEYINPUT33), .ZN(n770) );
  NOR2_X1 U856 ( .A1(n770), .A2(n769), .ZN(n772) );
  XOR2_X1 U857 ( .A(G1981), .B(G305), .Z(n967) );
  INV_X1 U858 ( .A(n967), .ZN(n771) );
  NOR2_X1 U859 ( .A1(n772), .A2(n771), .ZN(n773) );
  OR2_X1 U860 ( .A1(n774), .A2(n773), .ZN(n796) );
  XOR2_X1 U861 ( .A(KEYINPUT94), .B(G1991), .Z(n940) );
  NAND2_X1 U862 ( .A1(G119), .A2(n891), .ZN(n776) );
  NAND2_X1 U863 ( .A1(G107), .A2(n892), .ZN(n775) );
  NAND2_X1 U864 ( .A1(n776), .A2(n775), .ZN(n780) );
  NAND2_X1 U865 ( .A1(G131), .A2(n886), .ZN(n778) );
  NAND2_X1 U866 ( .A1(G95), .A2(n887), .ZN(n777) );
  NAND2_X1 U867 ( .A1(n778), .A2(n777), .ZN(n779) );
  NOR2_X1 U868 ( .A1(n780), .A2(n779), .ZN(n781) );
  XOR2_X1 U869 ( .A(KEYINPUT93), .B(n781), .Z(n873) );
  NOR2_X1 U870 ( .A1(n940), .A2(n873), .ZN(n791) );
  NAND2_X1 U871 ( .A1(G105), .A2(n887), .ZN(n782) );
  XNOR2_X1 U872 ( .A(n782), .B(KEYINPUT38), .ZN(n789) );
  NAND2_X1 U873 ( .A1(G117), .A2(n892), .ZN(n784) );
  NAND2_X1 U874 ( .A1(G141), .A2(n886), .ZN(n783) );
  NAND2_X1 U875 ( .A1(n784), .A2(n783), .ZN(n787) );
  NAND2_X1 U876 ( .A1(G129), .A2(n891), .ZN(n785) );
  XNOR2_X1 U877 ( .A(KEYINPUT95), .B(n785), .ZN(n786) );
  NOR2_X1 U878 ( .A1(n787), .A2(n786), .ZN(n788) );
  NAND2_X1 U879 ( .A1(n789), .A2(n788), .ZN(n874) );
  AND2_X1 U880 ( .A1(n874), .A2(G1996), .ZN(n790) );
  NOR2_X1 U881 ( .A1(n791), .A2(n790), .ZN(n923) );
  NOR2_X1 U882 ( .A1(n793), .A2(n792), .ZN(n822) );
  XOR2_X1 U883 ( .A(n822), .B(KEYINPUT96), .Z(n794) );
  NOR2_X1 U884 ( .A1(n923), .A2(n794), .ZN(n815) );
  INV_X1 U885 ( .A(n815), .ZN(n795) );
  NAND2_X1 U886 ( .A1(n796), .A2(n795), .ZN(n810) );
  XNOR2_X1 U887 ( .A(G2067), .B(KEYINPUT37), .ZN(n797) );
  XOR2_X1 U888 ( .A(n797), .B(KEYINPUT91), .Z(n820) );
  NAND2_X1 U889 ( .A1(G128), .A2(n891), .ZN(n799) );
  NAND2_X1 U890 ( .A1(G116), .A2(n892), .ZN(n798) );
  NAND2_X1 U891 ( .A1(n799), .A2(n798), .ZN(n800) );
  XNOR2_X1 U892 ( .A(n800), .B(KEYINPUT35), .ZN(n805) );
  NAND2_X1 U893 ( .A1(G140), .A2(n886), .ZN(n802) );
  NAND2_X1 U894 ( .A1(G104), .A2(n887), .ZN(n801) );
  NAND2_X1 U895 ( .A1(n802), .A2(n801), .ZN(n803) );
  XOR2_X1 U896 ( .A(KEYINPUT34), .B(n803), .Z(n804) );
  NAND2_X1 U897 ( .A1(n805), .A2(n804), .ZN(n806) );
  XOR2_X1 U898 ( .A(n806), .B(KEYINPUT36), .Z(n898) );
  OR2_X1 U899 ( .A1(n820), .A2(n898), .ZN(n807) );
  XNOR2_X1 U900 ( .A(n807), .B(KEYINPUT92), .ZN(n931) );
  XOR2_X1 U901 ( .A(G1986), .B(G290), .Z(n974) );
  NAND2_X1 U902 ( .A1(n931), .A2(n974), .ZN(n808) );
  AND2_X1 U903 ( .A1(n808), .A2(n822), .ZN(n809) );
  NOR2_X1 U904 ( .A1(n810), .A2(n809), .ZN(n811) );
  NAND2_X1 U905 ( .A1(n812), .A2(n811), .ZN(n825) );
  NOR2_X1 U906 ( .A1(G1996), .A2(n874), .ZN(n912) );
  AND2_X1 U907 ( .A1(n940), .A2(n873), .ZN(n921) );
  NOR2_X1 U908 ( .A1(G1986), .A2(G290), .ZN(n813) );
  NOR2_X1 U909 ( .A1(n921), .A2(n813), .ZN(n814) );
  NOR2_X1 U910 ( .A1(n815), .A2(n814), .ZN(n816) );
  XNOR2_X1 U911 ( .A(n816), .B(KEYINPUT104), .ZN(n817) );
  NOR2_X1 U912 ( .A1(n912), .A2(n817), .ZN(n818) );
  XNOR2_X1 U913 ( .A(KEYINPUT39), .B(n818), .ZN(n819) );
  NAND2_X1 U914 ( .A1(n819), .A2(n931), .ZN(n821) );
  NAND2_X1 U915 ( .A1(n898), .A2(n820), .ZN(n917) );
  NAND2_X1 U916 ( .A1(n821), .A2(n917), .ZN(n823) );
  NAND2_X1 U917 ( .A1(n823), .A2(n822), .ZN(n824) );
  NAND2_X1 U918 ( .A1(n825), .A2(n824), .ZN(n827) );
  XOR2_X1 U919 ( .A(KEYINPUT105), .B(KEYINPUT40), .Z(n826) );
  XNOR2_X1 U920 ( .A(n827), .B(n826), .ZN(G329) );
  NAND2_X1 U921 ( .A1(n828), .A2(G2106), .ZN(n829) );
  XNOR2_X1 U922 ( .A(n829), .B(KEYINPUT106), .ZN(G217) );
  AND2_X1 U923 ( .A1(G15), .A2(G2), .ZN(n830) );
  NAND2_X1 U924 ( .A1(G661), .A2(n830), .ZN(G259) );
  NAND2_X1 U925 ( .A1(G3), .A2(G1), .ZN(n832) );
  NAND2_X1 U926 ( .A1(n832), .A2(n831), .ZN(n833) );
  XOR2_X1 U927 ( .A(KEYINPUT107), .B(n833), .Z(G188) );
  INV_X1 U929 ( .A(G120), .ZN(G236) );
  INV_X1 U930 ( .A(G96), .ZN(G221) );
  INV_X1 U931 ( .A(G69), .ZN(G235) );
  NOR2_X1 U932 ( .A1(n835), .A2(n834), .ZN(G325) );
  INV_X1 U933 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U934 ( .A(G286), .B(n836), .ZN(n838) );
  XNOR2_X1 U935 ( .A(G171), .B(n970), .ZN(n837) );
  XNOR2_X1 U936 ( .A(n838), .B(n837), .ZN(n839) );
  XNOR2_X1 U937 ( .A(n839), .B(n980), .ZN(n840) );
  NOR2_X1 U938 ( .A1(G37), .A2(n840), .ZN(G397) );
  XNOR2_X1 U939 ( .A(G1961), .B(G2474), .ZN(n850) );
  XOR2_X1 U940 ( .A(G1981), .B(G1971), .Z(n842) );
  XNOR2_X1 U941 ( .A(G1966), .B(G1956), .ZN(n841) );
  XNOR2_X1 U942 ( .A(n842), .B(n841), .ZN(n846) );
  XOR2_X1 U943 ( .A(G1976), .B(G1986), .Z(n844) );
  XNOR2_X1 U944 ( .A(G1996), .B(G1991), .ZN(n843) );
  XNOR2_X1 U945 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U946 ( .A(n846), .B(n845), .Z(n848) );
  XNOR2_X1 U947 ( .A(KEYINPUT108), .B(KEYINPUT41), .ZN(n847) );
  XNOR2_X1 U948 ( .A(n848), .B(n847), .ZN(n849) );
  XNOR2_X1 U949 ( .A(n850), .B(n849), .ZN(G229) );
  XOR2_X1 U950 ( .A(G2100), .B(G2096), .Z(n852) );
  XNOR2_X1 U951 ( .A(KEYINPUT42), .B(G2678), .ZN(n851) );
  XNOR2_X1 U952 ( .A(n852), .B(n851), .ZN(n856) );
  XOR2_X1 U953 ( .A(KEYINPUT43), .B(G2090), .Z(n854) );
  XNOR2_X1 U954 ( .A(G2067), .B(G2072), .ZN(n853) );
  XNOR2_X1 U955 ( .A(n854), .B(n853), .ZN(n855) );
  XOR2_X1 U956 ( .A(n856), .B(n855), .Z(n858) );
  XNOR2_X1 U957 ( .A(G2078), .B(G2084), .ZN(n857) );
  XNOR2_X1 U958 ( .A(n858), .B(n857), .ZN(G227) );
  NAND2_X1 U959 ( .A1(G124), .A2(n891), .ZN(n859) );
  XOR2_X1 U960 ( .A(KEYINPUT109), .B(n859), .Z(n860) );
  XNOR2_X1 U961 ( .A(n860), .B(KEYINPUT44), .ZN(n862) );
  NAND2_X1 U962 ( .A1(G112), .A2(n892), .ZN(n861) );
  NAND2_X1 U963 ( .A1(n862), .A2(n861), .ZN(n866) );
  NAND2_X1 U964 ( .A1(G136), .A2(n886), .ZN(n864) );
  NAND2_X1 U965 ( .A1(G100), .A2(n887), .ZN(n863) );
  NAND2_X1 U966 ( .A1(n864), .A2(n863), .ZN(n865) );
  NOR2_X1 U967 ( .A1(n866), .A2(n865), .ZN(G162) );
  XOR2_X1 U968 ( .A(KEYINPUT112), .B(KEYINPUT113), .Z(n868) );
  XNOR2_X1 U969 ( .A(G160), .B(KEYINPUT48), .ZN(n867) );
  XNOR2_X1 U970 ( .A(n868), .B(n867), .ZN(n869) );
  XNOR2_X1 U971 ( .A(KEYINPUT46), .B(n869), .ZN(n871) );
  XNOR2_X1 U972 ( .A(n918), .B(KEYINPUT111), .ZN(n870) );
  XNOR2_X1 U973 ( .A(n871), .B(n870), .ZN(n872) );
  XOR2_X1 U974 ( .A(n872), .B(G162), .Z(n876) );
  XOR2_X1 U975 ( .A(n874), .B(n873), .Z(n875) );
  XNOR2_X1 U976 ( .A(n876), .B(n875), .ZN(n885) );
  NAND2_X1 U977 ( .A1(G130), .A2(n891), .ZN(n878) );
  NAND2_X1 U978 ( .A1(G118), .A2(n892), .ZN(n877) );
  NAND2_X1 U979 ( .A1(n878), .A2(n877), .ZN(n883) );
  NAND2_X1 U980 ( .A1(G142), .A2(n886), .ZN(n880) );
  NAND2_X1 U981 ( .A1(G106), .A2(n887), .ZN(n879) );
  NAND2_X1 U982 ( .A1(n880), .A2(n879), .ZN(n881) );
  XOR2_X1 U983 ( .A(KEYINPUT45), .B(n881), .Z(n882) );
  NOR2_X1 U984 ( .A1(n883), .A2(n882), .ZN(n884) );
  XOR2_X1 U985 ( .A(n885), .B(n884), .Z(n900) );
  NAND2_X1 U986 ( .A1(G139), .A2(n886), .ZN(n889) );
  NAND2_X1 U987 ( .A1(G103), .A2(n887), .ZN(n888) );
  NAND2_X1 U988 ( .A1(n889), .A2(n888), .ZN(n890) );
  XNOR2_X1 U989 ( .A(KEYINPUT110), .B(n890), .ZN(n897) );
  NAND2_X1 U990 ( .A1(G127), .A2(n891), .ZN(n894) );
  NAND2_X1 U991 ( .A1(G115), .A2(n892), .ZN(n893) );
  NAND2_X1 U992 ( .A1(n894), .A2(n893), .ZN(n895) );
  XOR2_X1 U993 ( .A(KEYINPUT47), .B(n895), .Z(n896) );
  NOR2_X1 U994 ( .A1(n897), .A2(n896), .ZN(n924) );
  XOR2_X1 U995 ( .A(n898), .B(n924), .Z(n899) );
  XNOR2_X1 U996 ( .A(n900), .B(n899), .ZN(n901) );
  XOR2_X1 U997 ( .A(n901), .B(G164), .Z(n902) );
  NOR2_X1 U998 ( .A1(G37), .A2(n902), .ZN(G395) );
  NOR2_X1 U999 ( .A1(G401), .A2(n909), .ZN(n906) );
  NOR2_X1 U1000 ( .A1(G229), .A2(G227), .ZN(n903) );
  XNOR2_X1 U1001 ( .A(KEYINPUT49), .B(n903), .ZN(n904) );
  NOR2_X1 U1002 ( .A1(G397), .A2(n904), .ZN(n905) );
  NAND2_X1 U1003 ( .A1(n906), .A2(n905), .ZN(n907) );
  NOR2_X1 U1004 ( .A1(n907), .A2(G395), .ZN(n908) );
  XNOR2_X1 U1005 ( .A(n908), .B(KEYINPUT114), .ZN(G308) );
  INV_X1 U1006 ( .A(G308), .ZN(G225) );
  INV_X1 U1007 ( .A(n909), .ZN(G319) );
  INV_X1 U1008 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1009 ( .A(KEYINPUT51), .B(KEYINPUT117), .Z(n910) );
  XNOR2_X1 U1010 ( .A(KEYINPUT116), .B(n910), .ZN(n915) );
  XNOR2_X1 U1011 ( .A(G2090), .B(G162), .ZN(n911) );
  XNOR2_X1 U1012 ( .A(n911), .B(KEYINPUT115), .ZN(n913) );
  NOR2_X1 U1013 ( .A1(n913), .A2(n912), .ZN(n914) );
  XOR2_X1 U1014 ( .A(n915), .B(n914), .Z(n916) );
  NAND2_X1 U1015 ( .A1(n917), .A2(n916), .ZN(n933) );
  XNOR2_X1 U1016 ( .A(G160), .B(G2084), .ZN(n919) );
  NAND2_X1 U1017 ( .A1(n919), .A2(n918), .ZN(n920) );
  NOR2_X1 U1018 ( .A1(n921), .A2(n920), .ZN(n922) );
  NAND2_X1 U1019 ( .A1(n923), .A2(n922), .ZN(n929) );
  XOR2_X1 U1020 ( .A(G2072), .B(n924), .Z(n926) );
  XOR2_X1 U1021 ( .A(G164), .B(G2078), .Z(n925) );
  NOR2_X1 U1022 ( .A1(n926), .A2(n925), .ZN(n927) );
  XOR2_X1 U1023 ( .A(KEYINPUT50), .B(n927), .Z(n928) );
  NOR2_X1 U1024 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1025 ( .A1(n931), .A2(n930), .ZN(n932) );
  NOR2_X1 U1026 ( .A1(n933), .A2(n932), .ZN(n934) );
  XOR2_X1 U1027 ( .A(KEYINPUT52), .B(n934), .Z(n935) );
  NOR2_X1 U1028 ( .A1(KEYINPUT55), .A2(n935), .ZN(n936) );
  XOR2_X1 U1029 ( .A(KEYINPUT118), .B(n936), .Z(n937) );
  NAND2_X1 U1030 ( .A1(G29), .A2(n937), .ZN(n938) );
  XOR2_X1 U1031 ( .A(KEYINPUT119), .B(n938), .Z(n1019) );
  XOR2_X1 U1032 ( .A(G2072), .B(G33), .Z(n939) );
  NAND2_X1 U1033 ( .A1(n939), .A2(G28), .ZN(n951) );
  XNOR2_X1 U1034 ( .A(KEYINPUT120), .B(n940), .ZN(n941) );
  XNOR2_X1 U1035 ( .A(n941), .B(G25), .ZN(n949) );
  XOR2_X1 U1036 ( .A(G2067), .B(G26), .Z(n944) );
  XNOR2_X1 U1037 ( .A(n942), .B(G32), .ZN(n943) );
  NAND2_X1 U1038 ( .A1(n944), .A2(n943), .ZN(n947) );
  XNOR2_X1 U1039 ( .A(G27), .B(n945), .ZN(n946) );
  NOR2_X1 U1040 ( .A1(n947), .A2(n946), .ZN(n948) );
  NAND2_X1 U1041 ( .A1(n949), .A2(n948), .ZN(n950) );
  NOR2_X1 U1042 ( .A1(n951), .A2(n950), .ZN(n952) );
  XOR2_X1 U1043 ( .A(KEYINPUT53), .B(n952), .Z(n956) );
  XNOR2_X1 U1044 ( .A(KEYINPUT54), .B(G34), .ZN(n953) );
  XNOR2_X1 U1045 ( .A(n953), .B(KEYINPUT121), .ZN(n954) );
  XNOR2_X1 U1046 ( .A(G2084), .B(n954), .ZN(n955) );
  NAND2_X1 U1047 ( .A1(n956), .A2(n955), .ZN(n958) );
  XNOR2_X1 U1048 ( .A(G35), .B(G2090), .ZN(n957) );
  NOR2_X1 U1049 ( .A1(n958), .A2(n957), .ZN(n959) );
  XOR2_X1 U1050 ( .A(KEYINPUT55), .B(n959), .Z(n960) );
  NOR2_X1 U1051 ( .A1(G29), .A2(n960), .ZN(n1015) );
  XNOR2_X1 U1052 ( .A(G16), .B(KEYINPUT56), .ZN(n986) );
  XNOR2_X1 U1053 ( .A(G166), .B(G1971), .ZN(n965) );
  NAND2_X1 U1054 ( .A1(n753), .A2(n962), .ZN(n963) );
  XOR2_X1 U1055 ( .A(KEYINPUT122), .B(n963), .Z(n964) );
  NAND2_X1 U1056 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1057 ( .A(n966), .B(KEYINPUT123), .ZN(n984) );
  XNOR2_X1 U1058 ( .A(G1966), .B(G168), .ZN(n968) );
  NAND2_X1 U1059 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1060 ( .A(KEYINPUT57), .B(n969), .ZN(n979) );
  XNOR2_X1 U1061 ( .A(n970), .B(G1348), .ZN(n972) );
  XNOR2_X1 U1062 ( .A(G171), .B(G1961), .ZN(n971) );
  NAND2_X1 U1063 ( .A1(n972), .A2(n971), .ZN(n977) );
  XNOR2_X1 U1064 ( .A(n973), .B(G1956), .ZN(n975) );
  NAND2_X1 U1065 ( .A1(n975), .A2(n974), .ZN(n976) );
  NOR2_X1 U1066 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1067 ( .A1(n979), .A2(n978), .ZN(n982) );
  XNOR2_X1 U1068 ( .A(G1341), .B(n980), .ZN(n981) );
  NOR2_X1 U1069 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1070 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1071 ( .A1(n986), .A2(n985), .ZN(n1013) );
  INV_X1 U1072 ( .A(G16), .ZN(n1011) );
  XNOR2_X1 U1073 ( .A(G1341), .B(G19), .ZN(n988) );
  XNOR2_X1 U1074 ( .A(G1981), .B(G6), .ZN(n987) );
  NOR2_X1 U1075 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1076 ( .A(KEYINPUT124), .B(n989), .ZN(n992) );
  XNOR2_X1 U1077 ( .A(n990), .B(G20), .ZN(n991) );
  NAND2_X1 U1078 ( .A1(n992), .A2(n991), .ZN(n995) );
  XOR2_X1 U1079 ( .A(KEYINPUT59), .B(G1348), .Z(n993) );
  XNOR2_X1 U1080 ( .A(G4), .B(n993), .ZN(n994) );
  NOR2_X1 U1081 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1082 ( .A(KEYINPUT60), .B(n996), .ZN(n1000) );
  XNOR2_X1 U1083 ( .A(G1966), .B(G21), .ZN(n998) );
  XNOR2_X1 U1084 ( .A(G1961), .B(G5), .ZN(n997) );
  NOR2_X1 U1085 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1086 ( .A1(n1000), .A2(n999), .ZN(n1008) );
  XNOR2_X1 U1087 ( .A(G1986), .B(G24), .ZN(n1002) );
  XNOR2_X1 U1088 ( .A(G23), .B(G1976), .ZN(n1001) );
  NOR2_X1 U1089 ( .A1(n1002), .A2(n1001), .ZN(n1005) );
  XNOR2_X1 U1090 ( .A(G1971), .B(KEYINPUT125), .ZN(n1003) );
  XNOR2_X1 U1091 ( .A(n1003), .B(G22), .ZN(n1004) );
  NAND2_X1 U1092 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XNOR2_X1 U1093 ( .A(KEYINPUT58), .B(n1006), .ZN(n1007) );
  NOR2_X1 U1094 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1095 ( .A(KEYINPUT61), .B(n1009), .ZN(n1010) );
  NAND2_X1 U1096 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1097 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NOR2_X1 U1098 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1099 ( .A1(G11), .A2(n1016), .ZN(n1017) );
  XOR2_X1 U1100 ( .A(KEYINPUT126), .B(n1017), .Z(n1018) );
  NAND2_X1 U1101 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1102 ( .A(n1020), .B(KEYINPUT127), .ZN(n1021) );
  XNOR2_X1 U1103 ( .A(KEYINPUT62), .B(n1021), .ZN(G311) );
  INV_X1 U1104 ( .A(G311), .ZN(G150) );
endmodule

