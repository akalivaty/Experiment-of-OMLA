

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773;

  XNOR2_X1 U380 ( .A(n495), .B(n494), .ZN(n529) );
  NAND2_X1 U381 ( .A1(n770), .A2(KEYINPUT44), .ZN(n649) );
  XNOR2_X1 U382 ( .A(n415), .B(G953), .ZN(n498) );
  NOR2_X1 U383 ( .A1(n658), .A2(n747), .ZN(n453) );
  XNOR2_X2 U384 ( .A(n541), .B(n497), .ZN(n570) );
  INV_X2 U385 ( .A(KEYINPUT68), .ZN(n490) );
  XNOR2_X2 U386 ( .A(n596), .B(n595), .ZN(n626) );
  NAND2_X2 U387 ( .A1(n386), .A2(n384), .ZN(n596) );
  XNOR2_X2 U388 ( .A(n620), .B(n392), .ZN(n470) );
  XNOR2_X2 U389 ( .A(n591), .B(n590), .ZN(n771) );
  XNOR2_X2 U390 ( .A(n458), .B(n363), .ZN(n641) );
  NAND2_X2 U391 ( .A1(n412), .A2(n411), .ZN(n522) );
  XNOR2_X1 U392 ( .A(n381), .B(n367), .ZN(n768) );
  AND2_X1 U393 ( .A1(n717), .A2(n653), .ZN(n479) );
  NAND2_X1 U394 ( .A1(n753), .A2(n652), .ZN(n717) );
  NOR2_X1 U395 ( .A1(n427), .A2(n425), .ZN(n489) );
  AND2_X1 U396 ( .A1(n615), .A2(n589), .ZN(n674) );
  NAND2_X1 U397 ( .A1(n623), .A2(n400), .ZN(n639) );
  NAND2_X2 U398 ( .A1(n375), .A2(n372), .ZN(n644) );
  AND2_X1 U399 ( .A1(n388), .A2(n387), .ZN(n386) );
  XNOR2_X1 U400 ( .A(n532), .B(n531), .ZN(n594) );
  XNOR2_X1 U401 ( .A(n477), .B(n504), .ZN(n759) );
  XOR2_X1 U402 ( .A(G113), .B(G116), .Z(n495) );
  XNOR2_X1 U403 ( .A(n649), .B(KEYINPUT95), .ZN(n357) );
  INV_X1 U404 ( .A(n697), .ZN(n358) );
  XNOR2_X1 U405 ( .A(n649), .B(KEYINPUT95), .ZN(n428) );
  XNOR2_X2 U406 ( .A(n541), .B(n488), .ZN(n726) );
  INV_X1 U407 ( .A(KEYINPUT96), .ZN(n472) );
  XNOR2_X1 U408 ( .A(n441), .B(G146), .ZN(n525) );
  INV_X1 U409 ( .A(G125), .ZN(n441) );
  XNOR2_X1 U410 ( .A(n408), .B(KEYINPUT70), .ZN(n437) );
  INV_X1 U411 ( .A(G131), .ZN(n408) );
  OR2_X1 U412 ( .A1(G237), .A2(G902), .ZN(n533) );
  AND2_X1 U413 ( .A1(n519), .A2(n520), .ZN(n609) );
  XNOR2_X1 U414 ( .A(n525), .B(n459), .ZN(n556) );
  XNOR2_X1 U415 ( .A(KEYINPUT10), .B(KEYINPUT69), .ZN(n459) );
  NAND2_X1 U416 ( .A1(n543), .A2(n374), .ZN(n385) );
  OR2_X1 U417 ( .A1(n570), .A2(n373), .ZN(n372) );
  AND2_X1 U418 ( .A1(n377), .A2(n376), .ZN(n375) );
  NAND2_X1 U419 ( .A1(G472), .A2(n374), .ZN(n373) );
  XNOR2_X1 U420 ( .A(n644), .B(KEYINPUT6), .ZN(n444) );
  INV_X1 U421 ( .A(n639), .ZN(n619) );
  OR2_X1 U422 ( .A1(n742), .A2(G902), .ZN(n458) );
  NAND2_X1 U423 ( .A1(n359), .A2(n647), .ZN(n394) );
  OR2_X1 U424 ( .A1(n661), .A2(n361), .ZN(n457) );
  XNOR2_X1 U425 ( .A(n525), .B(n526), .ZN(n468) );
  XNOR2_X1 U426 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n526) );
  NOR2_X1 U427 ( .A1(G953), .A2(G237), .ZN(n512) );
  NOR2_X1 U428 ( .A1(n772), .A2(n484), .ZN(n483) );
  INV_X1 U429 ( .A(n769), .ZN(n484) );
  XNOR2_X1 U430 ( .A(n409), .B(n437), .ZN(n477) );
  XNOR2_X1 U431 ( .A(n522), .B(n410), .ZN(n409) );
  XNOR2_X1 U432 ( .A(G137), .B(KEYINPUT72), .ZN(n410) );
  XNOR2_X1 U433 ( .A(n476), .B(G128), .ZN(n521) );
  INV_X1 U434 ( .A(G143), .ZN(n476) );
  XNOR2_X1 U435 ( .A(G140), .B(KEYINPUT71), .ZN(n555) );
  NOR2_X1 U436 ( .A1(n653), .A2(n655), .ZN(n532) );
  XNOR2_X1 U437 ( .A(n451), .B(n487), .ZN(n540) );
  XNOR2_X1 U438 ( .A(n527), .B(n528), .ZN(n451) );
  INV_X1 U439 ( .A(KEYINPUT80), .ZN(n528) );
  XNOR2_X1 U440 ( .A(G128), .B(G137), .ZN(n557) );
  XNOR2_X1 U441 ( .A(KEYINPUT100), .B(KEYINPUT23), .ZN(n559) );
  XNOR2_X1 U442 ( .A(n556), .B(n555), .ZN(n758) );
  XNOR2_X1 U443 ( .A(n516), .B(n447), .ZN(n733) );
  XNOR2_X1 U444 ( .A(n556), .B(n515), .ZN(n447) );
  XNOR2_X1 U445 ( .A(n405), .B(KEYINPUT39), .ZN(n383) );
  NAND2_X1 U446 ( .A1(n413), .A2(n402), .ZN(n405) );
  AND2_X1 U447 ( .A1(n403), .A2(n406), .ZN(n402) );
  NOR2_X1 U448 ( .A1(n686), .A2(n404), .ZN(n403) );
  AND2_X1 U449 ( .A1(n593), .A2(n445), .ZN(n602) );
  AND2_X1 U450 ( .A1(n444), .A2(n687), .ZN(n445) );
  BUF_X1 U451 ( .A(n594), .Z(n414) );
  XNOR2_X1 U452 ( .A(n461), .B(n460), .ZN(n623) );
  INV_X1 U453 ( .A(KEYINPUT22), .ZN(n460) );
  NAND2_X1 U454 ( .A1(n619), .A2(n618), .ZN(n620) );
  NAND2_X1 U455 ( .A1(n771), .A2(KEYINPUT46), .ZN(n431) );
  NAND2_X1 U456 ( .A1(n394), .A2(KEYINPUT47), .ZN(n393) );
  INV_X1 U457 ( .A(KEYINPUT73), .ZN(n599) );
  NAND2_X1 U458 ( .A1(n389), .A2(G902), .ZN(n387) );
  NAND2_X1 U459 ( .A1(n570), .A2(n378), .ZN(n377) );
  NAND2_X1 U460 ( .A1(n378), .A2(G902), .ZN(n376) );
  XOR2_X1 U461 ( .A(KEYINPUT101), .B(KEYINPUT20), .Z(n546) );
  XOR2_X1 U462 ( .A(KEYINPUT5), .B(G101), .Z(n493) );
  XNOR2_X1 U463 ( .A(G101), .B(G110), .ZN(n527) );
  NAND2_X1 U464 ( .A1(n457), .A2(KEYINPUT94), .ZN(n426) );
  NAND2_X1 U465 ( .A1(n416), .A2(KEYINPUT44), .ZN(n420) );
  AND2_X1 U466 ( .A1(n469), .A2(n474), .ZN(n473) );
  NAND2_X1 U467 ( .A1(n391), .A2(KEYINPUT96), .ZN(n474) );
  XOR2_X1 U468 ( .A(KEYINPUT104), .B(KEYINPUT12), .Z(n509) );
  XNOR2_X1 U469 ( .A(G104), .B(G122), .ZN(n508) );
  XOR2_X1 U470 ( .A(KEYINPUT11), .B(G140), .Z(n514) );
  XNOR2_X1 U471 ( .A(G143), .B(G113), .ZN(n446) );
  XOR2_X1 U472 ( .A(G902), .B(KEYINPUT15), .Z(n653) );
  XNOR2_X1 U473 ( .A(n466), .B(n749), .ZN(n655) );
  XNOR2_X1 U474 ( .A(n467), .B(n524), .ZN(n466) );
  XNOR2_X1 U475 ( .A(n523), .B(n468), .ZN(n467) );
  XNOR2_X1 U476 ( .A(n569), .B(n442), .ZN(n592) );
  INV_X1 U477 ( .A(KEYINPUT74), .ZN(n442) );
  XNOR2_X1 U478 ( .A(G119), .B(KEYINPUT3), .ZN(n494) );
  XNOR2_X1 U479 ( .A(n501), .B(n500), .ZN(n502) );
  INV_X1 U480 ( .A(KEYINPUT7), .ZN(n500) );
  XOR2_X1 U481 ( .A(G122), .B(KEYINPUT9), .Z(n501) );
  XNOR2_X1 U482 ( .A(G116), .B(G107), .ZN(n503) );
  XNOR2_X1 U483 ( .A(n521), .B(n475), .ZN(n504) );
  INV_X1 U484 ( .A(G134), .ZN(n475) );
  NOR2_X1 U485 ( .A1(n705), .A2(n399), .ZN(n706) );
  XNOR2_X1 U486 ( .A(n482), .B(n481), .ZN(n652) );
  INV_X1 U487 ( .A(KEYINPUT90), .ZN(n481) );
  NAND2_X1 U488 ( .A1(n438), .A2(KEYINPUT2), .ZN(n482) );
  XNOR2_X1 U489 ( .A(n580), .B(n407), .ZN(n413) );
  INV_X1 U490 ( .A(KEYINPUT30), .ZN(n407) );
  XNOR2_X1 U491 ( .A(n505), .B(G478), .ZN(n519) );
  INV_X1 U492 ( .A(n444), .ZN(n400) );
  NAND2_X1 U493 ( .A1(n732), .A2(G472), .ZN(n465) );
  INV_X1 U494 ( .A(n747), .ZN(n463) );
  INV_X1 U495 ( .A(KEYINPUT64), .ZN(n415) );
  XNOR2_X1 U496 ( .A(n397), .B(n540), .ZN(n749) );
  XNOR2_X1 U497 ( .A(n529), .B(n398), .ZN(n397) );
  XNOR2_X1 U498 ( .A(n485), .B(KEYINPUT79), .ZN(n398) );
  XNOR2_X1 U499 ( .A(KEYINPUT16), .B(G122), .ZN(n485) );
  XNOR2_X1 U500 ( .A(n401), .B(n564), .ZN(n742) );
  XNOR2_X1 U501 ( .A(n758), .B(n565), .ZN(n401) );
  XNOR2_X1 U502 ( .A(n419), .B(n417), .ZN(n740) );
  XNOR2_X1 U503 ( .A(n418), .B(n504), .ZN(n417) );
  NAND2_X1 U504 ( .A1(n563), .A2(G217), .ZN(n419) );
  XNOR2_X1 U505 ( .A(n502), .B(n503), .ZN(n418) );
  XNOR2_X1 U506 ( .A(n733), .B(n486), .ZN(n734) );
  BUF_X1 U507 ( .A(n732), .Z(n743) );
  NOR2_X1 U508 ( .A1(G952), .A2(n498), .ZN(n747) );
  XNOR2_X1 U509 ( .A(n380), .B(n379), .ZN(n597) );
  INV_X1 U510 ( .A(KEYINPUT36), .ZN(n379) );
  NAND2_X1 U511 ( .A1(n602), .A2(n414), .ZN(n380) );
  NOR2_X1 U512 ( .A1(n642), .A2(n399), .ZN(n643) );
  XNOR2_X1 U513 ( .A(n470), .B(G119), .ZN(n773) );
  OR2_X1 U514 ( .A1(n674), .A2(KEYINPUT87), .ZN(n359) );
  INV_X1 U515 ( .A(n520), .ZN(n584) );
  INV_X1 U516 ( .A(n668), .ZN(n391) );
  XOR2_X1 U517 ( .A(KEYINPUT25), .B(KEYINPUT102), .Z(n360) );
  INV_X1 U518 ( .A(n642), .ZN(n406) );
  AND2_X1 U519 ( .A1(n648), .A2(n647), .ZN(n361) );
  AND2_X1 U520 ( .A1(n636), .A2(n471), .ZN(n362) );
  XOR2_X1 U521 ( .A(n567), .B(n360), .Z(n363) );
  INV_X1 U522 ( .A(G902), .ZN(n374) );
  INV_X1 U523 ( .A(G472), .ZN(n378) );
  NAND2_X1 U524 ( .A1(n519), .A2(n584), .ZN(n678) );
  AND2_X1 U525 ( .A1(n668), .A2(n472), .ZN(n364) );
  AND2_X1 U526 ( .A1(n413), .A2(n406), .ZN(n365) );
  XOR2_X1 U527 ( .A(KEYINPUT98), .B(KEYINPUT0), .Z(n366) );
  INV_X1 U528 ( .A(KEYINPUT46), .ZN(n436) );
  XOR2_X1 U529 ( .A(KEYINPUT112), .B(KEYINPUT40), .Z(n367) );
  INV_X1 U530 ( .A(n681), .ZN(n382) );
  XOR2_X1 U531 ( .A(n570), .B(KEYINPUT62), .Z(n368) );
  XOR2_X1 U532 ( .A(n657), .B(n656), .Z(n369) );
  XOR2_X1 U533 ( .A(n599), .B(KEYINPUT48), .Z(n370) );
  XOR2_X1 U534 ( .A(n654), .B(KEYINPUT63), .Z(n371) );
  XNOR2_X2 U535 ( .A(n644), .B(n571), .ZN(n621) );
  AND2_X2 U536 ( .A1(n455), .A2(n479), .ZN(n732) );
  AND2_X1 U537 ( .A1(n396), .A2(n673), .ZN(n395) );
  NAND2_X1 U538 ( .A1(n383), .A2(n675), .ZN(n381) );
  XNOR2_X2 U539 ( .A(n635), .B(KEYINPUT35), .ZN(n770) );
  NAND2_X1 U540 ( .A1(n627), .A2(n444), .ZN(n628) );
  AND2_X2 U541 ( .A1(n626), .A2(n625), .ZN(n627) );
  NAND2_X1 U542 ( .A1(n424), .A2(n423), .ZN(n422) );
  AND2_X1 U543 ( .A1(n383), .A2(n382), .ZN(n600) );
  OR2_X1 U544 ( .A1(n726), .A2(n385), .ZN(n384) );
  NAND2_X1 U545 ( .A1(n726), .A2(n389), .ZN(n388) );
  INV_X1 U546 ( .A(n543), .ZN(n389) );
  NAND2_X1 U547 ( .A1(n390), .A2(n364), .ZN(n471) );
  INV_X1 U548 ( .A(n470), .ZN(n390) );
  OR2_X1 U549 ( .A1(n470), .A2(n391), .ZN(n416) );
  INV_X1 U550 ( .A(KEYINPUT32), .ZN(n392) );
  NAND2_X1 U551 ( .A1(n395), .A2(n393), .ZN(n449) );
  NAND2_X1 U552 ( .A1(n579), .A2(n578), .ZN(n396) );
  AND2_X1 U553 ( .A1(n627), .A2(n399), .ZN(n707) );
  INV_X1 U554 ( .A(n644), .ZN(n399) );
  INV_X1 U555 ( .A(n581), .ZN(n404) );
  NAND2_X1 U556 ( .A1(n490), .A2(KEYINPUT4), .ZN(n411) );
  NAND2_X1 U557 ( .A1(n491), .A2(KEYINPUT68), .ZN(n412) );
  NAND2_X1 U558 ( .A1(n498), .A2(G234), .ZN(n499) );
  INV_X1 U559 ( .A(n519), .ZN(n585) );
  NAND2_X1 U560 ( .A1(n609), .A2(n608), .ZN(n610) );
  NAND2_X1 U561 ( .A1(n420), .A2(n426), .ZN(n425) );
  NAND2_X1 U562 ( .A1(n422), .A2(n421), .ZN(n427) );
  NAND2_X1 U563 ( .A1(n357), .A2(KEYINPUT94), .ZN(n421) );
  NOR2_X1 U564 ( .A1(n457), .A2(KEYINPUT94), .ZN(n423) );
  INV_X1 U565 ( .A(n428), .ZN(n424) );
  NAND2_X1 U566 ( .A1(n768), .A2(KEYINPUT46), .ZN(n432) );
  NAND2_X1 U567 ( .A1(n448), .A2(n429), .ZN(n443) );
  NOR2_X1 U568 ( .A1(n433), .A2(n430), .ZN(n429) );
  NAND2_X1 U569 ( .A1(n432), .A2(n431), .ZN(n430) );
  NOR2_X1 U570 ( .A1(n434), .A2(n768), .ZN(n433) );
  NAND2_X1 U571 ( .A1(n435), .A2(n436), .ZN(n434) );
  INV_X1 U572 ( .A(n771), .ZN(n435) );
  XNOR2_X1 U573 ( .A(n437), .B(n446), .ZN(n511) );
  NAND2_X1 U574 ( .A1(n365), .A2(n581), .ZN(n583) );
  INV_X1 U575 ( .A(n439), .ZN(n438) );
  XNOR2_X2 U576 ( .A(n439), .B(KEYINPUT89), .ZN(n761) );
  NAND2_X1 U577 ( .A1(n601), .A2(n483), .ZN(n439) );
  NOR2_X1 U578 ( .A1(n449), .A2(n598), .ZN(n448) );
  INV_X1 U579 ( .A(KEYINPUT2), .ZN(n480) );
  NAND2_X1 U580 ( .A1(n732), .A2(G210), .ZN(n478) );
  NAND2_X1 U581 ( .A1(n617), .A2(n645), .ZN(n461) );
  XNOR2_X2 U582 ( .A(n452), .B(n366), .ZN(n645) );
  XNOR2_X2 U583 ( .A(n440), .B(KEYINPUT45), .ZN(n753) );
  NAND2_X1 U584 ( .A1(n489), .A2(n650), .ZN(n440) );
  XNOR2_X1 U585 ( .A(n465), .B(n368), .ZN(n464) );
  NAND2_X1 U586 ( .A1(n621), .A2(n592), .ZN(n573) );
  XNOR2_X1 U587 ( .A(n443), .B(n370), .ZN(n601) );
  XNOR2_X1 U588 ( .A(n478), .B(n369), .ZN(n658) );
  NAND2_X1 U589 ( .A1(n464), .A2(n463), .ZN(n462) );
  INV_X1 U590 ( .A(n641), .ZN(n699) );
  NAND2_X1 U591 ( .A1(n641), .A2(n568), .ZN(n569) );
  NAND2_X1 U592 ( .A1(n621), .A2(n687), .ZN(n580) );
  NOR2_X1 U593 ( .A1(n736), .A2(n747), .ZN(n738) );
  NAND2_X1 U594 ( .A1(n450), .A2(n697), .ZN(n640) );
  XNOR2_X1 U595 ( .A(n639), .B(KEYINPUT93), .ZN(n450) );
  NAND2_X1 U596 ( .A1(n615), .A2(n616), .ZN(n452) );
  XNOR2_X1 U597 ( .A(n453), .B(n660), .ZN(G51) );
  NAND2_X1 U598 ( .A1(n454), .A2(n753), .ZN(n456) );
  INV_X1 U599 ( .A(n651), .ZN(n454) );
  NAND2_X1 U600 ( .A1(n456), .A2(n480), .ZN(n455) );
  XNOR2_X1 U601 ( .A(n462), .B(n371), .ZN(G57) );
  NAND2_X1 U602 ( .A1(n470), .A2(KEYINPUT96), .ZN(n469) );
  NAND2_X1 U603 ( .A1(n473), .A2(n362), .ZN(n638) );
  XNOR2_X1 U604 ( .A(n638), .B(n637), .ZN(n650) );
  XNOR2_X1 U605 ( .A(n735), .B(n734), .ZN(n736) );
  XNOR2_X1 U606 ( .A(KEYINPUT125), .B(KEYINPUT59), .ZN(n486) );
  XOR2_X1 U607 ( .A(G107), .B(G104), .Z(n487) );
  XOR2_X1 U608 ( .A(n540), .B(n539), .Z(n488) );
  INV_X1 U609 ( .A(KEYINPUT77), .ZN(n637) );
  INV_X1 U610 ( .A(KEYINPUT76), .ZN(n542) );
  XNOR2_X1 U611 ( .A(n496), .B(n529), .ZN(n497) );
  XNOR2_X1 U612 ( .A(n542), .B(G469), .ZN(n543) );
  INV_X1 U613 ( .A(KEYINPUT108), .ZN(n571) );
  AND2_X1 U614 ( .A1(n358), .A2(n641), .ZN(n618) );
  XNOR2_X1 U615 ( .A(n530), .B(KEYINPUT86), .ZN(n531) );
  INV_X1 U616 ( .A(KEYINPUT4), .ZN(n491) );
  XNOR2_X2 U617 ( .A(n759), .B(G146), .ZN(n541) );
  NAND2_X1 U618 ( .A1(n512), .A2(G210), .ZN(n492) );
  XNOR2_X1 U619 ( .A(n493), .B(n492), .ZN(n496) );
  INV_X1 U620 ( .A(KEYINPUT87), .ZN(n576) );
  XOR2_X1 U621 ( .A(KEYINPUT8), .B(n499), .Z(n563) );
  NOR2_X1 U622 ( .A1(G902), .A2(n740), .ZN(n505) );
  XOR2_X1 U623 ( .A(KEYINPUT106), .B(KEYINPUT13), .Z(n507) );
  XNOR2_X1 U624 ( .A(KEYINPUT105), .B(G475), .ZN(n506) );
  XNOR2_X1 U625 ( .A(n507), .B(n506), .ZN(n518) );
  XNOR2_X1 U626 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U627 ( .A(n511), .B(n510), .ZN(n516) );
  NAND2_X1 U628 ( .A1(G214), .A2(n512), .ZN(n513) );
  XNOR2_X1 U629 ( .A(n514), .B(n513), .ZN(n515) );
  NOR2_X1 U630 ( .A1(G902), .A2(n733), .ZN(n517) );
  XOR2_X1 U631 ( .A(n518), .B(n517), .Z(n520) );
  NAND2_X1 U632 ( .A1(n585), .A2(n520), .ZN(n681) );
  NAND2_X1 U633 ( .A1(n678), .A2(n681), .ZN(n647) );
  XOR2_X1 U634 ( .A(n522), .B(n521), .Z(n524) );
  NAND2_X1 U635 ( .A1(G224), .A2(n498), .ZN(n523) );
  NAND2_X1 U636 ( .A1(G210), .A2(n533), .ZN(n530) );
  NAND2_X1 U637 ( .A1(G214), .A2(n533), .ZN(n687) );
  NAND2_X1 U638 ( .A1(n594), .A2(n687), .ZN(n536) );
  XNOR2_X1 U639 ( .A(KEYINPUT19), .B(KEYINPUT66), .ZN(n534) );
  XNOR2_X1 U640 ( .A(n534), .B(KEYINPUT82), .ZN(n535) );
  XNOR2_X1 U641 ( .A(n536), .B(n535), .ZN(n615) );
  XNOR2_X1 U642 ( .A(n555), .B(KEYINPUT83), .ZN(n538) );
  NAND2_X1 U643 ( .A1(G227), .A2(n498), .ZN(n537) );
  XNOR2_X1 U644 ( .A(n538), .B(n537), .ZN(n539) );
  INV_X1 U645 ( .A(n653), .ZN(n544) );
  NAND2_X1 U646 ( .A1(G234), .A2(n544), .ZN(n545) );
  XNOR2_X1 U647 ( .A(n546), .B(n545), .ZN(n566) );
  NAND2_X1 U648 ( .A1(n566), .A2(G221), .ZN(n547) );
  XOR2_X1 U649 ( .A(n547), .B(KEYINPUT21), .Z(n700) );
  NAND2_X1 U650 ( .A1(G234), .A2(G237), .ZN(n548) );
  XNOR2_X1 U651 ( .A(KEYINPUT14), .B(n548), .ZN(n550) );
  NAND2_X1 U652 ( .A1(G952), .A2(n550), .ZN(n715) );
  NOR2_X1 U653 ( .A1(n715), .A2(G953), .ZN(n549) );
  XNOR2_X1 U654 ( .A(n549), .B(KEYINPUT99), .ZN(n613) );
  NAND2_X1 U655 ( .A1(G902), .A2(n550), .ZN(n611) );
  NOR2_X1 U656 ( .A1(G900), .A2(n611), .ZN(n552) );
  INV_X1 U657 ( .A(n498), .ZN(n551) );
  NAND2_X1 U658 ( .A1(n552), .A2(n551), .ZN(n553) );
  NAND2_X1 U659 ( .A1(n613), .A2(n553), .ZN(n581) );
  NAND2_X1 U660 ( .A1(n700), .A2(n581), .ZN(n554) );
  XNOR2_X1 U661 ( .A(n554), .B(KEYINPUT75), .ZN(n568) );
  XOR2_X1 U662 ( .A(G110), .B(G119), .Z(n558) );
  XNOR2_X1 U663 ( .A(n558), .B(n557), .ZN(n562) );
  XOR2_X1 U664 ( .A(KEYINPUT88), .B(KEYINPUT24), .Z(n560) );
  XNOR2_X1 U665 ( .A(n560), .B(n559), .ZN(n561) );
  XOR2_X1 U666 ( .A(n562), .B(n561), .Z(n565) );
  NAND2_X1 U667 ( .A1(G221), .A2(n563), .ZN(n564) );
  NAND2_X1 U668 ( .A1(G217), .A2(n566), .ZN(n567) );
  XNOR2_X1 U669 ( .A(KEYINPUT111), .B(KEYINPUT28), .ZN(n572) );
  XNOR2_X1 U670 ( .A(n573), .B(n572), .ZN(n574) );
  AND2_X1 U671 ( .A1(n596), .A2(n574), .ZN(n589) );
  NAND2_X1 U672 ( .A1(n647), .A2(n674), .ZN(n575) );
  NAND2_X1 U673 ( .A1(n576), .A2(n575), .ZN(n579) );
  NAND2_X1 U674 ( .A1(KEYINPUT87), .A2(n674), .ZN(n577) );
  NAND2_X1 U675 ( .A1(n577), .A2(KEYINPUT47), .ZN(n578) );
  NAND2_X1 U676 ( .A1(n584), .A2(n585), .ZN(n632) );
  XOR2_X1 U677 ( .A(KEYINPUT103), .B(n700), .Z(n608) );
  NAND2_X1 U678 ( .A1(n699), .A2(n608), .ZN(n696) );
  INV_X1 U679 ( .A(n696), .ZN(n625) );
  NAND2_X1 U680 ( .A1(n625), .A2(n596), .ZN(n642) );
  NOR2_X1 U681 ( .A1(n632), .A2(n583), .ZN(n582) );
  NAND2_X1 U682 ( .A1(n582), .A2(n414), .ZN(n673) );
  INV_X1 U683 ( .A(n647), .ZN(n691) );
  INV_X1 U684 ( .A(n594), .ZN(n605) );
  XOR2_X1 U685 ( .A(n605), .B(KEYINPUT38), .Z(n686) );
  INV_X1 U686 ( .A(n609), .ZN(n689) );
  XNOR2_X1 U687 ( .A(n605), .B(KEYINPUT38), .ZN(n586) );
  NAND2_X1 U688 ( .A1(n586), .A2(n687), .ZN(n690) );
  NOR2_X1 U689 ( .A1(n689), .A2(n690), .ZN(n588) );
  XNOR2_X1 U690 ( .A(KEYINPUT113), .B(KEYINPUT41), .ZN(n587) );
  XNOR2_X1 U691 ( .A(n588), .B(n587), .ZN(n709) );
  NAND2_X1 U692 ( .A1(n709), .A2(n589), .ZN(n591) );
  XOR2_X1 U693 ( .A(KEYINPUT114), .B(KEYINPUT42), .Z(n590) );
  INV_X1 U694 ( .A(n678), .ZN(n675) );
  AND2_X1 U695 ( .A1(n592), .A2(n675), .ZN(n593) );
  XOR2_X1 U696 ( .A(KEYINPUT1), .B(KEYINPUT65), .Z(n595) );
  INV_X1 U697 ( .A(n626), .ZN(n697) );
  NAND2_X1 U698 ( .A1(n597), .A2(n358), .ZN(n685) );
  XOR2_X1 U699 ( .A(n685), .B(KEYINPUT92), .Z(n598) );
  XNOR2_X1 U700 ( .A(n600), .B(KEYINPUT115), .ZN(n769) );
  XOR2_X1 U701 ( .A(KEYINPUT43), .B(KEYINPUT109), .Z(n604) );
  NAND2_X1 U702 ( .A1(n602), .A2(n697), .ZN(n603) );
  XNOR2_X1 U703 ( .A(n604), .B(n603), .ZN(n606) );
  NAND2_X1 U704 ( .A1(n606), .A2(n605), .ZN(n607) );
  XOR2_X1 U705 ( .A(KEYINPUT110), .B(n607), .Z(n772) );
  XNOR2_X1 U706 ( .A(n761), .B(KEYINPUT81), .ZN(n651) );
  XNOR2_X1 U707 ( .A(KEYINPUT107), .B(n610), .ZN(n617) );
  INV_X1 U708 ( .A(n611), .ZN(n612) );
  INV_X1 U709 ( .A(G953), .ZN(n752) );
  NOR2_X1 U710 ( .A1(G898), .A2(n752), .ZN(n748) );
  NAND2_X1 U711 ( .A1(n612), .A2(n748), .ZN(n614) );
  NAND2_X1 U712 ( .A1(n614), .A2(n613), .ZN(n616) );
  OR2_X1 U713 ( .A1(n621), .A2(n626), .ZN(n622) );
  NOR2_X1 U714 ( .A1(n699), .A2(n622), .ZN(n624) );
  NAND2_X1 U715 ( .A1(n624), .A2(n623), .ZN(n668) );
  XNOR2_X2 U716 ( .A(n628), .B(KEYINPUT33), .ZN(n719) );
  NAND2_X1 U717 ( .A1(n719), .A2(n645), .ZN(n631) );
  XNOR2_X1 U718 ( .A(KEYINPUT78), .B(KEYINPUT34), .ZN(n629) );
  XNOR2_X1 U719 ( .A(n629), .B(KEYINPUT85), .ZN(n630) );
  XNOR2_X1 U720 ( .A(n631), .B(n630), .ZN(n634) );
  XOR2_X1 U721 ( .A(KEYINPUT84), .B(n632), .Z(n633) );
  NAND2_X1 U722 ( .A1(n634), .A2(n633), .ZN(n635) );
  NOR2_X1 U723 ( .A1(KEYINPUT44), .A2(n770), .ZN(n636) );
  NOR2_X1 U724 ( .A1(n641), .A2(n640), .ZN(n661) );
  NAND2_X1 U725 ( .A1(n645), .A2(n643), .ZN(n663) );
  NAND2_X1 U726 ( .A1(n645), .A2(n707), .ZN(n646) );
  XOR2_X1 U727 ( .A(KEYINPUT31), .B(n646), .Z(n680) );
  NAND2_X1 U728 ( .A1(n663), .A2(n680), .ZN(n648) );
  INV_X1 U729 ( .A(KEYINPUT116), .ZN(n654) );
  XOR2_X1 U730 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n657) );
  XNOR2_X1 U731 ( .A(n655), .B(KEYINPUT97), .ZN(n656) );
  INV_X1 U732 ( .A(KEYINPUT56), .ZN(n659) );
  XNOR2_X1 U733 ( .A(n659), .B(KEYINPUT91), .ZN(n660) );
  XOR2_X1 U734 ( .A(n661), .B(G101), .Z(G3) );
  NOR2_X1 U735 ( .A1(n678), .A2(n663), .ZN(n662) );
  XOR2_X1 U736 ( .A(G104), .B(n662), .Z(G6) );
  NOR2_X1 U737 ( .A1(n663), .A2(n681), .ZN(n667) );
  XOR2_X1 U738 ( .A(KEYINPUT117), .B(KEYINPUT26), .Z(n665) );
  XNOR2_X1 U739 ( .A(G107), .B(KEYINPUT27), .ZN(n664) );
  XNOR2_X1 U740 ( .A(n665), .B(n664), .ZN(n666) );
  XNOR2_X1 U741 ( .A(n667), .B(n666), .ZN(G9) );
  XNOR2_X1 U742 ( .A(G110), .B(KEYINPUT118), .ZN(n669) );
  XNOR2_X1 U743 ( .A(n669), .B(n668), .ZN(G12) );
  XOR2_X1 U744 ( .A(KEYINPUT119), .B(KEYINPUT29), .Z(n671) );
  NAND2_X1 U745 ( .A1(n674), .A2(n382), .ZN(n670) );
  XNOR2_X1 U746 ( .A(n671), .B(n670), .ZN(n672) );
  XOR2_X1 U747 ( .A(G128), .B(n672), .Z(G30) );
  XNOR2_X1 U748 ( .A(G143), .B(n673), .ZN(G45) );
  XNOR2_X1 U749 ( .A(G146), .B(KEYINPUT120), .ZN(n677) );
  NAND2_X1 U750 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U751 ( .A(n677), .B(n676), .ZN(G48) );
  NOR2_X1 U752 ( .A1(n678), .A2(n680), .ZN(n679) );
  XOR2_X1 U753 ( .A(G113), .B(n679), .Z(G15) );
  NOR2_X1 U754 ( .A1(n681), .A2(n680), .ZN(n683) );
  XNOR2_X1 U755 ( .A(G116), .B(KEYINPUT121), .ZN(n682) );
  XNOR2_X1 U756 ( .A(n683), .B(n682), .ZN(G18) );
  XOR2_X1 U757 ( .A(G125), .B(KEYINPUT37), .Z(n684) );
  XNOR2_X1 U758 ( .A(n685), .B(n684), .ZN(G27) );
  NOR2_X1 U759 ( .A1(n687), .A2(n586), .ZN(n688) );
  NOR2_X1 U760 ( .A1(n689), .A2(n688), .ZN(n693) );
  NOR2_X1 U761 ( .A1(n691), .A2(n690), .ZN(n692) );
  NOR2_X1 U762 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U763 ( .A(n694), .B(KEYINPUT123), .ZN(n695) );
  NAND2_X1 U764 ( .A1(n695), .A2(n719), .ZN(n712) );
  NAND2_X1 U765 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U766 ( .A(KEYINPUT50), .B(n698), .ZN(n704) );
  XOR2_X1 U767 ( .A(KEYINPUT49), .B(KEYINPUT122), .Z(n702) );
  OR2_X1 U768 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U769 ( .A(n702), .B(n701), .ZN(n703) );
  NAND2_X1 U770 ( .A1(n704), .A2(n703), .ZN(n705) );
  NOR2_X1 U771 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U772 ( .A(KEYINPUT51), .B(n708), .ZN(n710) );
  NAND2_X1 U773 ( .A1(n710), .A2(n709), .ZN(n711) );
  NAND2_X1 U774 ( .A1(n712), .A2(n711), .ZN(n713) );
  XOR2_X1 U775 ( .A(KEYINPUT52), .B(n713), .Z(n714) );
  NOR2_X1 U776 ( .A1(n715), .A2(n714), .ZN(n723) );
  NAND2_X1 U777 ( .A1(n753), .A2(n761), .ZN(n716) );
  NAND2_X1 U778 ( .A1(n716), .A2(n480), .ZN(n718) );
  NAND2_X1 U779 ( .A1(n718), .A2(n717), .ZN(n721) );
  NAND2_X1 U780 ( .A1(n719), .A2(n709), .ZN(n720) );
  NAND2_X1 U781 ( .A1(n721), .A2(n720), .ZN(n722) );
  NOR2_X1 U782 ( .A1(n723), .A2(n722), .ZN(n724) );
  NAND2_X1 U783 ( .A1(n752), .A2(n724), .ZN(n725) );
  XOR2_X1 U784 ( .A(KEYINPUT53), .B(n725), .Z(G75) );
  XOR2_X1 U785 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n728) );
  XNOR2_X1 U786 ( .A(n726), .B(KEYINPUT124), .ZN(n727) );
  XNOR2_X1 U787 ( .A(n728), .B(n727), .ZN(n730) );
  NAND2_X1 U788 ( .A1(n743), .A2(G469), .ZN(n729) );
  XNOR2_X1 U789 ( .A(n730), .B(n729), .ZN(n731) );
  NOR2_X1 U790 ( .A1(n747), .A2(n731), .ZN(G54) );
  NAND2_X1 U791 ( .A1(n732), .A2(G475), .ZN(n735) );
  XOR2_X1 U792 ( .A(KEYINPUT60), .B(KEYINPUT67), .Z(n737) );
  XNOR2_X1 U793 ( .A(n738), .B(n737), .ZN(G60) );
  NAND2_X1 U794 ( .A1(G478), .A2(n743), .ZN(n739) );
  XNOR2_X1 U795 ( .A(n740), .B(n739), .ZN(n741) );
  NOR2_X1 U796 ( .A1(n747), .A2(n741), .ZN(G63) );
  XNOR2_X1 U797 ( .A(n742), .B(KEYINPUT126), .ZN(n745) );
  NAND2_X1 U798 ( .A1(G217), .A2(n743), .ZN(n744) );
  XNOR2_X1 U799 ( .A(n745), .B(n744), .ZN(n746) );
  NOR2_X1 U800 ( .A1(n747), .A2(n746), .ZN(G66) );
  NOR2_X1 U801 ( .A1(n749), .A2(n748), .ZN(n757) );
  NAND2_X1 U802 ( .A1(G953), .A2(G224), .ZN(n750) );
  XNOR2_X1 U803 ( .A(KEYINPUT61), .B(n750), .ZN(n751) );
  NAND2_X1 U804 ( .A1(n751), .A2(G898), .ZN(n755) );
  NAND2_X1 U805 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U806 ( .A1(n755), .A2(n754), .ZN(n756) );
  XNOR2_X1 U807 ( .A(n757), .B(n756), .ZN(G69) );
  XNOR2_X1 U808 ( .A(n759), .B(n758), .ZN(n763) );
  INV_X1 U809 ( .A(n763), .ZN(n760) );
  XNOR2_X1 U810 ( .A(n761), .B(n760), .ZN(n762) );
  NAND2_X1 U811 ( .A1(n498), .A2(n762), .ZN(n767) );
  XNOR2_X1 U812 ( .A(G227), .B(n763), .ZN(n764) );
  NAND2_X1 U813 ( .A1(n764), .A2(G900), .ZN(n765) );
  NAND2_X1 U814 ( .A1(G953), .A2(n765), .ZN(n766) );
  NAND2_X1 U815 ( .A1(n767), .A2(n766), .ZN(G72) );
  XOR2_X1 U816 ( .A(n768), .B(G131), .Z(G33) );
  XNOR2_X1 U817 ( .A(G134), .B(n769), .ZN(G36) );
  XOR2_X1 U818 ( .A(n770), .B(G122), .Z(G24) );
  XOR2_X1 U819 ( .A(G137), .B(n771), .Z(G39) );
  XOR2_X1 U820 ( .A(G140), .B(n772), .Z(G42) );
  XNOR2_X1 U821 ( .A(KEYINPUT127), .B(n773), .ZN(G21) );
endmodule

