

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590;

  NOR2_X1 U325 ( .A1(n376), .A2(n582), .ZN(n377) );
  XNOR2_X1 U326 ( .A(n303), .B(n325), .ZN(n304) );
  XNOR2_X1 U327 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U328 ( .A(n297), .B(n296), .ZN(n299) );
  XNOR2_X1 U329 ( .A(n299), .B(n298), .ZN(n392) );
  XNOR2_X1 U330 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U331 ( .A(n450), .B(n449), .ZN(G1349GAT) );
  XOR2_X1 U332 ( .A(KEYINPUT31), .B(KEYINPUT32), .Z(n294) );
  NAND2_X1 U333 ( .A1(G230GAT), .A2(G233GAT), .ZN(n293) );
  XNOR2_X1 U334 ( .A(n294), .B(n293), .ZN(n295) );
  XNOR2_X1 U335 ( .A(KEYINPUT71), .B(n295), .ZN(n307) );
  XOR2_X1 U336 ( .A(KEYINPUT33), .B(KEYINPUT69), .Z(n301) );
  XNOR2_X1 U337 ( .A(G99GAT), .B(G85GAT), .ZN(n297) );
  INV_X1 U338 ( .A(G106GAT), .ZN(n296) );
  XOR2_X1 U339 ( .A(KEYINPUT70), .B(G92GAT), .Z(n298) );
  XOR2_X1 U340 ( .A(G57GAT), .B(KEYINPUT13), .Z(n364) );
  XNOR2_X1 U341 ( .A(n392), .B(n364), .ZN(n300) );
  XOR2_X1 U342 ( .A(n301), .B(n300), .Z(n305) );
  XOR2_X1 U343 ( .A(G120GAT), .B(G71GAT), .Z(n310) );
  XNOR2_X1 U344 ( .A(G78GAT), .B(G204GAT), .ZN(n302) );
  XNOR2_X1 U345 ( .A(n302), .B(G148GAT), .ZN(n419) );
  XNOR2_X1 U346 ( .A(n310), .B(n419), .ZN(n303) );
  XOR2_X1 U347 ( .A(G176GAT), .B(G64GAT), .Z(n325) );
  XNOR2_X1 U348 ( .A(n307), .B(n306), .ZN(n396) );
  XNOR2_X1 U349 ( .A(KEYINPUT41), .B(n396), .ZN(n549) );
  XNOR2_X1 U350 ( .A(KEYINPUT103), .B(n549), .ZN(n533) );
  XOR2_X1 U351 ( .A(G99GAT), .B(G134GAT), .Z(n309) );
  XNOR2_X1 U352 ( .A(G43GAT), .B(G190GAT), .ZN(n308) );
  XNOR2_X1 U353 ( .A(n309), .B(n308), .ZN(n324) );
  XOR2_X1 U354 ( .A(G15GAT), .B(G127GAT), .Z(n371) );
  XOR2_X1 U355 ( .A(n371), .B(n310), .Z(n312) );
  NAND2_X1 U356 ( .A1(G227GAT), .A2(G233GAT), .ZN(n311) );
  XNOR2_X1 U357 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U358 ( .A(G113GAT), .B(KEYINPUT0), .Z(n431) );
  XOR2_X1 U359 ( .A(n313), .B(n431), .Z(n322) );
  XOR2_X1 U360 ( .A(KEYINPUT81), .B(KEYINPUT82), .Z(n315) );
  XNOR2_X1 U361 ( .A(G169GAT), .B(G176GAT), .ZN(n314) );
  XNOR2_X1 U362 ( .A(n315), .B(n314), .ZN(n320) );
  XOR2_X1 U363 ( .A(G183GAT), .B(KEYINPUT17), .Z(n317) );
  XNOR2_X1 U364 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n316) );
  XNOR2_X1 U365 ( .A(n317), .B(n316), .ZN(n334) );
  XNOR2_X1 U366 ( .A(n334), .B(KEYINPUT83), .ZN(n318) );
  XNOR2_X1 U367 ( .A(n318), .B(KEYINPUT20), .ZN(n319) );
  XNOR2_X1 U368 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U369 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U370 ( .A(n324), .B(n323), .Z(n520) );
  INV_X1 U371 ( .A(n520), .ZN(n527) );
  XOR2_X1 U372 ( .A(G169GAT), .B(G8GAT), .Z(n343) );
  XNOR2_X1 U373 ( .A(n343), .B(n325), .ZN(n338) );
  XNOR2_X1 U374 ( .A(G36GAT), .B(G190GAT), .ZN(n326) );
  XNOR2_X1 U375 ( .A(n326), .B(G218GAT), .ZN(n381) );
  XOR2_X1 U376 ( .A(n381), .B(KEYINPUT88), .Z(n328) );
  NAND2_X1 U377 ( .A1(G226GAT), .A2(G233GAT), .ZN(n327) );
  XNOR2_X1 U378 ( .A(n328), .B(n327), .ZN(n332) );
  XOR2_X1 U379 ( .A(KEYINPUT89), .B(KEYINPUT76), .Z(n330) );
  XNOR2_X1 U380 ( .A(G204GAT), .B(G92GAT), .ZN(n329) );
  XNOR2_X1 U381 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U382 ( .A(n332), .B(n331), .Z(n336) );
  XNOR2_X1 U383 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n333) );
  XNOR2_X1 U384 ( .A(n333), .B(G211GAT), .ZN(n407) );
  XNOR2_X1 U385 ( .A(n334), .B(n407), .ZN(n335) );
  XNOR2_X1 U386 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U387 ( .A(n338), .B(n337), .Z(n517) );
  INV_X1 U388 ( .A(n517), .ZN(n489) );
  XOR2_X1 U389 ( .A(G22GAT), .B(G141GAT), .Z(n340) );
  XNOR2_X1 U390 ( .A(G113GAT), .B(G15GAT), .ZN(n339) );
  XNOR2_X1 U391 ( .A(n340), .B(n339), .ZN(n356) );
  XOR2_X1 U392 ( .A(G29GAT), .B(G43GAT), .Z(n342) );
  XNOR2_X1 U393 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n341) );
  XNOR2_X1 U394 ( .A(n342), .B(n341), .ZN(n382) );
  XOR2_X1 U395 ( .A(n343), .B(n382), .Z(n345) );
  XNOR2_X1 U396 ( .A(G36GAT), .B(G50GAT), .ZN(n344) );
  XNOR2_X1 U397 ( .A(n345), .B(n344), .ZN(n349) );
  XOR2_X1 U398 ( .A(KEYINPUT67), .B(KEYINPUT30), .Z(n347) );
  NAND2_X1 U399 ( .A1(G229GAT), .A2(G233GAT), .ZN(n346) );
  XNOR2_X1 U400 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U401 ( .A(n349), .B(n348), .Z(n354) );
  XOR2_X1 U402 ( .A(KEYINPUT29), .B(KEYINPUT68), .Z(n351) );
  XNOR2_X1 U403 ( .A(G197GAT), .B(G1GAT), .ZN(n350) );
  XNOR2_X1 U404 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U405 ( .A(n352), .B(KEYINPUT66), .ZN(n353) );
  XNOR2_X1 U406 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U407 ( .A(n356), .B(n355), .ZN(n531) );
  NOR2_X1 U408 ( .A1(n531), .A2(n549), .ZN(n357) );
  XNOR2_X1 U409 ( .A(n357), .B(KEYINPUT46), .ZN(n376) );
  XOR2_X1 U410 ( .A(KEYINPUT76), .B(G64GAT), .Z(n359) );
  XNOR2_X1 U411 ( .A(G78GAT), .B(G211GAT), .ZN(n358) );
  XNOR2_X1 U412 ( .A(n359), .B(n358), .ZN(n363) );
  XOR2_X1 U413 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n361) );
  XNOR2_X1 U414 ( .A(G1GAT), .B(G8GAT), .ZN(n360) );
  XNOR2_X1 U415 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U416 ( .A(n363), .B(n362), .ZN(n375) );
  XOR2_X1 U417 ( .A(G22GAT), .B(G155GAT), .Z(n410) );
  XOR2_X1 U418 ( .A(n364), .B(n410), .Z(n366) );
  XNOR2_X1 U419 ( .A(G183GAT), .B(G71GAT), .ZN(n365) );
  XNOR2_X1 U420 ( .A(n366), .B(n365), .ZN(n370) );
  XOR2_X1 U421 ( .A(KEYINPUT12), .B(KEYINPUT77), .Z(n368) );
  NAND2_X1 U422 ( .A1(G231GAT), .A2(G233GAT), .ZN(n367) );
  XNOR2_X1 U423 ( .A(n368), .B(n367), .ZN(n369) );
  XOR2_X1 U424 ( .A(n370), .B(n369), .Z(n373) );
  XNOR2_X1 U425 ( .A(n371), .B(KEYINPUT78), .ZN(n372) );
  XNOR2_X1 U426 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U427 ( .A(n375), .B(n374), .Z(n480) );
  INV_X1 U428 ( .A(n480), .ZN(n582) );
  XNOR2_X1 U429 ( .A(n377), .B(KEYINPUT112), .ZN(n393) );
  XOR2_X1 U430 ( .A(KEYINPUT65), .B(KEYINPUT72), .Z(n379) );
  NAND2_X1 U431 ( .A1(G232GAT), .A2(G233GAT), .ZN(n378) );
  XNOR2_X1 U432 ( .A(n379), .B(n378), .ZN(n380) );
  XOR2_X1 U433 ( .A(n380), .B(KEYINPUT9), .Z(n384) );
  XNOR2_X1 U434 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U435 ( .A(n384), .B(n383), .ZN(n388) );
  XOR2_X1 U436 ( .A(KEYINPUT11), .B(KEYINPUT10), .Z(n386) );
  XNOR2_X1 U437 ( .A(KEYINPUT64), .B(KEYINPUT74), .ZN(n385) );
  XNOR2_X1 U438 ( .A(n386), .B(n385), .ZN(n387) );
  XOR2_X1 U439 ( .A(n388), .B(n387), .Z(n390) );
  XOR2_X1 U440 ( .A(G50GAT), .B(G162GAT), .Z(n406) );
  XOR2_X1 U441 ( .A(G134GAT), .B(KEYINPUT73), .Z(n430) );
  XNOR2_X1 U442 ( .A(n406), .B(n430), .ZN(n389) );
  XNOR2_X1 U443 ( .A(n390), .B(n389), .ZN(n391) );
  XNOR2_X1 U444 ( .A(n392), .B(n391), .ZN(n560) );
  NAND2_X1 U445 ( .A1(n393), .A2(n560), .ZN(n394) );
  XNOR2_X1 U446 ( .A(n394), .B(KEYINPUT47), .ZN(n395) );
  XNOR2_X1 U447 ( .A(n395), .B(KEYINPUT113), .ZN(n402) );
  XNOR2_X1 U448 ( .A(KEYINPUT75), .B(n560), .ZN(n565) );
  XNOR2_X1 U449 ( .A(n565), .B(KEYINPUT97), .ZN(n397) );
  XNOR2_X1 U450 ( .A(n397), .B(KEYINPUT36), .ZN(n587) );
  NOR2_X1 U451 ( .A1(n587), .A2(n480), .ZN(n398) );
  XOR2_X1 U452 ( .A(KEYINPUT45), .B(n398), .Z(n399) );
  NOR2_X1 U453 ( .A1(n396), .A2(n399), .ZN(n400) );
  NAND2_X1 U454 ( .A1(n400), .A2(n531), .ZN(n401) );
  NAND2_X1 U455 ( .A1(n402), .A2(n401), .ZN(n404) );
  INV_X1 U456 ( .A(KEYINPUT48), .ZN(n403) );
  XNOR2_X1 U457 ( .A(n404), .B(n403), .ZN(n543) );
  NOR2_X1 U458 ( .A1(n489), .A2(n543), .ZN(n405) );
  XNOR2_X1 U459 ( .A(KEYINPUT54), .B(n405), .ZN(n571) );
  XOR2_X1 U460 ( .A(n407), .B(n406), .Z(n409) );
  NAND2_X1 U461 ( .A1(G228GAT), .A2(G233GAT), .ZN(n408) );
  XNOR2_X1 U462 ( .A(n409), .B(n408), .ZN(n411) );
  XOR2_X1 U463 ( .A(n411), .B(n410), .Z(n413) );
  XNOR2_X1 U464 ( .A(G218GAT), .B(G106GAT), .ZN(n412) );
  XNOR2_X1 U465 ( .A(n413), .B(n412), .ZN(n417) );
  XOR2_X1 U466 ( .A(KEYINPUT24), .B(KEYINPUT22), .Z(n415) );
  XNOR2_X1 U467 ( .A(KEYINPUT84), .B(KEYINPUT23), .ZN(n414) );
  XNOR2_X1 U468 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U469 ( .A(n417), .B(n416), .Z(n421) );
  XNOR2_X1 U470 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n418) );
  XNOR2_X1 U471 ( .A(n418), .B(KEYINPUT2), .ZN(n439) );
  XNOR2_X1 U472 ( .A(n439), .B(n419), .ZN(n420) );
  XNOR2_X1 U473 ( .A(n421), .B(n420), .ZN(n457) );
  XOR2_X1 U474 ( .A(KEYINPUT85), .B(G57GAT), .Z(n423) );
  XNOR2_X1 U475 ( .A(G1GAT), .B(G155GAT), .ZN(n422) );
  XNOR2_X1 U476 ( .A(n423), .B(n422), .ZN(n427) );
  XOR2_X1 U477 ( .A(G85GAT), .B(G148GAT), .Z(n425) );
  XNOR2_X1 U478 ( .A(G120GAT), .B(G127GAT), .ZN(n424) );
  XNOR2_X1 U479 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U480 ( .A(n427), .B(n426), .ZN(n443) );
  XOR2_X1 U481 ( .A(KEYINPUT5), .B(KEYINPUT87), .Z(n429) );
  XNOR2_X1 U482 ( .A(KEYINPUT4), .B(KEYINPUT86), .ZN(n428) );
  XNOR2_X1 U483 ( .A(n429), .B(n428), .ZN(n435) );
  XOR2_X1 U484 ( .A(n430), .B(G162GAT), .Z(n433) );
  XNOR2_X1 U485 ( .A(G29GAT), .B(n431), .ZN(n432) );
  XNOR2_X1 U486 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U487 ( .A(n435), .B(n434), .Z(n437) );
  NAND2_X1 U488 ( .A1(G225GAT), .A2(G233GAT), .ZN(n436) );
  XNOR2_X1 U489 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U490 ( .A(n438), .B(KEYINPUT6), .Z(n441) );
  XNOR2_X1 U491 ( .A(n439), .B(KEYINPUT1), .ZN(n440) );
  XNOR2_X1 U492 ( .A(n441), .B(n440), .ZN(n442) );
  XOR2_X1 U493 ( .A(n443), .B(n442), .Z(n515) );
  NOR2_X1 U494 ( .A1(n457), .A2(n515), .ZN(n444) );
  AND2_X1 U495 ( .A1(n571), .A2(n444), .ZN(n445) );
  XNOR2_X1 U496 ( .A(n445), .B(KEYINPUT55), .ZN(n446) );
  NOR2_X2 U497 ( .A1(n527), .A2(n446), .ZN(n566) );
  NAND2_X1 U498 ( .A1(n533), .A2(n566), .ZN(n450) );
  XOR2_X1 U499 ( .A(G176GAT), .B(KEYINPUT122), .Z(n448) );
  XNOR2_X1 U500 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n447) );
  INV_X1 U501 ( .A(n515), .ZN(n570) );
  XNOR2_X1 U502 ( .A(n457), .B(KEYINPUT28), .ZN(n522) );
  XOR2_X1 U503 ( .A(n517), .B(KEYINPUT27), .Z(n454) );
  OR2_X1 U504 ( .A1(n522), .A2(n454), .ZN(n451) );
  NOR2_X1 U505 ( .A1(n570), .A2(n451), .ZN(n529) );
  NAND2_X1 U506 ( .A1(n529), .A2(n527), .ZN(n452) );
  XOR2_X1 U507 ( .A(KEYINPUT90), .B(n452), .Z(n462) );
  NAND2_X1 U508 ( .A1(n527), .A2(n457), .ZN(n453) );
  XNOR2_X1 U509 ( .A(n453), .B(KEYINPUT26), .ZN(n573) );
  NOR2_X1 U510 ( .A1(n573), .A2(n454), .ZN(n545) );
  NOR2_X1 U511 ( .A1(n489), .A2(n527), .ZN(n455) );
  XOR2_X1 U512 ( .A(KEYINPUT91), .B(n455), .Z(n456) );
  NOR2_X1 U513 ( .A1(n457), .A2(n456), .ZN(n458) );
  XOR2_X1 U514 ( .A(KEYINPUT25), .B(n458), .Z(n459) );
  NOR2_X1 U515 ( .A1(n545), .A2(n459), .ZN(n460) );
  NOR2_X1 U516 ( .A1(n515), .A2(n460), .ZN(n461) );
  NOR2_X1 U517 ( .A1(n462), .A2(n461), .ZN(n479) );
  NOR2_X1 U518 ( .A1(n565), .A2(n480), .ZN(n464) );
  XNOR2_X1 U519 ( .A(KEYINPUT16), .B(KEYINPUT80), .ZN(n463) );
  XNOR2_X1 U520 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U521 ( .A(KEYINPUT79), .B(n465), .ZN(n466) );
  NOR2_X1 U522 ( .A1(n479), .A2(n466), .ZN(n499) );
  NOR2_X1 U523 ( .A1(n396), .A2(n531), .ZN(n484) );
  NAND2_X1 U524 ( .A1(n499), .A2(n484), .ZN(n467) );
  XOR2_X1 U525 ( .A(KEYINPUT92), .B(n467), .Z(n476) );
  NAND2_X1 U526 ( .A1(n476), .A2(n515), .ZN(n471) );
  XOR2_X1 U527 ( .A(KEYINPUT34), .B(KEYINPUT93), .Z(n469) );
  XNOR2_X1 U528 ( .A(G1GAT), .B(KEYINPUT94), .ZN(n468) );
  XNOR2_X1 U529 ( .A(n469), .B(n468), .ZN(n470) );
  XNOR2_X1 U530 ( .A(n471), .B(n470), .ZN(G1324GAT) );
  NAND2_X1 U531 ( .A1(n476), .A2(n517), .ZN(n472) );
  XNOR2_X1 U532 ( .A(n472), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U533 ( .A(KEYINPUT35), .B(KEYINPUT95), .Z(n474) );
  NAND2_X1 U534 ( .A1(n520), .A2(n476), .ZN(n473) );
  XNOR2_X1 U535 ( .A(n474), .B(n473), .ZN(n475) );
  XOR2_X1 U536 ( .A(G15GAT), .B(n475), .Z(G1326GAT) );
  NAND2_X1 U537 ( .A1(n476), .A2(n522), .ZN(n477) );
  XNOR2_X1 U538 ( .A(n477), .B(KEYINPUT96), .ZN(n478) );
  XNOR2_X1 U539 ( .A(G22GAT), .B(n478), .ZN(G1327GAT) );
  XNOR2_X1 U540 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n488) );
  XOR2_X1 U541 ( .A(KEYINPUT99), .B(KEYINPUT38), .Z(n486) );
  XNOR2_X1 U542 ( .A(KEYINPUT37), .B(KEYINPUT98), .ZN(n483) );
  NOR2_X1 U543 ( .A1(n587), .A2(n479), .ZN(n481) );
  NAND2_X1 U544 ( .A1(n481), .A2(n480), .ZN(n482) );
  XNOR2_X1 U545 ( .A(n483), .B(n482), .ZN(n512) );
  NAND2_X1 U546 ( .A1(n484), .A2(n512), .ZN(n485) );
  XNOR2_X1 U547 ( .A(n486), .B(n485), .ZN(n495) );
  NOR2_X1 U548 ( .A1(n570), .A2(n495), .ZN(n487) );
  XNOR2_X1 U549 ( .A(n488), .B(n487), .ZN(G1328GAT) );
  NOR2_X1 U550 ( .A1(n489), .A2(n495), .ZN(n490) );
  XOR2_X1 U551 ( .A(KEYINPUT100), .B(n490), .Z(n491) );
  XNOR2_X1 U552 ( .A(G36GAT), .B(n491), .ZN(G1329GAT) );
  NOR2_X1 U553 ( .A1(n495), .A2(n527), .ZN(n493) );
  XNOR2_X1 U554 ( .A(KEYINPUT40), .B(KEYINPUT101), .ZN(n492) );
  XNOR2_X1 U555 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U556 ( .A(G43GAT), .B(n494), .ZN(G1330GAT) );
  INV_X1 U557 ( .A(n522), .ZN(n496) );
  NOR2_X1 U558 ( .A1(n496), .A2(n495), .ZN(n497) );
  XOR2_X1 U559 ( .A(G50GAT), .B(n497), .Z(G1331GAT) );
  XOR2_X1 U560 ( .A(G57GAT), .B(KEYINPUT102), .Z(n502) );
  NAND2_X1 U561 ( .A1(n531), .A2(n533), .ZN(n498) );
  XOR2_X1 U562 ( .A(KEYINPUT104), .B(n498), .Z(n513) );
  NAND2_X1 U563 ( .A1(n513), .A2(n499), .ZN(n500) );
  XNOR2_X1 U564 ( .A(n500), .B(KEYINPUT105), .ZN(n509) );
  NAND2_X1 U565 ( .A1(n509), .A2(n515), .ZN(n501) );
  XNOR2_X1 U566 ( .A(n502), .B(n501), .ZN(n504) );
  XOR2_X1 U567 ( .A(KEYINPUT106), .B(KEYINPUT42), .Z(n503) );
  XNOR2_X1 U568 ( .A(n504), .B(n503), .ZN(G1332GAT) );
  XOR2_X1 U569 ( .A(G64GAT), .B(KEYINPUT107), .Z(n506) );
  NAND2_X1 U570 ( .A1(n509), .A2(n517), .ZN(n505) );
  XNOR2_X1 U571 ( .A(n506), .B(n505), .ZN(G1333GAT) );
  NAND2_X1 U572 ( .A1(n509), .A2(n520), .ZN(n507) );
  XNOR2_X1 U573 ( .A(n507), .B(KEYINPUT108), .ZN(n508) );
  XNOR2_X1 U574 ( .A(G71GAT), .B(n508), .ZN(G1334GAT) );
  XOR2_X1 U575 ( .A(G78GAT), .B(KEYINPUT43), .Z(n511) );
  NAND2_X1 U576 ( .A1(n509), .A2(n522), .ZN(n510) );
  XNOR2_X1 U577 ( .A(n511), .B(n510), .ZN(G1335GAT) );
  NAND2_X1 U578 ( .A1(n513), .A2(n512), .ZN(n514) );
  XNOR2_X1 U579 ( .A(n514), .B(KEYINPUT109), .ZN(n523) );
  NAND2_X1 U580 ( .A1(n515), .A2(n523), .ZN(n516) );
  XNOR2_X1 U581 ( .A(n516), .B(G85GAT), .ZN(G1336GAT) );
  NAND2_X1 U582 ( .A1(n517), .A2(n523), .ZN(n518) );
  XNOR2_X1 U583 ( .A(n518), .B(KEYINPUT110), .ZN(n519) );
  XNOR2_X1 U584 ( .A(G92GAT), .B(n519), .ZN(G1337GAT) );
  NAND2_X1 U585 ( .A1(n523), .A2(n520), .ZN(n521) );
  XNOR2_X1 U586 ( .A(n521), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U587 ( .A(KEYINPUT111), .B(KEYINPUT44), .Z(n525) );
  NAND2_X1 U588 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U589 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U590 ( .A(G106GAT), .B(n526), .ZN(G1339GAT) );
  NOR2_X1 U591 ( .A1(n527), .A2(n543), .ZN(n528) );
  NAND2_X1 U592 ( .A1(n529), .A2(n528), .ZN(n530) );
  XOR2_X1 U593 ( .A(KEYINPUT114), .B(n530), .Z(n539) );
  INV_X1 U594 ( .A(n531), .ZN(n574) );
  AND2_X1 U595 ( .A1(n539), .A2(n574), .ZN(n532) );
  XOR2_X1 U596 ( .A(G113GAT), .B(n532), .Z(G1340GAT) );
  XOR2_X1 U597 ( .A(G120GAT), .B(KEYINPUT49), .Z(n535) );
  NAND2_X1 U598 ( .A1(n533), .A2(n539), .ZN(n534) );
  XNOR2_X1 U599 ( .A(n535), .B(n534), .ZN(G1341GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT115), .B(KEYINPUT50), .Z(n537) );
  NAND2_X1 U601 ( .A1(n582), .A2(n539), .ZN(n536) );
  XNOR2_X1 U602 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U603 ( .A(G127GAT), .B(n538), .ZN(G1342GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT116), .B(KEYINPUT51), .Z(n541) );
  NAND2_X1 U605 ( .A1(n565), .A2(n539), .ZN(n540) );
  XNOR2_X1 U606 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U607 ( .A(G134GAT), .B(n542), .ZN(G1343GAT) );
  INV_X1 U608 ( .A(KEYINPUT117), .ZN(n547) );
  NOR2_X1 U609 ( .A1(n570), .A2(n543), .ZN(n544) );
  NAND2_X1 U610 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U611 ( .A(n547), .B(n546), .ZN(n559) );
  INV_X1 U612 ( .A(n559), .ZN(n556) );
  NAND2_X1 U613 ( .A1(n574), .A2(n556), .ZN(n548) );
  XNOR2_X1 U614 ( .A(G141GAT), .B(n548), .ZN(G1344GAT) );
  NOR2_X1 U615 ( .A1(n549), .A2(n559), .ZN(n551) );
  XNOR2_X1 U616 ( .A(KEYINPUT119), .B(KEYINPUT53), .ZN(n550) );
  XNOR2_X1 U617 ( .A(n551), .B(n550), .ZN(n553) );
  INV_X1 U618 ( .A(KEYINPUT118), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n553), .B(n552), .ZN(n555) );
  XNOR2_X1 U620 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n555), .B(n554), .ZN(G1345GAT) );
  NAND2_X1 U622 ( .A1(n556), .A2(n582), .ZN(n557) );
  XNOR2_X1 U623 ( .A(n557), .B(KEYINPUT120), .ZN(n558) );
  XNOR2_X1 U624 ( .A(G155GAT), .B(n558), .ZN(G1346GAT) );
  NOR2_X1 U625 ( .A1(n560), .A2(n559), .ZN(n562) );
  XNOR2_X1 U626 ( .A(G162GAT), .B(KEYINPUT121), .ZN(n561) );
  XNOR2_X1 U627 ( .A(n562), .B(n561), .ZN(G1347GAT) );
  NAND2_X1 U628 ( .A1(n566), .A2(n574), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n563), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U630 ( .A1(n566), .A2(n582), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n564), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U632 ( .A1(n566), .A2(n565), .ZN(n568) );
  XOR2_X1 U633 ( .A(KEYINPUT123), .B(KEYINPUT58), .Z(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n569), .B(G190GAT), .ZN(G1351GAT) );
  NAND2_X1 U636 ( .A1(n571), .A2(n570), .ZN(n572) );
  NOR2_X1 U637 ( .A1(n573), .A2(n572), .ZN(n585) );
  NAND2_X1 U638 ( .A1(n585), .A2(n574), .ZN(n578) );
  XOR2_X1 U639 ( .A(KEYINPUT60), .B(KEYINPUT124), .Z(n576) );
  XNOR2_X1 U640 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U642 ( .A(n578), .B(n577), .ZN(G1352GAT) );
  XOR2_X1 U643 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n580) );
  NAND2_X1 U644 ( .A1(n585), .A2(n396), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(n581) );
  XOR2_X1 U646 ( .A(G204GAT), .B(n581), .Z(G1353GAT) );
  NAND2_X1 U647 ( .A1(n585), .A2(n582), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n583), .B(KEYINPUT126), .ZN(n584) );
  XNOR2_X1 U649 ( .A(G211GAT), .B(n584), .ZN(G1354GAT) );
  INV_X1 U650 ( .A(n585), .ZN(n586) );
  NOR2_X1 U651 ( .A1(n587), .A2(n586), .ZN(n589) );
  XNOR2_X1 U652 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n588) );
  XNOR2_X1 U653 ( .A(n589), .B(n588), .ZN(n590) );
  XNOR2_X1 U654 ( .A(G218GAT), .B(n590), .ZN(G1355GAT) );
endmodule

