//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 0 1 1 0 1 1 1 0 1 1 0 0 1 1 1 1 1 0 1 1 0 0 1 1 0 1 0 0 1 1 1 0 1 0 0 0 1 1 1 0 1 1 0 1 1 1 1 1 1 0 1 1 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:52 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n746, new_n747, new_n748, new_n749,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n762, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n805, new_n806, new_n807, new_n808, new_n809, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n860, new_n861, new_n863,
    new_n864, new_n865, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n917, new_n918, new_n920, new_n921, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n936, new_n937, new_n938, new_n939, new_n940, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n972,
    new_n973, new_n974, new_n975, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n983, new_n984;
  XOR2_X1   g000(.A(G15gat), .B(G43gat), .Z(new_n202));
  XNOR2_X1  g001(.A(G71gat), .B(G99gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT25), .ZN(new_n206));
  NAND2_X1  g005(.A1(G169gat), .A2(G176gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(KEYINPUT23), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n208), .B1(G169gat), .B2(G176gat), .ZN(new_n209));
  INV_X1    g008(.A(G169gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(KEYINPUT64), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT64), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(G169gat), .ZN(new_n213));
  INV_X1    g012(.A(G176gat), .ZN(new_n214));
  NAND4_X1  g013(.A1(new_n211), .A2(new_n213), .A3(KEYINPUT23), .A4(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n209), .A2(new_n215), .ZN(new_n216));
  AND3_X1   g015(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(G183gat), .A2(G190gat), .ZN(new_n218));
  OAI21_X1  g017(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n217), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n206), .B1(new_n216), .B2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT65), .ZN(new_n222));
  NOR2_X1   g021(.A1(G169gat), .A2(G176gat), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n206), .B1(new_n223), .B2(KEYINPUT23), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n209), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n222), .B1(new_n225), .B2(new_n220), .ZN(new_n226));
  MUX2_X1   g025(.A(KEYINPUT24), .B(new_n219), .S(new_n218), .Z(new_n227));
  NAND4_X1  g026(.A1(new_n227), .A2(KEYINPUT65), .A3(new_n209), .A4(new_n224), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n221), .A2(new_n226), .A3(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT26), .ZN(new_n230));
  AND3_X1   g029(.A1(new_n223), .A2(KEYINPUT66), .A3(new_n230), .ZN(new_n231));
  AOI22_X1  g030(.A1(new_n223), .A2(KEYINPUT66), .B1(new_n207), .B2(new_n230), .ZN(new_n232));
  XNOR2_X1  g031(.A(KEYINPUT27), .B(G183gat), .ZN(new_n233));
  INV_X1    g032(.A(G190gat), .ZN(new_n234));
  AND3_X1   g033(.A1(new_n233), .A2(KEYINPUT28), .A3(new_n234), .ZN(new_n235));
  AOI21_X1  g034(.A(KEYINPUT28), .B1(new_n233), .B2(new_n234), .ZN(new_n236));
  OAI221_X1 g035(.A(new_n218), .B1(new_n231), .B2(new_n232), .C1(new_n235), .C2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n229), .A2(new_n237), .ZN(new_n238));
  XOR2_X1   g037(.A(G127gat), .B(G134gat), .Z(new_n239));
  XNOR2_X1  g038(.A(G113gat), .B(G120gat), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n239), .B1(new_n240), .B2(KEYINPUT1), .ZN(new_n241));
  XOR2_X1   g040(.A(G113gat), .B(G120gat), .Z(new_n242));
  XNOR2_X1  g041(.A(G127gat), .B(G134gat), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT1), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n242), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  AND2_X1   g044(.A1(new_n241), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n238), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(G227gat), .ZN(new_n248));
  INV_X1    g047(.A(G233gat), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n241), .A2(new_n245), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n229), .A2(new_n251), .A3(new_n237), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n247), .A2(new_n250), .A3(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT32), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(KEYINPUT33), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n205), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n254), .B1(new_n204), .B2(KEYINPUT33), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n253), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n258), .A2(KEYINPUT67), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT67), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n253), .A2(new_n260), .A3(new_n257), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n256), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n250), .B1(new_n247), .B2(new_n252), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT34), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(KEYINPUT68), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT68), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n263), .A2(new_n267), .A3(new_n264), .ZN(new_n268));
  OR2_X1    g067(.A1(new_n263), .A2(new_n264), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n262), .A2(new_n266), .A3(new_n268), .A4(new_n269), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n266), .A2(new_n269), .A3(new_n268), .ZN(new_n271));
  INV_X1    g070(.A(new_n261), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n260), .B1(new_n253), .B2(new_n257), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n271), .B1(new_n274), .B2(new_n256), .ZN(new_n275));
  AND3_X1   g074(.A1(new_n270), .A2(new_n275), .A3(KEYINPUT36), .ZN(new_n276));
  AOI21_X1  g075(.A(KEYINPUT36), .B1(new_n270), .B2(new_n275), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT79), .ZN(new_n279));
  NAND2_X1  g078(.A1(G155gat), .A2(G162gat), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  NOR2_X1   g080(.A1(G155gat), .A2(G162gat), .ZN(new_n282));
  OAI21_X1  g081(.A(KEYINPUT77), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(G155gat), .ZN(new_n284));
  INV_X1    g083(.A(G162gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT77), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n286), .A2(new_n287), .A3(new_n280), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n283), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(G148gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(KEYINPUT76), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT76), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(G148gat), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n291), .A2(new_n293), .A3(G141gat), .ZN(new_n294));
  INV_X1    g093(.A(G141gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(G148gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n280), .A2(KEYINPUT2), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n289), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  AND2_X1   g098(.A1(KEYINPUT74), .A2(KEYINPUT2), .ZN(new_n300));
  NOR2_X1   g099(.A1(KEYINPUT74), .A2(KEYINPUT2), .ZN(new_n301));
  OAI21_X1  g100(.A(KEYINPUT75), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT74), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT2), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT75), .ZN(new_n306));
  NAND2_X1  g105(.A1(KEYINPUT74), .A2(KEYINPUT2), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n305), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n290), .A2(G141gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n296), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n302), .A2(new_n308), .A3(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT73), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n282), .A2(new_n312), .ZN(new_n313));
  OAI21_X1  g112(.A(KEYINPUT73), .B1(G155gat), .B2(G162gat), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n281), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n311), .A2(new_n315), .ZN(new_n316));
  XOR2_X1   g115(.A(KEYINPUT78), .B(KEYINPUT3), .Z(new_n317));
  NAND3_X1  g116(.A1(new_n299), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(new_n251), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT3), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n320), .B1(new_n299), .B2(new_n316), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n279), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  AOI22_X1  g121(.A1(new_n294), .A2(new_n296), .B1(KEYINPUT2), .B2(new_n280), .ZN(new_n323));
  AOI22_X1  g122(.A1(new_n289), .A2(new_n323), .B1(new_n311), .B2(new_n315), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n246), .B1(new_n324), .B2(new_n317), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n299), .A2(new_n316), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(KEYINPUT3), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n325), .A2(KEYINPUT79), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n322), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT81), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n330), .B1(new_n326), .B2(new_n251), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n324), .A2(KEYINPUT81), .A3(new_n246), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n331), .A2(KEYINPUT4), .A3(new_n332), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n326), .A2(new_n251), .ZN(new_n334));
  XNOR2_X1  g133(.A(KEYINPUT80), .B(KEYINPUT4), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n333), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT5), .ZN(new_n338));
  NAND2_X1  g137(.A1(G225gat), .A2(G233gat), .ZN(new_n339));
  NAND4_X1  g138(.A1(new_n329), .A2(new_n337), .A3(new_n338), .A4(new_n339), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n334), .A2(new_n335), .ZN(new_n341));
  AOI21_X1  g140(.A(KEYINPUT4), .B1(new_n331), .B2(new_n332), .ZN(new_n342));
  OAI211_X1 g141(.A(new_n329), .B(new_n339), .C1(new_n341), .C2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT83), .ZN(new_n344));
  NOR3_X1   g143(.A1(new_n324), .A2(new_n246), .A3(KEYINPUT82), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT82), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n346), .B1(new_n326), .B2(new_n251), .ZN(new_n347));
  OAI211_X1 g146(.A(new_n331), .B(new_n332), .C1(new_n345), .C2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(new_n339), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n338), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  AND3_X1   g149(.A1(new_n343), .A2(new_n344), .A3(new_n350), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n344), .B1(new_n343), .B2(new_n350), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n340), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  XNOR2_X1  g152(.A(G1gat), .B(G29gat), .ZN(new_n354));
  XNOR2_X1  g153(.A(new_n354), .B(KEYINPUT0), .ZN(new_n355));
  XNOR2_X1  g154(.A(G57gat), .B(G85gat), .ZN(new_n356));
  XOR2_X1   g155(.A(new_n355), .B(new_n356), .Z(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n353), .A2(KEYINPUT6), .A3(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT6), .ZN(new_n360));
  INV_X1    g159(.A(new_n340), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n339), .B1(new_n342), .B2(new_n341), .ZN(new_n362));
  NOR3_X1   g161(.A1(new_n319), .A2(new_n279), .A3(new_n321), .ZN(new_n363));
  AOI21_X1  g162(.A(KEYINPUT79), .B1(new_n325), .B2(new_n327), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n362), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n348), .A2(new_n349), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(KEYINPUT5), .ZN(new_n368));
  OAI21_X1  g167(.A(KEYINPUT83), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n343), .A2(new_n344), .A3(new_n350), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n361), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n360), .B1(new_n371), .B2(new_n357), .ZN(new_n372));
  OAI211_X1 g171(.A(new_n357), .B(new_n340), .C1(new_n351), .C2(new_n352), .ZN(new_n373));
  INV_X1    g172(.A(new_n373), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n359), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  XOR2_X1   g174(.A(G211gat), .B(G218gat), .Z(new_n376));
  INV_X1    g175(.A(KEYINPUT70), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT69), .ZN(new_n379));
  XNOR2_X1  g178(.A(G211gat), .B(G218gat), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(KEYINPUT70), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n378), .A2(new_n379), .A3(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT22), .ZN(new_n383));
  INV_X1    g182(.A(G211gat), .ZN(new_n384));
  INV_X1    g183(.A(G218gat), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n383), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(G204gat), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(G197gat), .ZN(new_n388));
  INV_X1    g187(.A(G197gat), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(G204gat), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n386), .A2(new_n388), .A3(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n382), .A2(new_n392), .ZN(new_n393));
  NAND4_X1  g192(.A1(new_n378), .A2(new_n379), .A3(new_n391), .A4(new_n381), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g194(.A(KEYINPUT29), .B1(new_n229), .B2(new_n237), .ZN(new_n396));
  NAND2_X1  g195(.A1(G226gat), .A2(G233gat), .ZN(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n397), .B1(new_n229), .B2(new_n237), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n395), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n400), .ZN(new_n402));
  INV_X1    g201(.A(new_n395), .ZN(new_n403));
  OAI211_X1 g202(.A(new_n402), .B(new_n403), .C1(new_n398), .C2(new_n396), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n401), .A2(new_n404), .ZN(new_n405));
  XNOR2_X1  g204(.A(G8gat), .B(G36gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(G64gat), .B(G92gat), .ZN(new_n407));
  XNOR2_X1  g206(.A(new_n406), .B(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n405), .A2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT30), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n410), .A2(KEYINPUT72), .A3(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT72), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n408), .B1(new_n401), .B2(new_n404), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n413), .B1(new_n414), .B2(KEYINPUT30), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n412), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n405), .A2(KEYINPUT30), .A3(new_n409), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n401), .A2(new_n408), .A3(new_n404), .ZN(new_n418));
  AND3_X1   g217(.A1(new_n417), .A2(KEYINPUT71), .A3(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(KEYINPUT71), .B1(new_n417), .B2(new_n418), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n416), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n375), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(G228gat), .A2(G233gat), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT29), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n395), .B1(new_n426), .B2(new_n318), .ZN(new_n427));
  AOI21_X1  g226(.A(KEYINPUT3), .B1(new_n395), .B2(new_n426), .ZN(new_n428));
  OAI22_X1  g227(.A1(new_n427), .A2(KEYINPUT85), .B1(new_n428), .B2(new_n324), .ZN(new_n429));
  AND2_X1   g228(.A1(new_n427), .A2(KEYINPUT85), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n425), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n378), .A2(new_n381), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n432), .B(new_n391), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n317), .B1(new_n433), .B2(KEYINPUT29), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(new_n326), .ZN(new_n435));
  INV_X1    g234(.A(new_n427), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n435), .A2(new_n424), .A3(new_n436), .ZN(new_n437));
  XNOR2_X1  g236(.A(G78gat), .B(G106gat), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n438), .B(KEYINPUT84), .ZN(new_n439));
  XNOR2_X1  g238(.A(KEYINPUT31), .B(G50gat), .ZN(new_n440));
  XNOR2_X1  g239(.A(new_n439), .B(new_n440), .ZN(new_n441));
  XNOR2_X1  g240(.A(new_n441), .B(G22gat), .ZN(new_n442));
  AND3_X1   g241(.A1(new_n431), .A2(new_n437), .A3(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n442), .B1(new_n431), .B2(new_n437), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(KEYINPUT86), .ZN(new_n447));
  OR3_X1    g246(.A1(new_n443), .A2(new_n444), .A3(KEYINPUT86), .ZN(new_n448));
  AND2_X1   g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n278), .B1(new_n423), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n417), .A2(new_n418), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n416), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n353), .A2(new_n358), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n339), .B1(new_n329), .B2(new_n337), .ZN(new_n455));
  OAI21_X1  g254(.A(KEYINPUT39), .B1(new_n348), .B2(new_n349), .ZN(new_n456));
  OR2_X1    g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT39), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n455), .A2(new_n458), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n457), .A2(KEYINPUT40), .A3(new_n357), .A4(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT40), .ZN(new_n461));
  INV_X1    g260(.A(new_n459), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n357), .B1(new_n455), .B2(new_n456), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n461), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n453), .A2(new_n454), .A3(new_n460), .A4(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT88), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT37), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n466), .B1(new_n405), .B2(new_n467), .ZN(new_n468));
  AOI211_X1 g267(.A(KEYINPUT88), .B(KEYINPUT37), .C1(new_n401), .C2(new_n404), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n401), .A2(KEYINPUT37), .A3(new_n404), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(new_n408), .ZN(new_n472));
  OAI21_X1  g271(.A(KEYINPUT38), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n471), .A2(KEYINPUT87), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT87), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n401), .A2(new_n404), .A3(new_n475), .A4(KEYINPUT37), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n409), .A2(KEYINPUT38), .ZN(new_n478));
  OAI211_X1 g277(.A(new_n477), .B(new_n478), .C1(new_n468), .C2(new_n469), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n473), .A2(new_n410), .A3(new_n479), .ZN(new_n480));
  OAI211_X1 g279(.A(new_n445), .B(new_n465), .C1(new_n375), .C2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n450), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n445), .A2(new_n270), .A3(new_n275), .ZN(new_n483));
  INV_X1    g282(.A(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT35), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n451), .B1(new_n415), .B2(new_n412), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n375), .A2(new_n484), .A3(new_n485), .A4(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n454), .A2(new_n360), .A3(new_n373), .ZN(new_n488));
  AOI211_X1 g287(.A(new_n483), .B(new_n421), .C1(new_n488), .C2(new_n359), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n487), .B1(new_n489), .B2(new_n485), .ZN(new_n490));
  AND2_X1   g289(.A1(new_n482), .A2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT92), .ZN(new_n492));
  XNOR2_X1  g291(.A(G15gat), .B(G22gat), .ZN(new_n493));
  OR2_X1    g292(.A1(new_n493), .A2(G1gat), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT16), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n493), .B1(new_n495), .B2(G1gat), .ZN(new_n496));
  INV_X1    g295(.A(G8gat), .ZN(new_n497));
  OR2_X1    g296(.A1(new_n497), .A2(KEYINPUT91), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n494), .A2(new_n496), .A3(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n499), .A2(KEYINPUT91), .A3(new_n497), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n497), .A2(KEYINPUT91), .ZN(new_n501));
  NAND4_X1  g300(.A1(new_n494), .A2(new_n496), .A3(new_n498), .A4(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n492), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT14), .ZN(new_n505));
  INV_X1    g304(.A(G29gat), .ZN(new_n506));
  INV_X1    g305(.A(G36gat), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n505), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  OAI21_X1  g307(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n509));
  AOI22_X1  g308(.A1(new_n508), .A2(new_n509), .B1(G29gat), .B2(G36gat), .ZN(new_n510));
  XNOR2_X1  g309(.A(G43gat), .B(G50gat), .ZN(new_n511));
  AOI22_X1  g310(.A1(new_n510), .A2(KEYINPUT90), .B1(KEYINPUT15), .B2(new_n511), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n510), .B1(KEYINPUT15), .B2(new_n511), .ZN(new_n513));
  OR2_X1    g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n512), .A2(new_n513), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(new_n516), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n500), .A2(new_n492), .A3(new_n502), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n504), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(G229gat), .A2(G233gat), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n516), .B(KEYINPUT17), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n500), .A2(new_n502), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  OAI211_X1 g322(.A(new_n519), .B(new_n520), .C1(new_n521), .C2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT18), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n517), .A2(KEYINPUT17), .ZN(new_n527));
  AND3_X1   g326(.A1(new_n514), .A2(KEYINPUT17), .A3(new_n515), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n522), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n529), .A2(KEYINPUT18), .A3(new_n519), .A4(new_n520), .ZN(new_n530));
  AND2_X1   g329(.A1(new_n526), .A2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(new_n518), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n516), .B1(new_n532), .B2(new_n503), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(new_n519), .ZN(new_n534));
  XOR2_X1   g333(.A(new_n520), .B(KEYINPUT13), .Z(new_n535));
  AOI21_X1  g334(.A(KEYINPUT93), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT93), .ZN(new_n537));
  INV_X1    g336(.A(new_n535), .ZN(new_n538));
  AOI211_X1 g337(.A(new_n537), .B(new_n538), .C1(new_n533), .C2(new_n519), .ZN(new_n539));
  OR2_X1    g338(.A1(new_n536), .A2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT94), .ZN(new_n541));
  XOR2_X1   g340(.A(G113gat), .B(G141gat), .Z(new_n542));
  XNOR2_X1  g341(.A(new_n542), .B(KEYINPUT11), .ZN(new_n543));
  XOR2_X1   g342(.A(new_n543), .B(KEYINPUT89), .Z(new_n544));
  XNOR2_X1  g343(.A(G169gat), .B(G197gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n544), .B(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n546), .B(KEYINPUT12), .ZN(new_n547));
  NAND4_X1  g346(.A1(new_n531), .A2(new_n540), .A3(new_n541), .A4(new_n547), .ZN(new_n548));
  OAI211_X1 g347(.A(new_n526), .B(new_n530), .C1(new_n536), .C2(new_n539), .ZN(new_n549));
  INV_X1    g348(.A(new_n547), .ZN(new_n550));
  OAI21_X1  g349(.A(KEYINPUT94), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n549), .A2(new_n550), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  XOR2_X1   g354(.A(G183gat), .B(G211gat), .Z(new_n556));
  OR2_X1    g355(.A1(G57gat), .A2(G64gat), .ZN(new_n557));
  NAND2_X1  g356(.A1(G57gat), .A2(G64gat), .ZN(new_n558));
  INV_X1    g357(.A(G71gat), .ZN(new_n559));
  INV_X1    g358(.A(G78gat), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  OAI211_X1 g360(.A(new_n557), .B(new_n558), .C1(new_n561), .C2(KEYINPUT9), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT95), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NOR2_X1   g363(.A1(G71gat), .A2(G78gat), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n561), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  OAI211_X1 g366(.A(new_n562), .B(new_n563), .C1(new_n561), .C2(new_n565), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n569), .A2(KEYINPUT21), .ZN(new_n570));
  NAND2_X1  g369(.A1(G231gat), .A2(G233gat), .ZN(new_n571));
  XOR2_X1   g370(.A(new_n570), .B(new_n571), .Z(new_n572));
  XNOR2_X1  g371(.A(G127gat), .B(G155gat), .ZN(new_n573));
  OR2_X1    g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n572), .A2(new_n573), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  XOR2_X1   g375(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  AOI22_X1  g377(.A1(new_n504), .A2(new_n518), .B1(KEYINPUT21), .B2(new_n569), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n577), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n574), .A2(new_n575), .A3(new_n581), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n578), .A2(new_n580), .A3(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n580), .B1(new_n578), .B2(new_n582), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n556), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n578), .A2(new_n582), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(new_n579), .ZN(new_n588));
  INV_X1    g387(.A(new_n556), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n588), .A2(new_n583), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n586), .A2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n593));
  NAND2_X1  g392(.A1(G99gat), .A2(G106gat), .ZN(new_n594));
  INV_X1    g393(.A(G85gat), .ZN(new_n595));
  INV_X1    g394(.A(G92gat), .ZN(new_n596));
  AOI22_X1  g395(.A1(KEYINPUT8), .A2(new_n594), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT7), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n598), .B1(new_n595), .B2(new_n596), .ZN(new_n599));
  NAND3_X1  g398(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n597), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(G99gat), .B(G106gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n593), .B1(new_n516), .B2(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(KEYINPUT96), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n604), .B1(new_n527), .B2(new_n528), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(G190gat), .B(G218gat), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  AOI21_X1  g409(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n609), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n606), .A2(new_n607), .A3(new_n613), .ZN(new_n614));
  AND3_X1   g413(.A1(new_n610), .A2(new_n612), .A3(new_n614), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n612), .B1(new_n610), .B2(new_n614), .ZN(new_n616));
  XOR2_X1   g415(.A(G134gat), .B(G162gat), .Z(new_n617));
  OR3_X1    g416(.A1(new_n615), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n617), .B1(new_n615), .B2(new_n616), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n592), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n569), .A2(KEYINPUT97), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT97), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n567), .A2(new_n623), .A3(new_n568), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n622), .A2(new_n603), .A3(new_n624), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n604), .A2(KEYINPUT97), .A3(new_n569), .ZN(new_n626));
  AOI21_X1  g425(.A(KEYINPUT10), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  AND3_X1   g426(.A1(new_n569), .A2(new_n603), .A3(KEYINPUT10), .ZN(new_n628));
  OR2_X1    g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(G230gat), .A2(G233gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(KEYINPUT98), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n625), .A2(new_n626), .ZN(new_n633));
  OR2_X1    g432(.A1(new_n633), .A2(new_n630), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(G120gat), .B(G148gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(G176gat), .B(G204gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n635), .A2(new_n638), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n630), .B1(new_n627), .B2(new_n628), .ZN(new_n640));
  INV_X1    g439(.A(new_n638), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n640), .A2(new_n634), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n639), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n621), .A2(new_n644), .ZN(new_n645));
  NOR3_X1   g444(.A1(new_n491), .A2(new_n555), .A3(new_n645), .ZN(new_n646));
  NOR3_X1   g445(.A1(new_n371), .A2(new_n360), .A3(new_n357), .ZN(new_n647));
  AOI21_X1  g446(.A(KEYINPUT6), .B1(new_n353), .B2(new_n358), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n647), .B1(new_n373), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n650), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g450(.A1(new_n646), .A2(new_n453), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n652), .A2(G8gat), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n653), .A2(KEYINPUT42), .ZN(new_n654));
  XNOR2_X1  g453(.A(KEYINPUT16), .B(G8gat), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  MUX2_X1   g455(.A(new_n654), .B(KEYINPUT42), .S(new_n656), .Z(G1325gat));
  INV_X1    g456(.A(new_n646), .ZN(new_n658));
  INV_X1    g457(.A(new_n278), .ZN(new_n659));
  OAI21_X1  g458(.A(G15gat), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n270), .A2(new_n275), .ZN(new_n661));
  OR2_X1    g460(.A1(new_n661), .A2(G15gat), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n660), .B1(new_n658), .B2(new_n662), .ZN(G1326gat));
  NAND2_X1  g462(.A1(new_n646), .A2(new_n449), .ZN(new_n664));
  XNOR2_X1  g463(.A(KEYINPUT43), .B(G22gat), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n664), .B(new_n665), .ZN(G1327gat));
  NOR2_X1   g465(.A1(new_n591), .A2(new_n643), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n667), .A2(new_n620), .ZN(new_n668));
  XOR2_X1   g467(.A(new_n668), .B(KEYINPUT99), .Z(new_n669));
  NOR2_X1   g468(.A1(new_n491), .A2(new_n555), .ZN(new_n670));
  AND2_X1   g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n671), .A2(new_n506), .A3(new_n649), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(KEYINPUT45), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n421), .B1(new_n488), .B2(new_n359), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n447), .A2(new_n448), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n659), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  OAI211_X1 g475(.A(new_n460), .B(new_n464), .C1(new_n371), .C2(new_n357), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n445), .B1(new_n677), .B2(new_n486), .ZN(new_n678));
  INV_X1    g477(.A(new_n480), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n678), .B1(new_n679), .B2(new_n649), .ZN(new_n680));
  OAI21_X1  g479(.A(KEYINPUT102), .B1(new_n676), .B2(new_n680), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n449), .B1(new_n649), .B2(new_n421), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT102), .ZN(new_n683));
  NAND4_X1  g482(.A1(new_n682), .A2(new_n481), .A3(new_n683), .A4(new_n659), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n681), .A2(new_n490), .A3(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT103), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT44), .ZN(new_n687));
  NAND4_X1  g486(.A1(new_n685), .A2(new_n686), .A3(new_n687), .A4(new_n620), .ZN(new_n688));
  INV_X1    g487(.A(new_n620), .ZN(new_n689));
  OAI21_X1  g488(.A(KEYINPUT44), .B1(new_n491), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n685), .A2(new_n687), .A3(new_n620), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(KEYINPUT103), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n554), .A2(KEYINPUT100), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT100), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n552), .A2(new_n697), .A3(new_n553), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(new_n667), .ZN(new_n701));
  XOR2_X1   g500(.A(new_n701), .B(KEYINPUT101), .Z(new_n702));
  NAND2_X1  g501(.A1(new_n695), .A2(new_n702), .ZN(new_n703));
  OAI21_X1  g502(.A(G29gat), .B1(new_n703), .B2(new_n375), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n673), .A2(new_n704), .ZN(G1328gat));
  NAND3_X1  g504(.A1(new_n671), .A2(new_n507), .A3(new_n453), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT104), .ZN(new_n707));
  OR3_X1    g506(.A1(new_n706), .A2(new_n707), .A3(KEYINPUT46), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n707), .B1(new_n706), .B2(KEYINPUT46), .ZN(new_n709));
  AOI22_X1  g508(.A1(new_n708), .A2(new_n709), .B1(KEYINPUT46), .B2(new_n706), .ZN(new_n710));
  OAI21_X1  g509(.A(G36gat), .B1(new_n703), .B2(new_n486), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(G1329gat));
  INV_X1    g511(.A(G43gat), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n669), .A2(new_n670), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n713), .B1(new_n714), .B2(new_n661), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n659), .A2(new_n713), .ZN(new_n716));
  INV_X1    g515(.A(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n715), .B1(new_n703), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(KEYINPUT47), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT47), .ZN(new_n720));
  OAI211_X1 g519(.A(new_n720), .B(new_n715), .C1(new_n703), .C2(new_n717), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n719), .A2(new_n721), .ZN(G1330gat));
  OAI21_X1  g521(.A(G50gat), .B1(new_n703), .B2(new_n445), .ZN(new_n723));
  OR2_X1    g522(.A1(new_n675), .A2(G50gat), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n671), .A2(KEYINPUT105), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT105), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n714), .A2(new_n726), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n724), .B1(new_n725), .B2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT48), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n723), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n695), .A2(new_n449), .A3(new_n702), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n728), .B1(new_n732), .B2(G50gat), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n731), .B1(KEYINPUT48), .B2(new_n733), .ZN(G1331gat));
  NAND3_X1  g533(.A1(new_n621), .A2(new_n643), .A3(new_n699), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(KEYINPUT106), .ZN(new_n736));
  INV_X1    g535(.A(new_n685), .ZN(new_n737));
  OAI21_X1  g536(.A(KEYINPUT107), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT106), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n735), .B(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT107), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n740), .A2(new_n741), .A3(new_n685), .ZN(new_n742));
  AND2_X1   g541(.A1(new_n738), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(new_n649), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g544(.A(new_n486), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n743), .A2(new_n746), .ZN(new_n747));
  NOR2_X1   g546(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(KEYINPUT108), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n747), .B(new_n749), .ZN(G1333gat));
  XNOR2_X1  g549(.A(new_n661), .B(KEYINPUT109), .ZN(new_n751));
  INV_X1    g550(.A(new_n751), .ZN(new_n752));
  NAND4_X1  g551(.A1(new_n738), .A2(new_n742), .A3(new_n559), .A4(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n738), .A2(new_n742), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n754), .A2(new_n659), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n753), .B1(new_n755), .B2(new_n559), .ZN(new_n756));
  XOR2_X1   g555(.A(KEYINPUT110), .B(KEYINPUT50), .Z(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(new_n757), .ZN(new_n759));
  OAI211_X1 g558(.A(new_n753), .B(new_n759), .C1(new_n755), .C2(new_n559), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n758), .A2(new_n760), .ZN(G1334gat));
  NOR2_X1   g560(.A1(new_n754), .A2(new_n675), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(new_n560), .ZN(G1335gat));
  NAND3_X1  g562(.A1(new_n649), .A2(new_n595), .A3(new_n643), .ZN(new_n764));
  INV_X1    g563(.A(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT51), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT112), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n684), .A2(new_n490), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n683), .B1(new_n450), .B2(new_n481), .ZN(new_n769));
  OAI211_X1 g568(.A(new_n767), .B(new_n620), .C1(new_n768), .C2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n699), .A2(new_n592), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n771), .B(KEYINPUT111), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n767), .B1(new_n685), .B2(new_n620), .ZN(new_n774));
  OAI211_X1 g573(.A(KEYINPUT113), .B(new_n766), .C1(new_n773), .C2(new_n774), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n620), .B1(new_n768), .B2(new_n769), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(KEYINPUT112), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n777), .A2(KEYINPUT51), .A3(new_n772), .A4(new_n770), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n775), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n777), .A2(new_n772), .A3(new_n770), .ZN(new_n780));
  AOI21_X1  g579(.A(KEYINPUT113), .B1(new_n780), .B2(new_n766), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n765), .B1(new_n779), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n772), .A2(new_n643), .ZN(new_n783));
  INV_X1    g582(.A(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(new_n694), .ZN(new_n785));
  OAI211_X1 g584(.A(new_n649), .B(new_n784), .C1(new_n785), .C2(new_n691), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(G85gat), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n782), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(KEYINPUT114), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT114), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n782), .A2(new_n790), .A3(new_n787), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n789), .A2(new_n791), .ZN(G1336gat));
  NAND3_X1  g591(.A1(new_n695), .A2(new_n453), .A3(new_n784), .ZN(new_n793));
  AOI21_X1  g592(.A(KEYINPUT52), .B1(new_n793), .B2(G92gat), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n644), .A2(new_n486), .A3(G92gat), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n795), .B1(new_n779), .B2(new_n781), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n783), .B1(new_n692), .B2(new_n694), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n596), .B1(new_n798), .B2(new_n453), .ZN(new_n799));
  INV_X1    g598(.A(new_n795), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n780), .A2(new_n766), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n800), .B1(new_n801), .B2(new_n778), .ZN(new_n802));
  OAI21_X1  g601(.A(KEYINPUT52), .B1(new_n799), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n797), .A2(new_n803), .ZN(G1337gat));
  NAND2_X1  g603(.A1(new_n798), .A2(new_n278), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(G99gat), .ZN(new_n806));
  NOR3_X1   g605(.A1(new_n644), .A2(new_n661), .A3(G99gat), .ZN(new_n807));
  XNOR2_X1  g606(.A(new_n807), .B(KEYINPUT115), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n808), .B1(new_n779), .B2(new_n781), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n806), .A2(new_n809), .ZN(G1338gat));
  NAND3_X1  g609(.A1(new_n695), .A2(new_n446), .A3(new_n784), .ZN(new_n811));
  AOI21_X1  g610(.A(KEYINPUT53), .B1(new_n811), .B2(G106gat), .ZN(new_n812));
  NOR3_X1   g611(.A1(new_n644), .A2(G106gat), .A3(new_n445), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n813), .B1(new_n779), .B2(new_n781), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(G106gat), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n816), .B1(new_n798), .B2(new_n449), .ZN(new_n817));
  INV_X1    g616(.A(new_n813), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n818), .B1(new_n801), .B2(new_n778), .ZN(new_n819));
  OAI21_X1  g618(.A(KEYINPUT53), .B1(new_n817), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n815), .A2(new_n820), .ZN(G1339gat));
  NAND2_X1  g620(.A1(new_n649), .A2(new_n486), .ZN(new_n822));
  OAI211_X1 g621(.A(KEYINPUT54), .B(new_n640), .C1(new_n629), .C2(new_n631), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT54), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n629), .A2(new_n824), .A3(new_n631), .ZN(new_n825));
  AND3_X1   g624(.A1(new_n823), .A2(new_n638), .A3(new_n825), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n826), .A2(KEYINPUT55), .ZN(new_n827));
  INV_X1    g626(.A(new_n827), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n823), .A2(KEYINPUT55), .A3(new_n638), .A4(new_n825), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(new_n642), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(KEYINPUT116), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT116), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n829), .A2(new_n832), .A3(new_n642), .ZN(new_n833));
  AND3_X1   g632(.A1(new_n828), .A2(new_n831), .A3(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n696), .A2(new_n834), .A3(new_n698), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n520), .B1(new_n529), .B2(new_n519), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT117), .ZN(new_n837));
  NOR3_X1   g636(.A1(new_n534), .A2(new_n837), .A3(new_n535), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n837), .B1(new_n534), .B2(new_n535), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(new_n546), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n552), .A2(new_n842), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n843), .A2(new_n644), .ZN(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n620), .B1(new_n835), .B2(new_n845), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n620), .A2(new_n552), .A3(new_n834), .A4(new_n842), .ZN(new_n847));
  INV_X1    g646(.A(new_n847), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n592), .B1(new_n846), .B2(new_n848), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n621), .A2(new_n644), .A3(new_n699), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n822), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  AND2_X1   g650(.A1(new_n851), .A2(new_n484), .ZN(new_n852));
  AOI21_X1  g651(.A(G113gat), .B1(new_n852), .B2(new_n700), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n449), .A2(new_n661), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n851), .A2(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(G113gat), .ZN(new_n856));
  NOR3_X1   g655(.A1(new_n855), .A2(new_n856), .A3(new_n555), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n853), .A2(new_n857), .ZN(G1340gat));
  AOI21_X1  g657(.A(G120gat), .B1(new_n852), .B2(new_n643), .ZN(new_n859));
  INV_X1    g658(.A(G120gat), .ZN(new_n860));
  NOR3_X1   g659(.A1(new_n855), .A2(new_n860), .A3(new_n644), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n859), .A2(new_n861), .ZN(G1341gat));
  INV_X1    g661(.A(G127gat), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n852), .A2(new_n863), .A3(new_n591), .ZN(new_n864));
  OAI21_X1  g663(.A(G127gat), .B1(new_n855), .B2(new_n592), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(G1342gat));
  AND2_X1   g665(.A1(new_n851), .A2(new_n620), .ZN(new_n867));
  INV_X1    g666(.A(G134gat), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n867), .A2(new_n868), .A3(new_n484), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT56), .ZN(new_n870));
  AND2_X1   g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n869), .A2(new_n870), .ZN(new_n872));
  AND2_X1   g671(.A1(new_n867), .A2(new_n854), .ZN(new_n873));
  OAI22_X1  g672(.A1(new_n871), .A2(new_n872), .B1(new_n868), .B2(new_n873), .ZN(G1343gat));
  AOI21_X1  g673(.A(new_n445), .B1(new_n849), .B2(new_n850), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT57), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n659), .A2(new_n649), .A3(new_n486), .ZN(new_n878));
  XOR2_X1   g677(.A(new_n878), .B(KEYINPUT118), .Z(new_n879));
  INV_X1    g678(.A(new_n850), .ZN(new_n880));
  AOI211_X1 g679(.A(new_n830), .B(new_n827), .C1(new_n552), .C2(new_n553), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n689), .B1(new_n881), .B2(new_n844), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n591), .B1(new_n882), .B2(new_n847), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n449), .B1(new_n880), .B2(new_n883), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n879), .B1(new_n884), .B2(KEYINPUT57), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n877), .A2(new_n885), .A3(new_n700), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(G141gat), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n278), .A2(new_n445), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n555), .A2(G141gat), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n851), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n887), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n891), .A2(KEYINPUT119), .A3(KEYINPUT58), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT119), .ZN(new_n893));
  AND2_X1   g692(.A1(new_n851), .A2(new_n888), .ZN(new_n894));
  AOI22_X1  g693(.A1(new_n886), .A2(G141gat), .B1(new_n894), .B2(new_n889), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT58), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n893), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  XNOR2_X1  g696(.A(new_n890), .B(KEYINPUT120), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n877), .A2(new_n885), .ZN(new_n899));
  OAI21_X1  g698(.A(G141gat), .B1(new_n899), .B2(new_n555), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n898), .A2(new_n896), .A3(new_n900), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n892), .A2(new_n897), .A3(new_n901), .ZN(G1344gat));
  AND2_X1   g701(.A1(new_n291), .A2(new_n293), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n894), .A2(new_n903), .A3(new_n643), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(KEYINPUT121), .ZN(new_n905));
  OR2_X1    g704(.A1(new_n904), .A2(KEYINPUT121), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n899), .A2(new_n644), .ZN(new_n907));
  NOR3_X1   g706(.A1(new_n907), .A2(KEYINPUT59), .A3(new_n903), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT59), .ZN(new_n909));
  OR2_X1    g708(.A1(new_n875), .A2(new_n876), .ZN(new_n910));
  INV_X1    g709(.A(new_n879), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n645), .A2(new_n554), .ZN(new_n912));
  OAI211_X1 g711(.A(new_n876), .B(new_n449), .C1(new_n912), .C2(new_n883), .ZN(new_n913));
  NAND4_X1  g712(.A1(new_n910), .A2(new_n643), .A3(new_n911), .A4(new_n913), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n909), .B1(new_n914), .B2(G148gat), .ZN(new_n915));
  OAI211_X1 g714(.A(new_n905), .B(new_n906), .C1(new_n908), .C2(new_n915), .ZN(G1345gat));
  OAI21_X1  g715(.A(G155gat), .B1(new_n899), .B2(new_n592), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n894), .A2(new_n284), .A3(new_n591), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(G1346gat));
  OAI21_X1  g718(.A(G162gat), .B1(new_n899), .B2(new_n689), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n894), .A2(new_n285), .A3(new_n620), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(G1347gat));
  NAND2_X1  g721(.A1(new_n849), .A2(new_n850), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n649), .A2(new_n486), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n925), .A2(new_n484), .ZN(new_n926));
  NAND4_X1  g725(.A1(new_n926), .A2(new_n211), .A3(new_n213), .A4(new_n700), .ZN(new_n927));
  XNOR2_X1  g726(.A(new_n924), .B(KEYINPUT122), .ZN(new_n928));
  AND3_X1   g727(.A1(new_n928), .A2(new_n675), .A3(new_n752), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n923), .A2(new_n929), .ZN(new_n930));
  OAI21_X1  g729(.A(G169gat), .B1(new_n930), .B2(new_n555), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n927), .A2(new_n931), .ZN(G1348gat));
  NAND3_X1  g731(.A1(new_n926), .A2(new_n214), .A3(new_n643), .ZN(new_n933));
  OAI21_X1  g732(.A(G176gat), .B1(new_n930), .B2(new_n644), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(new_n934), .ZN(G1349gat));
  NAND4_X1  g734(.A1(new_n925), .A2(new_n233), .A3(new_n484), .A4(new_n591), .ZN(new_n936));
  OAI21_X1  g735(.A(G183gat), .B1(new_n930), .B2(new_n592), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT60), .ZN(new_n938));
  AOI22_X1  g737(.A1(new_n936), .A2(new_n937), .B1(KEYINPUT123), .B2(new_n938), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n938), .A2(KEYINPUT123), .ZN(new_n940));
  XNOR2_X1  g739(.A(new_n939), .B(new_n940), .ZN(G1350gat));
  INV_X1    g740(.A(new_n698), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n697), .B1(new_n552), .B2(new_n553), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n828), .A2(new_n831), .A3(new_n833), .ZN(new_n944));
  NOR3_X1   g743(.A1(new_n942), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n689), .B1(new_n945), .B2(new_n844), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n591), .B1(new_n946), .B2(new_n847), .ZN(new_n947));
  OAI211_X1 g746(.A(new_n620), .B(new_n929), .C1(new_n947), .C2(new_n880), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT61), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n948), .A2(new_n949), .A3(G190gat), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT124), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND4_X1  g751(.A1(new_n948), .A2(KEYINPUT124), .A3(new_n949), .A4(G190gat), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n948), .A2(G190gat), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n954), .A2(KEYINPUT61), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n952), .A2(new_n953), .A3(new_n955), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n926), .A2(new_n234), .A3(new_n620), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT125), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n956), .A2(new_n957), .A3(KEYINPUT125), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n960), .A2(new_n961), .ZN(G1351gat));
  AND2_X1   g761(.A1(new_n925), .A2(new_n888), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n963), .A2(new_n389), .A3(new_n700), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n928), .A2(new_n659), .ZN(new_n965));
  INV_X1    g764(.A(new_n965), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n910), .A2(new_n913), .A3(new_n966), .ZN(new_n967));
  OAI21_X1  g766(.A(KEYINPUT126), .B1(new_n967), .B2(new_n555), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n968), .A2(G197gat), .ZN(new_n969));
  NOR3_X1   g768(.A1(new_n967), .A2(KEYINPUT126), .A3(new_n555), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n964), .B1(new_n969), .B2(new_n970), .ZN(G1352gat));
  AND4_X1   g770(.A1(new_n387), .A2(new_n925), .A3(new_n643), .A4(new_n888), .ZN(new_n972));
  AND2_X1   g771(.A1(new_n972), .A2(KEYINPUT62), .ZN(new_n973));
  NOR2_X1   g772(.A1(new_n972), .A2(KEYINPUT62), .ZN(new_n974));
  AND4_X1   g773(.A1(new_n643), .A2(new_n910), .A3(new_n913), .A4(new_n966), .ZN(new_n975));
  OAI22_X1  g774(.A1(new_n973), .A2(new_n974), .B1(new_n387), .B2(new_n975), .ZN(G1353gat));
  NAND3_X1  g775(.A1(new_n963), .A2(new_n384), .A3(new_n591), .ZN(new_n977));
  NAND4_X1  g776(.A1(new_n910), .A2(new_n591), .A3(new_n913), .A4(new_n966), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n978), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n979));
  INV_X1    g778(.A(new_n979), .ZN(new_n980));
  AOI21_X1  g779(.A(KEYINPUT63), .B1(new_n978), .B2(G211gat), .ZN(new_n981));
  OAI21_X1  g780(.A(new_n977), .B1(new_n980), .B2(new_n981), .ZN(G1354gat));
  OAI21_X1  g781(.A(G218gat), .B1(new_n967), .B2(new_n689), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n963), .A2(new_n385), .A3(new_n620), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n983), .A2(new_n984), .ZN(G1355gat));
endmodule


