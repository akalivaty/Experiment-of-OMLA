

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731;

  XNOR2_X1 U365 ( .A(n406), .B(G101), .ZN(n408) );
  INV_X2 U366 ( .A(G953), .ZN(n710) );
  OR2_X2 U367 ( .A1(n615), .A2(n600), .ZN(n393) );
  XNOR2_X2 U368 ( .A(n508), .B(KEYINPUT33), .ZN(n687) );
  NAND2_X2 U369 ( .A1(n514), .A2(n579), .ZN(n500) );
  XNOR2_X2 U370 ( .A(n457), .B(n456), .ZN(n514) );
  XNOR2_X1 U371 ( .A(n582), .B(n421), .ZN(n571) );
  NOR2_X1 U372 ( .A1(n527), .A2(n526), .ZN(n577) );
  INV_X1 U373 ( .A(G125), .ZN(n400) );
  AND2_X1 U374 ( .A1(n597), .A2(n596), .ZN(n603) );
  NOR2_X1 U375 ( .A1(n376), .A2(n375), .ZN(n566) );
  AND2_X1 U376 ( .A1(n594), .A2(n577), .ZN(n558) );
  NOR2_X1 U377 ( .A1(n570), .A2(n559), .ZN(n557) );
  NAND2_X1 U378 ( .A1(n571), .A2(n426), .ZN(n429) );
  XNOR2_X1 U379 ( .A(n397), .B(KEYINPUT77), .ZN(n396) );
  XNOR2_X1 U380 ( .A(n395), .B(n352), .ZN(n394) );
  XNOR2_X1 U381 ( .A(n577), .B(n576), .ZN(n651) );
  NAND2_X1 U382 ( .A1(n588), .A2(n677), .ZN(n582) );
  XNOR2_X1 U383 ( .A(n629), .B(n632), .ZN(n633) );
  XNOR2_X1 U384 ( .A(n440), .B(n363), .ZN(n527) );
  XOR2_X1 U385 ( .A(KEYINPUT59), .B(n623), .Z(n624) );
  XNOR2_X1 U386 ( .A(n496), .B(n399), .ZN(n716) );
  XNOR2_X1 U387 ( .A(G143), .B(G128), .ZN(n448) );
  NOR2_X2 U388 ( .A1(n389), .A2(n613), .ZN(n353) );
  XNOR2_X1 U389 ( .A(n575), .B(n358), .ZN(n357) );
  INV_X1 U390 ( .A(KEYINPUT47), .ZN(n358) );
  NOR2_X1 U391 ( .A1(n731), .A2(n730), .ZN(n567) );
  XNOR2_X1 U392 ( .A(n437), .B(KEYINPUT10), .ZN(n720) );
  NOR2_X1 U393 ( .A1(n374), .A2(n348), .ZN(n372) );
  XNOR2_X1 U394 ( .A(n567), .B(KEYINPUT46), .ZN(n371) );
  NAND2_X1 U395 ( .A1(n357), .A2(n356), .ZN(n374) );
  INV_X1 U396 ( .A(KEYINPUT48), .ZN(n370) );
  XNOR2_X1 U397 ( .A(n360), .B(n359), .ZN(n530) );
  BUF_X1 U398 ( .A(n604), .Z(n701) );
  NOR2_X1 U399 ( .A1(n681), .A2(n383), .ZN(n382) );
  INV_X1 U400 ( .A(n677), .ZN(n383) );
  XNOR2_X1 U401 ( .A(n588), .B(KEYINPUT38), .ZN(n559) );
  XOR2_X1 U402 ( .A(KEYINPUT68), .B(KEYINPUT8), .Z(n441) );
  XNOR2_X1 U403 ( .A(G119), .B(G128), .ZN(n490) );
  XNOR2_X1 U404 ( .A(G113), .B(G143), .ZN(n432) );
  XNOR2_X1 U405 ( .A(KEYINPUT69), .B(G131), .ZN(n468) );
  XNOR2_X1 U406 ( .A(n431), .B(KEYINPUT97), .ZN(n362) );
  XOR2_X1 U407 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n430) );
  INV_X1 U408 ( .A(KEYINPUT41), .ZN(n378) );
  NAND2_X1 U409 ( .A1(n381), .A2(n678), .ZN(n380) );
  AND2_X1 U410 ( .A1(n382), .A2(KEYINPUT41), .ZN(n381) );
  NOR2_X1 U411 ( .A1(n580), .A2(n579), .ZN(n585) );
  NAND2_X1 U412 ( .A1(n651), .A2(n578), .ZN(n580) );
  INV_X1 U413 ( .A(KEYINPUT108), .ZN(n581) );
  NAND2_X1 U414 ( .A1(n499), .A2(n350), .ZN(n387) );
  XNOR2_X1 U415 ( .A(n439), .B(KEYINPUT13), .ZN(n363) );
  INV_X1 U416 ( .A(G475), .ZN(n439) );
  NOR2_X1 U417 ( .A1(n716), .A2(G902), .ZN(n497) );
  INV_X1 U418 ( .A(n647), .ZN(n356) );
  INV_X1 U419 ( .A(KEYINPUT103), .ZN(n359) );
  NAND2_X1 U420 ( .A1(n678), .A2(n677), .ZN(n682) );
  XNOR2_X1 U421 ( .A(G101), .B(G146), .ZN(n461) );
  XNOR2_X1 U422 ( .A(KEYINPUT4), .B(G137), .ZN(n467) );
  NOR2_X1 U423 ( .A1(G953), .A2(G237), .ZN(n458) );
  INV_X1 U424 ( .A(G146), .ZN(n476) );
  NAND2_X1 U425 ( .A1(G234), .A2(G237), .ZN(n422) );
  XNOR2_X1 U426 ( .A(n361), .B(n370), .ZN(n597) );
  INV_X1 U427 ( .A(n660), .ZN(n595) );
  NAND2_X1 U428 ( .A1(n504), .A2(n392), .ZN(n518) );
  INV_X1 U429 ( .A(n661), .ZN(n392) );
  AND2_X1 U430 ( .A1(n562), .A2(n560), .ZN(n398) );
  NAND2_X1 U431 ( .A1(n668), .A2(n677), .ZN(n395) );
  INV_X1 U432 ( .A(G237), .ZN(n417) );
  NOR2_X1 U433 ( .A1(n562), .A2(n561), .ZN(n578) );
  XOR2_X1 U434 ( .A(KEYINPUT76), .B(G110), .Z(n407) );
  XOR2_X1 U435 ( .A(KEYINPUT9), .B(G122), .Z(n446) );
  XNOR2_X1 U436 ( .A(G116), .B(G107), .ZN(n445) );
  XNOR2_X1 U437 ( .A(KEYINPUT16), .B(G122), .ZN(n414) );
  NAND2_X1 U438 ( .A1(n351), .A2(n345), .ZN(n696) );
  NAND2_X1 U439 ( .A1(n539), .A2(n538), .ZN(n540) );
  INV_X1 U440 ( .A(n720), .ZN(n399) );
  NAND2_X1 U441 ( .A1(n369), .A2(n602), .ZN(n368) );
  XNOR2_X1 U442 ( .A(n362), .B(n430), .ZN(n435) );
  AND2_X1 U443 ( .A1(n379), .A2(n378), .ZN(n375) );
  XNOR2_X1 U444 ( .A(n585), .B(n581), .ZN(n583) );
  XNOR2_X1 U445 ( .A(n390), .B(n512), .ZN(n613) );
  NAND2_X1 U446 ( .A1(n386), .A2(n385), .ZN(n384) );
  NOR2_X1 U447 ( .A1(n499), .A2(n350), .ZN(n385) );
  NOR2_X1 U448 ( .A1(n573), .A2(n572), .ZN(n648) );
  XNOR2_X1 U449 ( .A(n525), .B(n524), .ZN(n654) );
  INV_X1 U450 ( .A(KEYINPUT105), .ZN(n576) );
  XNOR2_X1 U451 ( .A(n355), .B(n354), .ZN(n516) );
  INV_X1 U452 ( .A(KEYINPUT87), .ZN(n354) );
  INV_X1 U453 ( .A(n504), .ZN(n662) );
  AND2_X1 U454 ( .A1(n380), .A2(n349), .ZN(n345) );
  AND2_X1 U455 ( .A1(n388), .A2(n387), .ZN(n346) );
  XOR2_X1 U456 ( .A(G104), .B(G122), .Z(n347) );
  AND2_X1 U457 ( .A1(n373), .A2(n504), .ZN(n348) );
  OR2_X1 U458 ( .A1(n382), .A2(KEYINPUT41), .ZN(n349) );
  XOR2_X1 U459 ( .A(KEYINPUT65), .B(KEYINPUT32), .Z(n350) );
  OR2_X1 U460 ( .A1(n678), .A2(KEYINPUT41), .ZN(n351) );
  XNOR2_X1 U461 ( .A(KEYINPUT30), .B(KEYINPUT107), .ZN(n352) );
  NAND2_X1 U462 ( .A1(n346), .A2(n384), .ZN(n622) );
  XNOR2_X1 U463 ( .A(n353), .B(KEYINPUT44), .ZN(n531) );
  NAND2_X1 U464 ( .A1(n514), .A2(n513), .ZN(n355) );
  NOR2_X1 U465 ( .A1(n620), .A2(n529), .ZN(n360) );
  NAND2_X1 U466 ( .A1(n622), .A2(n644), .ZN(n389) );
  XNOR2_X1 U467 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U468 ( .A(n495), .B(n494), .ZN(n496) );
  NAND2_X1 U469 ( .A1(n372), .A2(n371), .ZN(n361) );
  INV_X1 U470 ( .A(n364), .ZN(n705) );
  AND2_X4 U471 ( .A1(n367), .A2(n364), .ZN(n715) );
  NAND2_X1 U472 ( .A1(n701), .A2(n365), .ZN(n364) );
  XNOR2_X1 U473 ( .A(n366), .B(KEYINPUT85), .ZN(n365) );
  NAND2_X1 U474 ( .A1(n603), .A2(KEYINPUT2), .ZN(n366) );
  XNOR2_X2 U475 ( .A(n368), .B(KEYINPUT64), .ZN(n367) );
  NAND2_X1 U476 ( .A1(n599), .A2(n604), .ZN(n369) );
  XNOR2_X1 U477 ( .A(n584), .B(KEYINPUT36), .ZN(n373) );
  NAND2_X1 U478 ( .A1(n377), .A2(n380), .ZN(n376) );
  INV_X1 U479 ( .A(n573), .ZN(n377) );
  NAND2_X1 U480 ( .A1(n678), .A2(n382), .ZN(n379) );
  NAND2_X1 U481 ( .A1(n396), .A2(n394), .ZN(n570) );
  NAND2_X1 U482 ( .A1(n398), .A2(n564), .ZN(n397) );
  INV_X1 U483 ( .A(n500), .ZN(n386) );
  XNOR2_X1 U484 ( .A(n510), .B(n509), .ZN(n391) );
  NAND2_X1 U485 ( .A1(n500), .A2(n350), .ZN(n388) );
  NAND2_X1 U486 ( .A1(n391), .A2(n568), .ZN(n390) );
  XNOR2_X2 U487 ( .A(n564), .B(n485), .ZN(n504) );
  XNOR2_X2 U488 ( .A(n484), .B(G469), .ZN(n564) );
  XNOR2_X2 U489 ( .A(n393), .B(n419), .ZN(n588) );
  XNOR2_X1 U490 ( .A(n416), .B(n542), .ZN(n615) );
  XNOR2_X2 U491 ( .A(n473), .B(G472), .ZN(n668) );
  XNOR2_X2 U492 ( .A(n400), .B(G146), .ZN(n436) );
  NOR2_X1 U493 ( .A1(n729), .A2(n595), .ZN(n596) );
  XNOR2_X1 U494 ( .A(n603), .B(KEYINPUT83), .ZN(n700) );
  NOR2_X1 U495 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U496 ( .A(n535), .B(n534), .ZN(n539) );
  INV_X1 U497 ( .A(KEYINPUT39), .ZN(n556) );
  INV_X1 U498 ( .A(KEYINPUT126), .ZN(n546) );
  XNOR2_X1 U499 ( .A(n557), .B(n556), .ZN(n594) );
  INV_X1 U500 ( .A(KEYINPUT63), .ZN(n611) );
  XNOR2_X1 U501 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U502 ( .A(n549), .B(n548), .ZN(G69) );
  XOR2_X1 U503 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n403) );
  NAND2_X1 U504 ( .A1(G224), .A2(n710), .ZN(n401) );
  XNOR2_X1 U505 ( .A(n401), .B(KEYINPUT4), .ZN(n402) );
  XNOR2_X1 U506 ( .A(n403), .B(n402), .ZN(n405) );
  XNOR2_X1 U507 ( .A(n436), .B(n448), .ZN(n404) );
  XNOR2_X1 U508 ( .A(n405), .B(n404), .ZN(n409) );
  XNOR2_X2 U509 ( .A(G107), .B(G104), .ZN(n406) );
  XNOR2_X2 U510 ( .A(n408), .B(n407), .ZN(n541) );
  XNOR2_X2 U511 ( .A(n541), .B(KEYINPUT72), .ZN(n481) );
  XNOR2_X1 U512 ( .A(n481), .B(n409), .ZN(n416) );
  XNOR2_X1 U513 ( .A(G119), .B(G116), .ZN(n411) );
  XNOR2_X1 U514 ( .A(G113), .B(KEYINPUT71), .ZN(n410) );
  XNOR2_X1 U515 ( .A(n411), .B(n410), .ZN(n413) );
  XNOR2_X1 U516 ( .A(KEYINPUT90), .B(KEYINPUT3), .ZN(n412) );
  XNOR2_X1 U517 ( .A(n413), .B(n412), .ZN(n465) );
  XNOR2_X1 U518 ( .A(n414), .B(KEYINPUT74), .ZN(n415) );
  XNOR2_X1 U519 ( .A(n465), .B(n415), .ZN(n542) );
  XNOR2_X1 U520 ( .A(G902), .B(KEYINPUT15), .ZN(n598) );
  INV_X1 U521 ( .A(n598), .ZN(n600) );
  INV_X1 U522 ( .A(G902), .ZN(n472) );
  NAND2_X1 U523 ( .A1(n472), .A2(n417), .ZN(n420) );
  NAND2_X1 U524 ( .A1(n420), .A2(G210), .ZN(n418) );
  XNOR2_X1 U525 ( .A(n418), .B(KEYINPUT91), .ZN(n419) );
  NAND2_X1 U526 ( .A1(n420), .A2(G214), .ZN(n677) );
  XNOR2_X1 U527 ( .A(KEYINPUT78), .B(KEYINPUT19), .ZN(n421) );
  XNOR2_X1 U528 ( .A(n422), .B(KEYINPUT14), .ZN(n423) );
  NAND2_X1 U529 ( .A1(G952), .A2(n423), .ZN(n693) );
  NOR2_X1 U530 ( .A1(G953), .A2(n693), .ZN(n553) );
  OR2_X1 U531 ( .A1(n710), .A2(G898), .ZN(n544) );
  NAND2_X1 U532 ( .A1(G902), .A2(n423), .ZN(n550) );
  NOR2_X1 U533 ( .A1(n544), .A2(n550), .ZN(n424) );
  OR2_X1 U534 ( .A1(n553), .A2(n424), .ZN(n425) );
  XNOR2_X1 U535 ( .A(n425), .B(KEYINPUT92), .ZN(n426) );
  INV_X1 U536 ( .A(KEYINPUT88), .ZN(n427) );
  XNOR2_X1 U537 ( .A(n427), .B(KEYINPUT0), .ZN(n428) );
  XNOR2_X2 U538 ( .A(n429), .B(n428), .ZN(n523) );
  NAND2_X1 U539 ( .A1(G214), .A2(n458), .ZN(n431) );
  XNOR2_X1 U540 ( .A(n347), .B(n432), .ZN(n433) );
  XNOR2_X1 U541 ( .A(n433), .B(n468), .ZN(n434) );
  XNOR2_X1 U542 ( .A(n435), .B(n434), .ZN(n438) );
  XNOR2_X1 U543 ( .A(n436), .B(G140), .ZN(n437) );
  XNOR2_X1 U544 ( .A(n438), .B(n720), .ZN(n623) );
  NOR2_X1 U545 ( .A1(G902), .A2(n623), .ZN(n440) );
  XOR2_X1 U546 ( .A(KEYINPUT98), .B(KEYINPUT7), .Z(n444) );
  NAND2_X1 U547 ( .A1(G234), .A2(n710), .ZN(n442) );
  XNOR2_X1 U548 ( .A(n442), .B(n441), .ZN(n489) );
  NAND2_X1 U549 ( .A1(G217), .A2(n489), .ZN(n443) );
  XNOR2_X1 U550 ( .A(n444), .B(n443), .ZN(n451) );
  XNOR2_X1 U551 ( .A(n446), .B(n445), .ZN(n449) );
  INV_X1 U552 ( .A(G134), .ZN(n447) );
  XNOR2_X1 U553 ( .A(n448), .B(n447), .ZN(n470) );
  XNOR2_X1 U554 ( .A(n449), .B(n470), .ZN(n450) );
  XNOR2_X1 U555 ( .A(n451), .B(n450), .ZN(n713) );
  NAND2_X1 U556 ( .A1(n713), .A2(n472), .ZN(n452) );
  XNOR2_X1 U557 ( .A(n452), .B(G478), .ZN(n526) );
  INV_X1 U558 ( .A(n526), .ZN(n511) );
  NAND2_X1 U559 ( .A1(n527), .A2(n511), .ZN(n681) );
  NAND2_X1 U560 ( .A1(n598), .A2(G234), .ZN(n453) );
  XNOR2_X1 U561 ( .A(n453), .B(KEYINPUT20), .ZN(n486) );
  AND2_X1 U562 ( .A1(n486), .A2(G221), .ZN(n454) );
  XNOR2_X1 U563 ( .A(n454), .B(KEYINPUT21), .ZN(n665) );
  INV_X1 U564 ( .A(n665), .ZN(n555) );
  NOR2_X1 U565 ( .A1(n681), .A2(n555), .ZN(n455) );
  NAND2_X1 U566 ( .A1(n523), .A2(n455), .ZN(n457) );
  XNOR2_X1 U567 ( .A(KEYINPUT73), .B(KEYINPUT22), .ZN(n456) );
  XOR2_X1 U568 ( .A(KEYINPUT95), .B(KEYINPUT5), .Z(n460) );
  NAND2_X1 U569 ( .A1(n458), .A2(G210), .ZN(n459) );
  XNOR2_X1 U570 ( .A(n460), .B(n459), .ZN(n464) );
  XOR2_X1 U571 ( .A(KEYINPUT75), .B(KEYINPUT94), .Z(n462) );
  XNOR2_X1 U572 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U573 ( .A(n464), .B(n463), .ZN(n466) );
  XNOR2_X1 U574 ( .A(n466), .B(n465), .ZN(n471) );
  XNOR2_X1 U575 ( .A(n468), .B(n467), .ZN(n469) );
  XNOR2_X1 U576 ( .A(n470), .B(n469), .ZN(n482) );
  XNOR2_X1 U577 ( .A(n471), .B(n482), .ZN(n606) );
  NAND2_X1 U578 ( .A1(n606), .A2(n472), .ZN(n473) );
  INV_X1 U579 ( .A(KEYINPUT101), .ZN(n474) );
  XNOR2_X1 U580 ( .A(n474), .B(KEYINPUT6), .ZN(n475) );
  XNOR2_X1 U581 ( .A(n668), .B(n475), .ZN(n579) );
  NAND2_X1 U582 ( .A1(n710), .A2(G227), .ZN(n477) );
  XNOR2_X1 U583 ( .A(n477), .B(n476), .ZN(n479) );
  XNOR2_X1 U584 ( .A(KEYINPUT80), .B(G140), .ZN(n478) );
  XNOR2_X1 U585 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U586 ( .A(n481), .B(n480), .ZN(n483) );
  XNOR2_X1 U587 ( .A(n482), .B(KEYINPUT93), .ZN(n721) );
  XNOR2_X1 U588 ( .A(n483), .B(n721), .ZN(n628) );
  OR2_X2 U589 ( .A1(n628), .A2(G902), .ZN(n484) );
  XNOR2_X1 U590 ( .A(KEYINPUT66), .B(KEYINPUT1), .ZN(n485) );
  XOR2_X1 U591 ( .A(KEYINPUT25), .B(KEYINPUT79), .Z(n488) );
  NAND2_X1 U592 ( .A1(G217), .A2(n486), .ZN(n487) );
  XNOR2_X1 U593 ( .A(n488), .B(n487), .ZN(n498) );
  NAND2_X1 U594 ( .A1(n489), .A2(G221), .ZN(n495) );
  XOR2_X1 U595 ( .A(G110), .B(G137), .Z(n491) );
  XNOR2_X1 U596 ( .A(n491), .B(n490), .ZN(n493) );
  XOR2_X1 U597 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n492) );
  XNOR2_X2 U598 ( .A(n498), .B(n497), .ZN(n562) );
  XNOR2_X1 U599 ( .A(n562), .B(KEYINPUT102), .ZN(n664) );
  INV_X1 U600 ( .A(n664), .ZN(n515) );
  NAND2_X1 U601 ( .A1(n504), .A2(n515), .ZN(n499) );
  INV_X1 U602 ( .A(n668), .ZN(n517) );
  INV_X1 U603 ( .A(n562), .ZN(n501) );
  NAND2_X1 U604 ( .A1(n517), .A2(n501), .ZN(n502) );
  NOR2_X1 U605 ( .A1(n504), .A2(n502), .ZN(n503) );
  NAND2_X1 U606 ( .A1(n514), .A2(n503), .ZN(n644) );
  NAND2_X1 U607 ( .A1(n665), .A2(n562), .ZN(n661) );
  INV_X1 U608 ( .A(KEYINPUT104), .ZN(n505) );
  XNOR2_X1 U609 ( .A(n518), .B(n505), .ZN(n507) );
  INV_X1 U610 ( .A(n579), .ZN(n506) );
  NAND2_X1 U611 ( .A1(n507), .A2(n506), .ZN(n508) );
  NAND2_X1 U612 ( .A1(n687), .A2(n523), .ZN(n510) );
  XNOR2_X1 U613 ( .A(KEYINPUT81), .B(KEYINPUT34), .ZN(n509) );
  NOR2_X1 U614 ( .A1(n527), .A2(n511), .ZN(n568) );
  XNOR2_X1 U615 ( .A(KEYINPUT86), .B(KEYINPUT35), .ZN(n512) );
  AND2_X1 U616 ( .A1(n579), .A2(n662), .ZN(n513) );
  NOR2_X1 U617 ( .A1(n516), .A2(n515), .ZN(n620) );
  XOR2_X1 U618 ( .A(KEYINPUT31), .B(KEYINPUT96), .Z(n520) );
  NOR2_X1 U619 ( .A1(n518), .A2(n517), .ZN(n671) );
  NAND2_X1 U620 ( .A1(n523), .A2(n671), .ZN(n519) );
  XOR2_X1 U621 ( .A(n520), .B(n519), .Z(n653) );
  NOR2_X1 U622 ( .A1(n668), .A2(n661), .ZN(n521) );
  AND2_X1 U623 ( .A1(n564), .A2(n521), .ZN(n522) );
  AND2_X1 U624 ( .A1(n523), .A2(n522), .ZN(n639) );
  NOR2_X1 U625 ( .A1(n653), .A2(n639), .ZN(n528) );
  INV_X1 U626 ( .A(KEYINPUT99), .ZN(n525) );
  AND2_X1 U627 ( .A1(n527), .A2(n526), .ZN(n524) );
  XNOR2_X1 U628 ( .A(KEYINPUT100), .B(n654), .ZN(n593) );
  NOR2_X1 U629 ( .A1(n593), .A2(n577), .ZN(n683) );
  NOR2_X1 U630 ( .A1(n528), .A2(n683), .ZN(n529) );
  NAND2_X1 U631 ( .A1(n531), .A2(n530), .ZN(n533) );
  XNOR2_X1 U632 ( .A(KEYINPUT84), .B(KEYINPUT45), .ZN(n532) );
  XNOR2_X2 U633 ( .A(n533), .B(n532), .ZN(n604) );
  NAND2_X1 U634 ( .A1(n701), .A2(n710), .ZN(n535) );
  INV_X1 U635 ( .A(KEYINPUT123), .ZN(n534) );
  NAND2_X1 U636 ( .A1(G953), .A2(G224), .ZN(n536) );
  XNOR2_X1 U637 ( .A(KEYINPUT61), .B(n536), .ZN(n537) );
  NAND2_X1 U638 ( .A1(n537), .A2(G898), .ZN(n538) );
  XNOR2_X1 U639 ( .A(n540), .B(KEYINPUT124), .ZN(n549) );
  XNOR2_X1 U640 ( .A(n541), .B(KEYINPUT125), .ZN(n543) );
  XNOR2_X1 U641 ( .A(n543), .B(n542), .ZN(n545) );
  NAND2_X1 U642 ( .A1(n545), .A2(n544), .ZN(n547) );
  OR2_X1 U643 ( .A1(n710), .A2(n550), .ZN(n551) );
  NOR2_X1 U644 ( .A1(n551), .A2(G900), .ZN(n552) );
  NOR2_X1 U645 ( .A1(n553), .A2(n552), .ZN(n554) );
  NOR2_X1 U646 ( .A1(n555), .A2(n554), .ZN(n560) );
  XNOR2_X1 U647 ( .A(n558), .B(KEYINPUT40), .ZN(n731) );
  INV_X1 U648 ( .A(n559), .ZN(n678) );
  XOR2_X1 U649 ( .A(n560), .B(KEYINPUT70), .Z(n561) );
  AND2_X1 U650 ( .A1(n668), .A2(n578), .ZN(n563) );
  XNOR2_X1 U651 ( .A(KEYINPUT28), .B(n563), .ZN(n565) );
  NAND2_X1 U652 ( .A1(n565), .A2(n564), .ZN(n573) );
  XNOR2_X1 U653 ( .A(n566), .B(KEYINPUT42), .ZN(n730) );
  NAND2_X1 U654 ( .A1(n568), .A2(n588), .ZN(n569) );
  NOR2_X1 U655 ( .A1(n570), .A2(n569), .ZN(n647) );
  INV_X1 U656 ( .A(n683), .ZN(n574) );
  INV_X1 U657 ( .A(n571), .ZN(n572) );
  NAND2_X1 U658 ( .A1(n574), .A2(n648), .ZN(n575) );
  AND2_X1 U659 ( .A1(n585), .A2(n677), .ZN(n586) );
  NAND2_X1 U660 ( .A1(n586), .A2(n662), .ZN(n587) );
  XNOR2_X1 U661 ( .A(n587), .B(KEYINPUT43), .ZN(n590) );
  INV_X1 U662 ( .A(n588), .ZN(n589) );
  NAND2_X1 U663 ( .A1(n590), .A2(n589), .ZN(n592) );
  INV_X1 U664 ( .A(KEYINPUT106), .ZN(n591) );
  XNOR2_X1 U665 ( .A(n592), .B(n591), .ZN(n729) );
  NAND2_X1 U666 ( .A1(n594), .A2(n593), .ZN(n660) );
  NOR2_X1 U667 ( .A1(n700), .A2(n598), .ZN(n599) );
  NAND2_X1 U668 ( .A1(n600), .A2(KEYINPUT2), .ZN(n601) );
  XOR2_X1 U669 ( .A(KEYINPUT67), .B(n601), .Z(n602) );
  NAND2_X1 U670 ( .A1(n715), .A2(G472), .ZN(n608) );
  XNOR2_X1 U671 ( .A(KEYINPUT89), .B(KEYINPUT62), .ZN(n605) );
  XNOR2_X1 U672 ( .A(n606), .B(n605), .ZN(n607) );
  XNOR2_X1 U673 ( .A(n608), .B(n607), .ZN(n610) );
  INV_X1 U674 ( .A(G952), .ZN(n609) );
  AND2_X1 U675 ( .A1(n609), .A2(G953), .ZN(n719) );
  NOR2_X2 U676 ( .A1(n610), .A2(n719), .ZN(n612) );
  XNOR2_X1 U677 ( .A(n612), .B(n611), .ZN(G57) );
  XOR2_X1 U678 ( .A(n613), .B(G122), .Z(G24) );
  NAND2_X1 U679 ( .A1(n715), .A2(G210), .ZN(n617) );
  XOR2_X1 U680 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n614) );
  XNOR2_X1 U681 ( .A(n615), .B(n614), .ZN(n616) );
  XNOR2_X1 U682 ( .A(n617), .B(n616), .ZN(n618) );
  NOR2_X2 U683 ( .A1(n618), .A2(n719), .ZN(n619) );
  XNOR2_X1 U684 ( .A(n619), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U685 ( .A(G101), .B(KEYINPUT109), .ZN(n621) );
  XNOR2_X1 U686 ( .A(n620), .B(n621), .ZN(G3) );
  XNOR2_X1 U687 ( .A(n622), .B(G119), .ZN(G21) );
  NAND2_X1 U688 ( .A1(n715), .A2(G475), .ZN(n625) );
  XNOR2_X1 U689 ( .A(n625), .B(n624), .ZN(n626) );
  NOR2_X2 U690 ( .A1(n626), .A2(n719), .ZN(n627) );
  XNOR2_X1 U691 ( .A(n627), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U692 ( .A1(n715), .A2(G469), .ZN(n634) );
  BUF_X1 U693 ( .A(n628), .Z(n629) );
  XNOR2_X1 U694 ( .A(KEYINPUT121), .B(KEYINPUT57), .ZN(n631) );
  XNOR2_X1 U695 ( .A(KEYINPUT58), .B(KEYINPUT120), .ZN(n630) );
  XNOR2_X1 U696 ( .A(n631), .B(n630), .ZN(n632) );
  XNOR2_X1 U697 ( .A(n634), .B(n633), .ZN(n635) );
  NOR2_X2 U698 ( .A1(n635), .A2(n719), .ZN(n636) );
  XNOR2_X1 U699 ( .A(n636), .B(KEYINPUT122), .ZN(G54) );
  NAND2_X1 U700 ( .A1(n639), .A2(n651), .ZN(n637) );
  XNOR2_X1 U701 ( .A(n637), .B(KEYINPUT110), .ZN(n638) );
  XNOR2_X1 U702 ( .A(G104), .B(n638), .ZN(G6) );
  XOR2_X1 U703 ( .A(KEYINPUT111), .B(KEYINPUT26), .Z(n641) );
  NAND2_X1 U704 ( .A1(n639), .A2(n654), .ZN(n640) );
  XNOR2_X1 U705 ( .A(n641), .B(n640), .ZN(n643) );
  XOR2_X1 U706 ( .A(G107), .B(KEYINPUT27), .Z(n642) );
  XNOR2_X1 U707 ( .A(n643), .B(n642), .ZN(G9) );
  XNOR2_X1 U708 ( .A(G110), .B(n644), .ZN(G12) );
  XOR2_X1 U709 ( .A(G128), .B(KEYINPUT29), .Z(n646) );
  NAND2_X1 U710 ( .A1(n648), .A2(n654), .ZN(n645) );
  XNOR2_X1 U711 ( .A(n646), .B(n645), .ZN(G30) );
  XOR2_X1 U712 ( .A(G143), .B(n647), .Z(G45) );
  NAND2_X1 U713 ( .A1(n648), .A2(n651), .ZN(n649) );
  XNOR2_X1 U714 ( .A(n649), .B(KEYINPUT112), .ZN(n650) );
  XNOR2_X1 U715 ( .A(G146), .B(n650), .ZN(G48) );
  NAND2_X1 U716 ( .A1(n653), .A2(n651), .ZN(n652) );
  XNOR2_X1 U717 ( .A(n652), .B(G113), .ZN(G15) );
  XOR2_X1 U718 ( .A(G116), .B(KEYINPUT113), .Z(n656) );
  NAND2_X1 U719 ( .A1(n654), .A2(n653), .ZN(n655) );
  XNOR2_X1 U720 ( .A(n656), .B(n655), .ZN(G18) );
  XNOR2_X1 U721 ( .A(n348), .B(KEYINPUT114), .ZN(n657) );
  XNOR2_X1 U722 ( .A(n657), .B(KEYINPUT37), .ZN(n658) );
  XNOR2_X1 U723 ( .A(G125), .B(n658), .ZN(G27) );
  XOR2_X1 U724 ( .A(G134), .B(KEYINPUT115), .Z(n659) );
  XNOR2_X1 U725 ( .A(n660), .B(n659), .ZN(G36) );
  INV_X1 U726 ( .A(n696), .ZN(n676) );
  NAND2_X1 U727 ( .A1(n662), .A2(n661), .ZN(n663) );
  XNOR2_X1 U728 ( .A(n663), .B(KEYINPUT50), .ZN(n670) );
  NOR2_X1 U729 ( .A1(n665), .A2(n664), .ZN(n666) );
  XOR2_X1 U730 ( .A(KEYINPUT49), .B(n666), .Z(n667) );
  NOR2_X1 U731 ( .A1(n668), .A2(n667), .ZN(n669) );
  NAND2_X1 U732 ( .A1(n670), .A2(n669), .ZN(n673) );
  INV_X1 U733 ( .A(n671), .ZN(n672) );
  NAND2_X1 U734 ( .A1(n673), .A2(n672), .ZN(n674) );
  XOR2_X1 U735 ( .A(KEYINPUT51), .B(n674), .Z(n675) );
  NAND2_X1 U736 ( .A1(n676), .A2(n675), .ZN(n690) );
  NOR2_X1 U737 ( .A1(n678), .A2(n677), .ZN(n679) );
  XNOR2_X1 U738 ( .A(n679), .B(KEYINPUT116), .ZN(n680) );
  NOR2_X1 U739 ( .A1(n681), .A2(n680), .ZN(n685) );
  NOR2_X1 U740 ( .A1(n683), .A2(n682), .ZN(n684) );
  NOR2_X1 U741 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U742 ( .A(n686), .B(KEYINPUT117), .ZN(n688) );
  NAND2_X1 U743 ( .A1(n688), .A2(n687), .ZN(n689) );
  NAND2_X1 U744 ( .A1(n690), .A2(n689), .ZN(n692) );
  XOR2_X1 U745 ( .A(KEYINPUT52), .B(KEYINPUT118), .Z(n691) );
  XNOR2_X1 U746 ( .A(n692), .B(n691), .ZN(n694) );
  NOR2_X1 U747 ( .A1(n694), .A2(n693), .ZN(n698) );
  INV_X1 U748 ( .A(n687), .ZN(n695) );
  NOR2_X1 U749 ( .A1(n696), .A2(n695), .ZN(n697) );
  NOR2_X1 U750 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U751 ( .A(n699), .B(KEYINPUT119), .ZN(n708) );
  INV_X1 U752 ( .A(n700), .ZN(n702) );
  NAND2_X1 U753 ( .A1(n702), .A2(n701), .ZN(n704) );
  XOR2_X1 U754 ( .A(KEYINPUT2), .B(KEYINPUT82), .Z(n703) );
  AND2_X1 U755 ( .A1(n704), .A2(n703), .ZN(n706) );
  NOR2_X1 U756 ( .A1(n706), .A2(n705), .ZN(n707) );
  NOR2_X1 U757 ( .A1(n708), .A2(n707), .ZN(n709) );
  NAND2_X1 U758 ( .A1(n710), .A2(n709), .ZN(n711) );
  XOR2_X1 U759 ( .A(KEYINPUT53), .B(n711), .Z(G75) );
  NAND2_X1 U760 ( .A1(n715), .A2(G478), .ZN(n712) );
  XOR2_X1 U761 ( .A(n713), .B(n712), .Z(n714) );
  NOR2_X1 U762 ( .A1(n719), .A2(n714), .ZN(G63) );
  NAND2_X1 U763 ( .A1(n715), .A2(G217), .ZN(n717) );
  XNOR2_X1 U764 ( .A(n717), .B(n716), .ZN(n718) );
  NOR2_X1 U765 ( .A1(n719), .A2(n718), .ZN(G66) );
  XNOR2_X1 U766 ( .A(n721), .B(n720), .ZN(n724) );
  XNOR2_X1 U767 ( .A(n700), .B(n724), .ZN(n722) );
  NOR2_X1 U768 ( .A1(G953), .A2(n722), .ZN(n723) );
  XNOR2_X1 U769 ( .A(n723), .B(KEYINPUT127), .ZN(n728) );
  XOR2_X1 U770 ( .A(G227), .B(n724), .Z(n725) );
  NAND2_X1 U771 ( .A1(n725), .A2(G900), .ZN(n726) );
  NAND2_X1 U772 ( .A1(n726), .A2(G953), .ZN(n727) );
  NAND2_X1 U773 ( .A1(n728), .A2(n727), .ZN(G72) );
  XOR2_X1 U774 ( .A(G140), .B(n729), .Z(G42) );
  XOR2_X1 U775 ( .A(G137), .B(n730), .Z(G39) );
  XOR2_X1 U776 ( .A(n731), .B(G131), .Z(G33) );
endmodule

