//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 1 1 0 0 1 1 1 0 1 0 1 0 0 0 1 1 1 1 0 0 0 1 1 1 1 1 0 1 1 1 0 1 1 1 1 0 0 0 1 0 0 1 0 0 1 0 0 0 0 0 1 0 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:44 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n594, new_n595,
    new_n597, new_n598, new_n599, new_n600, new_n601, new_n602, new_n603,
    new_n604, new_n605, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n630, new_n631, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n640, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n689,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n862, new_n863,
    new_n864, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G143), .ZN(new_n189));
  INV_X1    g003(.A(G143), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G146), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT1), .ZN(new_n192));
  NAND4_X1  g006(.A1(new_n189), .A2(new_n191), .A3(new_n192), .A4(G128), .ZN(new_n193));
  INV_X1    g007(.A(G128), .ZN(new_n194));
  AOI21_X1  g008(.A(new_n194), .B1(new_n189), .B2(KEYINPUT1), .ZN(new_n195));
  XNOR2_X1  g009(.A(G143), .B(G146), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n193), .B1(new_n195), .B2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT11), .ZN(new_n198));
  INV_X1    g012(.A(G134), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n198), .B1(new_n199), .B2(G137), .ZN(new_n200));
  INV_X1    g014(.A(G137), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n201), .A2(KEYINPUT11), .A3(G134), .ZN(new_n202));
  INV_X1    g016(.A(G131), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n199), .A2(G137), .ZN(new_n204));
  NAND4_X1  g018(.A1(new_n200), .A2(new_n202), .A3(new_n203), .A4(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(new_n204), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n199), .A2(G137), .ZN(new_n207));
  OAI21_X1  g021(.A(G131), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n197), .A2(new_n205), .A3(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(KEYINPUT64), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT30), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n200), .A2(new_n204), .A3(new_n202), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G131), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(new_n205), .ZN(new_n214));
  AND2_X1   g028(.A1(KEYINPUT0), .A2(G128), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n189), .A2(new_n191), .A3(new_n215), .ZN(new_n216));
  XNOR2_X1  g030(.A(KEYINPUT0), .B(G128), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n216), .B1(new_n196), .B2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n214), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT64), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n197), .A2(new_n221), .A3(new_n205), .A4(new_n208), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n210), .A2(new_n211), .A3(new_n220), .A4(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT65), .ZN(new_n224));
  AND3_X1   g038(.A1(new_n214), .A2(new_n224), .A3(new_n219), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n224), .B1(new_n214), .B2(new_n219), .ZN(new_n226));
  INV_X1    g040(.A(new_n209), .ZN(new_n227));
  NOR3_X1   g041(.A1(new_n225), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n223), .B1(new_n228), .B2(new_n211), .ZN(new_n229));
  XNOR2_X1  g043(.A(G116), .B(G119), .ZN(new_n230));
  XNOR2_X1  g044(.A(KEYINPUT2), .B(G113), .ZN(new_n231));
  XNOR2_X1  g045(.A(new_n230), .B(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n229), .A2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT31), .ZN(new_n235));
  AND2_X1   g049(.A1(new_n209), .A2(new_n232), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n220), .A2(KEYINPUT65), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n214), .A2(new_n224), .A3(new_n219), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n236), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT66), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n225), .A2(new_n226), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n242), .A2(KEYINPUT66), .A3(new_n236), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(G237), .ZN(new_n245));
  INV_X1    g059(.A(G953), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n245), .A2(new_n246), .A3(G210), .ZN(new_n247));
  XNOR2_X1  g061(.A(new_n247), .B(G101), .ZN(new_n248));
  XNOR2_X1  g062(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n249));
  XNOR2_X1  g063(.A(new_n248), .B(new_n249), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n234), .A2(new_n235), .A3(new_n244), .A4(new_n250), .ZN(new_n251));
  AOI21_X1  g065(.A(KEYINPUT28), .B1(new_n236), .B2(new_n220), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n210), .A2(new_n220), .A3(new_n222), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(new_n233), .ZN(new_n254));
  AOI21_X1  g068(.A(KEYINPUT66), .B1(new_n242), .B2(new_n236), .ZN(new_n255));
  AND4_X1   g069(.A1(KEYINPUT66), .A2(new_n236), .A3(new_n237), .A4(new_n238), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n254), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n252), .B1(new_n257), .B2(KEYINPUT28), .ZN(new_n258));
  XNOR2_X1  g072(.A(new_n250), .B(KEYINPUT68), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n251), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n234), .A2(new_n244), .A3(new_n250), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(KEYINPUT31), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT67), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n261), .A2(KEYINPUT67), .A3(KEYINPUT31), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n260), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NOR2_X1   g080(.A1(G472), .A2(G902), .ZN(new_n267));
  XOR2_X1   g081(.A(new_n267), .B(KEYINPUT69), .Z(new_n268));
  OAI21_X1  g082(.A(new_n187), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT71), .ZN(new_n270));
  INV_X1    g084(.A(new_n268), .ZN(new_n271));
  AND3_X1   g085(.A1(new_n261), .A2(KEYINPUT67), .A3(KEYINPUT31), .ZN(new_n272));
  AOI21_X1  g086(.A(KEYINPUT67), .B1(new_n261), .B2(KEYINPUT31), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  OAI211_X1 g088(.A(KEYINPUT32), .B(new_n271), .C1(new_n274), .C2(new_n260), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n269), .A2(new_n270), .A3(new_n275), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n266), .A2(new_n268), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n277), .A2(KEYINPUT71), .A3(KEYINPUT32), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n234), .A2(new_n244), .ZN(new_n280));
  INV_X1    g094(.A(new_n250), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(new_n252), .ZN(new_n283));
  AOI22_X1  g097(.A1(new_n241), .A2(new_n243), .B1(new_n233), .B2(new_n253), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT28), .ZN(new_n285));
  OAI211_X1 g099(.A(new_n283), .B(new_n259), .C1(new_n284), .C2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT29), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n282), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(KEYINPUT70), .ZN(new_n289));
  INV_X1    g103(.A(G902), .ZN(new_n290));
  OAI22_X1  g104(.A1(new_n255), .A2(new_n256), .B1(new_n232), .B2(new_n228), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n252), .B1(new_n291), .B2(KEYINPUT28), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n292), .A2(KEYINPUT29), .A3(new_n250), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT70), .ZN(new_n294));
  NAND4_X1  g108(.A1(new_n282), .A2(new_n286), .A3(new_n294), .A4(new_n287), .ZN(new_n295));
  NAND4_X1  g109(.A1(new_n289), .A2(new_n290), .A3(new_n293), .A4(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(G472), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n279), .A2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT81), .ZN(new_n299));
  INV_X1    g113(.A(G104), .ZN(new_n300));
  OAI21_X1  g114(.A(KEYINPUT3), .B1(new_n300), .B2(G107), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT3), .ZN(new_n302));
  INV_X1    g116(.A(G107), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n302), .A2(new_n303), .A3(G104), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n300), .A2(G107), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n301), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(G101), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n299), .B1(new_n307), .B2(KEYINPUT4), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT4), .ZN(new_n309));
  NAND4_X1  g123(.A1(new_n306), .A2(KEYINPUT81), .A3(new_n309), .A4(G101), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  XNOR2_X1  g125(.A(KEYINPUT80), .B(G101), .ZN(new_n312));
  NAND4_X1  g126(.A1(new_n312), .A2(new_n305), .A3(new_n301), .A4(new_n304), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n307), .A2(KEYINPUT4), .A3(new_n313), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n311), .A2(new_n233), .A3(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT5), .ZN(new_n316));
  INV_X1    g130(.A(G119), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n316), .A2(new_n317), .A3(G116), .ZN(new_n318));
  XNOR2_X1  g132(.A(new_n318), .B(KEYINPUT85), .ZN(new_n319));
  INV_X1    g133(.A(new_n230), .ZN(new_n320));
  OAI211_X1 g134(.A(new_n319), .B(G113), .C1(new_n316), .C2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(new_n305), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n300), .A2(G107), .ZN(new_n323));
  OAI21_X1  g137(.A(G101), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n313), .A2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  OR2_X1    g140(.A1(new_n320), .A2(new_n231), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n321), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n315), .A2(new_n328), .ZN(new_n329));
  XOR2_X1   g143(.A(G110), .B(G122), .Z(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT6), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT86), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n334), .B1(new_n329), .B2(new_n330), .ZN(new_n335));
  INV_X1    g149(.A(new_n330), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n315), .A2(KEYINPUT86), .A3(new_n336), .A4(new_n328), .ZN(new_n337));
  AOI22_X1  g151(.A1(new_n335), .A2(new_n337), .B1(new_n330), .B2(new_n329), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n333), .B1(new_n338), .B2(new_n332), .ZN(new_n339));
  OR2_X1    g153(.A1(new_n197), .A2(G125), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n218), .A2(G125), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(G224), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n343), .A2(G953), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n342), .B(new_n344), .ZN(new_n345));
  AOI21_X1  g159(.A(G902), .B1(new_n339), .B2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT7), .ZN(new_n347));
  INV_X1    g161(.A(new_n344), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n347), .B1(new_n348), .B2(KEYINPUT88), .ZN(new_n349));
  OR2_X1    g163(.A1(new_n348), .A2(KEYINPUT88), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n340), .A2(new_n341), .A3(new_n349), .A4(new_n350), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n342), .B1(new_n347), .B2(new_n344), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n351), .B1(new_n352), .B2(KEYINPUT87), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n353), .B1(KEYINPUT87), .B2(new_n352), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n335), .A2(new_n337), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n321), .A2(new_n327), .ZN(new_n356));
  XNOR2_X1  g170(.A(new_n356), .B(new_n326), .ZN(new_n357));
  XNOR2_X1  g171(.A(new_n330), .B(KEYINPUT8), .ZN(new_n358));
  OAI211_X1 g172(.A(new_n354), .B(new_n355), .C1(new_n357), .C2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n346), .A2(new_n359), .ZN(new_n360));
  OAI21_X1  g174(.A(G210), .B1(G237), .B2(G902), .ZN(new_n361));
  XOR2_X1   g175(.A(new_n361), .B(KEYINPUT89), .Z(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n360), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(G952), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n365), .A2(G953), .ZN(new_n366));
  NAND2_X1  g180(.A1(G234), .A2(G237), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  XOR2_X1   g182(.A(KEYINPUT21), .B(G898), .Z(new_n369));
  NAND3_X1  g183(.A1(new_n367), .A2(G902), .A3(G953), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n368), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  XNOR2_X1  g185(.A(new_n371), .B(KEYINPUT97), .ZN(new_n372));
  OAI21_X1  g186(.A(G214), .B1(G237), .B2(G902), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n346), .A2(new_n362), .A3(new_n359), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n364), .A2(new_n372), .A3(new_n373), .A4(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(G478), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n376), .A2(KEYINPUT15), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT96), .ZN(new_n378));
  INV_X1    g192(.A(G116), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n379), .A2(KEYINPUT14), .A3(G122), .ZN(new_n380));
  XNOR2_X1  g194(.A(G116), .B(G122), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  OAI211_X1 g196(.A(G107), .B(new_n380), .C1(new_n382), .C2(KEYINPUT14), .ZN(new_n383));
  XNOR2_X1  g197(.A(G128), .B(G143), .ZN(new_n384));
  XNOR2_X1  g198(.A(new_n384), .B(KEYINPUT95), .ZN(new_n385));
  AND2_X1   g199(.A1(new_n385), .A2(new_n199), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n385), .A2(new_n199), .ZN(new_n387));
  OAI221_X1 g201(.A(new_n383), .B1(G107), .B2(new_n382), .C1(new_n386), .C2(new_n387), .ZN(new_n388));
  XOR2_X1   g202(.A(KEYINPUT9), .B(G234), .Z(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  XNOR2_X1  g204(.A(KEYINPUT72), .B(G217), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  NOR3_X1   g206(.A1(new_n390), .A2(G953), .A3(new_n392), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n199), .B1(new_n384), .B2(KEYINPUT13), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n190), .A2(G128), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n394), .B1(KEYINPUT13), .B2(new_n395), .ZN(new_n396));
  OR2_X1    g210(.A1(new_n396), .A2(KEYINPUT94), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n385), .A2(new_n199), .ZN(new_n398));
  XNOR2_X1  g212(.A(new_n381), .B(new_n303), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n396), .A2(KEYINPUT94), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n397), .A2(new_n398), .A3(new_n399), .A4(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n388), .A2(new_n393), .A3(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n393), .B1(new_n388), .B2(new_n401), .ZN(new_n404));
  OAI211_X1 g218(.A(new_n378), .B(new_n290), .C1(new_n403), .C2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n388), .A2(new_n401), .ZN(new_n407));
  INV_X1    g221(.A(new_n393), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(new_n402), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n378), .B1(new_n410), .B2(new_n290), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n377), .B1(new_n406), .B2(new_n411), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n412), .B1(new_n377), .B2(new_n411), .ZN(new_n413));
  NOR2_X1   g227(.A1(G475), .A2(G902), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT93), .ZN(new_n415));
  XNOR2_X1  g229(.A(G125), .B(G140), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT19), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  XNOR2_X1  g232(.A(new_n416), .B(KEYINPUT74), .ZN(new_n419));
  AOI211_X1 g233(.A(G146), .B(new_n418), .C1(new_n419), .C2(new_n417), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT16), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(G125), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n422), .A2(G140), .ZN(new_n423));
  AOI211_X1 g237(.A(new_n188), .B(new_n423), .C1(KEYINPUT16), .C2(new_n416), .ZN(new_n424));
  OAI21_X1  g238(.A(KEYINPUT91), .B1(new_n420), .B2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT91), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n423), .B1(new_n416), .B2(KEYINPUT16), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(G146), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n419), .A2(new_n417), .ZN(new_n429));
  INV_X1    g243(.A(new_n418), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  OAI211_X1 g245(.A(new_n426), .B(new_n428), .C1(new_n431), .C2(G146), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n245), .A2(new_n246), .A3(G214), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n190), .A2(KEYINPUT90), .ZN(new_n434));
  OR2_X1    g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  OR2_X1    g249(.A1(new_n190), .A2(KEYINPUT90), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n436), .A2(new_n433), .A3(new_n434), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(new_n203), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n435), .A2(new_n437), .A3(G131), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n425), .A2(new_n432), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n419), .A2(new_n188), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n443), .B1(new_n188), .B2(new_n416), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT18), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n438), .B1(new_n445), .B2(new_n203), .ZN(new_n446));
  OAI211_X1 g260(.A(new_n444), .B(new_n446), .C1(new_n445), .C2(new_n440), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n442), .A2(new_n447), .ZN(new_n448));
  XNOR2_X1  g262(.A(G113), .B(G122), .ZN(new_n449));
  XNOR2_X1  g263(.A(new_n449), .B(new_n300), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n448), .A2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT92), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT17), .ZN(new_n454));
  OR3_X1    g268(.A1(new_n440), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n427), .A2(G146), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n456), .A2(new_n424), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n439), .A2(new_n454), .A3(new_n440), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n453), .B1(new_n440), .B2(new_n454), .ZN(new_n459));
  NAND4_X1  g273(.A1(new_n455), .A2(new_n457), .A3(new_n458), .A4(new_n459), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n447), .A2(new_n450), .A3(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n415), .B1(new_n452), .B2(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n450), .B1(new_n442), .B2(new_n447), .ZN(new_n463));
  INV_X1    g277(.A(new_n461), .ZN(new_n464));
  NOR3_X1   g278(.A1(new_n463), .A2(KEYINPUT93), .A3(new_n464), .ZN(new_n465));
  OAI211_X1 g279(.A(KEYINPUT20), .B(new_n414), .C1(new_n462), .C2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT20), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n463), .A2(new_n464), .ZN(new_n468));
  INV_X1    g282(.A(new_n414), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n450), .B1(new_n447), .B2(new_n460), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n290), .B1(new_n464), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(G475), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n466), .A2(new_n470), .A3(new_n473), .ZN(new_n474));
  NOR3_X1   g288(.A1(new_n375), .A2(new_n413), .A3(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT23), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n476), .B1(new_n317), .B2(G128), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n194), .A2(KEYINPUT23), .A3(G119), .ZN(new_n478));
  OAI211_X1 g292(.A(new_n477), .B(new_n478), .C1(G119), .C2(new_n194), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(G110), .ZN(new_n480));
  XOR2_X1   g294(.A(KEYINPUT24), .B(G110), .Z(new_n481));
  XNOR2_X1  g295(.A(G119), .B(G128), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  OAI211_X1 g297(.A(new_n480), .B(new_n483), .C1(new_n456), .C2(new_n424), .ZN(new_n484));
  XNOR2_X1  g298(.A(KEYINPUT73), .B(G110), .ZN(new_n485));
  OAI22_X1  g299(.A1(new_n479), .A2(new_n485), .B1(new_n482), .B2(new_n481), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n443), .A2(new_n428), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  XNOR2_X1  g302(.A(KEYINPUT22), .B(G137), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n246), .A2(G221), .A3(G234), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n489), .B(new_n490), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n491), .B(KEYINPUT75), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n488), .A2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT76), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n484), .A2(new_n491), .A3(new_n487), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n488), .A2(KEYINPUT76), .A3(new_n492), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n495), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n392), .B1(G234), .B2(new_n290), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n500), .A2(G902), .ZN(new_n501));
  XOR2_X1   g315(.A(new_n501), .B(KEYINPUT77), .Z(new_n502));
  NAND2_X1  g316(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n503), .B(KEYINPUT78), .ZN(new_n504));
  OAI21_X1  g318(.A(KEYINPUT25), .B1(new_n498), .B2(G902), .ZN(new_n505));
  AND3_X1   g319(.A1(new_n488), .A2(KEYINPUT76), .A3(new_n492), .ZN(new_n506));
  AOI21_X1  g320(.A(KEYINPUT76), .B1(new_n488), .B2(new_n492), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT25), .ZN(new_n509));
  NAND4_X1  g323(.A1(new_n508), .A2(new_n509), .A3(new_n290), .A4(new_n496), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n505), .A2(new_n500), .A3(new_n510), .ZN(new_n511));
  AND2_X1   g325(.A1(new_n504), .A2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n311), .A2(new_n219), .A3(new_n314), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(KEYINPUT82), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT82), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n311), .A2(new_n516), .A3(new_n219), .A4(new_n314), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n196), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n189), .A2(KEYINPUT83), .A3(KEYINPUT1), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(G128), .ZN(new_n521));
  AOI21_X1  g335(.A(KEYINPUT83), .B1(new_n189), .B2(KEYINPUT1), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n519), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n325), .B1(new_n523), .B2(new_n193), .ZN(new_n524));
  OR2_X1    g338(.A1(new_n524), .A2(KEYINPUT10), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n326), .A2(KEYINPUT10), .A3(new_n197), .ZN(new_n526));
  XOR2_X1   g340(.A(new_n214), .B(KEYINPUT84), .Z(new_n527));
  NAND4_X1  g341(.A1(new_n518), .A2(new_n525), .A3(new_n526), .A4(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n246), .A2(G227), .ZN(new_n529));
  XNOR2_X1  g343(.A(new_n529), .B(G140), .ZN(new_n530));
  XNOR2_X1  g344(.A(KEYINPUT79), .B(G110), .ZN(new_n531));
  XNOR2_X1  g345(.A(new_n530), .B(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  AND2_X1   g347(.A1(new_n528), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n518), .A2(new_n525), .A3(new_n526), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(new_n214), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n326), .A2(new_n197), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n214), .B1(new_n537), .B2(new_n524), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT12), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n538), .B(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n528), .A2(new_n540), .ZN(new_n541));
  AOI22_X1  g355(.A1(new_n534), .A2(new_n536), .B1(new_n541), .B2(new_n532), .ZN(new_n542));
  OAI21_X1  g356(.A(G469), .B1(new_n542), .B2(G902), .ZN(new_n543));
  INV_X1    g357(.A(G469), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n533), .B1(new_n536), .B2(new_n528), .ZN(new_n545));
  AND3_X1   g359(.A1(new_n528), .A2(new_n533), .A3(new_n540), .ZN(new_n546));
  OAI211_X1 g360(.A(new_n544), .B(new_n290), .C1(new_n545), .C2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n543), .A2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(G221), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n549), .B1(new_n389), .B2(new_n290), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n513), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n298), .A2(new_n475), .A3(new_n553), .ZN(new_n554));
  XOR2_X1   g368(.A(new_n554), .B(new_n312), .Z(G3));
  NOR2_X1   g369(.A1(new_n266), .A2(G902), .ZN(new_n556));
  INV_X1    g370(.A(G472), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n558), .A2(new_n277), .ZN(new_n559));
  INV_X1    g373(.A(new_n375), .ZN(new_n560));
  AND3_X1   g374(.A1(new_n553), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n410), .A2(KEYINPUT33), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT33), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n409), .A2(new_n563), .A3(new_n402), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n562), .A2(G478), .A3(new_n564), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n376), .A2(new_n290), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n410), .A2(new_n376), .A3(new_n290), .ZN(new_n568));
  AND3_X1   g382(.A1(new_n565), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n474), .A2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n561), .A2(new_n571), .ZN(new_n572));
  XOR2_X1   g386(.A(KEYINPUT34), .B(G104), .Z(new_n573));
  XNOR2_X1  g387(.A(new_n572), .B(new_n573), .ZN(G6));
  OR2_X1    g388(.A1(new_n462), .A2(new_n465), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n467), .B1(new_n576), .B2(new_n469), .ZN(new_n577));
  AND2_X1   g391(.A1(new_n466), .A2(new_n473), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(new_n413), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n561), .A2(new_n581), .ZN(new_n582));
  XOR2_X1   g396(.A(KEYINPUT35), .B(G107), .Z(new_n583));
  XNOR2_X1  g397(.A(new_n582), .B(new_n583), .ZN(G9));
  INV_X1    g398(.A(KEYINPUT98), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n488), .B(new_n585), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n492), .A2(KEYINPUT36), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n586), .B(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(new_n502), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(new_n511), .ZN(new_n590));
  XOR2_X1   g404(.A(new_n590), .B(KEYINPUT99), .Z(new_n591));
  NOR2_X1   g405(.A1(new_n591), .A2(new_n552), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n475), .A2(new_n592), .A3(new_n559), .ZN(new_n593));
  XOR2_X1   g407(.A(KEYINPUT37), .B(G110), .Z(new_n594));
  XNOR2_X1  g408(.A(new_n594), .B(KEYINPUT100), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n593), .B(new_n595), .ZN(G12));
  NAND2_X1  g410(.A1(new_n364), .A2(new_n374), .ZN(new_n597));
  INV_X1    g411(.A(new_n373), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  XOR2_X1   g413(.A(new_n368), .B(KEYINPUT102), .Z(new_n600));
  INV_X1    g414(.A(new_n370), .ZN(new_n601));
  XOR2_X1   g415(.A(KEYINPUT101), .B(G900), .Z(new_n602));
  AOI21_X1  g416(.A(new_n600), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NOR3_X1   g417(.A1(new_n579), .A2(new_n580), .A3(new_n603), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n298), .A2(new_n599), .A3(new_n592), .A4(new_n604), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n605), .B(G128), .ZN(G30));
  INV_X1    g420(.A(KEYINPUT38), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n597), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n364), .A2(KEYINPUT38), .A3(new_n374), .ZN(new_n609));
  AND2_X1   g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(new_n552), .ZN(new_n611));
  XOR2_X1   g425(.A(new_n603), .B(KEYINPUT39), .Z(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT40), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n611), .A2(KEYINPUT40), .A3(new_n612), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n610), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n590), .B(KEYINPUT99), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n474), .A2(new_n413), .A3(new_n373), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT103), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n620), .B(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n261), .ZN(new_n623));
  INV_X1    g437(.A(new_n259), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n623), .B1(new_n291), .B2(new_n624), .ZN(new_n625));
  OAI21_X1  g439(.A(G472), .B1(new_n625), .B2(G902), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n279), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n617), .A2(new_n622), .A3(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(G143), .ZN(G45));
  NOR2_X1   g443(.A1(new_n570), .A2(new_n603), .ZN(new_n630));
  NAND4_X1  g444(.A1(new_n298), .A2(new_n599), .A3(new_n592), .A4(new_n630), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n631), .B(G146), .ZN(G48));
  OAI21_X1  g446(.A(new_n290), .B1(new_n545), .B2(new_n546), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(G469), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n634), .A2(new_n551), .A3(new_n547), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n375), .A2(new_n635), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n298), .A2(new_n512), .A3(new_n571), .A4(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(KEYINPUT41), .B(G113), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(G15));
  NAND4_X1  g453(.A1(new_n298), .A2(new_n512), .A3(new_n581), .A4(new_n636), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(G116), .ZN(G18));
  INV_X1    g455(.A(new_n635), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n298), .A2(new_n475), .A3(new_n618), .A4(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(G119), .ZN(G21));
  OAI21_X1  g458(.A(KEYINPUT105), .B1(new_n556), .B2(new_n557), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT104), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n292), .B(new_n646), .ZN(new_n647));
  OAI211_X1 g461(.A(new_n251), .B(new_n262), .C1(new_n647), .C2(new_n259), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(new_n271), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT105), .ZN(new_n650));
  OAI211_X1 g464(.A(new_n650), .B(G472), .C1(new_n266), .C2(G902), .ZN(new_n651));
  AND3_X1   g465(.A1(new_n645), .A2(new_n649), .A3(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n372), .ZN(new_n653));
  NOR3_X1   g467(.A1(new_n597), .A2(new_n619), .A3(new_n653), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n652), .A2(new_n512), .A3(new_n642), .A4(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(G122), .ZN(G24));
  NOR3_X1   g470(.A1(new_n597), .A2(new_n598), .A3(new_n635), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n652), .A2(new_n618), .A3(new_n630), .A4(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(KEYINPUT106), .B(G125), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G27));
  INV_X1    g474(.A(new_n603), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n571), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n662), .A2(KEYINPUT42), .ZN(new_n663));
  INV_X1    g477(.A(new_n547), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n536), .A2(new_n528), .A3(new_n533), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n541), .A2(new_n532), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n665), .A2(new_n666), .A3(G469), .ZN(new_n667));
  NAND2_X1  g481(.A1(G469), .A2(G902), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  OAI21_X1  g483(.A(KEYINPUT107), .B1(new_n664), .B2(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT107), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n543), .A2(new_n671), .A3(new_n547), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n670), .A2(new_n551), .A3(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n374), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n362), .B1(new_n346), .B2(new_n359), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n373), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n298), .A2(new_n663), .A3(new_n677), .A4(new_n512), .ZN(new_n678));
  NOR3_X1   g492(.A1(new_n664), .A2(new_n669), .A3(KEYINPUT107), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n671), .B1(new_n543), .B2(new_n547), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n598), .B1(new_n364), .B2(new_n374), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n681), .A2(new_n630), .A3(new_n551), .A4(new_n682), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n297), .A2(new_n275), .A3(new_n269), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(new_n512), .ZN(new_n685));
  OAI21_X1  g499(.A(KEYINPUT42), .B1(new_n683), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n678), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(new_n203), .ZN(G33));
  NAND4_X1  g502(.A1(new_n298), .A2(new_n512), .A3(new_n677), .A4(new_n604), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G134), .ZN(G36));
  NAND4_X1  g504(.A1(new_n578), .A2(KEYINPUT43), .A3(new_n470), .A4(new_n569), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n569), .A2(new_n470), .A3(new_n466), .A4(new_n473), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT43), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT109), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n591), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n691), .A2(new_n694), .A3(KEYINPUT109), .ZN(new_n698));
  INV_X1    g512(.A(new_n559), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n697), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT44), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n702), .A2(new_n676), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n542), .A2(KEYINPUT45), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n665), .A2(new_n666), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT45), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n704), .A2(new_n707), .A3(G469), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(new_n668), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT46), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n664), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n708), .A2(KEYINPUT46), .A3(new_n668), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n713), .A2(new_n551), .A3(new_n612), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(KEYINPUT108), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT108), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n713), .A2(new_n716), .A3(new_n551), .A4(new_n612), .ZN(new_n717));
  AOI22_X1  g531(.A1(new_n715), .A2(new_n717), .B1(new_n700), .B2(new_n701), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n703), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G137), .ZN(G39));
  INV_X1    g534(.A(KEYINPUT47), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n709), .A2(new_n710), .ZN(new_n722));
  AND3_X1   g536(.A1(new_n722), .A2(new_n547), .A3(new_n712), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n721), .B1(new_n723), .B2(new_n550), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n713), .A2(KEYINPUT47), .A3(new_n551), .ZN(new_n725));
  AOI211_X1 g539(.A(new_n662), .B(new_n676), .C1(new_n724), .C2(new_n725), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n298), .A2(new_n512), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G140), .ZN(G42));
  NAND2_X1  g543(.A1(new_n365), .A2(new_n246), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n611), .A2(new_n618), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n731), .B1(new_n279), .B2(new_n297), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n579), .A2(new_n603), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n732), .A2(new_n580), .A3(new_n733), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n645), .A2(new_n618), .A3(new_n649), .A4(new_n651), .ZN(new_n735));
  INV_X1    g549(.A(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(new_n673), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n736), .A2(new_n630), .A3(new_n737), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n676), .B1(new_n734), .B2(new_n738), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n637), .A2(new_n643), .A3(new_n593), .A4(new_n655), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n678), .A2(new_n689), .A3(new_n686), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n570), .B1(new_n580), .B2(new_n474), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n553), .A2(new_n559), .A3(new_n560), .A4(new_n742), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n640), .A2(new_n554), .A3(new_n743), .ZN(new_n744));
  NOR4_X1   g558(.A1(new_n739), .A2(new_n740), .A3(new_n741), .A4(new_n744), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n605), .A2(new_n631), .A3(new_n658), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT52), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n673), .B1(new_n279), .B2(new_n626), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n589), .A2(new_n511), .A3(new_n661), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT110), .ZN(new_n750));
  AND2_X1   g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n749), .A2(new_n750), .ZN(new_n752));
  NOR4_X1   g566(.A1(new_n597), .A2(new_n619), .A3(new_n751), .A4(new_n752), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n747), .B1(new_n748), .B2(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(new_n754), .ZN(new_n755));
  OAI21_X1  g569(.A(KEYINPUT111), .B1(new_n746), .B2(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n627), .A2(new_n753), .A3(new_n737), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n605), .A2(new_n631), .A3(new_n658), .A4(new_n757), .ZN(new_n758));
  XOR2_X1   g572(.A(KEYINPUT112), .B(KEYINPUT52), .Z(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  OAI211_X1 g574(.A(new_n732), .B(new_n599), .C1(new_n604), .C2(new_n630), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT111), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n761), .A2(new_n762), .A3(new_n658), .A4(new_n754), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n756), .A2(new_n760), .A3(new_n763), .ZN(new_n764));
  AOI21_X1  g578(.A(KEYINPUT53), .B1(new_n745), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n758), .A2(new_n747), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n761), .A2(new_n658), .A3(new_n754), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NOR3_X1   g582(.A1(new_n740), .A2(new_n741), .A3(new_n744), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n734), .A2(new_n738), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(new_n682), .ZN(new_n771));
  XOR2_X1   g585(.A(KEYINPUT113), .B(KEYINPUT53), .Z(new_n772));
  AND4_X1   g586(.A1(new_n768), .A2(new_n769), .A3(new_n771), .A4(new_n772), .ZN(new_n773));
  OAI21_X1  g587(.A(KEYINPUT54), .B1(new_n765), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(KEYINPUT114), .ZN(new_n775));
  INV_X1    g589(.A(new_n772), .ZN(new_n776));
  AND2_X1   g590(.A1(new_n766), .A2(new_n767), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n740), .A2(new_n744), .ZN(new_n778));
  INV_X1    g592(.A(new_n741), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n778), .A2(new_n771), .A3(new_n779), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n776), .B1(new_n777), .B2(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT54), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n745), .A2(new_n764), .A3(KEYINPUT53), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n781), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT114), .ZN(new_n785));
  OAI211_X1 g599(.A(new_n785), .B(KEYINPUT54), .C1(new_n765), .C2(new_n773), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n775), .A2(new_n784), .A3(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT51), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT115), .ZN(new_n789));
  AOI21_X1  g603(.A(KEYINPUT47), .B1(new_n713), .B2(new_n551), .ZN(new_n790));
  AOI211_X1 g604(.A(new_n721), .B(new_n550), .C1(new_n711), .C2(new_n712), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n789), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n724), .A2(KEYINPUT115), .A3(new_n725), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n634), .A2(new_n550), .A3(new_n547), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n792), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n695), .A2(new_n600), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n645), .A2(new_n512), .A3(new_n649), .A4(new_n651), .ZN(new_n797));
  NOR3_X1   g611(.A1(new_n796), .A2(new_n797), .A3(new_n676), .ZN(new_n798));
  AND2_X1   g612(.A1(new_n795), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n682), .A2(new_n642), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(KEYINPUT116), .ZN(new_n801));
  INV_X1    g615(.A(new_n796), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n803), .A2(new_n736), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n627), .A2(new_n513), .ZN(new_n805));
  INV_X1    g619(.A(new_n368), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n474), .A2(new_n569), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n801), .A2(new_n805), .A3(new_n806), .A4(new_n807), .ZN(new_n808));
  NOR3_X1   g622(.A1(new_n796), .A2(new_n797), .A3(new_n373), .ZN(new_n809));
  AND3_X1   g623(.A1(new_n608), .A2(new_n609), .A3(new_n642), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT50), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  AOI21_X1  g627(.A(KEYINPUT50), .B1(new_n809), .B2(new_n810), .ZN(new_n814));
  OAI211_X1 g628(.A(new_n804), .B(new_n808), .C1(new_n813), .C2(new_n814), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n788), .B1(new_n799), .B2(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n803), .A2(new_n512), .A3(new_n684), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(KEYINPUT48), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n801), .A2(new_n805), .A3(new_n806), .A4(new_n571), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n802), .A2(new_n512), .A3(new_n652), .A4(new_n657), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n819), .A2(new_n366), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n821), .A2(KEYINPUT117), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT117), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n819), .A2(new_n823), .A3(new_n366), .A4(new_n820), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  XNOR2_X1  g639(.A(new_n811), .B(new_n812), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n724), .A2(new_n725), .A3(new_n794), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n788), .B1(new_n827), .B2(new_n798), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n826), .A2(new_n804), .A3(new_n808), .A4(new_n828), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n816), .A2(new_n818), .A3(new_n825), .A4(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n830), .A2(KEYINPUT118), .ZN(new_n831));
  AND2_X1   g645(.A1(new_n829), .A2(new_n825), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT118), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n832), .A2(new_n833), .A3(new_n818), .A4(new_n816), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n831), .A2(new_n834), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n730), .B1(new_n787), .B2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(new_n627), .ZN(new_n837));
  NOR4_X1   g651(.A1(new_n513), .A2(new_n692), .A3(new_n598), .A4(new_n550), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n634), .A2(new_n547), .ZN(new_n839));
  XOR2_X1   g653(.A(new_n839), .B(KEYINPUT49), .Z(new_n840));
  NAND4_X1  g654(.A1(new_n837), .A2(new_n610), .A3(new_n838), .A4(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n836), .A2(new_n841), .ZN(G75));
  INV_X1    g656(.A(KEYINPUT56), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n781), .A2(new_n783), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(G902), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n843), .B1(new_n845), .B2(new_n363), .ZN(new_n846));
  XNOR2_X1  g660(.A(new_n339), .B(new_n345), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n847), .B(KEYINPUT55), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n246), .A2(G952), .ZN(new_n850));
  INV_X1    g664(.A(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(new_n848), .ZN(new_n852));
  OAI211_X1 g666(.A(new_n843), .B(new_n852), .C1(new_n845), .C2(new_n363), .ZN(new_n853));
  AND3_X1   g667(.A1(new_n849), .A2(new_n851), .A3(new_n853), .ZN(G51));
  XOR2_X1   g668(.A(new_n668), .B(KEYINPUT57), .Z(new_n855));
  AND3_X1   g669(.A1(new_n781), .A2(new_n782), .A3(new_n783), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n782), .B1(new_n781), .B2(new_n783), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n855), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n858), .B1(new_n545), .B2(new_n546), .ZN(new_n859));
  OR2_X1    g673(.A1(new_n845), .A2(new_n708), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n850), .B1(new_n859), .B2(new_n860), .ZN(G54));
  NAND4_X1  g675(.A1(new_n844), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n862));
  AND2_X1   g676(.A1(new_n862), .A2(new_n576), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n862), .A2(new_n576), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n863), .A2(new_n864), .A3(new_n850), .ZN(G60));
  NAND2_X1  g679(.A1(new_n562), .A2(new_n564), .ZN(new_n866));
  INV_X1    g680(.A(new_n866), .ZN(new_n867));
  XNOR2_X1  g681(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n868));
  XNOR2_X1  g682(.A(new_n567), .B(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n870), .B1(new_n856), .B2(new_n857), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n871), .A2(new_n851), .ZN(new_n872));
  INV_X1    g686(.A(new_n869), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n787), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n872), .B1(new_n874), .B2(new_n867), .ZN(G63));
  NAND2_X1  g689(.A1(G217), .A2(G902), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n876), .B(KEYINPUT60), .ZN(new_n877));
  INV_X1    g691(.A(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n844), .A2(new_n878), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n850), .B1(new_n879), .B2(new_n498), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n877), .B1(new_n781), .B2(new_n783), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n588), .B(KEYINPUT120), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT121), .ZN(new_n884));
  OAI211_X1 g698(.A(new_n880), .B(new_n883), .C1(new_n884), .C2(KEYINPUT61), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT61), .ZN(new_n886));
  OAI211_X1 g700(.A(new_n884), .B(new_n851), .C1(new_n881), .C2(new_n499), .ZN(new_n887));
  INV_X1    g701(.A(new_n883), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n851), .B1(new_n881), .B2(new_n499), .ZN(new_n889));
  OAI211_X1 g703(.A(new_n886), .B(new_n887), .C1(new_n888), .C2(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n885), .A2(new_n890), .ZN(G66));
  INV_X1    g705(.A(new_n369), .ZN(new_n892));
  OAI21_X1  g706(.A(G953), .B1(new_n892), .B2(new_n343), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n893), .B1(new_n778), .B2(G953), .ZN(new_n894));
  INV_X1    g708(.A(new_n339), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n895), .B1(G898), .B2(new_n246), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n896), .B(KEYINPUT122), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n894), .B(new_n897), .ZN(G69));
  XOR2_X1   g712(.A(new_n229), .B(new_n431), .Z(new_n899));
  AOI21_X1  g713(.A(new_n246), .B1(G227), .B2(G900), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n628), .A2(new_n658), .A3(new_n761), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT62), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n901), .B(new_n902), .ZN(new_n903));
  AOI22_X1  g717(.A1(new_n718), .A2(new_n703), .B1(new_n726), .B2(new_n727), .ZN(new_n904));
  AND3_X1   g718(.A1(new_n742), .A2(new_n611), .A3(new_n612), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n905), .A2(new_n298), .A3(new_n512), .A4(new_n682), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n903), .A2(new_n904), .A3(new_n906), .ZN(new_n907));
  AOI211_X1 g721(.A(new_n899), .B(new_n900), .C1(new_n907), .C2(new_n246), .ZN(new_n908));
  XOR2_X1   g722(.A(new_n741), .B(KEYINPUT123), .Z(new_n909));
  AOI21_X1  g723(.A(new_n685), .B1(new_n715), .B2(new_n717), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n597), .A2(new_n619), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n746), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n909), .A2(new_n904), .A3(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT124), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n909), .A2(new_n904), .A3(KEYINPUT124), .A4(new_n912), .ZN(new_n916));
  AND2_X1   g730(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(new_n900), .ZN(new_n918));
  XNOR2_X1  g732(.A(KEYINPUT125), .B(G900), .ZN(new_n919));
  OAI22_X1  g733(.A1(new_n917), .A2(G953), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n908), .B1(new_n920), .B2(new_n899), .ZN(G72));
  NAND2_X1  g735(.A1(G472), .A2(G902), .ZN(new_n922));
  XOR2_X1   g736(.A(new_n922), .B(KEYINPUT63), .Z(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(KEYINPUT126), .ZN(new_n924));
  INV_X1    g738(.A(new_n778), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n924), .B1(new_n907), .B2(new_n925), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n926), .A2(new_n250), .A3(new_n280), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n282), .A2(new_n261), .ZN(new_n928));
  OAI211_X1 g742(.A(new_n923), .B(new_n928), .C1(new_n765), .C2(new_n773), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n927), .A2(new_n851), .A3(new_n929), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n915), .A2(new_n778), .A3(new_n916), .ZN(new_n931));
  AOI211_X1 g745(.A(new_n250), .B(new_n280), .C1(new_n931), .C2(new_n924), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n930), .A2(new_n932), .ZN(G57));
endmodule


