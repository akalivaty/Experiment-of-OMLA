//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 1 0 0 0 1 0 0 0 0 1 0 1 0 1 0 1 0 1 1 1 1 1 1 0 0 1 0 0 0 0 0 0 0 1 1 0 1 1 0 1 0 1 0 1 0 0 0 0 0 1 0 0 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:58 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n723, new_n725, new_n726, new_n727,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n736,
    new_n737, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n757, new_n758, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020;
  INV_X1    g000(.A(G119), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G128), .ZN(new_n188));
  INV_X1    g002(.A(G128), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G119), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT24), .B(G110), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT23), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n190), .A2(new_n194), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n189), .A2(KEYINPUT23), .A3(G119), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n195), .A2(new_n196), .A3(new_n188), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n193), .B1(new_n197), .B2(G110), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT76), .ZN(new_n199));
  XNOR2_X1  g013(.A(new_n198), .B(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G140), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G125), .ZN(new_n202));
  INV_X1    g016(.A(G125), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G140), .ZN(new_n204));
  NAND4_X1  g018(.A1(new_n202), .A2(new_n204), .A3(KEYINPUT74), .A4(KEYINPUT16), .ZN(new_n205));
  AND3_X1   g019(.A1(new_n202), .A2(new_n204), .A3(KEYINPUT16), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT74), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n207), .B1(new_n202), .B2(KEYINPUT16), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n205), .B1(new_n206), .B2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G146), .ZN(new_n210));
  INV_X1    g024(.A(G146), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n202), .A2(new_n204), .A3(new_n211), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n200), .A2(new_n210), .A3(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n197), .A2(KEYINPUT72), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT72), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n195), .A2(new_n196), .A3(new_n215), .A4(new_n188), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n214), .A2(G110), .A3(new_n216), .ZN(new_n217));
  XOR2_X1   g031(.A(new_n217), .B(KEYINPUT73), .Z(new_n218));
  INV_X1    g032(.A(KEYINPUT75), .ZN(new_n219));
  OAI211_X1 g033(.A(new_n211), .B(new_n205), .C1(new_n206), .C2(new_n208), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n210), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  OR3_X1    g035(.A1(new_n209), .A2(new_n219), .A3(G146), .ZN(new_n222));
  OR2_X1    g036(.A1(new_n191), .A2(new_n192), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n213), .B1(new_n218), .B2(new_n224), .ZN(new_n225));
  XNOR2_X1  g039(.A(KEYINPUT22), .B(G137), .ZN(new_n226));
  INV_X1    g040(.A(G953), .ZN(new_n227));
  AND3_X1   g041(.A1(new_n227), .A2(G221), .A3(G234), .ZN(new_n228));
  XOR2_X1   g042(.A(new_n226), .B(new_n228), .Z(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n225), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(G902), .ZN(new_n232));
  XNOR2_X1  g046(.A(new_n217), .B(KEYINPUT73), .ZN(new_n233));
  NAND4_X1  g047(.A1(new_n233), .A2(new_n222), .A3(new_n221), .A4(new_n223), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n234), .A2(new_n213), .A3(new_n229), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n231), .A2(new_n232), .A3(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT25), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n231), .A2(KEYINPUT25), .A3(new_n235), .A4(new_n232), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(G217), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n241), .B1(G234), .B2(new_n232), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  AND2_X1   g057(.A1(new_n231), .A2(new_n235), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n242), .A2(G902), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n243), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT71), .ZN(new_n248));
  NOR2_X1   g062(.A1(G472), .A2(G902), .ZN(new_n249));
  NOR2_X1   g063(.A1(G237), .A2(G953), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(G210), .ZN(new_n251));
  XNOR2_X1  g065(.A(new_n251), .B(KEYINPUT27), .ZN(new_n252));
  XNOR2_X1  g066(.A(KEYINPUT26), .B(G101), .ZN(new_n253));
  XNOR2_X1  g067(.A(new_n252), .B(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT11), .ZN(new_n255));
  INV_X1    g069(.A(G134), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n255), .B1(new_n256), .B2(G137), .ZN(new_n257));
  INV_X1    g071(.A(G137), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n258), .A2(KEYINPUT11), .A3(G134), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n256), .A2(G137), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n257), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G131), .ZN(new_n262));
  INV_X1    g076(.A(G131), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n257), .A2(new_n259), .A3(new_n263), .A4(new_n260), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n211), .A2(G143), .ZN(new_n266));
  INV_X1    g080(.A(G143), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G146), .ZN(new_n268));
  AND2_X1   g082(.A1(KEYINPUT0), .A2(G128), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n266), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  XNOR2_X1  g084(.A(G143), .B(G146), .ZN(new_n271));
  XNOR2_X1  g085(.A(KEYINPUT0), .B(G128), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n270), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n265), .A2(new_n274), .ZN(new_n275));
  XNOR2_X1  g089(.A(G116), .B(G119), .ZN(new_n276));
  XNOR2_X1  g090(.A(KEYINPUT2), .B(G113), .ZN(new_n277));
  XNOR2_X1  g091(.A(new_n276), .B(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n266), .A2(new_n268), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n266), .A2(KEYINPUT1), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n279), .A2(new_n280), .A3(G128), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT64), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n282), .A2(new_n258), .A3(G134), .ZN(new_n283));
  OAI21_X1  g097(.A(KEYINPUT64), .B1(new_n256), .B2(G137), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n258), .A2(G134), .ZN(new_n285));
  OAI211_X1 g099(.A(G131), .B(new_n283), .C1(new_n284), .C2(new_n285), .ZN(new_n286));
  OAI211_X1 g100(.A(new_n266), .B(new_n268), .C1(KEYINPUT1), .C2(new_n189), .ZN(new_n287));
  NAND4_X1  g101(.A1(new_n281), .A2(new_n286), .A3(new_n264), .A4(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n275), .A2(new_n278), .A3(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT66), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n275), .A2(new_n288), .ZN(new_n291));
  INV_X1    g105(.A(new_n276), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(new_n277), .ZN(new_n293));
  XOR2_X1   g107(.A(KEYINPUT2), .B(G113), .Z(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(new_n276), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n290), .B1(new_n291), .B2(new_n296), .ZN(new_n297));
  AOI211_X1 g111(.A(KEYINPUT66), .B(new_n278), .C1(new_n275), .C2(new_n288), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n289), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(KEYINPUT28), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT28), .ZN(new_n301));
  AND3_X1   g115(.A1(new_n289), .A2(KEYINPUT67), .A3(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(KEYINPUT67), .B1(new_n289), .B2(new_n301), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n254), .B1(new_n300), .B2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(new_n288), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n273), .B1(new_n264), .B2(new_n262), .ZN(new_n307));
  NOR3_X1   g121(.A1(new_n306), .A2(new_n307), .A3(KEYINPUT30), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT30), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n309), .B1(new_n275), .B2(new_n288), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n296), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  XNOR2_X1  g125(.A(KEYINPUT65), .B(KEYINPUT31), .ZN(new_n312));
  NAND4_X1  g126(.A1(new_n311), .A2(new_n289), .A3(new_n254), .A4(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(KEYINPUT30), .B1(new_n306), .B2(new_n307), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n275), .A2(new_n309), .A3(new_n288), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n278), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(new_n289), .ZN(new_n317));
  INV_X1    g131(.A(new_n254), .ZN(new_n318));
  NOR3_X1   g132(.A1(new_n316), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT31), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n313), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n249), .B1(new_n305), .B2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT68), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  OAI211_X1 g138(.A(KEYINPUT68), .B(new_n249), .C1(new_n305), .C2(new_n321), .ZN(new_n325));
  XOR2_X1   g139(.A(KEYINPUT69), .B(KEYINPUT32), .Z(new_n326));
  AND3_X1   g140(.A1(new_n324), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n296), .B1(new_n306), .B2(new_n307), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(KEYINPUT66), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n291), .A2(new_n290), .A3(new_n296), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n317), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  OAI211_X1 g145(.A(new_n304), .B(new_n254), .C1(new_n331), .C2(new_n301), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n318), .B1(new_n316), .B2(new_n317), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT29), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n332), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n328), .A2(new_n289), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(KEYINPUT28), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n318), .A2(new_n334), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n304), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  AND2_X1   g153(.A1(new_n339), .A2(new_n232), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n335), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(G472), .ZN(new_n342));
  AND2_X1   g156(.A1(new_n249), .A2(KEYINPUT32), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n343), .B1(new_n305), .B2(new_n321), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(KEYINPUT70), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT70), .ZN(new_n346));
  OAI211_X1 g160(.A(new_n346), .B(new_n343), .C1(new_n305), .C2(new_n321), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n342), .A2(new_n345), .A3(new_n347), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n248), .B1(new_n327), .B2(new_n348), .ZN(new_n349));
  AND2_X1   g163(.A1(new_n345), .A2(new_n347), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n324), .A2(new_n325), .A3(new_n326), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n350), .A2(new_n351), .A3(KEYINPUT71), .A4(new_n342), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n247), .B1(new_n349), .B2(new_n352), .ZN(new_n353));
  XNOR2_X1  g167(.A(G110), .B(G122), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(G104), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(G107), .ZN(new_n357));
  OR2_X1    g171(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n358));
  INV_X1    g172(.A(G107), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(G104), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n357), .B1(new_n358), .B2(new_n360), .ZN(new_n361));
  NOR2_X1   g175(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n356), .A2(G107), .ZN(new_n363));
  NAND2_X1  g177(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n362), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  OAI21_X1  g179(.A(G101), .B1(new_n361), .B2(new_n365), .ZN(new_n366));
  AND2_X1   g180(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n358), .B1(new_n360), .B2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(G101), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n363), .A2(new_n362), .ZN(new_n370));
  NAND4_X1  g184(.A1(new_n368), .A2(new_n369), .A3(new_n357), .A4(new_n370), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n366), .A2(KEYINPUT4), .A3(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT81), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT4), .ZN(new_n374));
  OAI211_X1 g188(.A(new_n374), .B(G101), .C1(new_n361), .C2(new_n365), .ZN(new_n375));
  NAND4_X1  g189(.A1(new_n372), .A2(new_n373), .A3(new_n296), .A4(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(G113), .ZN(new_n377));
  XOR2_X1   g191(.A(KEYINPUT82), .B(KEYINPUT5), .Z(new_n378));
  INV_X1    g192(.A(G116), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n379), .A2(G119), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n377), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  XNOR2_X1  g195(.A(KEYINPUT82), .B(KEYINPUT5), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n276), .A2(new_n382), .ZN(new_n383));
  AOI22_X1  g197(.A1(new_n381), .A2(new_n383), .B1(new_n276), .B2(new_n294), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n360), .A2(new_n357), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(G101), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n384), .A2(new_n371), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n376), .A2(new_n387), .ZN(new_n388));
  AND2_X1   g202(.A1(new_n296), .A2(new_n375), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n373), .B1(new_n389), .B2(new_n372), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n355), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n372), .A2(new_n296), .A3(new_n375), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(KEYINPUT81), .ZN(new_n393));
  NAND4_X1  g207(.A1(new_n393), .A2(new_n354), .A3(new_n387), .A4(new_n376), .ZN(new_n394));
  NAND4_X1  g208(.A1(new_n391), .A2(new_n394), .A3(KEYINPUT83), .A4(KEYINPUT6), .ZN(new_n395));
  AND3_X1   g209(.A1(new_n391), .A2(KEYINPUT6), .A3(new_n394), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT6), .ZN(new_n397));
  OAI211_X1 g211(.A(new_n397), .B(new_n355), .C1(new_n388), .C2(new_n390), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT83), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n395), .B1(new_n396), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n281), .A2(new_n287), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(new_n203), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT85), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n403), .B(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n273), .A2(G125), .ZN(new_n406));
  XNOR2_X1  g220(.A(new_n406), .B(KEYINPUT84), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n227), .A2(G224), .ZN(new_n409));
  XNOR2_X1  g223(.A(new_n408), .B(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n401), .A2(new_n411), .ZN(new_n412));
  XOR2_X1   g226(.A(new_n354), .B(KEYINPUT8), .Z(new_n413));
  NAND2_X1  g227(.A1(new_n371), .A2(new_n386), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n413), .B1(new_n384), .B2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT5), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n381), .B1(new_n416), .B2(new_n292), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(new_n295), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT86), .ZN(new_n419));
  XNOR2_X1  g233(.A(new_n418), .B(new_n419), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n415), .B1(new_n420), .B2(new_n414), .ZN(new_n421));
  NAND4_X1  g235(.A1(new_n405), .A2(KEYINPUT7), .A3(new_n409), .A4(new_n407), .ZN(new_n422));
  AND3_X1   g236(.A1(new_n421), .A2(new_n394), .A3(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT87), .ZN(new_n424));
  OR2_X1    g238(.A1(new_n405), .A2(new_n424), .ZN(new_n425));
  AOI22_X1  g239(.A1(new_n405), .A2(new_n424), .B1(G125), .B2(new_n273), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT7), .ZN(new_n427));
  OR2_X1    g241(.A1(new_n427), .A2(KEYINPUT88), .ZN(new_n428));
  AOI22_X1  g242(.A1(KEYINPUT88), .A2(new_n427), .B1(new_n227), .B2(G224), .ZN(new_n429));
  AOI22_X1  g243(.A1(new_n425), .A2(new_n426), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  AOI21_X1  g245(.A(G902), .B1(new_n423), .B2(new_n431), .ZN(new_n432));
  OAI21_X1  g246(.A(G210), .B1(G237), .B2(G902), .ZN(new_n433));
  XOR2_X1   g247(.A(new_n433), .B(KEYINPUT89), .Z(new_n434));
  NAND3_X1  g248(.A1(new_n412), .A2(new_n432), .A3(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(new_n434), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n391), .A2(KEYINPUT6), .A3(new_n394), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n437), .A2(new_n399), .A3(new_n398), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n410), .B1(new_n438), .B2(new_n395), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n421), .A2(new_n394), .A3(new_n422), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n232), .B1(new_n440), .B2(new_n430), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n436), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  OAI21_X1  g256(.A(G214), .B1(G237), .B2(G902), .ZN(new_n443));
  XNOR2_X1  g257(.A(new_n443), .B(KEYINPUT80), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n435), .A2(new_n442), .A3(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(G469), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n371), .A2(new_n287), .A3(new_n281), .A4(new_n386), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  AOI22_X1  g262(.A1(new_n371), .A2(new_n386), .B1(new_n287), .B2(new_n281), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n265), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT12), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(new_n265), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n414), .A2(new_n402), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n453), .B1(new_n454), .B2(new_n447), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(KEYINPUT12), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n452), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n372), .A2(new_n274), .A3(new_n375), .ZN(new_n458));
  INV_X1    g272(.A(new_n402), .ZN(new_n459));
  NAND4_X1  g273(.A1(new_n459), .A2(KEYINPUT10), .A3(new_n371), .A4(new_n386), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT10), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n447), .A2(new_n461), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n458), .A2(new_n453), .A3(new_n460), .A4(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n457), .A2(new_n463), .ZN(new_n464));
  XNOR2_X1  g278(.A(G110), .B(G140), .ZN(new_n465));
  INV_X1    g279(.A(G227), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n466), .A2(G953), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n465), .B(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n464), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n458), .A2(new_n462), .A3(new_n460), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(new_n265), .ZN(new_n471));
  INV_X1    g285(.A(new_n468), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n471), .A2(new_n463), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n469), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n446), .B1(new_n474), .B2(new_n232), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n455), .A2(KEYINPUT12), .ZN(new_n476));
  AOI211_X1 g290(.A(new_n451), .B(new_n453), .C1(new_n454), .C2(new_n447), .ZN(new_n477));
  OAI211_X1 g291(.A(new_n463), .B(new_n472), .C1(new_n476), .C2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT78), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n457), .A2(KEYINPUT78), .A3(new_n463), .A4(new_n472), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n471), .A2(new_n463), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(new_n468), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n480), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n484), .A2(new_n446), .A3(new_n232), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT79), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n484), .A2(KEYINPUT79), .A3(new_n446), .A4(new_n232), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n475), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT92), .ZN(new_n490));
  AND3_X1   g304(.A1(new_n202), .A2(new_n204), .A3(KEYINPUT19), .ZN(new_n491));
  AOI21_X1  g305(.A(KEYINPUT19), .B1(new_n202), .B2(new_n204), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n211), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(KEYINPUT91), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT19), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n203), .A2(G140), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n201), .A2(G125), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n202), .A2(new_n204), .A3(KEYINPUT19), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT91), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n500), .A2(new_n501), .A3(new_n211), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n494), .A2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(G237), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n504), .A2(new_n227), .A3(G214), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n505), .A2(new_n267), .ZN(new_n506));
  AOI21_X1  g320(.A(G143), .B1(new_n250), .B2(G214), .ZN(new_n507));
  OAI21_X1  g321(.A(G131), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n505), .A2(new_n267), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n250), .A2(G143), .A3(G214), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n509), .A2(new_n263), .A3(new_n510), .ZN(new_n511));
  AOI22_X1  g325(.A1(new_n209), .A2(G146), .B1(new_n508), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n509), .A2(new_n510), .ZN(new_n513));
  NAND2_X1  g327(.A1(KEYINPUT18), .A2(G131), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  OAI21_X1  g329(.A(KEYINPUT90), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT90), .ZN(new_n517));
  NAND4_X1  g331(.A1(new_n509), .A2(new_n517), .A3(new_n510), .A4(new_n514), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  OAI21_X1  g333(.A(G146), .B1(new_n496), .B2(new_n497), .ZN(new_n520));
  AOI22_X1  g334(.A1(new_n513), .A2(new_n515), .B1(new_n520), .B2(new_n212), .ZN(new_n521));
  AOI22_X1  g335(.A1(new_n503), .A2(new_n512), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  XNOR2_X1  g336(.A(G113), .B(G122), .ZN(new_n523));
  XNOR2_X1  g337(.A(new_n523), .B(new_n356), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n490), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n519), .A2(new_n521), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n501), .B1(new_n500), .B2(new_n211), .ZN(new_n527));
  AOI211_X1 g341(.A(KEYINPUT91), .B(G146), .C1(new_n498), .C2(new_n499), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n508), .A2(new_n511), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n210), .A2(new_n530), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n526), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(new_n524), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n532), .A2(KEYINPUT92), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n525), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n221), .A2(new_n222), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n513), .A2(KEYINPUT17), .A3(G131), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n537), .B1(new_n530), .B2(KEYINPUT17), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n536), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n540), .A2(new_n524), .A3(new_n526), .ZN(new_n541));
  AOI21_X1  g355(.A(KEYINPUT94), .B1(new_n535), .B2(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n538), .B1(new_n222), .B2(new_n221), .ZN(new_n543));
  INV_X1    g357(.A(new_n526), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  AOI22_X1  g359(.A1(new_n525), .A2(new_n534), .B1(new_n545), .B2(new_n524), .ZN(new_n546));
  NOR2_X1   g360(.A1(G475), .A2(G902), .ZN(new_n547));
  XNOR2_X1  g361(.A(new_n547), .B(KEYINPUT93), .ZN(new_n548));
  OAI22_X1  g362(.A1(new_n542), .A2(KEYINPUT20), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(KEYINPUT92), .B1(new_n532), .B2(new_n533), .ZN(new_n550));
  NOR3_X1   g364(.A1(new_n522), .A2(new_n490), .A3(new_n524), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n541), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT20), .ZN(new_n553));
  INV_X1    g367(.A(new_n548), .ZN(new_n554));
  NAND4_X1  g368(.A1(new_n552), .A2(KEYINPUT94), .A3(new_n553), .A4(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n549), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n227), .A2(G952), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n557), .B1(G234), .B2(G237), .ZN(new_n558));
  AOI211_X1 g372(.A(new_n232), .B(new_n227), .C1(G234), .C2(G237), .ZN(new_n559));
  XNOR2_X1  g373(.A(KEYINPUT21), .B(G898), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT97), .ZN(new_n563));
  OAI22_X1  g377(.A1(new_n563), .A2(KEYINPUT13), .B1(new_n267), .B2(G128), .ZN(new_n564));
  AND2_X1   g378(.A1(new_n563), .A2(KEYINPUT13), .ZN(new_n565));
  OAI21_X1  g379(.A(G134), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  XNOR2_X1  g380(.A(G128), .B(G143), .ZN(new_n567));
  XOR2_X1   g381(.A(new_n566), .B(new_n567), .Z(new_n568));
  OR2_X1    g382(.A1(KEYINPUT96), .A2(G122), .ZN(new_n569));
  NAND2_X1  g383(.A1(KEYINPUT96), .A2(G122), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n379), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(G122), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n572), .A2(G116), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n574), .A2(new_n359), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n359), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n568), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  XOR2_X1   g392(.A(new_n573), .B(KEYINPUT14), .Z(new_n579));
  OAI21_X1  g393(.A(G107), .B1(new_n579), .B2(new_n571), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n567), .B(new_n256), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n580), .A2(new_n576), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n578), .A2(new_n582), .ZN(new_n583));
  XNOR2_X1  g397(.A(KEYINPUT9), .B(G234), .ZN(new_n584));
  NOR3_X1   g398(.A1(new_n584), .A2(new_n241), .A3(G953), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n578), .A2(new_n582), .A3(new_n585), .ZN(new_n588));
  AOI21_X1  g402(.A(G902), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(G478), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n590), .A2(KEYINPUT15), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n589), .B(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n524), .B1(new_n540), .B2(new_n526), .ZN(new_n593));
  NOR3_X1   g407(.A1(new_n543), .A2(new_n533), .A3(new_n544), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n232), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(KEYINPUT95), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n533), .B1(new_n543), .B2(new_n544), .ZN(new_n597));
  AOI21_X1  g411(.A(G902), .B1(new_n541), .B2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT95), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n596), .A2(G475), .A3(new_n600), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n556), .A2(new_n562), .A3(new_n592), .A4(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(G221), .ZN(new_n603));
  INV_X1    g417(.A(new_n584), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n603), .B1(new_n604), .B2(new_n232), .ZN(new_n605));
  NOR4_X1   g419(.A1(new_n445), .A2(new_n489), .A3(new_n602), .A4(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n353), .A2(new_n606), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(G101), .ZN(G3));
  NOR2_X1   g422(.A1(new_n489), .A2(new_n605), .ZN(new_n609));
  INV_X1    g423(.A(new_n247), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n324), .A2(new_n325), .ZN(new_n611));
  INV_X1    g425(.A(G472), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n232), .B1(new_n305), .B2(new_n321), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT98), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n612), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n613), .A2(KEYINPUT98), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n611), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n609), .A2(new_n610), .A3(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n587), .A2(new_n588), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(KEYINPUT33), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT33), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n587), .A2(new_n623), .A3(new_n588), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n622), .A2(G478), .A3(new_n624), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n590), .A2(new_n232), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n626), .B1(new_n589), .B2(new_n590), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n628), .B1(new_n556), .B2(new_n601), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n435), .A2(new_n442), .A3(new_n443), .ZN(new_n631));
  NOR3_X1   g445(.A1(new_n630), .A2(new_n631), .A3(new_n561), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n620), .A2(new_n632), .ZN(new_n633));
  XOR2_X1   g447(.A(KEYINPUT34), .B(G104), .Z(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G6));
  XOR2_X1   g449(.A(new_n589), .B(new_n591), .Z(new_n636));
  AND3_X1   g450(.A1(new_n435), .A2(new_n442), .A3(new_n443), .ZN(new_n637));
  OAI21_X1  g451(.A(G475), .B1(new_n598), .B2(new_n599), .ZN(new_n638));
  AOI211_X1 g452(.A(KEYINPUT95), .B(G902), .C1(new_n541), .C2(new_n597), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n553), .B1(new_n546), .B2(new_n548), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n552), .A2(KEYINPUT20), .A3(new_n554), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n561), .B(KEYINPUT99), .ZN(new_n645));
  AND4_X1   g459(.A1(new_n636), .A2(new_n637), .A3(new_n644), .A4(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n620), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(KEYINPUT100), .ZN(new_n648));
  XNOR2_X1  g462(.A(KEYINPUT35), .B(G107), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G9));
  NOR2_X1   g464(.A1(new_n230), .A2(KEYINPUT36), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT101), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n234), .A2(new_n653), .A3(new_n213), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n653), .B1(new_n234), .B2(new_n213), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n652), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n225), .A2(KEYINPUT101), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n658), .A2(new_n651), .A3(new_n654), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(new_n245), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n243), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n606), .A2(new_n618), .A3(new_n662), .ZN(new_n663));
  XOR2_X1   g477(.A(KEYINPUT37), .B(G110), .Z(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G12));
  NAND2_X1  g479(.A1(new_n349), .A2(new_n352), .ZN(new_n666));
  AND2_X1   g480(.A1(new_n641), .A2(new_n642), .ZN(new_n667));
  XOR2_X1   g481(.A(new_n558), .B(KEYINPUT103), .Z(new_n668));
  OR2_X1    g482(.A1(KEYINPUT102), .A2(G900), .ZN(new_n669));
  NAND2_X1  g483(.A1(KEYINPUT102), .A2(G900), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n559), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n667), .A2(new_n636), .A3(new_n601), .A4(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT104), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n644), .A2(KEYINPUT104), .A3(new_n636), .A4(new_n672), .ZN(new_n676));
  AND3_X1   g490(.A1(new_n675), .A2(new_n637), .A3(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(new_n475), .ZN(new_n678));
  AOI22_X1  g492(.A1(new_n478), .A2(new_n479), .B1(new_n482), .B2(new_n468), .ZN(new_n679));
  AOI21_X1  g493(.A(G902), .B1(new_n679), .B2(new_n481), .ZN(new_n680));
  AOI21_X1  g494(.A(KEYINPUT79), .B1(new_n680), .B2(new_n446), .ZN(new_n681));
  INV_X1    g495(.A(new_n488), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n678), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n605), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n683), .A2(new_n684), .A3(new_n662), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n666), .A2(new_n677), .A3(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G128), .ZN(G30));
  XNOR2_X1  g502(.A(new_n672), .B(KEYINPUT39), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n609), .A2(new_n689), .ZN(new_n690));
  AND2_X1   g504(.A1(new_n690), .A2(KEYINPUT40), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n690), .A2(KEYINPUT40), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n435), .A2(new_n442), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(KEYINPUT38), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n318), .B1(new_n311), .B2(new_n289), .ZN(new_n695));
  OAI21_X1  g509(.A(new_n232), .B1(new_n336), .B2(new_n254), .ZN(new_n696));
  OAI21_X1  g510(.A(G472), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(KEYINPUT105), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n350), .A2(new_n351), .A3(new_n698), .ZN(new_n699));
  AOI22_X1  g513(.A1(new_n240), .A2(new_n242), .B1(new_n660), .B2(new_n245), .ZN(new_n700));
  INV_X1    g514(.A(G475), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n701), .B1(new_n595), .B2(KEYINPUT95), .ZN(new_n702));
  AOI22_X1  g516(.A1(new_n549), .A2(new_n555), .B1(new_n702), .B2(new_n600), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n703), .A2(new_n592), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n699), .A2(new_n443), .A3(new_n700), .A4(new_n704), .ZN(new_n705));
  NOR4_X1   g519(.A1(new_n691), .A2(new_n692), .A3(new_n694), .A4(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(new_n267), .ZN(G45));
  INV_X1    g521(.A(KEYINPUT106), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n708), .B1(new_n629), .B2(new_n672), .ZN(new_n709));
  INV_X1    g523(.A(new_n672), .ZN(new_n710));
  NOR4_X1   g524(.A1(new_n703), .A2(KEYINPUT106), .A3(new_n628), .A4(new_n710), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n666), .A2(new_n712), .A3(new_n686), .A4(new_n637), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G146), .ZN(G48));
  NAND2_X1  g528(.A1(new_n487), .A2(new_n488), .ZN(new_n715));
  OR2_X1    g529(.A1(new_n680), .A2(new_n446), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n715), .A2(new_n684), .A3(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n353), .A2(new_n632), .A3(new_n718), .ZN(new_n719));
  XOR2_X1   g533(.A(KEYINPUT41), .B(G113), .Z(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(KEYINPUT107), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n719), .B(new_n721), .ZN(G15));
  NAND3_X1  g536(.A1(new_n353), .A2(new_n646), .A3(new_n718), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G116), .ZN(G18));
  NOR2_X1   g538(.A1(new_n717), .A2(new_n631), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n602), .A2(new_n700), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n666), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G119), .ZN(G21));
  NOR3_X1   g542(.A1(new_n631), .A2(new_n592), .A3(new_n703), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n254), .B1(new_n304), .B2(new_n337), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n249), .B1(new_n321), .B2(new_n730), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n731), .B1(new_n614), .B2(new_n612), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n247), .A2(new_n732), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n729), .A2(new_n718), .A3(new_n645), .A4(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G122), .ZN(G24));
  NOR2_X1   g549(.A1(new_n700), .A2(new_n732), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n712), .A2(new_n725), .A3(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G125), .ZN(G27));
  INV_X1    g552(.A(new_n443), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n739), .B1(new_n435), .B2(new_n442), .ZN(new_n740));
  AND3_X1   g554(.A1(new_n740), .A2(new_n683), .A3(new_n684), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n666), .A2(new_n712), .A3(new_n610), .A4(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT108), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT42), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n353), .A2(KEYINPUT108), .A3(new_n712), .A4(new_n741), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n744), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(new_n322), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n344), .B1(new_n748), .B2(KEYINPUT32), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT109), .ZN(new_n750));
  OR2_X1    g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  AOI22_X1  g565(.A1(new_n749), .A2(new_n750), .B1(G472), .B2(new_n341), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n247), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n753), .A2(KEYINPUT42), .A3(new_n712), .A4(new_n741), .ZN(new_n754));
  AND2_X1   g568(.A1(new_n747), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(new_n263), .ZN(G33));
  AND2_X1   g570(.A1(new_n675), .A2(new_n676), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n666), .A2(new_n610), .A3(new_n757), .A4(new_n741), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G134), .ZN(G36));
  AND2_X1   g573(.A1(new_n469), .A2(new_n473), .ZN(new_n760));
  OR2_X1    g574(.A1(new_n760), .A2(KEYINPUT45), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(KEYINPUT45), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n761), .A2(G469), .A3(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(G469), .A2(G902), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT46), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n763), .A2(KEYINPUT46), .A3(new_n764), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n767), .A2(new_n715), .A3(new_n768), .ZN(new_n769));
  AND3_X1   g583(.A1(new_n769), .A2(new_n684), .A3(new_n689), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n618), .A2(new_n700), .ZN(new_n771));
  INV_X1    g585(.A(new_n628), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n703), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(KEYINPUT43), .ZN(new_n774));
  OR2_X1    g588(.A1(new_n773), .A2(KEYINPUT43), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n771), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT44), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n770), .A2(new_n778), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n740), .B1(new_n776), .B2(new_n777), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT110), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  OAI211_X1 g596(.A(KEYINPUT110), .B(new_n740), .C1(new_n776), .C2(new_n777), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n779), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(new_n258), .ZN(G39));
  NAND2_X1  g599(.A1(new_n769), .A2(new_n684), .ZN(new_n786));
  XNOR2_X1  g600(.A(KEYINPUT111), .B(KEYINPUT47), .ZN(new_n787));
  INV_X1    g601(.A(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT47), .ZN(new_n790));
  OAI211_X1 g604(.A(new_n769), .B(new_n684), .C1(KEYINPUT111), .C2(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n712), .A2(new_n247), .A3(new_n740), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n792), .A2(new_n666), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n789), .A2(new_n791), .A3(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(G140), .ZN(G42));
  XNOR2_X1  g609(.A(new_n557), .B(KEYINPUT119), .ZN(new_n796));
  INV_X1    g610(.A(new_n558), .ZN(new_n797));
  NOR3_X1   g611(.A1(new_n699), .A2(new_n247), .A3(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(new_n740), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n799), .A2(new_n717), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n775), .A2(new_n774), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n802), .A2(new_n668), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n803), .A2(new_n733), .ZN(new_n804));
  INV_X1    g618(.A(new_n725), .ZN(new_n805));
  OAI221_X1 g619(.A(new_n796), .B1(new_n801), .B2(new_n630), .C1(new_n804), .C2(new_n805), .ZN(new_n806));
  AND2_X1   g620(.A1(new_n803), .A2(new_n800), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(new_n753), .ZN(new_n808));
  OR2_X1    g622(.A1(new_n808), .A2(KEYINPUT48), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(KEYINPUT48), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n806), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT51), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n789), .A2(new_n791), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n715), .A2(new_n605), .A3(new_n716), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n804), .A2(new_n799), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n812), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n548), .B1(new_n535), .B2(new_n541), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT94), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n552), .A2(new_n819), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n818), .B1(new_n820), .B2(new_n553), .ZN(new_n821));
  INV_X1    g635(.A(new_n555), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n601), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n801), .A2(new_n823), .A3(new_n772), .ZN(new_n824));
  OR2_X1    g638(.A1(new_n824), .A2(KEYINPUT118), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n807), .A2(new_n736), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n824), .A2(KEYINPUT118), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n817), .A2(new_n825), .A3(new_n826), .A4(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n694), .A2(new_n739), .A3(new_n718), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT116), .ZN(new_n830));
  OR2_X1    g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n829), .A2(new_n830), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n831), .A2(new_n733), .A3(new_n832), .A4(new_n803), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n833), .B(KEYINPUT50), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n811), .B1(new_n828), .B2(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT117), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT50), .ZN(new_n838));
  XNOR2_X1  g652(.A(new_n833), .B(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n839), .A2(KEYINPUT117), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n825), .A2(new_n826), .A3(new_n827), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n813), .A2(KEYINPUT115), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT115), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n789), .A2(new_n843), .A3(new_n791), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n842), .A2(new_n844), .A3(new_n814), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n841), .B1(new_n845), .B2(new_n816), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n837), .A2(new_n840), .A3(new_n846), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n835), .B1(new_n847), .B2(new_n812), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n723), .A2(new_n719), .A3(new_n727), .A4(new_n734), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n849), .B1(new_n747), .B2(new_n754), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n662), .A2(new_n710), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n729), .A2(new_n609), .A3(new_n699), .A4(new_n851), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n713), .A2(new_n687), .A3(new_n737), .A4(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT52), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n685), .B1(new_n349), .B2(new_n352), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n823), .A2(new_n772), .A3(new_n672), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n857), .A2(KEYINPUT106), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n629), .A2(new_n708), .A3(new_n672), .ZN(new_n859));
  AND3_X1   g673(.A1(new_n858), .A2(new_n859), .A3(new_n736), .ZN(new_n860));
  AOI22_X1  g674(.A1(new_n856), .A2(new_n677), .B1(new_n860), .B2(new_n725), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n861), .A2(KEYINPUT52), .A3(new_n713), .A4(new_n852), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n855), .A2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT112), .ZN(new_n864));
  AND3_X1   g678(.A1(new_n606), .A2(new_n666), .A3(new_n610), .ZN(new_n865));
  INV_X1    g679(.A(new_n445), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n703), .A2(new_n592), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n823), .A2(new_n628), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n866), .A2(new_n867), .A3(new_n645), .A4(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n445), .A2(new_n602), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n870), .A2(new_n609), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n618), .A2(new_n662), .ZN(new_n872));
  OAI22_X1  g686(.A1(new_n619), .A2(new_n869), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n864), .B1(new_n865), .B2(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n868), .A2(new_n867), .A3(new_n645), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n875), .A2(new_n445), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n876), .A2(new_n610), .A3(new_n609), .A4(new_n618), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n607), .A2(new_n663), .A3(new_n877), .A4(KEYINPUT112), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n874), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n860), .A2(new_n741), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n758), .A2(new_n880), .ZN(new_n881));
  AND4_X1   g695(.A1(new_n592), .A2(new_n662), .A3(new_n644), .A4(new_n672), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n666), .A2(new_n741), .A3(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT113), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n666), .A2(KEYINPUT113), .A3(new_n741), .A4(new_n882), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n881), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n850), .A2(new_n863), .A3(new_n879), .A4(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT53), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  AND2_X1   g704(.A1(new_n879), .A2(new_n887), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n891), .A2(KEYINPUT53), .A3(new_n850), .A4(new_n863), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n893), .A2(KEYINPUT54), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n889), .B1(new_n874), .B2(new_n878), .ZN(new_n895));
  AND4_X1   g709(.A1(new_n850), .A2(new_n863), .A3(new_n895), .A4(new_n887), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT114), .ZN(new_n897));
  AOI22_X1  g711(.A1(new_n896), .A2(new_n897), .B1(new_n888), .B2(new_n889), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT54), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n850), .A2(new_n863), .A3(new_n895), .A4(new_n887), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(KEYINPUT114), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n898), .A2(new_n899), .A3(new_n901), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n848), .A2(new_n894), .A3(new_n902), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n903), .B1(G952), .B2(G953), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n715), .A2(new_n716), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n905), .B(KEYINPUT49), .Z(new_n906));
  NAND3_X1  g720(.A1(new_n610), .A2(new_n684), .A3(new_n444), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n907), .A2(new_n699), .A3(new_n773), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n906), .A2(new_n908), .A3(new_n694), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n904), .A2(new_n909), .ZN(G75));
  AND3_X1   g724(.A1(new_n879), .A2(new_n887), .A3(KEYINPUT53), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n911), .A2(new_n897), .A3(new_n850), .A4(new_n863), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n890), .A2(new_n912), .A3(new_n901), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n913), .A2(G902), .A3(new_n434), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT56), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n401), .B(new_n410), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n916), .B(KEYINPUT55), .ZN(new_n917));
  AND3_X1   g731(.A1(new_n914), .A2(new_n915), .A3(new_n917), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n917), .B1(new_n914), .B2(new_n915), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n227), .A2(G952), .ZN(new_n920));
  NOR3_X1   g734(.A1(new_n918), .A2(new_n919), .A3(new_n920), .ZN(G51));
  XOR2_X1   g735(.A(new_n764), .B(KEYINPUT57), .Z(new_n922));
  AOI21_X1  g736(.A(new_n899), .B1(new_n898), .B2(new_n901), .ZN(new_n923));
  AND4_X1   g737(.A1(new_n899), .A2(new_n890), .A3(new_n912), .A4(new_n901), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n922), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n925), .A2(new_n484), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n913), .A2(G902), .ZN(new_n927));
  OR2_X1    g741(.A1(new_n927), .A2(new_n763), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n920), .B1(new_n926), .B2(new_n928), .ZN(G54));
  INV_X1    g743(.A(KEYINPUT121), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n232), .B1(new_n898), .B2(new_n901), .ZN(new_n931));
  NAND2_X1  g745(.A1(KEYINPUT58), .A2(G475), .ZN(new_n932));
  XOR2_X1   g746(.A(new_n932), .B(KEYINPUT120), .Z(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n552), .B1(new_n931), .B2(new_n934), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n546), .A2(new_n933), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n913), .A2(G902), .A3(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(new_n920), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n930), .B1(new_n935), .B2(new_n939), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n546), .B1(new_n927), .B2(new_n933), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n941), .A2(KEYINPUT121), .A3(new_n938), .A4(new_n937), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n940), .A2(new_n942), .ZN(G60));
  NAND2_X1  g757(.A1(new_n622), .A2(new_n624), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n902), .A2(new_n894), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n626), .B(KEYINPUT59), .Z(new_n946));
  AOI21_X1  g760(.A(new_n944), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n944), .A2(new_n946), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n913), .A2(KEYINPUT54), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n948), .B1(new_n949), .B2(new_n902), .ZN(new_n950));
  NOR3_X1   g764(.A1(new_n947), .A2(new_n920), .A3(new_n950), .ZN(G63));
  NAND2_X1  g765(.A1(G217), .A2(G902), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n952), .B(KEYINPUT122), .Z(new_n953));
  XOR2_X1   g767(.A(new_n953), .B(KEYINPUT60), .Z(new_n954));
  NAND3_X1  g768(.A1(new_n913), .A2(new_n660), .A3(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(new_n954), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n956), .B1(new_n898), .B2(new_n901), .ZN(new_n957));
  OAI211_X1 g771(.A(new_n938), .B(new_n955), .C1(new_n957), .C2(new_n244), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT61), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n913), .A2(new_n954), .ZN(new_n961));
  INV_X1    g775(.A(new_n244), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n920), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n963), .A2(KEYINPUT61), .A3(new_n955), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n960), .A2(new_n964), .ZN(G66));
  INV_X1    g779(.A(new_n849), .ZN(new_n966));
  AOI21_X1  g780(.A(G953), .B1(new_n879), .B2(new_n966), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n967), .B(KEYINPUT123), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT124), .ZN(new_n969));
  INV_X1    g783(.A(G224), .ZN(new_n970));
  OAI21_X1  g784(.A(G953), .B1(new_n560), .B2(new_n970), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n968), .A2(new_n969), .A3(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(new_n972), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n969), .B1(new_n968), .B2(new_n971), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(new_n401), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n976), .B1(G898), .B2(new_n227), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n975), .B(new_n977), .ZN(G69));
  NAND2_X1  g792(.A1(G900), .A2(G953), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n769), .A2(new_n684), .A3(new_n689), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n753), .A2(new_n729), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n982), .B(KEYINPUT126), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n794), .A2(new_n758), .ZN(new_n984));
  NOR3_X1   g798(.A1(new_n983), .A2(new_n755), .A3(new_n984), .ZN(new_n985));
  INV_X1    g799(.A(KEYINPUT125), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n861), .A2(new_n713), .ZN(new_n987));
  OR3_X1    g801(.A1(new_n784), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n986), .B1(new_n784), .B2(new_n987), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n985), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n979), .B1(new_n990), .B2(G953), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n314), .A2(new_n315), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n992), .B(new_n500), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n991), .A2(new_n993), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n227), .B1(G227), .B2(G900), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n995), .B(KEYINPUT127), .ZN(new_n996));
  INV_X1    g810(.A(new_n996), .ZN(new_n997));
  OR2_X1    g811(.A1(new_n706), .A2(new_n987), .ZN(new_n998));
  OR2_X1    g812(.A1(new_n998), .A2(KEYINPUT62), .ZN(new_n999));
  INV_X1    g813(.A(new_n784), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n998), .A2(KEYINPUT62), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n740), .A2(new_n867), .A3(new_n868), .ZN(new_n1002));
  NOR2_X1   g816(.A1(new_n690), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1003), .A2(new_n353), .ZN(new_n1004));
  AND2_X1   g818(.A1(new_n794), .A2(new_n1004), .ZN(new_n1005));
  NAND4_X1  g819(.A1(new_n999), .A2(new_n1000), .A3(new_n1001), .A4(new_n1005), .ZN(new_n1006));
  NOR2_X1   g820(.A1(new_n993), .A2(G953), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  AND3_X1   g822(.A1(new_n994), .A2(new_n997), .A3(new_n1008), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n997), .B1(new_n994), .B2(new_n1008), .ZN(new_n1010));
  NOR2_X1   g824(.A1(new_n1009), .A2(new_n1010), .ZN(G72));
  INV_X1    g825(.A(new_n319), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1012), .A2(new_n333), .ZN(new_n1013));
  NAND2_X1  g827(.A1(G472), .A2(G902), .ZN(new_n1014));
  XOR2_X1   g828(.A(new_n1014), .B(KEYINPUT63), .Z(new_n1015));
  OAI21_X1  g829(.A(new_n938), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1016));
  AND3_X1   g830(.A1(new_n893), .A2(new_n1015), .A3(new_n1013), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n879), .A2(new_n966), .ZN(new_n1018));
  AOI211_X1 g832(.A(new_n1018), .B(new_n1013), .C1(new_n1006), .C2(new_n254), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n990), .A2(new_n318), .ZN(new_n1020));
  AOI211_X1 g834(.A(new_n1016), .B(new_n1017), .C1(new_n1019), .C2(new_n1020), .ZN(G57));
endmodule


