//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 1 0 1 1 0 1 0 1 1 1 1 1 1 1 0 0 0 1 0 1 0 1 1 0 0 1 0 1 1 1 0 1 0 0 0 1 1 1 1 0 0 1 0 0 0 0 1 0 0 0 1 0 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:59 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n534,
    new_n535, new_n536, new_n537, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n547, new_n548, new_n549, new_n550, new_n551, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n566, new_n567, new_n568, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n612, new_n613, new_n616, new_n618, new_n619,
    new_n620, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1139, new_n1140, new_n1142, new_n1143,
    new_n1144, new_n1145;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT64), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT65), .Z(new_n459));
  AOI21_X1  g034(.A(new_n459), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n463), .A2(new_n465), .A3(G125), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n461), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND4_X1  g043(.A1(new_n463), .A2(new_n465), .A3(G137), .A4(new_n461), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n461), .A2(G101), .A3(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n468), .A2(new_n471), .ZN(G160));
  NOR2_X1   g047(.A1(G100), .A2(G2105), .ZN(new_n473));
  XOR2_X1   g048(.A(new_n473), .B(KEYINPUT67), .Z(new_n474));
  OAI21_X1  g049(.A(G2104), .B1(new_n461), .B2(G112), .ZN(new_n475));
  INV_X1    g050(.A(G124), .ZN(new_n476));
  XNOR2_X1  g051(.A(KEYINPUT3), .B(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G2105), .ZN(new_n478));
  OAI22_X1  g053(.A1(new_n474), .A2(new_n475), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n477), .A2(new_n461), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT66), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n480), .B(new_n481), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n479), .B1(new_n482), .B2(G136), .ZN(G162));
  NAND4_X1  g058(.A1(new_n463), .A2(new_n465), .A3(G138), .A4(new_n461), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(KEYINPUT4), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT4), .ZN(new_n486));
  NAND4_X1  g061(.A1(new_n477), .A2(new_n486), .A3(G138), .A4(new_n461), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  NAND4_X1  g063(.A1(new_n463), .A2(new_n465), .A3(G126), .A4(G2105), .ZN(new_n489));
  OR2_X1    g064(.A1(G102), .A2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(G114), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G2105), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n490), .A2(new_n492), .A3(G2104), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n489), .A2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT68), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n489), .A2(KEYINPUT68), .A3(new_n493), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n488), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(G164));
  INV_X1    g074(.A(KEYINPUT5), .ZN(new_n500));
  INV_X1    g075(.A(G543), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n500), .B1(new_n501), .B2(KEYINPUT70), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT70), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n503), .A2(KEYINPUT5), .A3(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G62), .ZN(new_n506));
  NAND2_X1  g081(.A1(G75), .A2(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G651), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G50), .ZN(new_n511));
  INV_X1    g086(.A(G651), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n512), .A2(KEYINPUT6), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT6), .ZN(new_n514));
  OAI21_X1  g089(.A(KEYINPUT69), .B1(new_n514), .B2(G651), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT69), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n516), .A2(new_n512), .A3(KEYINPUT6), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n513), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G543), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n505), .ZN(new_n520));
  INV_X1    g095(.A(G88), .ZN(new_n521));
  OAI22_X1  g096(.A1(new_n511), .A2(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  OR2_X1    g097(.A1(new_n510), .A2(new_n522), .ZN(G303));
  INV_X1    g098(.A(G303), .ZN(G166));
  AND2_X1   g099(.A1(new_n518), .A2(new_n505), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(G89), .ZN(new_n526));
  AOI211_X1 g101(.A(new_n501), .B(new_n513), .C1(new_n515), .C2(new_n517), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G51), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n505), .A2(G63), .A3(G651), .ZN(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n530), .B(KEYINPUT7), .ZN(new_n531));
  NAND4_X1  g106(.A1(new_n526), .A2(new_n528), .A3(new_n529), .A4(new_n531), .ZN(new_n532));
  XOR2_X1   g107(.A(new_n532), .B(KEYINPUT71), .Z(G168));
  AOI22_X1  g108(.A1(new_n505), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n534));
  OR2_X1    g109(.A1(new_n534), .A2(new_n512), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n525), .A2(G90), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n527), .A2(G52), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(G301));
  INV_X1    g113(.A(G301), .ZN(G171));
  AOI22_X1  g114(.A1(new_n505), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n540), .A2(new_n512), .ZN(new_n541));
  XOR2_X1   g116(.A(new_n541), .B(KEYINPUT72), .Z(new_n542));
  AOI22_X1  g117(.A1(new_n525), .A2(G81), .B1(new_n527), .B2(G43), .ZN(new_n543));
  AND2_X1   g118(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G860), .ZN(G153));
  NAND4_X1  g120(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND3_X1  g121(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n547));
  NAND2_X1  g122(.A1(G1), .A2(G3), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(KEYINPUT8), .ZN(new_n549));
  OR2_X1    g124(.A1(new_n548), .A2(KEYINPUT8), .ZN(new_n550));
  AOI21_X1  g125(.A(new_n547), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT73), .ZN(G188));
  INV_X1    g127(.A(G53), .ZN(new_n553));
  OR3_X1    g128(.A1(new_n519), .A2(KEYINPUT9), .A3(new_n553), .ZN(new_n554));
  OAI21_X1  g129(.A(KEYINPUT9), .B1(new_n519), .B2(new_n553), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n505), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n557));
  OR2_X1    g132(.A1(new_n557), .A2(new_n512), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT74), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n525), .A2(new_n559), .A3(G91), .ZN(new_n560));
  INV_X1    g135(.A(G91), .ZN(new_n561));
  OAI21_X1  g136(.A(KEYINPUT74), .B1(new_n520), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n556), .A2(new_n558), .A3(new_n563), .ZN(G299));
  INV_X1    g139(.A(G168), .ZN(G286));
  NAND2_X1  g140(.A1(new_n525), .A2(G87), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n527), .A2(G49), .ZN(new_n567));
  OAI21_X1  g142(.A(G651), .B1(new_n505), .B2(G74), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(G288));
  NAND3_X1  g144(.A1(new_n518), .A2(G48), .A3(G543), .ZN(new_n570));
  AND3_X1   g145(.A1(new_n503), .A2(KEYINPUT5), .A3(G543), .ZN(new_n571));
  AOI21_X1  g146(.A(KEYINPUT5), .B1(new_n503), .B2(G543), .ZN(new_n572));
  OAI21_X1  g147(.A(G61), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(G73), .A2(G543), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n512), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT75), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n570), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n515), .A2(new_n517), .ZN(new_n578));
  INV_X1    g153(.A(new_n513), .ZN(new_n579));
  NAND4_X1  g154(.A1(new_n578), .A2(new_n505), .A3(G86), .A4(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT76), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(G61), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n583), .B1(new_n502), .B2(new_n504), .ZN(new_n584));
  INV_X1    g159(.A(new_n574), .ZN(new_n585));
  OAI211_X1 g160(.A(new_n576), .B(G651), .C1(new_n584), .C2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n582), .A2(new_n586), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n577), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n525), .A2(KEYINPUT76), .A3(G86), .ZN(new_n589));
  AND2_X1   g164(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(G305));
  AOI22_X1  g166(.A1(new_n505), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n592));
  OR2_X1    g167(.A1(new_n592), .A2(KEYINPUT77), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(KEYINPUT77), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n593), .A2(G651), .A3(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT78), .ZN(new_n596));
  OR2_X1    g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n525), .A2(G85), .B1(new_n527), .B2(G47), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n595), .A2(new_n596), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(G290));
  NAND2_X1  g175(.A1(G301), .A2(G868), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n525), .A2(G92), .ZN(new_n602));
  XOR2_X1   g177(.A(KEYINPUT79), .B(KEYINPUT10), .Z(new_n603));
  XNOR2_X1  g178(.A(new_n602), .B(new_n603), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n505), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n605));
  NOR2_X1   g180(.A1(new_n605), .A2(new_n512), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n606), .B1(G54), .B2(new_n527), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n604), .A2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n601), .B1(new_n609), .B2(G868), .ZN(G284));
  OAI21_X1  g185(.A(new_n601), .B1(new_n609), .B2(G868), .ZN(G321));
  INV_X1    g186(.A(G868), .ZN(new_n612));
  NAND2_X1  g187(.A1(G299), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n613), .B1(G168), .B2(new_n612), .ZN(G297));
  OAI21_X1  g189(.A(new_n613), .B1(G168), .B2(new_n612), .ZN(G280));
  INV_X1    g190(.A(G559), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n609), .B1(new_n616), .B2(G860), .ZN(G148));
  NAND2_X1  g192(.A1(new_n609), .A2(new_n616), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT80), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n619), .A2(G868), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n620), .B1(G868), .B2(new_n544), .ZN(G323));
  XNOR2_X1  g196(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g197(.A1(new_n482), .A2(G135), .ZN(new_n623));
  INV_X1    g198(.A(G123), .ZN(new_n624));
  OAI21_X1  g199(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n625));
  NOR2_X1   g200(.A1(new_n461), .A2(G111), .ZN(new_n626));
  OAI221_X1 g201(.A(new_n623), .B1(new_n624), .B2(new_n478), .C1(new_n625), .C2(new_n626), .ZN(new_n627));
  INV_X1    g202(.A(KEYINPUT81), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(G2096), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n461), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(KEYINPUT12), .Z(new_n632));
  XNOR2_X1  g207(.A(KEYINPUT13), .B(G2100), .ZN(new_n633));
  OR2_X1    g208(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n632), .A2(new_n633), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n630), .A2(new_n634), .A3(new_n635), .ZN(G156));
  XNOR2_X1  g211(.A(KEYINPUT15), .B(G2435), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT82), .B(G2438), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(G2427), .B(G2430), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n641), .A2(KEYINPUT14), .ZN(new_n642));
  XOR2_X1   g217(.A(KEYINPUT83), .B(KEYINPUT16), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2451), .B(G2454), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G2443), .B(G2446), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(KEYINPUT84), .B(KEYINPUT85), .Z(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  INV_X1    g226(.A(new_n647), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n646), .B(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n653), .A2(new_n649), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1341), .B(G1348), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n651), .A2(new_n654), .A3(new_n656), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n658), .A2(G14), .A3(new_n659), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(G401));
  XOR2_X1   g236(.A(G2084), .B(G2090), .Z(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(G2067), .B(G2678), .Z(new_n664));
  OR2_X1    g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n663), .A2(new_n664), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n665), .A2(new_n666), .A3(KEYINPUT17), .ZN(new_n667));
  INV_X1    g242(.A(KEYINPUT18), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(G2072), .B(G2078), .Z(new_n670));
  AOI21_X1  g245(.A(new_n670), .B1(new_n665), .B2(KEYINPUT18), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n669), .B(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(G2096), .B(G2100), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT86), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n672), .B(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(G227));
  XNOR2_X1  g251(.A(G1971), .B(G1976), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT19), .ZN(new_n678));
  XOR2_X1   g253(.A(G1956), .B(G2474), .Z(new_n679));
  XOR2_X1   g254(.A(G1961), .B(G1966), .Z(new_n680));
  NAND2_X1  g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(new_n682), .B(KEYINPUT20), .Z(new_n683));
  NOR2_X1   g258(.A1(new_n679), .A2(new_n680), .ZN(new_n684));
  INV_X1    g259(.A(new_n681), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n684), .B1(new_n678), .B2(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(KEYINPUT87), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n678), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n686), .B(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n683), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT88), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1991), .B(G1996), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1981), .B(G1986), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n691), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n696));
  XOR2_X1   g271(.A(new_n695), .B(new_n696), .Z(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(G229));
  NOR2_X1   g273(.A1(G6), .A2(G16), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n699), .B1(new_n590), .B2(G16), .ZN(new_n700));
  XOR2_X1   g275(.A(KEYINPUT32), .B(G1981), .Z(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(G16), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n703), .A2(G22), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(G166), .B2(new_n703), .ZN(new_n705));
  INV_X1    g280(.A(G1971), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  NOR2_X1   g282(.A1(G16), .A2(G23), .ZN(new_n708));
  INV_X1    g283(.A(G288), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n708), .B1(new_n709), .B2(G16), .ZN(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT33), .B(G1976), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  NAND3_X1  g287(.A1(new_n702), .A2(new_n707), .A3(new_n712), .ZN(new_n713));
  OR2_X1    g288(.A1(new_n713), .A2(KEYINPUT34), .ZN(new_n714));
  AOI21_X1  g289(.A(KEYINPUT89), .B1(new_n713), .B2(KEYINPUT34), .ZN(new_n715));
  OR2_X1    g290(.A1(G95), .A2(G2105), .ZN(new_n716));
  OAI211_X1 g291(.A(new_n716), .B(G2104), .C1(G107), .C2(new_n461), .ZN(new_n717));
  INV_X1    g292(.A(G119), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n480), .B(KEYINPUT66), .ZN(new_n719));
  INV_X1    g294(.A(G131), .ZN(new_n720));
  OAI221_X1 g295(.A(new_n717), .B1(new_n718), .B2(new_n478), .C1(new_n719), .C2(new_n720), .ZN(new_n721));
  MUX2_X1   g296(.A(G25), .B(new_n721), .S(G29), .Z(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT35), .B(G1991), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n722), .B(new_n723), .Z(new_n724));
  NOR2_X1   g299(.A1(G16), .A2(G24), .ZN(new_n725));
  INV_X1    g300(.A(G290), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n725), .B1(new_n726), .B2(G16), .ZN(new_n727));
  INV_X1    g302(.A(G1986), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  NAND4_X1  g304(.A1(new_n714), .A2(new_n715), .A3(new_n724), .A4(new_n729), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT36), .ZN(new_n731));
  NAND3_X1  g306(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT26), .Z(new_n733));
  NAND3_X1  g308(.A1(new_n461), .A2(G105), .A3(G2104), .ZN(new_n734));
  INV_X1    g309(.A(G129), .ZN(new_n735));
  OAI211_X1 g310(.A(new_n733), .B(new_n734), .C1(new_n478), .C2(new_n735), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(new_n482), .B2(G141), .ZN(new_n737));
  OR2_X1    g312(.A1(new_n737), .A2(KEYINPUT92), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n737), .A2(KEYINPUT92), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n741), .A2(G29), .ZN(new_n742));
  INV_X1    g317(.A(KEYINPUT93), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(G29), .B2(G32), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(KEYINPUT93), .B2(new_n742), .ZN(new_n746));
  XOR2_X1   g321(.A(KEYINPUT27), .B(G1996), .Z(new_n747));
  XNOR2_X1  g322(.A(new_n746), .B(new_n747), .ZN(new_n748));
  OR2_X1    g323(.A1(G29), .A2(G33), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(KEYINPUT25), .Z(new_n751));
  AOI22_X1  g326(.A1(new_n477), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n752));
  INV_X1    g327(.A(G139), .ZN(new_n753));
  OAI221_X1 g328(.A(new_n751), .B1(new_n461), .B2(new_n752), .C1(new_n719), .C2(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(G29), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n749), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(G2072), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT28), .ZN(new_n759));
  INV_X1    g334(.A(G26), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n759), .B1(new_n760), .B2(G29), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n760), .A2(G29), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n482), .A2(G140), .ZN(new_n763));
  INV_X1    g338(.A(G128), .ZN(new_n764));
  OAI21_X1  g339(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n461), .A2(G116), .ZN(new_n766));
  OAI221_X1 g341(.A(new_n763), .B1(new_n764), .B2(new_n478), .C1(new_n765), .C2(new_n766), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n762), .B1(new_n767), .B2(G29), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n761), .B1(new_n768), .B2(new_n759), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n758), .B1(new_n769), .B2(G2067), .ZN(new_n770));
  OAI211_X1 g345(.A(new_n748), .B(new_n770), .C1(G2067), .C2(new_n769), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n703), .A2(G19), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(new_n544), .B2(new_n703), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n773), .A2(G1341), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n756), .A2(new_n757), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n773), .A2(G1341), .ZN(new_n776));
  NOR2_X1   g351(.A1(G168), .A2(new_n703), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(new_n703), .B2(G21), .ZN(new_n778));
  INV_X1    g353(.A(G1966), .ZN(new_n779));
  OAI211_X1 g354(.A(new_n775), .B(new_n776), .C1(new_n778), .C2(new_n779), .ZN(new_n780));
  NOR3_X1   g355(.A1(new_n771), .A2(new_n774), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n703), .A2(G4), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(new_n609), .B2(new_n703), .ZN(new_n783));
  INV_X1    g358(.A(G1348), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(G299), .A2(G16), .ZN(new_n786));
  NAND3_X1  g361(.A1(new_n703), .A2(KEYINPUT23), .A3(G20), .ZN(new_n787));
  INV_X1    g362(.A(KEYINPUT23), .ZN(new_n788));
  INV_X1    g363(.A(G20), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n788), .B1(new_n789), .B2(G16), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n786), .A2(new_n787), .A3(new_n790), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(G1956), .Z(new_n792));
  INV_X1    g367(.A(G1961), .ZN(new_n793));
  NAND2_X1  g368(.A1(G171), .A2(G16), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(G5), .B2(G16), .ZN(new_n795));
  OAI211_X1 g370(.A(new_n785), .B(new_n792), .C1(new_n793), .C2(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n778), .A2(new_n779), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n795), .A2(new_n793), .ZN(new_n798));
  NOR2_X1   g373(.A1(G164), .A2(new_n755), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n799), .B1(G27), .B2(new_n755), .ZN(new_n800));
  INV_X1    g375(.A(G2078), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n797), .A2(new_n798), .A3(new_n802), .ZN(new_n803));
  NOR2_X1   g378(.A1(G29), .A2(G35), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n804), .B1(G162), .B2(G29), .ZN(new_n805));
  XNOR2_X1  g380(.A(KEYINPUT29), .B(G2090), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  XNOR2_X1  g382(.A(KEYINPUT31), .B(G11), .ZN(new_n808));
  XOR2_X1   g383(.A(KEYINPUT94), .B(KEYINPUT30), .Z(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(G28), .ZN(new_n810));
  OAI221_X1 g385(.A(new_n808), .B1(G29), .B2(new_n810), .C1(new_n800), .C2(new_n801), .ZN(new_n811));
  NOR4_X1   g386(.A1(new_n796), .A2(new_n803), .A3(new_n807), .A4(new_n811), .ZN(new_n812));
  AND3_X1   g387(.A1(new_n731), .A2(new_n781), .A3(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n629), .A2(G29), .ZN(new_n814));
  NAND2_X1  g389(.A1(G160), .A2(G29), .ZN(new_n815));
  XNOR2_X1  g390(.A(KEYINPUT90), .B(KEYINPUT24), .ZN(new_n816));
  XOR2_X1   g391(.A(new_n816), .B(G34), .Z(new_n817));
  OAI21_X1  g392(.A(new_n815), .B1(G29), .B2(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(new_n818), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n819), .A2(G2084), .ZN(new_n820));
  INV_X1    g395(.A(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n819), .A2(G2084), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT91), .ZN(new_n823));
  NAND4_X1  g398(.A1(new_n813), .A2(new_n814), .A3(new_n821), .A4(new_n823), .ZN(G150));
  INV_X1    g399(.A(G150), .ZN(G311));
  XNOR2_X1  g400(.A(KEYINPUT97), .B(G93), .ZN(new_n826));
  XNOR2_X1  g401(.A(KEYINPUT96), .B(G55), .ZN(new_n827));
  AOI22_X1  g402(.A1(new_n525), .A2(new_n826), .B1(new_n527), .B2(new_n827), .ZN(new_n828));
  AOI22_X1  g403(.A1(new_n505), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n829));
  XOR2_X1   g404(.A(new_n829), .B(KEYINPUT95), .Z(new_n830));
  OAI21_X1  g405(.A(new_n828), .B1(new_n830), .B2(new_n512), .ZN(new_n831));
  XNOR2_X1  g406(.A(KEYINPUT98), .B(G860), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n833), .B(KEYINPUT37), .Z(new_n834));
  XNOR2_X1  g409(.A(new_n544), .B(new_n831), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT39), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n609), .A2(G559), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT38), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n836), .B(new_n838), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n834), .B1(new_n839), .B2(new_n832), .ZN(G145));
  INV_X1    g415(.A(G37), .ZN(new_n841));
  OR2_X1    g416(.A1(G106), .A2(G2105), .ZN(new_n842));
  OAI211_X1 g417(.A(new_n842), .B(G2104), .C1(G118), .C2(new_n461), .ZN(new_n843));
  INV_X1    g418(.A(G130), .ZN(new_n844));
  INV_X1    g419(.A(G142), .ZN(new_n845));
  OAI221_X1 g420(.A(new_n843), .B1(new_n844), .B2(new_n478), .C1(new_n719), .C2(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n721), .B(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT99), .ZN(new_n848));
  INV_X1    g423(.A(new_n632), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n848), .B(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n740), .B(new_n767), .ZN(new_n851));
  INV_X1    g426(.A(new_n494), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n488), .A2(new_n852), .ZN(new_n853));
  XOR2_X1   g428(.A(new_n754), .B(new_n853), .Z(new_n854));
  XNOR2_X1  g429(.A(new_n851), .B(new_n854), .ZN(new_n855));
  OR3_X1    g430(.A1(new_n850), .A2(KEYINPUT101), .A3(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(new_n855), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n848), .B(new_n632), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n859), .A2(KEYINPUT101), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n850), .A2(new_n855), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n629), .B(G160), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(G162), .ZN(new_n863));
  NAND4_X1  g438(.A1(new_n856), .A2(new_n860), .A3(new_n861), .A4(new_n863), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n863), .B1(new_n859), .B2(new_n861), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT100), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  AOI211_X1 g442(.A(KEYINPUT100), .B(new_n863), .C1(new_n859), .C2(new_n861), .ZN(new_n868));
  OAI211_X1 g443(.A(new_n841), .B(new_n864), .C1(new_n867), .C2(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g445(.A(KEYINPUT104), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n831), .A2(new_n612), .ZN(new_n872));
  XNOR2_X1  g447(.A(G303), .B(G288), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(new_n590), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(G290), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT103), .ZN(new_n877));
  OR2_X1    g452(.A1(new_n877), .A2(KEYINPUT42), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(KEYINPUT42), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n876), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n875), .A2(new_n877), .A3(KEYINPUT42), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  XOR2_X1   g457(.A(new_n619), .B(new_n835), .Z(new_n883));
  INV_X1    g458(.A(KEYINPUT102), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n884), .B1(new_n609), .B2(G299), .ZN(new_n885));
  XOR2_X1   g460(.A(new_n608), .B(G299), .Z(new_n886));
  AOI21_X1  g461(.A(new_n885), .B1(new_n886), .B2(new_n884), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n883), .A2(new_n887), .ZN(new_n888));
  MUX2_X1   g463(.A(new_n886), .B(new_n887), .S(KEYINPUT41), .Z(new_n889));
  OAI211_X1 g464(.A(new_n882), .B(new_n888), .C1(new_n883), .C2(new_n889), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n888), .B1(new_n883), .B2(new_n889), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n891), .A2(new_n880), .A3(new_n881), .ZN(new_n892));
  AND2_X1   g467(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  OAI211_X1 g468(.A(new_n871), .B(new_n872), .C1(new_n893), .C2(new_n612), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n612), .B1(new_n890), .B2(new_n892), .ZN(new_n895));
  INV_X1    g470(.A(new_n872), .ZN(new_n896));
  OAI21_X1  g471(.A(KEYINPUT104), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n894), .A2(new_n897), .ZN(G295));
  OAI21_X1  g473(.A(new_n872), .B1(new_n893), .B2(new_n612), .ZN(G331));
  XNOR2_X1  g474(.A(G168), .B(G301), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n900), .B(new_n835), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n902), .A2(new_n887), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n903), .B1(new_n889), .B2(new_n902), .ZN(new_n904));
  AOI21_X1  g479(.A(G37), .B1(new_n904), .B2(new_n876), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n901), .A2(KEYINPUT41), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n876), .B1(new_n906), .B2(new_n887), .ZN(new_n907));
  INV_X1    g482(.A(new_n886), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n907), .B1(new_n908), .B2(new_n906), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n905), .A2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT43), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  OAI211_X1 g487(.A(new_n903), .B(new_n875), .C1(new_n889), .C2(new_n902), .ZN(new_n913));
  AOI21_X1  g488(.A(KEYINPUT43), .B1(new_n905), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g489(.A(KEYINPUT44), .B1(new_n912), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n910), .A2(new_n911), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT44), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n905), .A2(KEYINPUT43), .A3(new_n913), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n915), .A2(new_n919), .ZN(G397));
  NOR2_X1   g495(.A1(G290), .A2(G1986), .ZN(new_n921));
  AOI21_X1  g496(.A(G1384), .B1(new_n488), .B2(new_n852), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT45), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(KEYINPUT105), .B1(G160), .B2(G40), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT105), .ZN(new_n927));
  INV_X1    g502(.A(G40), .ZN(new_n928));
  NOR4_X1   g503(.A1(new_n468), .A2(new_n471), .A3(new_n927), .A4(new_n928), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n926), .A2(new_n929), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n925), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n921), .A2(new_n931), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n932), .B(KEYINPUT127), .ZN(new_n933));
  XOR2_X1   g508(.A(new_n933), .B(KEYINPUT48), .Z(new_n934));
  INV_X1    g509(.A(G1996), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n740), .B(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(G2067), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n767), .B(new_n937), .ZN(new_n938));
  AND2_X1   g513(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n721), .A2(new_n723), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n721), .A2(new_n723), .ZN(new_n941));
  INV_X1    g516(.A(new_n941), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n939), .A2(new_n940), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n934), .B1(new_n931), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n931), .A2(new_n935), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT46), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  XOR2_X1   g522(.A(new_n947), .B(KEYINPUT125), .Z(new_n948));
  NOR2_X1   g523(.A1(new_n945), .A2(new_n946), .ZN(new_n949));
  XOR2_X1   g524(.A(new_n949), .B(KEYINPUT126), .Z(new_n950));
  NAND2_X1  g525(.A1(new_n938), .A2(new_n741), .ZN(new_n951));
  AOI211_X1 g526(.A(new_n948), .B(new_n950), .C1(new_n931), .C2(new_n951), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n952), .B(KEYINPUT47), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n939), .A2(new_n941), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n954), .B1(G2067), .B2(new_n767), .ZN(new_n955));
  AOI211_X1 g530(.A(new_n944), .B(new_n953), .C1(new_n931), .C2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT123), .ZN(new_n957));
  OAI22_X1  g532(.A1(new_n926), .A2(new_n929), .B1(new_n922), .B2(KEYINPUT45), .ZN(new_n958));
  INV_X1    g533(.A(G1384), .ZN(new_n959));
  AND3_X1   g534(.A1(new_n498), .A2(KEYINPUT45), .A3(new_n959), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n779), .B1(new_n958), .B2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT110), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  OR2_X1    g538(.A1(new_n923), .A2(KEYINPUT50), .ZN(new_n964));
  NOR3_X1   g539(.A1(new_n468), .A2(new_n471), .A3(new_n928), .ZN(new_n965));
  XNOR2_X1  g540(.A(new_n965), .B(KEYINPUT105), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n498), .A2(new_n959), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(KEYINPUT50), .ZN(new_n968));
  INV_X1    g543(.A(G2084), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n964), .A2(new_n966), .A3(new_n968), .A4(new_n969), .ZN(new_n970));
  OAI211_X1 g545(.A(KEYINPUT110), .B(new_n779), .C1(new_n958), .C2(new_n960), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n963), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(KEYINPUT119), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT119), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n963), .A2(new_n974), .A3(new_n970), .A4(new_n971), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n973), .A2(G168), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(G8), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n973), .A2(KEYINPUT51), .A3(new_n975), .ZN(new_n978));
  INV_X1    g553(.A(G8), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT51), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n972), .A2(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n979), .B1(new_n981), .B2(G168), .ZN(new_n982));
  AOI22_X1  g557(.A1(new_n977), .A2(KEYINPUT51), .B1(new_n978), .B2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT62), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n957), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT52), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n922), .B1(new_n926), .B2(new_n929), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(G8), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT107), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n987), .A2(KEYINPUT107), .A3(G8), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n709), .A2(G1976), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n986), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(G1981), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n588), .A2(KEYINPUT109), .A3(new_n995), .A4(new_n589), .ZN(new_n996));
  AOI22_X1  g571(.A1(new_n575), .A2(new_n576), .B1(new_n581), .B2(new_n580), .ZN(new_n997));
  OAI21_X1  g572(.A(G651), .B1(new_n584), .B2(new_n585), .ZN(new_n998));
  AOI22_X1  g573(.A1(new_n998), .A2(KEYINPUT75), .B1(new_n527), .B2(G48), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n997), .A2(new_n999), .A3(new_n995), .A4(new_n589), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT109), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n996), .A2(new_n1002), .ZN(new_n1003));
  AND2_X1   g578(.A1(new_n570), .A2(new_n580), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n995), .B1(new_n1004), .B2(new_n998), .ZN(new_n1005));
  INV_X1    g580(.A(new_n1005), .ZN(new_n1006));
  AOI21_X1  g581(.A(KEYINPUT49), .B1(new_n1003), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT49), .ZN(new_n1008));
  AOI211_X1 g583(.A(new_n1008), .B(new_n1005), .C1(new_n996), .C2(new_n1002), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n994), .B1(new_n1010), .B2(new_n992), .ZN(new_n1011));
  NAND2_X1  g586(.A1(G303), .A2(G8), .ZN(new_n1012));
  XOR2_X1   g587(.A(new_n1012), .B(KEYINPUT55), .Z(new_n1013));
  INV_X1    g588(.A(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n923), .A2(KEYINPUT50), .ZN(new_n1015));
  OAI211_X1 g590(.A(new_n966), .B(new_n1015), .C1(KEYINPUT50), .C2(new_n967), .ZN(new_n1016));
  AOI21_X1  g591(.A(KEYINPUT45), .B1(new_n498), .B2(new_n959), .ZN(new_n1017));
  AOI211_X1 g592(.A(new_n924), .B(G1384), .C1(new_n488), .C2(new_n852), .ZN(new_n1018));
  NOR3_X1   g593(.A1(new_n930), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1019));
  OAI22_X1  g594(.A1(new_n1016), .A2(G2090), .B1(new_n1019), .B2(G1971), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(G8), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1014), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT106), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1023), .B1(new_n1019), .B2(G1971), .ZN(new_n1024));
  INV_X1    g599(.A(G2090), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n964), .A2(new_n966), .A3(new_n968), .A4(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n967), .A2(new_n924), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1018), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n966), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1029), .A2(KEYINPUT106), .A3(new_n706), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1024), .A2(new_n1026), .A3(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1031), .A2(new_n1013), .A3(G8), .ZN(new_n1032));
  XNOR2_X1  g607(.A(KEYINPUT108), .B(G1976), .ZN(new_n1033));
  AOI21_X1  g608(.A(KEYINPUT52), .B1(G288), .B2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n992), .A2(new_n993), .A3(new_n1034), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n1011), .A2(new_n1022), .A3(new_n1032), .A4(new_n1035), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1036), .B1(new_n983), .B2(new_n984), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT53), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1038), .B1(new_n1029), .B2(G2078), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n964), .A2(new_n966), .A3(new_n968), .ZN(new_n1040));
  XNOR2_X1  g615(.A(KEYINPUT120), .B(G1961), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  OR2_X1    g617(.A1(new_n958), .A2(new_n960), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1038), .A2(G2078), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1044), .ZN(new_n1045));
  OAI211_X1 g620(.A(new_n1039), .B(new_n1042), .C1(new_n1043), .C2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(G171), .ZN(new_n1047));
  XNOR2_X1  g622(.A(new_n1047), .B(KEYINPUT121), .ZN(new_n1048));
  AND2_X1   g623(.A1(new_n982), .A2(new_n978), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n980), .B1(new_n976), .B2(G8), .ZN(new_n1050));
  OAI211_X1 g625(.A(KEYINPUT123), .B(KEYINPUT62), .C1(new_n1049), .C2(new_n1050), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n985), .A2(new_n1037), .A3(new_n1048), .A4(new_n1051), .ZN(new_n1052));
  XNOR2_X1  g627(.A(KEYINPUT112), .B(G1956), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1016), .A2(new_n1053), .ZN(new_n1054));
  XNOR2_X1  g629(.A(KEYINPUT56), .B(G2072), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1019), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1054), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT57), .ZN(new_n1058));
  XNOR2_X1  g633(.A(G299), .B(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1057), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1040), .A2(new_n784), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n966), .A2(new_n937), .A3(new_n922), .ZN(new_n1063));
  AND2_X1   g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1061), .B1(new_n608), .B2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1059), .A2(new_n1054), .A3(new_n1056), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(KEYINPUT113), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT113), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1059), .A2(new_n1054), .A3(new_n1068), .A4(new_n1056), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1065), .A2(new_n1067), .A3(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1067), .A2(new_n1069), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT61), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1061), .A2(KEYINPUT61), .A3(new_n1066), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT60), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1064), .A2(new_n1075), .A3(new_n609), .ZN(new_n1076));
  AND3_X1   g651(.A1(new_n1062), .A2(new_n608), .A3(new_n1063), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n608), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1078));
  OAI21_X1  g653(.A(KEYINPUT60), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1073), .A2(new_n1074), .A3(new_n1076), .A4(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(new_n544), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1081), .A2(KEYINPUT117), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT114), .ZN(new_n1083));
  NOR3_X1   g658(.A1(new_n1029), .A2(new_n1083), .A3(G1996), .ZN(new_n1084));
  AOI21_X1  g659(.A(KEYINPUT114), .B1(new_n1019), .B2(new_n935), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  XOR2_X1   g661(.A(KEYINPUT115), .B(KEYINPUT58), .Z(new_n1087));
  XNOR2_X1  g662(.A(new_n1087), .B(G1341), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n987), .A2(new_n1088), .ZN(new_n1089));
  XNOR2_X1  g664(.A(new_n1089), .B(KEYINPUT116), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1082), .B1(new_n1086), .B2(new_n1090), .ZN(new_n1091));
  XOR2_X1   g666(.A(KEYINPUT118), .B(KEYINPUT59), .Z(new_n1092));
  INV_X1    g667(.A(new_n1092), .ZN(new_n1093));
  XNOR2_X1  g668(.A(new_n1091), .B(new_n1093), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1070), .B1(new_n1080), .B2(new_n1094), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n925), .A2(new_n1028), .A3(new_n965), .A4(new_n1044), .ZN(new_n1096));
  XNOR2_X1  g671(.A(new_n1096), .B(KEYINPUT122), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1097), .A2(new_n1039), .A3(new_n1042), .ZN(new_n1098));
  AND2_X1   g673(.A1(new_n1098), .A2(G171), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT54), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1046), .A2(G171), .ZN(new_n1101));
  NOR3_X1   g676(.A1(new_n1099), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n983), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1036), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1098), .A2(G171), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1100), .B1(new_n1048), .B2(new_n1105), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1095), .A2(new_n1103), .A3(new_n1104), .A4(new_n1106), .ZN(new_n1107));
  AND2_X1   g682(.A1(new_n1011), .A2(new_n1035), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1032), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1003), .A2(new_n1006), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(new_n1008), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1003), .A2(KEYINPUT49), .A3(new_n1006), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1111), .A2(new_n992), .A3(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(G1976), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1113), .A2(new_n1114), .A3(new_n709), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(new_n1003), .ZN(new_n1116));
  AOI22_X1  g691(.A1(new_n1108), .A2(new_n1109), .B1(new_n1116), .B2(new_n992), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n972), .A2(G8), .A3(G168), .ZN(new_n1118));
  OAI21_X1  g693(.A(KEYINPUT111), .B1(new_n1036), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(new_n994), .ZN(new_n1120));
  AND4_X1   g695(.A1(new_n1032), .A2(new_n1120), .A3(new_n1113), .A4(new_n1035), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT111), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1118), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1121), .A2(new_n1122), .A3(new_n1022), .A4(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT63), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1119), .A2(new_n1124), .A3(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1031), .A2(G8), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1125), .B1(new_n1127), .B2(new_n1014), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1121), .A2(new_n1123), .A3(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1126), .A2(new_n1129), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1052), .A2(new_n1107), .A3(new_n1117), .A4(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(new_n943), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1132), .B1(new_n728), .B2(new_n726), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n931), .B1(new_n1133), .B2(new_n921), .ZN(new_n1134));
  AND3_X1   g709(.A1(new_n1131), .A2(KEYINPUT124), .A3(new_n1134), .ZN(new_n1135));
  AOI21_X1  g710(.A(KEYINPUT124), .B1(new_n1131), .B2(new_n1134), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n956), .B1(new_n1135), .B2(new_n1136), .ZN(G329));
  assign    G231 = 1'b0;
  NAND4_X1  g712(.A1(new_n916), .A2(G319), .A3(new_n869), .A4(new_n918), .ZN(new_n1139));
  NAND3_X1  g713(.A1(new_n660), .A2(new_n675), .A3(new_n697), .ZN(new_n1140));
  NOR2_X1   g714(.A1(new_n1139), .A2(new_n1140), .ZN(G308));
  AOI21_X1  g715(.A(KEYINPUT43), .B1(new_n905), .B2(new_n909), .ZN(new_n1142));
  AND2_X1   g716(.A1(new_n905), .A2(new_n913), .ZN(new_n1143));
  AOI21_X1  g717(.A(new_n1142), .B1(KEYINPUT43), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g718(.A(new_n1140), .ZN(new_n1145));
  NAND4_X1  g719(.A1(new_n1144), .A2(new_n1145), .A3(G319), .A4(new_n869), .ZN(G225));
endmodule


