

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586;

  XOR2_X1 U324 ( .A(n309), .B(n308), .Z(n521) );
  XNOR2_X1 U325 ( .A(n457), .B(KEYINPUT96), .ZN(n459) );
  XOR2_X1 U326 ( .A(n295), .B(G134GAT), .Z(n292) );
  INV_X1 U327 ( .A(n469), .ZN(n458) );
  OR2_X1 U328 ( .A1(n459), .A2(n458), .ZN(n460) );
  XNOR2_X1 U329 ( .A(KEYINPUT120), .B(KEYINPUT54), .ZN(n446) );
  XNOR2_X1 U330 ( .A(n447), .B(n446), .ZN(n448) );
  XOR2_X1 U331 ( .A(n555), .B(KEYINPUT36), .Z(n584) );
  NOR2_X1 U332 ( .A1(n530), .A2(n450), .ZN(n565) );
  XOR2_X1 U333 ( .A(KEYINPUT107), .B(n515), .Z(n523) );
  XNOR2_X1 U334 ( .A(n451), .B(G190GAT), .ZN(n452) );
  XNOR2_X1 U335 ( .A(n453), .B(n452), .ZN(G1351GAT) );
  XOR2_X1 U336 ( .A(KEYINPUT0), .B(G127GAT), .Z(n337) );
  XOR2_X1 U337 ( .A(G120GAT), .B(n337), .Z(n294) );
  XOR2_X1 U338 ( .A(G99GAT), .B(G71GAT), .Z(n369) );
  XNOR2_X1 U339 ( .A(G113GAT), .B(n369), .ZN(n293) );
  XNOR2_X1 U340 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U341 ( .A(G176GAT), .B(KEYINPUT84), .Z(n297) );
  XNOR2_X1 U342 ( .A(G169GAT), .B(G15GAT), .ZN(n296) );
  XNOR2_X1 U343 ( .A(n297), .B(n296), .ZN(n298) );
  XNOR2_X1 U344 ( .A(G43GAT), .B(n298), .ZN(n299) );
  XNOR2_X1 U345 ( .A(n292), .B(n299), .ZN(n303) );
  XOR2_X1 U346 ( .A(KEYINPUT20), .B(KEYINPUT82), .Z(n301) );
  NAND2_X1 U347 ( .A1(G227GAT), .A2(G233GAT), .ZN(n300) );
  XNOR2_X1 U348 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U349 ( .A(n303), .B(n302), .Z(n309) );
  XNOR2_X1 U350 ( .A(KEYINPUT81), .B(KEYINPUT18), .ZN(n304) );
  XNOR2_X1 U351 ( .A(n304), .B(KEYINPUT17), .ZN(n305) );
  XOR2_X1 U352 ( .A(n305), .B(KEYINPUT19), .Z(n307) );
  XNOR2_X1 U353 ( .A(G183GAT), .B(G190GAT), .ZN(n306) );
  XNOR2_X1 U354 ( .A(n307), .B(n306), .ZN(n354) );
  XNOR2_X1 U355 ( .A(n354), .B(KEYINPUT83), .ZN(n308) );
  INV_X1 U356 ( .A(n521), .ZN(n530) );
  XOR2_X1 U357 ( .A(KEYINPUT88), .B(KEYINPUT87), .Z(n311) );
  XNOR2_X1 U358 ( .A(KEYINPUT23), .B(KEYINPUT22), .ZN(n310) );
  XNOR2_X1 U359 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U360 ( .A(n312), .B(G148GAT), .Z(n314) );
  XOR2_X1 U361 ( .A(G141GAT), .B(G22GAT), .Z(n421) );
  XNOR2_X1 U362 ( .A(G50GAT), .B(n421), .ZN(n313) );
  XNOR2_X1 U363 ( .A(n314), .B(n313), .ZN(n320) );
  XOR2_X1 U364 ( .A(G155GAT), .B(KEYINPUT2), .Z(n316) );
  XNOR2_X1 U365 ( .A(G162GAT), .B(KEYINPUT3), .ZN(n315) );
  XNOR2_X1 U366 ( .A(n316), .B(n315), .ZN(n334) );
  XOR2_X1 U367 ( .A(G106GAT), .B(G78GAT), .Z(n368) );
  XOR2_X1 U368 ( .A(n334), .B(n368), .Z(n318) );
  NAND2_X1 U369 ( .A1(G228GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U370 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U371 ( .A(n320), .B(n319), .Z(n328) );
  XOR2_X1 U372 ( .A(KEYINPUT86), .B(G218GAT), .Z(n322) );
  XNOR2_X1 U373 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n321) );
  XNOR2_X1 U374 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U375 ( .A(G197GAT), .B(n323), .Z(n353) );
  XOR2_X1 U376 ( .A(G204GAT), .B(KEYINPUT85), .Z(n325) );
  XNOR2_X1 U377 ( .A(KEYINPUT89), .B(KEYINPUT24), .ZN(n324) );
  XNOR2_X1 U378 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U379 ( .A(n353), .B(n326), .ZN(n327) );
  XNOR2_X1 U380 ( .A(n328), .B(n327), .ZN(n469) );
  XOR2_X1 U381 ( .A(KEYINPUT90), .B(KEYINPUT92), .Z(n330) );
  NAND2_X1 U382 ( .A1(G225GAT), .A2(G233GAT), .ZN(n329) );
  XNOR2_X1 U383 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U384 ( .A(n331), .B(KEYINPUT5), .Z(n336) );
  XOR2_X1 U385 ( .A(G57GAT), .B(G85GAT), .Z(n333) );
  XNOR2_X1 U386 ( .A(G120GAT), .B(G148GAT), .ZN(n332) );
  XNOR2_X1 U387 ( .A(n333), .B(n332), .ZN(n361) );
  XNOR2_X1 U388 ( .A(n334), .B(n361), .ZN(n335) );
  XNOR2_X1 U389 ( .A(n336), .B(n335), .ZN(n341) );
  XOR2_X1 U390 ( .A(G134GAT), .B(KEYINPUT77), .Z(n391) );
  XOR2_X1 U391 ( .A(n337), .B(n391), .Z(n339) );
  XNOR2_X1 U392 ( .A(G29GAT), .B(G141GAT), .ZN(n338) );
  XNOR2_X1 U393 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U394 ( .A(n341), .B(n340), .Z(n346) );
  XOR2_X1 U395 ( .A(G113GAT), .B(G1GAT), .Z(n424) );
  XOR2_X1 U396 ( .A(KEYINPUT91), .B(KEYINPUT1), .Z(n343) );
  XNOR2_X1 U397 ( .A(KEYINPUT4), .B(KEYINPUT6), .ZN(n342) );
  XNOR2_X1 U398 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U399 ( .A(n424), .B(n344), .ZN(n345) );
  XNOR2_X1 U400 ( .A(n346), .B(n345), .ZN(n465) );
  XNOR2_X1 U401 ( .A(KEYINPUT93), .B(n465), .ZN(n468) );
  INV_X1 U402 ( .A(n468), .ZN(n516) );
  XNOR2_X1 U403 ( .A(G169GAT), .B(G36GAT), .ZN(n347) );
  XNOR2_X1 U404 ( .A(n347), .B(G8GAT), .ZN(n420) );
  XOR2_X1 U405 ( .A(KEYINPUT94), .B(n420), .Z(n349) );
  NAND2_X1 U406 ( .A1(G226GAT), .A2(G233GAT), .ZN(n348) );
  XNOR2_X1 U407 ( .A(n349), .B(n348), .ZN(n352) );
  XOR2_X1 U408 ( .A(G64GAT), .B(G92GAT), .Z(n351) );
  XNOR2_X1 U409 ( .A(G176GAT), .B(G204GAT), .ZN(n350) );
  XNOR2_X1 U410 ( .A(n351), .B(n350), .ZN(n360) );
  XOR2_X1 U411 ( .A(n352), .B(n360), .Z(n356) );
  XNOR2_X1 U412 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U413 ( .A(n356), .B(n355), .Z(n518) );
  XOR2_X1 U414 ( .A(KEYINPUT119), .B(n518), .Z(n445) );
  XOR2_X1 U415 ( .A(KEYINPUT31), .B(KEYINPUT32), .Z(n358) );
  NAND2_X1 U416 ( .A1(G230GAT), .A2(G233GAT), .ZN(n357) );
  XNOR2_X1 U417 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U418 ( .A(n359), .B(KEYINPUT13), .Z(n363) );
  XNOR2_X1 U419 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U420 ( .A(n363), .B(n362), .ZN(n367) );
  XOR2_X1 U421 ( .A(KEYINPUT73), .B(KEYINPUT33), .Z(n365) );
  XNOR2_X1 U422 ( .A(KEYINPUT71), .B(KEYINPUT72), .ZN(n364) );
  XNOR2_X1 U423 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U424 ( .A(n367), .B(n366), .Z(n371) );
  XNOR2_X1 U425 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U426 ( .A(n371), .B(n370), .Z(n454) );
  INV_X1 U427 ( .A(n454), .ZN(n574) );
  XOR2_X1 U428 ( .A(G78GAT), .B(G155GAT), .Z(n373) );
  XNOR2_X1 U429 ( .A(G22GAT), .B(G211GAT), .ZN(n372) );
  XNOR2_X1 U430 ( .A(n373), .B(n372), .ZN(n377) );
  XOR2_X1 U431 ( .A(G127GAT), .B(G71GAT), .Z(n375) );
  XNOR2_X1 U432 ( .A(G15GAT), .B(G183GAT), .ZN(n374) );
  XNOR2_X1 U433 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U434 ( .A(n377), .B(n376), .Z(n382) );
  XOR2_X1 U435 ( .A(KEYINPUT79), .B(KEYINPUT80), .Z(n379) );
  NAND2_X1 U436 ( .A1(G231GAT), .A2(G233GAT), .ZN(n378) );
  XNOR2_X1 U437 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U438 ( .A(KEYINPUT78), .B(n380), .ZN(n381) );
  XNOR2_X1 U439 ( .A(n382), .B(n381), .ZN(n390) );
  XOR2_X1 U440 ( .A(G64GAT), .B(G57GAT), .Z(n384) );
  XNOR2_X1 U441 ( .A(G1GAT), .B(G8GAT), .ZN(n383) );
  XNOR2_X1 U442 ( .A(n384), .B(n383), .ZN(n388) );
  XOR2_X1 U443 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n386) );
  XNOR2_X1 U444 ( .A(KEYINPUT13), .B(KEYINPUT12), .ZN(n385) );
  XNOR2_X1 U445 ( .A(n386), .B(n385), .ZN(n387) );
  XOR2_X1 U446 ( .A(n388), .B(n387), .Z(n389) );
  XOR2_X1 U447 ( .A(n390), .B(n389), .Z(n579) );
  INV_X1 U448 ( .A(n579), .ZN(n485) );
  XOR2_X1 U449 ( .A(KEYINPUT10), .B(n391), .Z(n393) );
  XNOR2_X1 U450 ( .A(G190GAT), .B(G218GAT), .ZN(n392) );
  XNOR2_X1 U451 ( .A(n393), .B(n392), .ZN(n412) );
  XOR2_X1 U452 ( .A(G92GAT), .B(KEYINPUT11), .Z(n395) );
  XNOR2_X1 U453 ( .A(G85GAT), .B(KEYINPUT66), .ZN(n394) );
  XNOR2_X1 U454 ( .A(n395), .B(n394), .ZN(n399) );
  XOR2_X1 U455 ( .A(KEYINPUT75), .B(G106GAT), .Z(n397) );
  XNOR2_X1 U456 ( .A(G99GAT), .B(G162GAT), .ZN(n396) );
  XNOR2_X1 U457 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U458 ( .A(n399), .B(n398), .Z(n408) );
  XNOR2_X1 U459 ( .A(G50GAT), .B(G43GAT), .ZN(n401) );
  XNOR2_X1 U460 ( .A(KEYINPUT7), .B(KEYINPUT68), .ZN(n400) );
  XNOR2_X1 U461 ( .A(n401), .B(n400), .ZN(n403) );
  XOR2_X1 U462 ( .A(KEYINPUT8), .B(G29GAT), .Z(n402) );
  XNOR2_X1 U463 ( .A(n403), .B(n402), .ZN(n430) );
  XOR2_X1 U464 ( .A(KEYINPUT9), .B(KEYINPUT76), .Z(n405) );
  XNOR2_X1 U465 ( .A(G36GAT), .B(KEYINPUT65), .ZN(n404) );
  XNOR2_X1 U466 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U467 ( .A(n430), .B(n406), .ZN(n407) );
  NAND2_X1 U468 ( .A1(n408), .A2(n407), .ZN(n410) );
  OR2_X1 U469 ( .A1(n408), .A2(n407), .ZN(n409) );
  NAND2_X1 U470 ( .A1(n410), .A2(n409), .ZN(n411) );
  XNOR2_X1 U471 ( .A(n412), .B(n411), .ZN(n414) );
  NAND2_X1 U472 ( .A1(G232GAT), .A2(G233GAT), .ZN(n413) );
  XNOR2_X2 U473 ( .A(n414), .B(n413), .ZN(n555) );
  NOR2_X1 U474 ( .A1(n485), .A2(n584), .ZN(n415) );
  XOR2_X1 U475 ( .A(n415), .B(KEYINPUT45), .Z(n416) );
  NOR2_X1 U476 ( .A1(n574), .A2(n416), .ZN(n417) );
  XNOR2_X1 U477 ( .A(n417), .B(KEYINPUT111), .ZN(n432) );
  XOR2_X1 U478 ( .A(KEYINPUT67), .B(KEYINPUT69), .Z(n419) );
  XNOR2_X1 U479 ( .A(KEYINPUT29), .B(KEYINPUT30), .ZN(n418) );
  XNOR2_X1 U480 ( .A(n419), .B(n418), .ZN(n429) );
  XOR2_X1 U481 ( .A(n421), .B(n420), .Z(n423) );
  NAND2_X1 U482 ( .A1(G229GAT), .A2(G233GAT), .ZN(n422) );
  XNOR2_X1 U483 ( .A(n423), .B(n422), .ZN(n425) );
  XOR2_X1 U484 ( .A(n425), .B(n424), .Z(n427) );
  XNOR2_X1 U485 ( .A(G197GAT), .B(G15GAT), .ZN(n426) );
  XNOR2_X1 U486 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U487 ( .A(n429), .B(n428), .Z(n431) );
  XNOR2_X1 U488 ( .A(n431), .B(n430), .ZN(n569) );
  INV_X1 U489 ( .A(n569), .ZN(n502) );
  XOR2_X1 U490 ( .A(KEYINPUT70), .B(n502), .Z(n557) );
  NOR2_X1 U491 ( .A1(n432), .A2(n557), .ZN(n434) );
  INV_X1 U492 ( .A(KEYINPUT112), .ZN(n433) );
  XNOR2_X1 U493 ( .A(n434), .B(n433), .ZN(n442) );
  XNOR2_X1 U494 ( .A(KEYINPUT41), .B(n454), .ZN(n549) );
  NAND2_X1 U495 ( .A1(n569), .A2(n549), .ZN(n435) );
  XNOR2_X1 U496 ( .A(n435), .B(KEYINPUT46), .ZN(n436) );
  XNOR2_X1 U497 ( .A(KEYINPUT110), .B(n436), .ZN(n438) );
  INV_X1 U498 ( .A(n555), .ZN(n437) );
  NAND2_X1 U499 ( .A1(n438), .A2(n437), .ZN(n439) );
  NOR2_X1 U500 ( .A1(n579), .A2(n439), .ZN(n440) );
  XNOR2_X1 U501 ( .A(KEYINPUT47), .B(n440), .ZN(n441) );
  NAND2_X1 U502 ( .A1(n442), .A2(n441), .ZN(n444) );
  XNOR2_X1 U503 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n443) );
  XNOR2_X1 U504 ( .A(n444), .B(n443), .ZN(n528) );
  NAND2_X1 U505 ( .A1(n445), .A2(n528), .ZN(n447) );
  NOR2_X1 U506 ( .A1(n516), .A2(n448), .ZN(n568) );
  AND2_X1 U507 ( .A1(n469), .A2(n568), .ZN(n449) );
  XNOR2_X1 U508 ( .A(n449), .B(KEYINPUT55), .ZN(n450) );
  NAND2_X1 U509 ( .A1(n565), .A2(n555), .ZN(n453) );
  XOR2_X1 U510 ( .A(KEYINPUT123), .B(KEYINPUT58), .Z(n451) );
  NAND2_X1 U511 ( .A1(n454), .A2(n557), .ZN(n455) );
  XNOR2_X1 U512 ( .A(n455), .B(KEYINPUT74), .ZN(n489) );
  NOR2_X1 U513 ( .A1(n555), .A2(n485), .ZN(n456) );
  XNOR2_X1 U514 ( .A(n456), .B(KEYINPUT16), .ZN(n474) );
  AND2_X1 U515 ( .A1(n521), .A2(n518), .ZN(n457) );
  XNOR2_X1 U516 ( .A(n460), .B(KEYINPUT25), .ZN(n463) );
  XOR2_X1 U517 ( .A(n518), .B(KEYINPUT27), .Z(n467) );
  NOR2_X1 U518 ( .A1(n521), .A2(n469), .ZN(n461) );
  XNOR2_X1 U519 ( .A(n461), .B(KEYINPUT26), .ZN(n567) );
  INV_X1 U520 ( .A(n567), .ZN(n547) );
  NOR2_X1 U521 ( .A1(n467), .A2(n547), .ZN(n462) );
  NOR2_X1 U522 ( .A1(n463), .A2(n462), .ZN(n464) );
  NOR2_X1 U523 ( .A1(n465), .A2(n464), .ZN(n466) );
  XNOR2_X1 U524 ( .A(n466), .B(KEYINPUT97), .ZN(n473) );
  NOR2_X1 U525 ( .A1(n468), .A2(n467), .ZN(n527) );
  XNOR2_X1 U526 ( .A(n469), .B(KEYINPUT28), .ZN(n482) );
  NAND2_X1 U527 ( .A1(n527), .A2(n482), .ZN(n470) );
  XNOR2_X1 U528 ( .A(KEYINPUT95), .B(n470), .ZN(n471) );
  NAND2_X1 U529 ( .A1(n471), .A2(n530), .ZN(n472) );
  NAND2_X1 U530 ( .A1(n473), .A2(n472), .ZN(n486) );
  NAND2_X1 U531 ( .A1(n474), .A2(n486), .ZN(n503) );
  NOR2_X1 U532 ( .A1(n489), .A2(n503), .ZN(n475) );
  XNOR2_X1 U533 ( .A(KEYINPUT98), .B(n475), .ZN(n483) );
  NAND2_X1 U534 ( .A1(n483), .A2(n516), .ZN(n476) );
  XNOR2_X1 U535 ( .A(n476), .B(KEYINPUT34), .ZN(n477) );
  XNOR2_X1 U536 ( .A(G1GAT), .B(n477), .ZN(G1324GAT) );
  NAND2_X1 U537 ( .A1(n483), .A2(n518), .ZN(n478) );
  XNOR2_X1 U538 ( .A(n478), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U539 ( .A(KEYINPUT35), .B(KEYINPUT99), .Z(n480) );
  NAND2_X1 U540 ( .A1(n483), .A2(n521), .ZN(n479) );
  XNOR2_X1 U541 ( .A(n480), .B(n479), .ZN(n481) );
  XOR2_X1 U542 ( .A(G15GAT), .B(n481), .Z(G1326GAT) );
  INV_X1 U543 ( .A(n482), .ZN(n533) );
  NAND2_X1 U544 ( .A1(n483), .A2(n533), .ZN(n484) );
  XNOR2_X1 U545 ( .A(n484), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U546 ( .A(G29GAT), .B(KEYINPUT39), .Z(n492) );
  NAND2_X1 U547 ( .A1(n486), .A2(n485), .ZN(n487) );
  NOR2_X1 U548 ( .A1(n584), .A2(n487), .ZN(n488) );
  XNOR2_X1 U549 ( .A(KEYINPUT37), .B(n488), .ZN(n514) );
  NOR2_X1 U550 ( .A1(n514), .A2(n489), .ZN(n490) );
  XNOR2_X1 U551 ( .A(n490), .B(KEYINPUT38), .ZN(n497) );
  NAND2_X1 U552 ( .A1(n516), .A2(n497), .ZN(n491) );
  XNOR2_X1 U553 ( .A(n492), .B(n491), .ZN(G1328GAT) );
  NAND2_X1 U554 ( .A1(n497), .A2(n518), .ZN(n493) );
  XNOR2_X1 U555 ( .A(n493), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U556 ( .A(KEYINPUT100), .B(KEYINPUT40), .Z(n495) );
  NAND2_X1 U557 ( .A1(n497), .A2(n521), .ZN(n494) );
  XNOR2_X1 U558 ( .A(n495), .B(n494), .ZN(n496) );
  XOR2_X1 U559 ( .A(G43GAT), .B(n496), .Z(G1330GAT) );
  XOR2_X1 U560 ( .A(G50GAT), .B(KEYINPUT101), .Z(n499) );
  NAND2_X1 U561 ( .A1(n533), .A2(n497), .ZN(n498) );
  XNOR2_X1 U562 ( .A(n499), .B(n498), .ZN(G1331GAT) );
  XNOR2_X1 U563 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n500) );
  XNOR2_X1 U564 ( .A(n500), .B(KEYINPUT103), .ZN(n501) );
  XOR2_X1 U565 ( .A(KEYINPUT104), .B(n501), .Z(n505) );
  XNOR2_X1 U566 ( .A(n549), .B(KEYINPUT102), .ZN(n560) );
  NAND2_X1 U567 ( .A1(n502), .A2(n560), .ZN(n513) );
  NOR2_X1 U568 ( .A1(n513), .A2(n503), .ZN(n509) );
  NAND2_X1 U569 ( .A1(n509), .A2(n516), .ZN(n504) );
  XNOR2_X1 U570 ( .A(n505), .B(n504), .ZN(G1332GAT) );
  XOR2_X1 U571 ( .A(G64GAT), .B(KEYINPUT105), .Z(n507) );
  NAND2_X1 U572 ( .A1(n509), .A2(n518), .ZN(n506) );
  XNOR2_X1 U573 ( .A(n507), .B(n506), .ZN(G1333GAT) );
  NAND2_X1 U574 ( .A1(n521), .A2(n509), .ZN(n508) );
  XNOR2_X1 U575 ( .A(n508), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U576 ( .A(KEYINPUT106), .B(KEYINPUT43), .Z(n511) );
  NAND2_X1 U577 ( .A1(n509), .A2(n533), .ZN(n510) );
  XNOR2_X1 U578 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U579 ( .A(G78GAT), .B(n512), .ZN(G1335GAT) );
  NOR2_X1 U580 ( .A1(n514), .A2(n513), .ZN(n515) );
  NAND2_X1 U581 ( .A1(n516), .A2(n523), .ZN(n517) );
  XNOR2_X1 U582 ( .A(G85GAT), .B(n517), .ZN(G1336GAT) );
  NAND2_X1 U583 ( .A1(n518), .A2(n523), .ZN(n519) );
  XNOR2_X1 U584 ( .A(n519), .B(KEYINPUT108), .ZN(n520) );
  XNOR2_X1 U585 ( .A(G92GAT), .B(n520), .ZN(G1337GAT) );
  NAND2_X1 U586 ( .A1(n521), .A2(n523), .ZN(n522) );
  XNOR2_X1 U587 ( .A(n522), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U588 ( .A(KEYINPUT44), .B(KEYINPUT109), .Z(n525) );
  NAND2_X1 U589 ( .A1(n523), .A2(n533), .ZN(n524) );
  XNOR2_X1 U590 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U591 ( .A(G106GAT), .B(n526), .ZN(G1339GAT) );
  XOR2_X1 U592 ( .A(G113GAT), .B(KEYINPUT115), .Z(n535) );
  NAND2_X1 U593 ( .A1(n528), .A2(n527), .ZN(n529) );
  XOR2_X1 U594 ( .A(KEYINPUT113), .B(n529), .Z(n546) );
  NOR2_X1 U595 ( .A1(n530), .A2(n546), .ZN(n531) );
  XOR2_X1 U596 ( .A(KEYINPUT114), .B(n531), .Z(n532) );
  NOR2_X1 U597 ( .A1(n533), .A2(n532), .ZN(n542) );
  NAND2_X1 U598 ( .A1(n542), .A2(n557), .ZN(n534) );
  XNOR2_X1 U599 ( .A(n535), .B(n534), .ZN(G1340GAT) );
  XOR2_X1 U600 ( .A(G120GAT), .B(KEYINPUT49), .Z(n537) );
  NAND2_X1 U601 ( .A1(n542), .A2(n560), .ZN(n536) );
  XNOR2_X1 U602 ( .A(n537), .B(n536), .ZN(G1341GAT) );
  XNOR2_X1 U603 ( .A(G127GAT), .B(KEYINPUT116), .ZN(n541) );
  XOR2_X1 U604 ( .A(KEYINPUT117), .B(KEYINPUT50), .Z(n539) );
  NAND2_X1 U605 ( .A1(n542), .A2(n579), .ZN(n538) );
  XNOR2_X1 U606 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U607 ( .A(n541), .B(n540), .ZN(G1342GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT118), .B(KEYINPUT51), .Z(n544) );
  NAND2_X1 U609 ( .A1(n542), .A2(n555), .ZN(n543) );
  XNOR2_X1 U610 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U611 ( .A(G134GAT), .B(n545), .ZN(G1343GAT) );
  NOR2_X1 U612 ( .A1(n547), .A2(n546), .ZN(n554) );
  NAND2_X1 U613 ( .A1(n554), .A2(n569), .ZN(n548) );
  XNOR2_X1 U614 ( .A(G141GAT), .B(n548), .ZN(G1344GAT) );
  XOR2_X1 U615 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n551) );
  NAND2_X1 U616 ( .A1(n554), .A2(n549), .ZN(n550) );
  XNOR2_X1 U617 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U618 ( .A(G148GAT), .B(n552), .ZN(G1345GAT) );
  NAND2_X1 U619 ( .A1(n554), .A2(n579), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n553), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U621 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U622 ( .A(n556), .B(G162GAT), .ZN(G1347GAT) );
  XOR2_X1 U623 ( .A(G169GAT), .B(KEYINPUT121), .Z(n559) );
  NAND2_X1 U624 ( .A1(n565), .A2(n557), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n559), .B(n558), .ZN(G1348GAT) );
  NAND2_X1 U626 ( .A1(n565), .A2(n560), .ZN(n562) );
  XOR2_X1 U627 ( .A(G176GAT), .B(KEYINPUT56), .Z(n561) );
  XNOR2_X1 U628 ( .A(n562), .B(n561), .ZN(n564) );
  XNOR2_X1 U629 ( .A(KEYINPUT57), .B(KEYINPUT122), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n564), .B(n563), .ZN(G1349GAT) );
  NAND2_X1 U631 ( .A1(n565), .A2(n579), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n566), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U633 ( .A1(n568), .A2(n567), .ZN(n583) );
  INV_X1 U634 ( .A(n583), .ZN(n580) );
  NAND2_X1 U635 ( .A1(n569), .A2(n580), .ZN(n573) );
  XOR2_X1 U636 ( .A(KEYINPUT59), .B(KEYINPUT124), .Z(n571) );
  XNOR2_X1 U637 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n570) );
  XNOR2_X1 U638 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n573), .B(n572), .ZN(G1352GAT) );
  XOR2_X1 U640 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n576) );
  NAND2_X1 U641 ( .A1(n580), .A2(n574), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n576), .B(n575), .ZN(n578) );
  XOR2_X1 U643 ( .A(G204GAT), .B(KEYINPUT125), .Z(n577) );
  XNOR2_X1 U644 ( .A(n578), .B(n577), .ZN(G1353GAT) );
  XOR2_X1 U645 ( .A(G211GAT), .B(KEYINPUT127), .Z(n582) );
  NAND2_X1 U646 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(G1354GAT) );
  NOR2_X1 U648 ( .A1(n584), .A2(n583), .ZN(n585) );
  XOR2_X1 U649 ( .A(KEYINPUT62), .B(n585), .Z(n586) );
  XNOR2_X1 U650 ( .A(G218GAT), .B(n586), .ZN(G1355GAT) );
endmodule

