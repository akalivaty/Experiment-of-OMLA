//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 0 0 1 1 0 0 1 1 0 0 1 1 0 0 1 0 0 0 1 0 1 0 1 1 1 1 1 1 0 1 1 0 0 0 1 1 0 0 0 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:26 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n739, new_n740, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n794, new_n795, new_n797, new_n798,
    new_n799, new_n801, new_n802, new_n803, new_n805, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n836, new_n837, new_n838,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n905, new_n906, new_n908, new_n909, new_n911, new_n912, new_n913,
    new_n914, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n997, new_n998, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1014, new_n1015,
    new_n1016, new_n1018, new_n1019, new_n1020, new_n1021, new_n1023,
    new_n1024, new_n1025, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1049, new_n1050, new_n1051;
  INV_X1    g000(.A(KEYINPUT12), .ZN(new_n202));
  XNOR2_X1  g001(.A(G113gat), .B(G141gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(G169gat), .B(G197gat), .ZN(new_n204));
  OR2_X1    g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(KEYINPUT89), .B(KEYINPUT11), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n203), .A2(new_n204), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n205), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  AOI21_X1  g008(.A(new_n206), .B1(new_n205), .B2(new_n207), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n202), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(new_n210), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n212), .A2(KEYINPUT12), .A3(new_n208), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT90), .ZN(new_n215));
  XNOR2_X1  g014(.A(new_n214), .B(new_n215), .ZN(new_n216));
  XOR2_X1   g015(.A(G43gat), .B(G50gat), .Z(new_n217));
  INV_X1    g016(.A(KEYINPUT15), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(G29gat), .ZN(new_n220));
  INV_X1    g019(.A(G36gat), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n220), .A2(new_n221), .A3(KEYINPUT14), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT14), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n223), .B1(G29gat), .B2(G36gat), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n222), .A2(new_n224), .A3(KEYINPUT91), .ZN(new_n225));
  NAND2_X1  g024(.A1(G29gat), .A2(G36gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  AOI21_X1  g026(.A(KEYINPUT91), .B1(new_n222), .B2(new_n224), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n219), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  OR2_X1    g028(.A1(G43gat), .A2(G50gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(G43gat), .A2(G50gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  AOI22_X1  g031(.A1(new_n232), .A2(KEYINPUT15), .B1(G29gat), .B2(G36gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n222), .A2(new_n224), .ZN(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n217), .A2(new_n218), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n233), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n229), .A2(new_n237), .A3(KEYINPUT17), .ZN(new_n238));
  INV_X1    g037(.A(G1gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(KEYINPUT16), .ZN(new_n240));
  INV_X1    g039(.A(G15gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(G22gat), .ZN(new_n242));
  INV_X1    g041(.A(G22gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(G15gat), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n240), .A2(new_n242), .A3(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  AOI21_X1  g045(.A(G1gat), .B1(new_n242), .B2(new_n244), .ZN(new_n247));
  OAI21_X1  g046(.A(G8gat), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n247), .ZN(new_n249));
  INV_X1    g048(.A(G8gat), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n249), .A2(new_n245), .A3(new_n250), .ZN(new_n251));
  AND2_X1   g050(.A1(new_n248), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT91), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n234), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n254), .A2(new_n225), .A3(new_n226), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n234), .B1(new_n218), .B2(new_n217), .ZN(new_n256));
  AOI22_X1  g055(.A1(new_n255), .A2(new_n219), .B1(new_n256), .B2(new_n233), .ZN(new_n257));
  XNOR2_X1  g056(.A(KEYINPUT92), .B(KEYINPUT17), .ZN(new_n258));
  OAI211_X1 g057(.A(new_n238), .B(new_n252), .C1(new_n257), .C2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(G229gat), .A2(G233gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n229), .A2(new_n237), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n248), .A2(new_n251), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n259), .A2(new_n260), .A3(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT18), .ZN(new_n265));
  AND2_X1   g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND4_X1  g065(.A1(new_n259), .A2(KEYINPUT18), .A3(new_n260), .A4(new_n263), .ZN(new_n267));
  XOR2_X1   g066(.A(new_n260), .B(KEYINPUT13), .Z(new_n268));
  INV_X1    g067(.A(new_n263), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n261), .A2(new_n262), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n268), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n267), .A2(new_n271), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n216), .B1(new_n266), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n264), .A2(new_n265), .ZN(new_n274));
  AND2_X1   g073(.A1(new_n211), .A2(new_n213), .ZN(new_n275));
  NAND4_X1  g074(.A1(new_n274), .A2(new_n271), .A3(new_n267), .A4(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n273), .A2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(G211gat), .B(G218gat), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(G218gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(KEYINPUT72), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT72), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(G218gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  AOI21_X1  g084(.A(KEYINPUT22), .B1(new_n285), .B2(G211gat), .ZN(new_n286));
  XOR2_X1   g085(.A(G197gat), .B(G204gat), .Z(new_n287));
  OAI21_X1  g086(.A(new_n280), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n287), .ZN(new_n289));
  XNOR2_X1  g088(.A(KEYINPUT72), .B(G218gat), .ZN(new_n290));
  INV_X1    g089(.A(G211gat), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  OAI211_X1 g091(.A(new_n279), .B(new_n289), .C1(new_n292), .C2(KEYINPUT22), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n288), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(G226gat), .ZN(new_n296));
  INV_X1    g095(.A(G233gat), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT25), .ZN(new_n299));
  NOR2_X1   g098(.A1(G169gat), .A2(G176gat), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT23), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  OAI21_X1  g101(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(G169gat), .A2(G176gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(KEYINPUT64), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT64), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n307), .A2(G169gat), .A3(G176gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n304), .A2(new_n309), .ZN(new_n310));
  NOR2_X1   g109(.A1(G183gat), .A2(G190gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(G183gat), .A2(G190gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(KEYINPUT24), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT24), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n314), .A2(G183gat), .A3(G190gat), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n311), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n299), .B1(new_n310), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n313), .A2(new_n315), .ZN(new_n318));
  XNOR2_X1  g117(.A(KEYINPUT65), .B(G190gat), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n318), .B1(new_n319), .B2(G183gat), .ZN(new_n320));
  AOI22_X1  g119(.A1(new_n303), .A2(new_n302), .B1(new_n306), .B2(new_n308), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n320), .A2(KEYINPUT25), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n317), .A2(new_n322), .ZN(new_n323));
  OAI21_X1  g122(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT26), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n300), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n309), .A2(new_n324), .A3(new_n326), .ZN(new_n327));
  XOR2_X1   g126(.A(KEYINPUT65), .B(G190gat), .Z(new_n328));
  XNOR2_X1  g127(.A(KEYINPUT27), .B(G183gat), .ZN(new_n329));
  AND3_X1   g128(.A1(new_n328), .A2(KEYINPUT28), .A3(new_n329), .ZN(new_n330));
  AOI21_X1  g129(.A(KEYINPUT28), .B1(new_n328), .B2(new_n329), .ZN(new_n331));
  OAI211_X1 g130(.A(new_n312), .B(new_n327), .C1(new_n330), .C2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n323), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT29), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n298), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT28), .ZN(new_n336));
  INV_X1    g135(.A(new_n329), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n336), .B1(new_n337), .B2(new_n319), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n328), .A2(KEYINPUT28), .A3(new_n329), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n327), .A2(new_n312), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  AOI22_X1  g141(.A1(new_n340), .A2(new_n342), .B1(new_n317), .B2(new_n322), .ZN(new_n343));
  INV_X1    g142(.A(new_n298), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n295), .B1(new_n335), .B2(new_n345), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n344), .B1(new_n343), .B2(KEYINPUT29), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n333), .A2(new_n298), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n347), .A2(new_n294), .A3(new_n348), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n346), .A2(new_n349), .A3(KEYINPUT73), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT73), .ZN(new_n351));
  OAI211_X1 g150(.A(new_n351), .B(new_n295), .C1(new_n335), .C2(new_n345), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n350), .A2(KEYINPUT37), .A3(new_n352), .ZN(new_n353));
  XNOR2_X1  g152(.A(G8gat), .B(G36gat), .ZN(new_n354));
  XNOR2_X1  g153(.A(G64gat), .B(G92gat), .ZN(new_n355));
  XOR2_X1   g154(.A(new_n354), .B(new_n355), .Z(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n353), .A2(KEYINPUT87), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n350), .A2(new_n352), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT37), .ZN(new_n360));
  AOI21_X1  g159(.A(KEYINPUT86), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT86), .ZN(new_n362));
  AOI211_X1 g161(.A(new_n362), .B(KEYINPUT37), .C1(new_n350), .C2(new_n352), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n358), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  AOI21_X1  g163(.A(KEYINPUT87), .B1(new_n353), .B2(new_n357), .ZN(new_n365));
  OAI21_X1  g164(.A(KEYINPUT38), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT88), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  OAI211_X1 g167(.A(KEYINPUT88), .B(KEYINPUT38), .C1(new_n364), .C2(new_n365), .ZN(new_n369));
  XOR2_X1   g168(.A(G1gat), .B(G29gat), .Z(new_n370));
  XNOR2_X1  g169(.A(new_n370), .B(KEYINPUT0), .ZN(new_n371));
  XNOR2_X1  g170(.A(G57gat), .B(G85gat), .ZN(new_n372));
  XNOR2_X1  g171(.A(new_n371), .B(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n373), .ZN(new_n374));
  XNOR2_X1  g173(.A(G127gat), .B(G134gat), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT66), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(G127gat), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n378), .A2(G134gat), .ZN(new_n379));
  INV_X1    g178(.A(G134gat), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n380), .A2(G127gat), .ZN(new_n381));
  OAI21_X1  g180(.A(KEYINPUT66), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(G113gat), .ZN(new_n383));
  INV_X1    g182(.A(G120gat), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT1), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n386), .B1(G113gat), .B2(G120gat), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n377), .A2(new_n382), .A3(new_n388), .ZN(new_n389));
  OAI211_X1 g188(.A(new_n375), .B(new_n376), .C1(new_n385), .C2(new_n387), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  OR2_X1    g190(.A1(KEYINPUT75), .A2(G141gat), .ZN(new_n392));
  NAND2_X1  g191(.A1(KEYINPUT75), .A2(G141gat), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n392), .A2(G148gat), .A3(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(G148gat), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(G141gat), .ZN(new_n396));
  NAND2_X1  g195(.A1(G155gat), .A2(G162gat), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT2), .ZN(new_n398));
  INV_X1    g197(.A(G155gat), .ZN(new_n399));
  INV_X1    g198(.A(G162gat), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n398), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  AOI22_X1  g200(.A1(new_n394), .A2(new_n396), .B1(new_n397), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n399), .A2(new_n400), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(new_n397), .ZN(new_n404));
  INV_X1    g203(.A(G141gat), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(G148gat), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n396), .A2(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n404), .B1(new_n398), .B2(new_n407), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n402), .A2(new_n408), .ZN(new_n409));
  AND3_X1   g208(.A1(new_n391), .A2(new_n409), .A3(KEYINPUT4), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT67), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n391), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n389), .A2(KEYINPUT67), .A3(new_n390), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n412), .A2(new_n409), .A3(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT4), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n410), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  OAI21_X1  g215(.A(KEYINPUT3), .B1(new_n402), .B2(new_n408), .ZN(new_n417));
  XNOR2_X1  g216(.A(G141gat), .B(G148gat), .ZN(new_n418));
  OAI211_X1 g217(.A(new_n397), .B(new_n403), .C1(new_n418), .C2(KEYINPUT2), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT3), .ZN(new_n420));
  INV_X1    g219(.A(new_n396), .ZN(new_n421));
  AND2_X1   g220(.A1(KEYINPUT75), .A2(G141gat), .ZN(new_n422));
  NOR2_X1   g221(.A1(KEYINPUT75), .A2(G141gat), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n421), .B1(new_n424), .B2(G148gat), .ZN(new_n425));
  AND2_X1   g224(.A1(new_n401), .A2(new_n397), .ZN(new_n426));
  OAI211_X1 g225(.A(new_n419), .B(new_n420), .C1(new_n425), .C2(new_n426), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n417), .A2(new_n427), .A3(new_n390), .A4(new_n389), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT5), .ZN(new_n429));
  NAND2_X1  g228(.A1(G225gat), .A2(G233gat), .ZN(new_n430));
  XOR2_X1   g229(.A(new_n430), .B(KEYINPUT76), .Z(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  AND3_X1   g231(.A1(new_n428), .A2(new_n429), .A3(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n374), .B1(new_n416), .B2(new_n433), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n412), .A2(KEYINPUT4), .A3(new_n409), .A4(new_n413), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n391), .A2(new_n409), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(new_n415), .ZN(new_n437));
  NAND4_X1  g236(.A1(new_n435), .A2(new_n432), .A3(new_n428), .A4(new_n437), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n419), .B1(new_n425), .B2(new_n426), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n439), .A2(new_n390), .A3(new_n389), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n436), .A2(new_n440), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n429), .B1(new_n441), .B2(new_n431), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n438), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n434), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(KEYINPUT77), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n416), .A2(new_n433), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n443), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(new_n374), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT6), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT77), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n434), .A2(new_n450), .A3(new_n443), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n445), .A2(new_n448), .A3(new_n449), .A4(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n373), .B1(new_n443), .B2(new_n446), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(KEYINPUT6), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n359), .A2(new_n356), .ZN(new_n455));
  AND3_X1   g254(.A1(new_n452), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  XOR2_X1   g255(.A(new_n356), .B(KEYINPUT74), .Z(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT85), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n347), .A2(new_n459), .A3(new_n348), .A4(new_n294), .ZN(new_n460));
  AND2_X1   g259(.A1(new_n460), .A2(KEYINPUT37), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n346), .A2(new_n349), .A3(KEYINPUT85), .ZN(new_n462));
  AOI211_X1 g261(.A(KEYINPUT38), .B(new_n458), .C1(new_n461), .C2(new_n462), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n463), .B1(new_n361), .B2(new_n363), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n456), .A2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n368), .A2(new_n369), .A3(new_n466), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n432), .B1(new_n416), .B2(new_n428), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT39), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(new_n373), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT84), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n472), .B1(new_n441), .B2(new_n431), .ZN(new_n473));
  NAND4_X1  g272(.A1(new_n436), .A2(new_n440), .A3(KEYINPUT84), .A4(new_n432), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n473), .A2(KEYINPUT39), .A3(new_n474), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n468), .A2(new_n475), .ZN(new_n476));
  OAI21_X1  g275(.A(KEYINPUT40), .B1(new_n471), .B2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(new_n476), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT40), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n478), .A2(new_n479), .A3(new_n373), .A4(new_n470), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n453), .B1(new_n477), .B2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT30), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n350), .A2(new_n352), .A3(new_n457), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n482), .B1(new_n455), .B2(new_n483), .ZN(new_n484));
  AOI21_X1  g283(.A(KEYINPUT30), .B1(new_n359), .B2(new_n356), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n481), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  XNOR2_X1  g285(.A(G78gat), .B(G106gat), .ZN(new_n487));
  XNOR2_X1  g286(.A(new_n487), .B(KEYINPUT80), .ZN(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  XNOR2_X1  g288(.A(KEYINPUT79), .B(KEYINPUT31), .ZN(new_n490));
  XNOR2_X1  g289(.A(new_n490), .B(G50gat), .ZN(new_n491));
  INV_X1    g290(.A(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT81), .ZN(new_n493));
  INV_X1    g292(.A(G228gat), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n494), .A2(new_n297), .ZN(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  AOI21_X1  g295(.A(KEYINPUT29), .B1(new_n409), .B2(new_n420), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n496), .B1(new_n497), .B2(new_n294), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n294), .A2(KEYINPUT82), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT82), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n334), .B1(new_n288), .B2(new_n500), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n420), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n498), .B1(new_n502), .B2(new_n439), .ZN(new_n503));
  AOI21_X1  g302(.A(KEYINPUT29), .B1(new_n288), .B2(new_n293), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n439), .B1(new_n504), .B2(KEYINPUT3), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(KEYINPUT83), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT83), .ZN(new_n507));
  OAI211_X1 g306(.A(new_n507), .B(new_n439), .C1(new_n504), .C2(KEYINPUT3), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n497), .A2(new_n294), .ZN(new_n509));
  INV_X1    g308(.A(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n506), .A2(new_n508), .A3(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n503), .B1(new_n495), .B2(new_n511), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n493), .B1(new_n512), .B2(new_n243), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n509), .B1(new_n505), .B2(KEYINPUT83), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n496), .B1(new_n514), .B2(new_n508), .ZN(new_n515));
  OAI21_X1  g314(.A(G22gat), .B1(new_n515), .B2(new_n503), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n492), .B1(new_n513), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n511), .A2(new_n495), .ZN(new_n518));
  INV_X1    g317(.A(new_n503), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n518), .A2(new_n243), .A3(new_n519), .ZN(new_n520));
  AND4_X1   g319(.A1(KEYINPUT81), .A2(new_n516), .A3(new_n520), .A4(new_n492), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n489), .B1(new_n517), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n516), .A2(new_n520), .A3(KEYINPUT81), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(new_n491), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n513), .A2(new_n492), .A3(new_n516), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n524), .A2(new_n525), .A3(new_n488), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n486), .A2(new_n522), .A3(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n467), .A2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT71), .ZN(new_n530));
  XNOR2_X1  g329(.A(G15gat), .B(G43gat), .ZN(new_n531));
  OR2_X1    g330(.A1(new_n531), .A2(KEYINPUT68), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(KEYINPUT68), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n534), .A2(G71gat), .ZN(new_n535));
  INV_X1    g334(.A(G71gat), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n532), .A2(new_n536), .A3(new_n533), .ZN(new_n537));
  AND3_X1   g336(.A1(new_n535), .A2(G99gat), .A3(new_n537), .ZN(new_n538));
  AOI21_X1  g337(.A(G99gat), .B1(new_n535), .B2(new_n537), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(G227gat), .A2(G233gat), .ZN(new_n541));
  INV_X1    g340(.A(new_n316), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(new_n321), .ZN(new_n543));
  AND3_X1   g342(.A1(new_n304), .A2(new_n309), .A3(KEYINPUT25), .ZN(new_n544));
  AOI22_X1  g343(.A1(new_n543), .A2(new_n299), .B1(new_n544), .B2(new_n320), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n341), .B1(new_n338), .B2(new_n339), .ZN(new_n546));
  AND3_X1   g345(.A1(new_n389), .A2(KEYINPUT67), .A3(new_n390), .ZN(new_n547));
  AOI21_X1  g346(.A(KEYINPUT67), .B1(new_n389), .B2(new_n390), .ZN(new_n548));
  OAI22_X1  g347(.A1(new_n545), .A2(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND4_X1  g348(.A1(new_n412), .A2(new_n323), .A3(new_n332), .A4(new_n413), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n541), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n540), .B1(new_n551), .B2(KEYINPUT33), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT32), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n549), .A2(new_n550), .ZN(new_n556));
  INV_X1    g355(.A(new_n541), .ZN(new_n557));
  AOI221_X4 g356(.A(new_n553), .B1(new_n540), .B2(KEYINPUT33), .C1(new_n556), .C2(new_n557), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n530), .B1(new_n555), .B2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n550), .ZN(new_n560));
  AOI22_X1  g359(.A1(new_n413), .A2(new_n412), .B1(new_n323), .B2(new_n332), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n557), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n562), .A2(KEYINPUT32), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT33), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n563), .A2(new_n565), .A3(new_n540), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n552), .A2(new_n554), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n566), .A2(KEYINPUT71), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n556), .A2(KEYINPUT70), .ZN(new_n569));
  AND2_X1   g368(.A1(KEYINPUT70), .A2(KEYINPUT34), .ZN(new_n570));
  OAI211_X1 g369(.A(new_n569), .B(new_n541), .C1(new_n556), .C2(new_n570), .ZN(new_n571));
  AND2_X1   g370(.A1(KEYINPUT69), .A2(KEYINPUT34), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n549), .A2(new_n541), .A3(new_n550), .ZN(new_n573));
  NOR2_X1   g372(.A1(KEYINPUT69), .A2(KEYINPUT34), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n572), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n571), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n559), .A2(new_n568), .A3(new_n576), .ZN(new_n577));
  AND2_X1   g376(.A1(new_n571), .A2(new_n575), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n578), .A2(KEYINPUT71), .A3(new_n566), .A4(new_n567), .ZN(new_n579));
  AND3_X1   g378(.A1(new_n577), .A2(KEYINPUT36), .A3(new_n579), .ZN(new_n580));
  AOI21_X1  g379(.A(KEYINPUT36), .B1(new_n577), .B2(new_n579), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n522), .A2(new_n526), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n451), .A2(new_n449), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n450), .B1(new_n434), .B2(new_n443), .ZN(new_n585));
  OAI21_X1  g384(.A(KEYINPUT78), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT78), .ZN(new_n587));
  NAND4_X1  g386(.A1(new_n445), .A2(new_n587), .A3(new_n449), .A4(new_n451), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n586), .A2(new_n448), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(new_n454), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n484), .A2(new_n485), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n583), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n529), .A2(new_n582), .A3(new_n593), .ZN(new_n594));
  AND2_X1   g393(.A1(new_n522), .A2(new_n526), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n455), .A2(new_n483), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n596), .A2(KEYINPUT30), .ZN(new_n597));
  INV_X1    g396(.A(new_n485), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  AND2_X1   g398(.A1(new_n452), .A2(new_n454), .ZN(new_n600));
  NOR3_X1   g399(.A1(new_n599), .A2(KEYINPUT35), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n577), .A2(new_n579), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n595), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n522), .A2(new_n526), .A3(new_n602), .ZN(new_n604));
  OAI21_X1  g403(.A(KEYINPUT35), .B1(new_n604), .B2(new_n592), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n278), .B1(new_n594), .B2(new_n606), .ZN(new_n607));
  AND2_X1   g406(.A1(G71gat), .A2(G78gat), .ZN(new_n608));
  NOR2_X1   g407(.A1(G71gat), .A2(G78gat), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(G57gat), .B(G64gat), .ZN(new_n611));
  AOI21_X1  g410(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n610), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(G57gat), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n614), .A2(G64gat), .ZN(new_n615));
  INV_X1    g414(.A(G64gat), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(G57gat), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(G71gat), .B(G78gat), .ZN(new_n619));
  INV_X1    g418(.A(new_n612), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n618), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  AND3_X1   g420(.A1(new_n613), .A2(new_n621), .A3(KEYINPUT93), .ZN(new_n622));
  AOI21_X1  g421(.A(KEYINPUT93), .B1(new_n613), .B2(new_n621), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT21), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(G127gat), .B(G155gat), .ZN(new_n627));
  OR2_X1    g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n626), .A2(new_n627), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n624), .A2(new_n625), .ZN(new_n631));
  NOR3_X1   g430(.A1(new_n631), .A2(KEYINPUT94), .A3(new_n262), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  OAI21_X1  g432(.A(KEYINPUT94), .B1(new_n631), .B2(new_n262), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n630), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n630), .A2(new_n633), .A3(new_n634), .ZN(new_n637));
  XNOR2_X1  g436(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n638));
  NAND2_X1  g437(.A1(G231gat), .A2(G233gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(G183gat), .B(G211gat), .ZN(new_n641));
  XOR2_X1   g440(.A(new_n640), .B(new_n641), .Z(new_n642));
  NAND3_X1  g441(.A1(new_n636), .A2(new_n637), .A3(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n642), .ZN(new_n644));
  INV_X1    g443(.A(new_n637), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n644), .B1(new_n645), .B2(new_n635), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n643), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(G92gat), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n649), .A2(KEYINPUT7), .A3(G85gat), .ZN(new_n650));
  NAND2_X1  g449(.A1(KEYINPUT7), .A2(G85gat), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n651), .A2(G92gat), .ZN(new_n652));
  NOR2_X1   g451(.A1(KEYINPUT7), .A2(G85gat), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n650), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(G99gat), .A2(G106gat), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n655), .A2(KEYINPUT95), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT95), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n657), .A2(G99gat), .A3(G106gat), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n656), .A2(new_n658), .A3(KEYINPUT8), .ZN(new_n659));
  XNOR2_X1  g458(.A(G99gat), .B(G106gat), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n654), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n660), .B1(new_n654), .B2(new_n659), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  OR2_X1    g463(.A1(new_n664), .A2(KEYINPUT96), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(KEYINPUT96), .ZN(new_n666));
  INV_X1    g465(.A(new_n258), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n261), .A2(new_n667), .ZN(new_n668));
  NAND4_X1  g467(.A1(new_n665), .A2(new_n666), .A3(new_n238), .A4(new_n668), .ZN(new_n669));
  AND2_X1   g468(.A1(G232gat), .A2(G233gat), .ZN(new_n670));
  AOI22_X1  g469(.A1(new_n261), .A2(new_n664), .B1(KEYINPUT41), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  XOR2_X1   g471(.A(G190gat), .B(G218gat), .Z(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n673), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n669), .A2(new_n671), .A3(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  XOR2_X1   g476(.A(G134gat), .B(G162gat), .Z(new_n678));
  NOR2_X1   g477(.A1(new_n670), .A2(KEYINPUT41), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XOR2_X1   g479(.A(new_n680), .B(KEYINPUT97), .Z(new_n681));
  NAND2_X1  g480(.A1(new_n677), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n680), .A2(KEYINPUT97), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n674), .A2(new_n683), .A3(new_n676), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(G230gat), .A2(G233gat), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n686), .B(KEYINPUT99), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  XOR2_X1   g487(.A(KEYINPUT98), .B(KEYINPUT10), .Z(new_n689));
  OAI22_X1  g488(.A1(new_n622), .A2(new_n623), .B1(new_n662), .B2(new_n663), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n654), .A2(new_n659), .ZN(new_n691));
  INV_X1    g490(.A(new_n660), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n613), .A2(new_n621), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n693), .A2(new_n694), .A3(new_n661), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n689), .B1(new_n690), .B2(new_n695), .ZN(new_n696));
  OAI21_X1  g495(.A(KEYINPUT10), .B1(new_n622), .B2(new_n623), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n693), .A2(new_n661), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n688), .B1(new_n696), .B2(new_n699), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n690), .A2(new_n687), .A3(new_n695), .ZN(new_n701));
  XNOR2_X1  g500(.A(G120gat), .B(G148gat), .ZN(new_n702));
  XNOR2_X1  g501(.A(G176gat), .B(G204gat), .ZN(new_n703));
  XOR2_X1   g502(.A(new_n702), .B(new_n703), .Z(new_n704));
  NAND3_X1  g503(.A1(new_n700), .A2(new_n701), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(KEYINPUT100), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT100), .ZN(new_n707));
  NAND4_X1  g506(.A1(new_n700), .A2(new_n707), .A3(new_n701), .A4(new_n704), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n700), .A2(new_n701), .ZN(new_n710));
  INV_X1    g509(.A(new_n704), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n709), .A2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(new_n713), .ZN(new_n714));
  NAND4_X1  g513(.A1(new_n648), .A2(KEYINPUT101), .A3(new_n685), .A4(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT101), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n685), .A2(new_n643), .A3(new_n646), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n716), .B1(new_n717), .B2(new_n713), .ZN(new_n718));
  AND2_X1   g517(.A1(new_n715), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n607), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n720), .A2(new_n590), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(new_n239), .ZN(G1324gat));
  INV_X1    g521(.A(new_n720), .ZN(new_n723));
  XOR2_X1   g522(.A(KEYINPUT16), .B(G8gat), .Z(new_n724));
  NAND3_X1  g523(.A1(new_n723), .A2(new_n599), .A3(new_n724), .ZN(new_n725));
  OAI21_X1  g524(.A(G8gat), .B1(new_n720), .B2(new_n591), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  MUX2_X1   g526(.A(new_n725), .B(new_n727), .S(KEYINPUT42), .Z(G1325gat));
  INV_X1    g527(.A(KEYINPUT102), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n729), .B1(new_n580), .B2(new_n581), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT36), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n602), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n577), .A2(KEYINPUT36), .A3(new_n579), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n732), .A2(KEYINPUT102), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n730), .A2(new_n734), .ZN(new_n735));
  OAI21_X1  g534(.A(G15gat), .B1(new_n720), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n602), .A2(new_n241), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n736), .B1(new_n720), .B2(new_n737), .ZN(G1326gat));
  NOR2_X1   g537(.A1(new_n720), .A2(new_n595), .ZN(new_n739));
  XOR2_X1   g538(.A(KEYINPUT43), .B(G22gat), .Z(new_n740));
  XNOR2_X1  g539(.A(new_n739), .B(new_n740), .ZN(G1327gat));
  INV_X1    g540(.A(new_n685), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n647), .A2(new_n742), .A3(new_n714), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(KEYINPUT103), .ZN(new_n744));
  AND2_X1   g543(.A1(new_n607), .A2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(new_n590), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n745), .A2(new_n220), .A3(new_n746), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(KEYINPUT45), .ZN(new_n748));
  NOR3_X1   g547(.A1(new_n580), .A2(new_n581), .A3(new_n729), .ZN(new_n749));
  AOI21_X1  g548(.A(KEYINPUT102), .B1(new_n732), .B2(new_n733), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n593), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n465), .B1(new_n366), .B2(new_n367), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n527), .B1(new_n752), .B2(new_n369), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n606), .B1(new_n751), .B2(new_n753), .ZN(new_n754));
  AOI21_X1  g553(.A(KEYINPUT44), .B1(new_n754), .B2(new_n742), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n742), .A2(KEYINPUT44), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n756), .B1(new_n594), .B2(new_n606), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  NOR3_X1   g557(.A1(new_n648), .A2(new_n278), .A3(new_n713), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  OAI21_X1  g559(.A(G29gat), .B1(new_n760), .B2(new_n590), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n748), .A2(new_n761), .ZN(G1328gat));
  NAND3_X1  g561(.A1(new_n745), .A2(new_n221), .A3(new_n599), .ZN(new_n763));
  AND2_X1   g562(.A1(KEYINPUT104), .A2(KEYINPUT46), .ZN(new_n764));
  NOR2_X1   g563(.A1(KEYINPUT104), .A2(KEYINPUT46), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n763), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  OAI21_X1  g565(.A(G36gat), .B1(new_n760), .B2(new_n591), .ZN(new_n767));
  OAI211_X1 g566(.A(new_n766), .B(new_n767), .C1(new_n764), .C2(new_n763), .ZN(G1329gat));
  INV_X1    g567(.A(KEYINPUT44), .ZN(new_n769));
  AOI22_X1  g568(.A1(new_n730), .A2(new_n734), .B1(new_n592), .B2(new_n583), .ZN(new_n770));
  AOI22_X1  g569(.A1(new_n529), .A2(new_n770), .B1(new_n605), .B2(new_n603), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n769), .B1(new_n771), .B2(new_n685), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n749), .A2(new_n750), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n593), .A2(new_n582), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n606), .B1(new_n753), .B2(new_n774), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n775), .A2(KEYINPUT44), .A3(new_n742), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n772), .A2(new_n773), .A3(new_n776), .A4(new_n759), .ZN(new_n777));
  AND2_X1   g576(.A1(new_n777), .A2(G43gat), .ZN(new_n778));
  INV_X1    g577(.A(new_n602), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n779), .A2(G43gat), .ZN(new_n780));
  AND2_X1   g579(.A1(new_n745), .A2(new_n780), .ZN(new_n781));
  OAI21_X1  g580(.A(KEYINPUT105), .B1(new_n778), .B2(new_n781), .ZN(new_n782));
  XNOR2_X1  g581(.A(new_n782), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g582(.A(G50gat), .B1(new_n760), .B2(new_n595), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT107), .ZN(new_n785));
  AOI21_X1  g584(.A(KEYINPUT48), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n595), .A2(G50gat), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n787), .B(KEYINPUT106), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n745), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n784), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n786), .A2(new_n790), .ZN(new_n791));
  OAI211_X1 g590(.A(new_n784), .B(new_n789), .C1(new_n785), .C2(KEYINPUT48), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(G1331gat));
  NOR4_X1   g592(.A1(new_n771), .A2(new_n277), .A3(new_n717), .A4(new_n714), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(new_n746), .ZN(new_n795));
  XNOR2_X1  g594(.A(new_n795), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g595(.A1(new_n794), .A2(new_n599), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n797), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n798));
  XOR2_X1   g597(.A(KEYINPUT49), .B(G64gat), .Z(new_n799));
  OAI21_X1  g598(.A(new_n798), .B1(new_n797), .B2(new_n799), .ZN(G1333gat));
  AOI21_X1  g599(.A(new_n536), .B1(new_n794), .B2(new_n773), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n779), .A2(G71gat), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n801), .B1(new_n794), .B2(new_n802), .ZN(new_n803));
  XNOR2_X1  g602(.A(new_n803), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g603(.A1(new_n794), .A2(new_n583), .ZN(new_n805));
  XNOR2_X1  g604(.A(new_n805), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g605(.A1(new_n647), .A2(new_n278), .ZN(new_n807));
  XOR2_X1   g606(.A(new_n807), .B(KEYINPUT108), .Z(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(new_n713), .ZN(new_n809));
  NOR3_X1   g608(.A1(new_n755), .A2(new_n757), .A3(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(new_n810), .ZN(new_n811));
  OAI21_X1  g610(.A(G85gat), .B1(new_n811), .B2(new_n590), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n529), .A2(new_n770), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n685), .B1(new_n813), .B2(new_n606), .ZN(new_n814));
  AOI21_X1  g613(.A(KEYINPUT51), .B1(new_n814), .B2(new_n808), .ZN(new_n815));
  AND4_X1   g614(.A1(KEYINPUT51), .A2(new_n754), .A3(new_n742), .A4(new_n808), .ZN(new_n816));
  OR2_X1    g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n590), .A2(G85gat), .A3(new_n714), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n812), .A2(new_n819), .ZN(G1336gat));
  OAI21_X1  g619(.A(KEYINPUT110), .B1(new_n811), .B2(new_n591), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT110), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n810), .A2(new_n822), .A3(new_n599), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n821), .A2(G92gat), .A3(new_n823), .ZN(new_n824));
  NOR3_X1   g623(.A1(new_n591), .A2(G92gat), .A3(new_n714), .ZN(new_n825));
  AOI21_X1  g624(.A(KEYINPUT52), .B1(new_n817), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n754), .A2(new_n742), .A3(new_n808), .ZN(new_n828));
  AND3_X1   g627(.A1(new_n828), .A2(KEYINPUT109), .A3(KEYINPUT51), .ZN(new_n829));
  AOI21_X1  g628(.A(KEYINPUT51), .B1(new_n828), .B2(KEYINPUT109), .ZN(new_n830));
  INV_X1    g629(.A(new_n825), .ZN(new_n831));
  NOR3_X1   g630(.A1(new_n829), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n649), .B1(new_n810), .B2(new_n599), .ZN(new_n833));
  OAI21_X1  g632(.A(KEYINPUT52), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n827), .A2(new_n834), .ZN(G1337gat));
  OAI21_X1  g634(.A(G99gat), .B1(new_n811), .B2(new_n735), .ZN(new_n836));
  NOR3_X1   g635(.A1(new_n779), .A2(G99gat), .A3(new_n714), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n817), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n836), .A2(new_n838), .ZN(G1338gat));
  NOR3_X1   g638(.A1(new_n595), .A2(G106gat), .A3(new_n714), .ZN(new_n840));
  INV_X1    g639(.A(new_n840), .ZN(new_n841));
  NOR3_X1   g640(.A1(new_n829), .A2(new_n830), .A3(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(new_n809), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n772), .A2(new_n583), .A3(new_n776), .A4(new_n843), .ZN(new_n844));
  AND2_X1   g643(.A1(new_n844), .A2(G106gat), .ZN(new_n845));
  OAI21_X1  g644(.A(KEYINPUT53), .B1(new_n842), .B2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT111), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n844), .A2(G106gat), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n840), .B1(new_n815), .B2(new_n816), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT53), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n849), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(KEYINPUT112), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT112), .ZN(new_n854));
  NAND4_X1  g653(.A1(new_n849), .A2(new_n850), .A3(new_n854), .A4(new_n851), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  OAI211_X1 g655(.A(KEYINPUT111), .B(KEYINPUT53), .C1(new_n842), .C2(new_n845), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n848), .A2(new_n856), .A3(new_n857), .ZN(G1339gat));
  NOR3_X1   g657(.A1(new_n717), .A2(new_n277), .A3(new_n713), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT55), .ZN(new_n860));
  INV_X1    g659(.A(new_n689), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT93), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n694), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n613), .A2(new_n621), .A3(KEYINPUT93), .ZN(new_n864));
  AOI22_X1  g663(.A1(new_n863), .A2(new_n864), .B1(new_n661), .B2(new_n693), .ZN(new_n865));
  INV_X1    g664(.A(new_n695), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n861), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  OAI211_X1 g666(.A(new_n664), .B(KEYINPUT10), .C1(new_n622), .C2(new_n623), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n867), .A2(new_n687), .A3(new_n868), .ZN(new_n869));
  AND3_X1   g668(.A1(new_n700), .A2(new_n869), .A3(KEYINPUT54), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT54), .ZN(new_n871));
  OAI211_X1 g670(.A(new_n871), .B(new_n688), .C1(new_n696), .C2(new_n699), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(new_n711), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n860), .B1(new_n870), .B2(new_n873), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n687), .B1(new_n867), .B2(new_n868), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n704), .B1(new_n875), .B2(new_n871), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n700), .A2(new_n869), .A3(KEYINPUT54), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n876), .A2(KEYINPUT55), .A3(new_n877), .ZN(new_n878));
  AND4_X1   g677(.A1(new_n277), .A2(new_n874), .A3(new_n709), .A4(new_n878), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n260), .B1(new_n259), .B2(new_n263), .ZN(new_n880));
  NOR3_X1   g679(.A1(new_n269), .A2(new_n270), .A3(new_n268), .ZN(new_n881));
  OAI22_X1  g680(.A1(new_n880), .A2(new_n881), .B1(new_n209), .B2(new_n210), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n276), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n883), .B1(new_n709), .B2(new_n712), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n685), .B1(new_n879), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n867), .A2(new_n868), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n871), .B1(new_n886), .B2(new_n688), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n873), .B1(new_n869), .B2(new_n887), .ZN(new_n888));
  AOI22_X1  g687(.A1(new_n888), .A2(KEYINPUT55), .B1(new_n706), .B2(new_n708), .ZN(new_n889));
  INV_X1    g688(.A(new_n883), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n742), .A2(new_n889), .A3(new_n890), .A4(new_n874), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n885), .A2(new_n891), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n859), .B1(new_n892), .B2(new_n647), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n893), .A2(new_n583), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n894), .A2(new_n746), .A3(new_n591), .A4(new_n602), .ZN(new_n895));
  NOR3_X1   g694(.A1(new_n895), .A2(new_n383), .A3(new_n278), .ZN(new_n896));
  INV_X1    g695(.A(new_n893), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(new_n746), .ZN(new_n898));
  INV_X1    g697(.A(new_n898), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n604), .A2(new_n599), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  INV_X1    g700(.A(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(new_n277), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n896), .B1(new_n903), .B2(new_n383), .ZN(G1340gat));
  NOR3_X1   g703(.A1(new_n895), .A2(new_n384), .A3(new_n714), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n902), .A2(new_n713), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n905), .B1(new_n906), .B2(new_n384), .ZN(G1341gat));
  OAI21_X1  g706(.A(G127gat), .B1(new_n895), .B2(new_n647), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n648), .A2(new_n378), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n908), .B1(new_n901), .B2(new_n909), .ZN(G1342gat));
  NAND3_X1  g709(.A1(new_n902), .A2(new_n380), .A3(new_n742), .ZN(new_n911));
  OR2_X1    g710(.A1(new_n911), .A2(KEYINPUT56), .ZN(new_n912));
  OAI21_X1  g711(.A(G134gat), .B1(new_n895), .B2(new_n685), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n911), .A2(KEYINPUT56), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(G1343gat));
  NOR2_X1   g714(.A1(new_n898), .A2(new_n599), .ZN(new_n916));
  OR3_X1    g715(.A1(new_n773), .A2(KEYINPUT116), .A3(new_n595), .ZN(new_n917));
  OAI21_X1  g716(.A(KEYINPUT116), .B1(new_n773), .B2(new_n595), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n278), .A2(G141gat), .ZN(new_n919));
  AND4_X1   g718(.A1(new_n916), .A2(new_n917), .A3(new_n918), .A4(new_n919), .ZN(new_n920));
  INV_X1    g719(.A(new_n920), .ZN(new_n921));
  INV_X1    g720(.A(new_n424), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n746), .A2(new_n591), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n773), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n583), .A2(KEYINPUT57), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n874), .A2(KEYINPUT113), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n876), .A2(new_n877), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT113), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n927), .A2(new_n928), .A3(new_n860), .ZN(new_n929));
  NAND4_X1  g728(.A1(new_n889), .A2(new_n926), .A3(new_n277), .A4(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(new_n884), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n742), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT114), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n891), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n928), .B1(new_n927), .B2(new_n860), .ZN(new_n935));
  AOI211_X1 g734(.A(KEYINPUT113), .B(KEYINPUT55), .C1(new_n876), .C2(new_n877), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  AND3_X1   g736(.A1(new_n277), .A2(new_n709), .A3(new_n878), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n884), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NOR3_X1   g738(.A1(new_n939), .A2(KEYINPUT114), .A3(new_n742), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n647), .B1(new_n934), .B2(new_n940), .ZN(new_n941));
  INV_X1    g740(.A(new_n859), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n925), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  AOI21_X1  g742(.A(KEYINPUT57), .B1(new_n897), .B2(new_n583), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n924), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n922), .B1(new_n945), .B2(new_n278), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT58), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n921), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT117), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT57), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n950), .B1(new_n893), .B2(new_n595), .ZN(new_n951));
  OAI21_X1  g750(.A(KEYINPUT114), .B1(new_n939), .B2(new_n742), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n926), .A2(new_n929), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n277), .A2(new_n709), .A3(new_n878), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n931), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n955), .A2(new_n933), .A3(new_n685), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n952), .A2(new_n891), .A3(new_n956), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n859), .B1(new_n957), .B2(new_n647), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n951), .B1(new_n958), .B2(new_n925), .ZN(new_n959));
  AND3_X1   g758(.A1(new_n959), .A2(KEYINPUT115), .A3(new_n924), .ZN(new_n960));
  AOI21_X1  g759(.A(KEYINPUT115), .B1(new_n959), .B2(new_n924), .ZN(new_n961));
  NOR3_X1   g760(.A1(new_n960), .A2(new_n961), .A3(new_n278), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n921), .B1(new_n962), .B2(new_n424), .ZN(new_n963));
  AOI21_X1  g762(.A(new_n949), .B1(new_n963), .B2(KEYINPUT58), .ZN(new_n964));
  INV_X1    g763(.A(KEYINPUT115), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n945), .A2(new_n965), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n959), .A2(KEYINPUT115), .A3(new_n924), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n966), .A2(new_n277), .A3(new_n967), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n920), .B1(new_n968), .B2(new_n922), .ZN(new_n969));
  NOR3_X1   g768(.A1(new_n969), .A2(KEYINPUT117), .A3(new_n947), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n948), .B1(new_n964), .B2(new_n970), .ZN(G1344gat));
  AND2_X1   g770(.A1(new_n917), .A2(new_n918), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n972), .A2(new_n916), .ZN(new_n973));
  NOR3_X1   g772(.A1(new_n973), .A2(G148gat), .A3(new_n714), .ZN(new_n974));
  XNOR2_X1  g773(.A(new_n974), .B(KEYINPUT118), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n891), .B1(new_n939), .B2(new_n742), .ZN(new_n976));
  INV_X1    g775(.A(KEYINPUT121), .ZN(new_n977));
  AOI21_X1  g776(.A(new_n648), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  OAI21_X1  g777(.A(new_n978), .B1(new_n977), .B2(new_n976), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n715), .A2(new_n718), .A3(new_n278), .ZN(new_n980));
  INV_X1    g779(.A(KEYINPUT120), .ZN(new_n981));
  XNOR2_X1  g780(.A(new_n980), .B(new_n981), .ZN(new_n982));
  AOI21_X1  g781(.A(new_n595), .B1(new_n979), .B2(new_n982), .ZN(new_n983));
  OAI22_X1  g782(.A1(new_n983), .A2(KEYINPUT57), .B1(new_n893), .B2(new_n925), .ZN(new_n984));
  NOR3_X1   g783(.A1(new_n773), .A2(new_n714), .A3(new_n923), .ZN(new_n985));
  NAND3_X1  g784(.A1(new_n984), .A2(KEYINPUT122), .A3(new_n985), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n986), .A2(G148gat), .ZN(new_n987));
  AOI21_X1  g786(.A(KEYINPUT122), .B1(new_n984), .B2(new_n985), .ZN(new_n988));
  OAI21_X1  g787(.A(KEYINPUT59), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  NOR2_X1   g788(.A1(new_n395), .A2(KEYINPUT59), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n966), .A2(new_n967), .ZN(new_n991));
  OAI21_X1  g790(.A(new_n990), .B1(new_n991), .B2(new_n714), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n992), .A2(KEYINPUT119), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n989), .A2(new_n993), .ZN(new_n994));
  NOR2_X1   g793(.A1(new_n992), .A2(KEYINPUT119), .ZN(new_n995));
  OAI21_X1  g794(.A(new_n975), .B1(new_n994), .B2(new_n995), .ZN(G1345gat));
  OAI21_X1  g795(.A(G155gat), .B1(new_n991), .B2(new_n647), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n648), .A2(new_n399), .ZN(new_n998));
  OAI21_X1  g797(.A(new_n997), .B1(new_n973), .B2(new_n998), .ZN(G1346gat));
  OAI21_X1  g798(.A(G162gat), .B1(new_n991), .B2(new_n685), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n742), .A2(new_n400), .ZN(new_n1001));
  OAI21_X1  g800(.A(new_n1000), .B1(new_n973), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g801(.A(KEYINPUT123), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  OAI211_X1 g803(.A(new_n1000), .B(KEYINPUT123), .C1(new_n973), .C2(new_n1001), .ZN(new_n1005));
  NAND2_X1  g804(.A1(new_n1004), .A2(new_n1005), .ZN(G1347gat));
  NOR3_X1   g805(.A1(new_n746), .A2(new_n779), .A3(new_n591), .ZN(new_n1007));
  NAND2_X1  g806(.A1(new_n894), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g807(.A(new_n1008), .ZN(new_n1009));
  AND3_X1   g808(.A1(new_n1009), .A2(G169gat), .A3(new_n277), .ZN(new_n1010));
  NOR4_X1   g809(.A1(new_n893), .A2(new_n746), .A3(new_n591), .A4(new_n604), .ZN(new_n1011));
  AOI21_X1  g810(.A(G169gat), .B1(new_n1011), .B2(new_n277), .ZN(new_n1012));
  NOR2_X1   g811(.A1(new_n1010), .A2(new_n1012), .ZN(G1348gat));
  OAI21_X1  g812(.A(G176gat), .B1(new_n1008), .B2(new_n714), .ZN(new_n1014));
  INV_X1    g813(.A(G176gat), .ZN(new_n1015));
  NAND3_X1  g814(.A1(new_n1011), .A2(new_n1015), .A3(new_n713), .ZN(new_n1016));
  NAND2_X1  g815(.A1(new_n1014), .A2(new_n1016), .ZN(G1349gat));
  NAND2_X1  g816(.A1(new_n1009), .A2(new_n648), .ZN(new_n1018));
  NOR2_X1   g817(.A1(new_n647), .A2(new_n337), .ZN(new_n1019));
  AOI22_X1  g818(.A1(new_n1018), .A2(G183gat), .B1(new_n1011), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g819(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n1021));
  XNOR2_X1  g820(.A(new_n1020), .B(new_n1021), .ZN(G1350gat));
  OAI21_X1  g821(.A(G190gat), .B1(new_n1008), .B2(new_n685), .ZN(new_n1023));
  XNOR2_X1  g822(.A(new_n1023), .B(KEYINPUT61), .ZN(new_n1024));
  NAND3_X1  g823(.A1(new_n1011), .A2(new_n328), .A3(new_n742), .ZN(new_n1025));
  NAND2_X1  g824(.A1(new_n1024), .A2(new_n1025), .ZN(G1351gat));
  NOR2_X1   g825(.A1(new_n893), .A2(new_n746), .ZN(new_n1027));
  AND4_X1   g826(.A1(new_n599), .A2(new_n1027), .A3(new_n583), .A4(new_n735), .ZN(new_n1028));
  AOI21_X1  g827(.A(G197gat), .B1(new_n1028), .B2(new_n277), .ZN(new_n1029));
  NAND3_X1  g828(.A1(new_n735), .A2(new_n590), .A3(new_n599), .ZN(new_n1030));
  XNOR2_X1  g829(.A(new_n1030), .B(KEYINPUT125), .ZN(new_n1031));
  AND3_X1   g830(.A1(new_n1031), .A2(G197gat), .A3(new_n277), .ZN(new_n1032));
  AOI21_X1  g831(.A(new_n1029), .B1(new_n1032), .B2(new_n984), .ZN(G1352gat));
  AOI21_X1  g832(.A(G204gat), .B1(KEYINPUT126), .B2(KEYINPUT62), .ZN(new_n1034));
  NAND3_X1  g833(.A1(new_n1028), .A2(new_n713), .A3(new_n1034), .ZN(new_n1035));
  NOR2_X1   g834(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n1036));
  XNOR2_X1  g835(.A(new_n1035), .B(new_n1036), .ZN(new_n1037));
  NAND3_X1  g836(.A1(new_n984), .A2(new_n713), .A3(new_n1031), .ZN(new_n1038));
  NAND2_X1  g837(.A1(new_n1038), .A2(G204gat), .ZN(new_n1039));
  NAND2_X1  g838(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g839(.A(KEYINPUT127), .ZN(new_n1041));
  XNOR2_X1  g840(.A(new_n1040), .B(new_n1041), .ZN(G1353gat));
  NAND3_X1  g841(.A1(new_n1028), .A2(new_n291), .A3(new_n648), .ZN(new_n1043));
  NOR2_X1   g842(.A1(new_n1030), .A2(new_n647), .ZN(new_n1044));
  NAND2_X1  g843(.A1(new_n984), .A2(new_n1044), .ZN(new_n1045));
  AND3_X1   g844(.A1(new_n1045), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1046));
  AOI21_X1  g845(.A(KEYINPUT63), .B1(new_n1045), .B2(G211gat), .ZN(new_n1047));
  OAI21_X1  g846(.A(new_n1043), .B1(new_n1046), .B2(new_n1047), .ZN(G1354gat));
  AOI21_X1  g847(.A(G218gat), .B1(new_n1028), .B2(new_n742), .ZN(new_n1049));
  AND2_X1   g848(.A1(new_n984), .A2(new_n1031), .ZN(new_n1050));
  NOR2_X1   g849(.A1(new_n685), .A2(new_n290), .ZN(new_n1051));
  AOI21_X1  g850(.A(new_n1049), .B1(new_n1050), .B2(new_n1051), .ZN(G1355gat));
endmodule


