//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 1 0 0 0 0 1 0 0 0 0 0 1 0 1 1 0 1 0 0 0 0 1 0 1 1 0 1 0 0 0 0 0 1 0 1 1 1 1 1 0 1 1 0 1 0 1 0 0 0 1 0 0 0 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n736, new_n737, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n767, new_n768, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n780, new_n781, new_n782, new_n783, new_n785, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n817,
    new_n818, new_n819, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n940, new_n941, new_n942, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n973, new_n974, new_n975, new_n976, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1003, new_n1004, new_n1005, new_n1006, new_n1008,
    new_n1009;
  INV_X1    g000(.A(KEYINPUT82), .ZN(new_n202));
  NOR2_X1   g001(.A1(G169gat), .A2(G176gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(G169gat), .A2(G176gat), .ZN(new_n204));
  AOI21_X1  g003(.A(new_n203), .B1(KEYINPUT23), .B2(new_n204), .ZN(new_n205));
  AND2_X1   g004(.A1(new_n203), .A2(KEYINPUT23), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(G183gat), .ZN(new_n208));
  INV_X1    g007(.A(G190gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND3_X1  g009(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  AOI21_X1  g011(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n213));
  OAI21_X1  g012(.A(KEYINPUT64), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(new_n213), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT64), .ZN(new_n216));
  NAND4_X1  g015(.A1(new_n215), .A2(new_n210), .A3(new_n216), .A4(new_n211), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n207), .A2(new_n214), .A3(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT25), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  XOR2_X1   g019(.A(KEYINPUT66), .B(KEYINPUT24), .Z(new_n221));
  INV_X1    g020(.A(KEYINPUT67), .ZN(new_n222));
  NAND2_X1  g021(.A1(G183gat), .A2(G190gat), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(KEYINPUT66), .B(KEYINPUT24), .ZN(new_n225));
  INV_X1    g024(.A(new_n223), .ZN(new_n226));
  OAI21_X1  g025(.A(KEYINPUT67), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n212), .B1(new_n224), .B2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT65), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n203), .A2(new_n229), .ZN(new_n230));
  OAI21_X1  g029(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n231));
  AND2_X1   g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(KEYINPUT23), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n205), .A2(new_n219), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n220), .B1(new_n228), .B2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT28), .ZN(new_n237));
  XNOR2_X1  g036(.A(KEYINPUT27), .B(G183gat), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT68), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n239), .B1(new_n208), .B2(KEYINPUT27), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(new_n209), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n237), .B1(new_n240), .B2(new_n242), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n238), .A2(KEYINPUT28), .A3(new_n209), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT26), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n230), .A2(new_n246), .A3(new_n231), .ZN(new_n247));
  INV_X1    g046(.A(new_n204), .ZN(new_n248));
  INV_X1    g047(.A(new_n203), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n248), .B1(new_n249), .B2(KEYINPUT26), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n226), .B1(new_n247), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n245), .A2(new_n251), .ZN(new_n252));
  AOI21_X1  g051(.A(KEYINPUT29), .B1(new_n236), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(G226gat), .A2(G233gat), .ZN(new_n254));
  XOR2_X1   g053(.A(new_n254), .B(KEYINPUT74), .Z(new_n255));
  OAI21_X1  g054(.A(KEYINPUT75), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT75), .ZN(new_n257));
  INV_X1    g056(.A(new_n255), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n224), .A2(new_n227), .ZN(new_n259));
  INV_X1    g058(.A(new_n212), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  AOI211_X1 g060(.A(new_n219), .B(new_n205), .C1(new_n232), .C2(KEYINPUT23), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  AOI22_X1  g062(.A1(new_n263), .A2(new_n220), .B1(new_n245), .B2(new_n251), .ZN(new_n264));
  OAI211_X1 g063(.A(new_n257), .B(new_n258), .C1(new_n264), .C2(KEYINPUT29), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n236), .A2(new_n252), .ZN(new_n266));
  INV_X1    g065(.A(new_n254), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n256), .A2(new_n265), .A3(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(G197gat), .B(G204gat), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT22), .ZN(new_n271));
  INV_X1    g070(.A(G211gat), .ZN(new_n272));
  INV_X1    g071(.A(G218gat), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n271), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n270), .A2(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(G211gat), .B(G218gat), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n276), .A2(new_n270), .A3(new_n274), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n280), .B(KEYINPUT73), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n202), .B1(new_n269), .B2(new_n281), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n258), .B1(new_n264), .B2(KEYINPUT29), .ZN(new_n283));
  AOI22_X1  g082(.A1(new_n283), .A2(KEYINPUT75), .B1(new_n267), .B2(new_n266), .ZN(new_n284));
  INV_X1    g083(.A(new_n281), .ZN(new_n285));
  NAND4_X1  g084(.A1(new_n284), .A2(KEYINPUT82), .A3(new_n265), .A4(new_n285), .ZN(new_n286));
  AOI22_X1  g085(.A1(new_n261), .A2(new_n262), .B1(new_n219), .B2(new_n218), .ZN(new_n287));
  INV_X1    g086(.A(new_n251), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n288), .B1(new_n243), .B2(new_n244), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n255), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n290), .B1(new_n253), .B2(new_n267), .ZN(new_n291));
  INV_X1    g090(.A(new_n280), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n282), .A2(new_n286), .A3(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(KEYINPUT37), .ZN(new_n295));
  XNOR2_X1  g094(.A(G8gat), .B(G36gat), .ZN(new_n296));
  XNOR2_X1  g095(.A(G64gat), .B(G92gat), .ZN(new_n297));
  XOR2_X1   g096(.A(new_n296), .B(new_n297), .Z(new_n298));
  NAND2_X1  g097(.A1(new_n269), .A2(new_n281), .ZN(new_n299));
  OAI211_X1 g098(.A(new_n290), .B(new_n280), .C1(new_n253), .C2(new_n267), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT37), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  AOI211_X1 g102(.A(KEYINPUT38), .B(new_n298), .C1(new_n299), .C2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n295), .A2(new_n304), .ZN(new_n305));
  XNOR2_X1  g104(.A(G1gat), .B(G29gat), .ZN(new_n306));
  XNOR2_X1  g105(.A(new_n306), .B(KEYINPUT0), .ZN(new_n307));
  XNOR2_X1  g106(.A(G57gat), .B(G85gat), .ZN(new_n308));
  XOR2_X1   g107(.A(new_n307), .B(new_n308), .Z(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT78), .ZN(new_n311));
  XNOR2_X1  g110(.A(G113gat), .B(G120gat), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n312), .A2(KEYINPUT1), .ZN(new_n313));
  XNOR2_X1  g112(.A(G127gat), .B(G134gat), .ZN(new_n314));
  OR2_X1    g113(.A1(KEYINPUT69), .A2(KEYINPUT1), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n313), .A2(new_n316), .ZN(new_n317));
  OAI211_X1 g116(.A(new_n314), .B(new_n315), .C1(new_n312), .C2(KEYINPUT1), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT77), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n317), .A2(KEYINPUT77), .A3(new_n318), .ZN(new_n322));
  XOR2_X1   g121(.A(G141gat), .B(G148gat), .Z(new_n323));
  NAND2_X1  g122(.A1(G155gat), .A2(G162gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(KEYINPUT2), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  NOR2_X1   g125(.A1(G155gat), .A2(G162gat), .ZN(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  AOI22_X1  g127(.A1(new_n324), .A2(new_n328), .B1(new_n325), .B2(KEYINPUT76), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n326), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(new_n324), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n331), .A2(new_n327), .ZN(new_n332));
  OAI211_X1 g131(.A(new_n323), .B(new_n325), .C1(new_n332), .C2(KEYINPUT76), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n330), .A2(new_n333), .A3(KEYINPUT3), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n321), .A2(new_n322), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n330), .A2(new_n333), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT3), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n311), .B1(new_n335), .B2(new_n339), .ZN(new_n340));
  AND3_X1   g139(.A1(new_n317), .A2(KEYINPUT77), .A3(new_n318), .ZN(new_n341));
  AOI21_X1  g140(.A(KEYINPUT77), .B1(new_n317), .B2(new_n318), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND4_X1  g142(.A1(new_n343), .A2(KEYINPUT78), .A3(new_n338), .A4(new_n334), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n340), .A2(new_n344), .ZN(new_n345));
  AOI22_X1  g144(.A1(new_n330), .A2(new_n333), .B1(new_n317), .B2(new_n318), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT80), .ZN(new_n347));
  XNOR2_X1  g146(.A(KEYINPUT79), .B(KEYINPUT4), .ZN(new_n348));
  AND3_X1   g147(.A1(new_n346), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n346), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(KEYINPUT4), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n347), .B1(new_n346), .B2(new_n348), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n349), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(G225gat), .A2(G233gat), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n355), .A2(KEYINPUT5), .ZN(new_n356));
  AND3_X1   g155(.A1(new_n345), .A2(new_n353), .A3(new_n356), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n336), .A2(KEYINPUT4), .A3(new_n319), .ZN(new_n358));
  INV_X1    g157(.A(new_n348), .ZN(new_n359));
  OAI211_X1 g158(.A(new_n358), .B(new_n354), .C1(new_n346), .C2(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n360), .B1(new_n340), .B2(new_n344), .ZN(new_n361));
  INV_X1    g160(.A(new_n336), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n346), .B1(new_n343), .B2(new_n362), .ZN(new_n363));
  OAI21_X1  g162(.A(KEYINPUT5), .B1(new_n363), .B2(new_n354), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n361), .A2(new_n364), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n310), .B1(new_n357), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n345), .A2(new_n353), .ZN(new_n367));
  INV_X1    g166(.A(new_n356), .ZN(new_n368));
  OAI221_X1 g167(.A(new_n309), .B1(new_n361), .B2(new_n364), .C1(new_n367), .C2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT6), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n366), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  OAI211_X1 g170(.A(KEYINPUT6), .B(new_n310), .C1(new_n357), .C2(new_n365), .ZN(new_n372));
  AND2_X1   g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n298), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n285), .B1(new_n284), .B2(new_n265), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n374), .B1(new_n375), .B2(new_n302), .ZN(new_n376));
  INV_X1    g175(.A(new_n300), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n377), .B1(new_n269), .B2(new_n281), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n378), .A2(new_n301), .ZN(new_n379));
  OAI21_X1  g178(.A(KEYINPUT38), .B1(new_n376), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n378), .A2(new_n298), .ZN(new_n381));
  NAND4_X1  g180(.A1(new_n305), .A2(new_n373), .A3(new_n380), .A4(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(G228gat), .ZN(new_n383));
  INV_X1    g182(.A(G233gat), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  AOI21_X1  g184(.A(KEYINPUT29), .B1(new_n278), .B2(new_n279), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT81), .ZN(new_n387));
  AND2_X1   g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n337), .B1(new_n386), .B2(new_n387), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n362), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT29), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n338), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(new_n292), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n385), .B1(new_n390), .B2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n281), .A2(new_n392), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n362), .B1(new_n386), .B2(KEYINPUT3), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n396), .A2(new_n385), .A3(new_n397), .ZN(new_n398));
  XOR2_X1   g197(.A(KEYINPUT31), .B(G50gat), .Z(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n395), .A2(new_n398), .A3(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n398), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n399), .B1(new_n402), .B2(new_n394), .ZN(new_n403));
  XNOR2_X1  g202(.A(G78gat), .B(G106gat), .ZN(new_n404));
  XNOR2_X1  g203(.A(new_n404), .B(G22gat), .ZN(new_n405));
  AND3_X1   g204(.A1(new_n401), .A2(new_n403), .A3(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n405), .B1(new_n401), .B2(new_n403), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT39), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n367), .A2(new_n409), .A3(new_n355), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n354), .B1(new_n345), .B2(new_n353), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n409), .B1(new_n363), .B2(new_n354), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  OAI211_X1 g212(.A(new_n410), .B(new_n309), .C1(new_n411), .C2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT40), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n310), .B1(new_n411), .B2(new_n409), .ZN(new_n417));
  OAI211_X1 g216(.A(new_n417), .B(KEYINPUT40), .C1(new_n411), .C2(new_n413), .ZN(new_n418));
  AND3_X1   g217(.A1(new_n416), .A2(new_n366), .A3(new_n418), .ZN(new_n419));
  AND2_X1   g218(.A1(new_n298), .A2(KEYINPUT30), .ZN(new_n420));
  AND3_X1   g219(.A1(new_n299), .A2(new_n300), .A3(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n298), .B1(new_n299), .B2(new_n300), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(KEYINPUT30), .B1(new_n378), .B2(new_n298), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n419), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n382), .A2(new_n408), .A3(new_n427), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n319), .B1(new_n287), .B2(new_n289), .ZN(new_n429));
  NAND2_X1  g228(.A1(G227gat), .A2(G233gat), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n319), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n236), .A2(new_n252), .A3(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n429), .A2(new_n431), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(KEYINPUT32), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT33), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  XOR2_X1   g236(.A(G15gat), .B(G43gat), .Z(new_n438));
  XNOR2_X1  g237(.A(G71gat), .B(G99gat), .ZN(new_n439));
  XNOR2_X1  g238(.A(new_n438), .B(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n435), .A2(new_n437), .A3(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(new_n440), .ZN(new_n442));
  OAI211_X1 g241(.A(new_n434), .B(KEYINPUT32), .C1(new_n436), .C2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT71), .ZN(new_n445));
  XNOR2_X1  g244(.A(KEYINPUT70), .B(KEYINPUT34), .ZN(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  AND2_X1   g246(.A1(new_n429), .A2(new_n433), .ZN(new_n448));
  OAI211_X1 g247(.A(new_n445), .B(new_n447), .C1(new_n448), .C2(new_n431), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n431), .B1(new_n429), .B2(new_n433), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT34), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  OAI21_X1  g251(.A(KEYINPUT71), .B1(new_n450), .B2(new_n446), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n449), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n444), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(KEYINPUT72), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT72), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n444), .A2(new_n454), .A3(new_n457), .ZN(new_n458));
  AND2_X1   g257(.A1(new_n453), .A2(new_n452), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n459), .A2(new_n441), .A3(new_n443), .A4(new_n449), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n456), .A2(KEYINPUT36), .A3(new_n458), .A4(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT36), .ZN(new_n462));
  INV_X1    g261(.A(new_n455), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n444), .A2(new_n454), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n462), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n371), .A2(new_n372), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n466), .A2(new_n423), .A3(new_n425), .ZN(new_n467));
  INV_X1    g266(.A(new_n408), .ZN(new_n468));
  AOI22_X1  g267(.A1(new_n461), .A2(new_n465), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n456), .A2(new_n408), .A3(new_n460), .A4(new_n458), .ZN(new_n470));
  OAI21_X1  g269(.A(KEYINPUT35), .B1(new_n470), .B2(new_n467), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n463), .A2(new_n464), .ZN(new_n472));
  NOR3_X1   g271(.A1(new_n424), .A2(new_n421), .A3(new_n422), .ZN(new_n473));
  NOR3_X1   g272(.A1(new_n406), .A2(new_n407), .A3(KEYINPUT35), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n472), .A2(new_n473), .A3(new_n466), .A4(new_n474), .ZN(new_n475));
  AOI22_X1  g274(.A1(new_n428), .A2(new_n469), .B1(new_n471), .B2(new_n475), .ZN(new_n476));
  XNOR2_X1  g275(.A(G113gat), .B(G141gat), .ZN(new_n477));
  XNOR2_X1  g276(.A(new_n477), .B(G197gat), .ZN(new_n478));
  XOR2_X1   g277(.A(KEYINPUT11), .B(G169gat), .Z(new_n479));
  XNOR2_X1  g278(.A(new_n478), .B(new_n479), .ZN(new_n480));
  XOR2_X1   g279(.A(new_n480), .B(KEYINPUT12), .Z(new_n481));
  INV_X1    g280(.A(G1gat), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(KEYINPUT16), .ZN(new_n483));
  INV_X1    g282(.A(G15gat), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(G22gat), .ZN(new_n485));
  INV_X1    g284(.A(G22gat), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(G15gat), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n483), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(G1gat), .B1(new_n485), .B2(new_n487), .ZN(new_n490));
  OAI21_X1  g289(.A(G8gat), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(G8gat), .ZN(new_n492));
  AND2_X1   g291(.A1(new_n485), .A2(new_n487), .ZN(new_n493));
  OAI211_X1 g292(.A(new_n492), .B(new_n488), .C1(new_n493), .C2(G1gat), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  OR2_X1    g295(.A1(G43gat), .A2(G50gat), .ZN(new_n497));
  NAND2_X1  g296(.A1(G43gat), .A2(G50gat), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n497), .A2(KEYINPUT83), .A3(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT83), .ZN(new_n500));
  AND2_X1   g299(.A1(G43gat), .A2(G50gat), .ZN(new_n501));
  NOR2_X1   g300(.A1(G43gat), .A2(G50gat), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n499), .A2(new_n503), .A3(KEYINPUT15), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT15), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n497), .A2(new_n505), .A3(new_n498), .ZN(new_n506));
  INV_X1    g305(.A(G29gat), .ZN(new_n507));
  INV_X1    g306(.A(G36gat), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n507), .A2(new_n508), .A3(KEYINPUT14), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT14), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n510), .B1(G29gat), .B2(G36gat), .ZN(new_n511));
  NAND2_X1  g310(.A1(G29gat), .A2(G36gat), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n509), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n504), .A2(new_n506), .A3(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT17), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n513), .A2(new_n499), .A3(new_n503), .A4(KEYINPUT15), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n516), .B1(new_n515), .B2(new_n517), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n496), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT18), .ZN(new_n522));
  NAND2_X1  g321(.A1(G229gat), .A2(G233gat), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  AND3_X1   g323(.A1(new_n499), .A2(new_n503), .A3(KEYINPUT15), .ZN(new_n525));
  NAND4_X1  g324(.A1(new_n506), .A2(new_n511), .A3(new_n509), .A4(new_n512), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n517), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  AOI211_X1 g326(.A(new_n522), .B(new_n524), .C1(new_n527), .C2(new_n495), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n521), .A2(KEYINPUT84), .A3(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT84), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n527), .A2(KEYINPUT17), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n495), .B1(new_n531), .B2(new_n518), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n527), .A2(new_n495), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n533), .A2(KEYINPUT18), .A3(new_n523), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n530), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  AND2_X1   g334(.A1(new_n529), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n533), .A2(new_n523), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n522), .B1(new_n532), .B2(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n527), .B(new_n495), .ZN(new_n539));
  XOR2_X1   g338(.A(new_n523), .B(KEYINPUT13), .Z(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n538), .A2(new_n541), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n481), .B1(new_n536), .B2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(new_n481), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n529), .A2(new_n535), .ZN(new_n545));
  NAND4_X1  g344(.A1(new_n544), .A2(new_n545), .A3(new_n538), .A4(new_n541), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n543), .A2(KEYINPUT85), .A3(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT85), .ZN(new_n548));
  OAI211_X1 g347(.A(new_n548), .B(new_n481), .C1(new_n536), .C2(new_n542), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n476), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT96), .ZN(new_n552));
  XNOR2_X1  g351(.A(G190gat), .B(G218gat), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT8), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n554), .B1(G99gat), .B2(G106gat), .ZN(new_n555));
  XNOR2_X1  g354(.A(KEYINPUT91), .B(G85gat), .ZN(new_n556));
  INV_X1    g355(.A(G92gat), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n555), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(G99gat), .A2(G106gat), .ZN(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  NOR2_X1   g359(.A1(G99gat), .A2(G106gat), .ZN(new_n561));
  OAI21_X1  g360(.A(KEYINPUT92), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  OR2_X1    g361(.A1(G99gat), .A2(G106gat), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT92), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n563), .A2(new_n564), .A3(new_n559), .ZN(new_n565));
  NAND2_X1  g364(.A1(G85gat), .A2(G92gat), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(KEYINPUT7), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT7), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n568), .A2(G85gat), .A3(G92gat), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  NAND4_X1  g369(.A1(new_n558), .A2(new_n562), .A3(new_n565), .A4(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(G85gat), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(KEYINPUT91), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT91), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n574), .A2(G85gat), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n573), .A2(new_n575), .A3(new_n557), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n559), .A2(KEYINPUT8), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n576), .A2(new_n570), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n565), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  AND3_X1   g379(.A1(new_n571), .A2(KEYINPUT93), .A3(new_n580), .ZN(new_n581));
  AOI21_X1  g380(.A(KEYINPUT93), .B1(new_n571), .B2(new_n580), .ZN(new_n582));
  OAI21_X1  g381(.A(KEYINPUT94), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n531), .A2(new_n518), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT93), .ZN(new_n585));
  AND2_X1   g384(.A1(new_n578), .A2(new_n579), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n578), .A2(new_n579), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n585), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT94), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n571), .A2(KEYINPUT93), .A3(new_n580), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  AND3_X1   g390(.A1(new_n583), .A2(new_n584), .A3(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n588), .A2(new_n527), .A3(new_n590), .ZN(new_n593));
  NAND2_X1  g392(.A1(G232gat), .A2(G233gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n594), .B(KEYINPUT90), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT41), .ZN(new_n596));
  OR2_X1    g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  OAI211_X1 g397(.A(KEYINPUT95), .B(new_n553), .C1(new_n592), .C2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n598), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n583), .A2(new_n591), .A3(new_n584), .ZN(new_n601));
  INV_X1    g400(.A(new_n553), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n600), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n595), .A2(new_n596), .ZN(new_n604));
  XNOR2_X1  g403(.A(G134gat), .B(G162gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n604), .B(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n599), .A2(new_n603), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n600), .A2(new_n601), .ZN(new_n609));
  AOI21_X1  g408(.A(KEYINPUT95), .B1(new_n609), .B2(new_n553), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n552), .B1(new_n608), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n609), .A2(new_n553), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT95), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  AND2_X1   g413(.A1(new_n603), .A2(new_n607), .ZN(new_n615));
  NAND4_X1  g414(.A1(new_n614), .A2(new_n615), .A3(KEYINPUT96), .A4(new_n599), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n612), .A2(new_n603), .ZN(new_n617));
  AOI22_X1  g416(.A1(new_n611), .A2(new_n616), .B1(new_n617), .B2(new_n606), .ZN(new_n618));
  INV_X1    g417(.A(G57gat), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n619), .A2(G64gat), .ZN(new_n620));
  INV_X1    g419(.A(G64gat), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n621), .A2(G57gat), .ZN(new_n622));
  OAI21_X1  g421(.A(KEYINPUT9), .B1(new_n620), .B2(new_n622), .ZN(new_n623));
  OR2_X1    g422(.A1(G71gat), .A2(G78gat), .ZN(new_n624));
  NAND2_X1  g423(.A1(G71gat), .A2(G78gat), .ZN(new_n625));
  AND2_X1   g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  OAI21_X1  g425(.A(KEYINPUT86), .B1(new_n619), .B2(G64gat), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT86), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n628), .A2(new_n621), .A3(G57gat), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n619), .A2(G64gat), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n627), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT9), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n625), .B1(new_n624), .B2(new_n632), .ZN(new_n633));
  AOI22_X1  g432(.A1(new_n623), .A2(new_n626), .B1(new_n631), .B2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT21), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  XOR2_X1   g436(.A(KEYINPUT89), .B(KEYINPUT19), .Z(new_n638));
  XNOR2_X1  g437(.A(new_n637), .B(new_n638), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n495), .B1(KEYINPUT21), .B2(new_n634), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n639), .B(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(G231gat), .A2(G233gat), .ZN(new_n642));
  XOR2_X1   g441(.A(new_n642), .B(KEYINPUT88), .Z(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(KEYINPUT87), .ZN(new_n644));
  XNOR2_X1  g443(.A(G127gat), .B(G155gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(KEYINPUT20), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n644), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(G183gat), .B(G211gat), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n641), .B(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n618), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(KEYINPUT97), .B(KEYINPUT10), .ZN(new_n653));
  AND3_X1   g452(.A1(new_n571), .A2(new_n634), .A3(new_n580), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n634), .B1(new_n571), .B2(new_n580), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n653), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  AND2_X1   g455(.A1(new_n634), .A2(KEYINPUT10), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n588), .A2(new_n590), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(G230gat), .A2(G233gat), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  OR3_X1    g460(.A1(new_n654), .A2(new_n655), .A3(new_n660), .ZN(new_n662));
  XNOR2_X1  g461(.A(G120gat), .B(G148gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(G176gat), .B(G204gat), .ZN(new_n664));
  XOR2_X1   g463(.A(new_n663), .B(new_n664), .Z(new_n665));
  AND3_X1   g464(.A1(new_n661), .A2(new_n662), .A3(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n661), .A2(new_n662), .ZN(new_n668));
  INV_X1    g467(.A(new_n665), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n652), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n551), .A2(new_n672), .ZN(new_n673));
  AND3_X1   g472(.A1(new_n371), .A2(new_n372), .A3(KEYINPUT98), .ZN(new_n674));
  AOI21_X1  g473(.A(KEYINPUT98), .B1(new_n371), .B2(new_n372), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n673), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g477(.A(KEYINPUT99), .B(G1gat), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n678), .B(new_n679), .ZN(G1324gat));
  NOR2_X1   g479(.A1(new_n673), .A2(new_n473), .ZN(new_n681));
  OR3_X1    g480(.A1(new_n681), .A2(KEYINPUT100), .A3(new_n492), .ZN(new_n682));
  OAI21_X1  g481(.A(KEYINPUT100), .B1(new_n681), .B2(new_n492), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT42), .ZN(new_n684));
  XOR2_X1   g483(.A(KEYINPUT16), .B(G8gat), .Z(new_n685));
  AOI21_X1  g484(.A(new_n684), .B1(new_n681), .B2(new_n685), .ZN(new_n686));
  AND3_X1   g485(.A1(new_n681), .A2(new_n684), .A3(new_n685), .ZN(new_n687));
  OAI211_X1 g486(.A(new_n682), .B(new_n683), .C1(new_n686), .C2(new_n687), .ZN(G1325gat));
  NAND2_X1  g487(.A1(new_n461), .A2(new_n465), .ZN(new_n689));
  OAI21_X1  g488(.A(G15gat), .B1(new_n673), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n472), .A2(new_n484), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n690), .B1(new_n673), .B2(new_n691), .ZN(G1326gat));
  OR3_X1    g491(.A1(new_n673), .A2(KEYINPUT101), .A3(new_n408), .ZN(new_n693));
  OAI21_X1  g492(.A(KEYINPUT101), .B1(new_n673), .B2(new_n408), .ZN(new_n694));
  XNOR2_X1  g493(.A(KEYINPUT43), .B(G22gat), .ZN(new_n695));
  AND3_X1   g494(.A1(new_n693), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n695), .B1(new_n693), .B2(new_n694), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n696), .A2(new_n697), .ZN(G1327gat));
  NAND2_X1  g497(.A1(new_n467), .A2(new_n468), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT38), .ZN(new_n700));
  OAI211_X1 g499(.A(new_n700), .B(new_n374), .C1(new_n375), .C2(new_n302), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n701), .B1(KEYINPUT37), .B2(new_n294), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n371), .A2(new_n372), .A3(new_n381), .ZN(new_n703));
  OAI21_X1  g502(.A(KEYINPUT37), .B1(new_n375), .B2(new_n377), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n298), .B1(new_n299), .B2(new_n303), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n700), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NOR3_X1   g505(.A1(new_n702), .A2(new_n703), .A3(new_n706), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n416), .A2(new_n366), .A3(new_n418), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n408), .B1(new_n473), .B2(new_n708), .ZN(new_n709));
  OAI211_X1 g508(.A(new_n689), .B(new_n699), .C1(new_n707), .C2(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n471), .A2(new_n475), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(new_n550), .ZN(new_n713));
  INV_X1    g512(.A(new_n671), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(new_n650), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n618), .A2(new_n715), .ZN(new_n716));
  XOR2_X1   g515(.A(new_n716), .B(KEYINPUT102), .Z(new_n717));
  AND3_X1   g516(.A1(new_n712), .A2(new_n713), .A3(new_n717), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n718), .A2(new_n507), .A3(new_n676), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n719), .B(KEYINPUT45), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT44), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n721), .B1(new_n476), .B2(new_n618), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n617), .A2(new_n606), .ZN(new_n723));
  AOI211_X1 g522(.A(new_n613), .B(new_n602), .C1(new_n600), .C2(new_n601), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n603), .A2(new_n607), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  AOI21_X1  g525(.A(KEYINPUT96), .B1(new_n726), .B2(new_n614), .ZN(new_n727));
  NOR3_X1   g526(.A1(new_n608), .A2(new_n552), .A3(new_n610), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n723), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n712), .A2(KEYINPUT44), .A3(new_n729), .ZN(new_n730));
  AND2_X1   g529(.A1(new_n722), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n715), .A2(new_n550), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(G29gat), .B1(new_n733), .B2(new_n677), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n720), .A2(new_n734), .ZN(G1328gat));
  NAND3_X1  g534(.A1(new_n718), .A2(new_n508), .A3(new_n426), .ZN(new_n736));
  XOR2_X1   g535(.A(KEYINPUT103), .B(KEYINPUT46), .Z(new_n737));
  XNOR2_X1  g536(.A(new_n736), .B(new_n737), .ZN(new_n738));
  OAI21_X1  g537(.A(G36gat), .B1(new_n733), .B2(new_n473), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(G1329gat));
  INV_X1    g539(.A(new_n689), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n722), .A2(new_n730), .A3(new_n741), .A4(new_n732), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT104), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(G43gat), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n742), .A2(new_n743), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n551), .A2(new_n717), .ZN(new_n748));
  INV_X1    g547(.A(new_n472), .ZN(new_n749));
  OR3_X1    g548(.A1(new_n748), .A2(G43gat), .A3(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(KEYINPUT47), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n742), .A2(G43gat), .ZN(new_n752));
  AND2_X1   g551(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  OAI22_X1  g552(.A1(new_n747), .A2(new_n751), .B1(new_n753), .B2(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g553(.A(KEYINPUT105), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n408), .B1(new_n718), .B2(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n748), .A2(KEYINPUT105), .ZN(new_n757));
  AOI21_X1  g556(.A(G50gat), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT48), .ZN(new_n760));
  AND2_X1   g559(.A1(new_n468), .A2(G50gat), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n731), .A2(new_n732), .A3(new_n761), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n759), .A2(new_n760), .A3(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(new_n762), .ZN(new_n764));
  OAI21_X1  g563(.A(KEYINPUT48), .B1(new_n764), .B2(new_n758), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n763), .A2(new_n765), .ZN(G1331gat));
  NOR4_X1   g565(.A1(new_n476), .A2(new_n713), .A3(new_n652), .A4(new_n714), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(new_n676), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g568(.A1(new_n378), .A2(new_n420), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n770), .B1(new_n298), .B2(new_n378), .ZN(new_n771));
  OAI21_X1  g570(.A(KEYINPUT106), .B1(new_n771), .B2(new_n424), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT106), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n423), .A2(new_n773), .A3(new_n425), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n767), .A2(new_n775), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n776), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n777));
  XOR2_X1   g576(.A(KEYINPUT49), .B(G64gat), .Z(new_n778));
  OAI21_X1  g577(.A(new_n777), .B1(new_n776), .B2(new_n778), .ZN(G1333gat));
  NAND2_X1  g578(.A1(new_n767), .A2(new_n741), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n749), .A2(G71gat), .ZN(new_n781));
  AOI22_X1  g580(.A1(new_n780), .A2(G71gat), .B1(new_n767), .B2(new_n781), .ZN(new_n782));
  XNOR2_X1  g581(.A(KEYINPUT107), .B(KEYINPUT50), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n782), .B(new_n783), .ZN(G1334gat));
  NAND2_X1  g583(.A1(new_n767), .A2(new_n468), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n785), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g585(.A1(new_n713), .A2(new_n651), .ZN(new_n787));
  INV_X1    g586(.A(new_n787), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n788), .A2(new_n714), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n731), .A2(new_n789), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n790), .A2(new_n677), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n712), .A2(new_n729), .A3(new_n787), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT51), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n618), .B1(new_n710), .B2(new_n711), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n795), .A2(KEYINPUT51), .A3(new_n787), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n676), .A2(new_n556), .A3(new_n671), .ZN(new_n799));
  OAI22_X1  g598(.A1(new_n791), .A2(new_n556), .B1(new_n798), .B2(new_n799), .ZN(G1336gat));
  NAND4_X1  g599(.A1(new_n722), .A2(new_n730), .A3(new_n426), .A4(new_n789), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(G92gat), .ZN(new_n802));
  INV_X1    g601(.A(new_n775), .ZN(new_n803));
  NOR3_X1   g602(.A1(new_n803), .A2(G92gat), .A3(new_n714), .ZN(new_n804));
  NOR4_X1   g603(.A1(new_n476), .A2(new_n793), .A3(new_n618), .A4(new_n788), .ZN(new_n805));
  AOI21_X1  g604(.A(KEYINPUT51), .B1(new_n795), .B2(new_n787), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n804), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n802), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(KEYINPUT52), .ZN(new_n809));
  AOI21_X1  g608(.A(KEYINPUT52), .B1(new_n797), .B2(new_n804), .ZN(new_n810));
  NAND4_X1  g609(.A1(new_n722), .A2(new_n730), .A3(new_n775), .A4(new_n789), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(G92gat), .ZN(new_n812));
  AOI21_X1  g611(.A(KEYINPUT108), .B1(new_n810), .B2(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT52), .ZN(new_n814));
  AND4_X1   g613(.A1(KEYINPUT108), .A2(new_n812), .A3(new_n814), .A4(new_n807), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n809), .B1(new_n813), .B2(new_n815), .ZN(G1337gat));
  XNOR2_X1  g615(.A(KEYINPUT109), .B(G99gat), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n817), .B1(new_n790), .B2(new_n689), .ZN(new_n818));
  OR3_X1    g617(.A1(new_n749), .A2(new_n714), .A3(new_n817), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n818), .B1(new_n798), .B2(new_n819), .ZN(G1338gat));
  NOR3_X1   g619(.A1(new_n408), .A2(G106gat), .A3(new_n714), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n797), .A2(new_n821), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n722), .A2(new_n730), .A3(new_n468), .A4(new_n789), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(G106gat), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n822), .A2(KEYINPUT110), .A3(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(KEYINPUT53), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT53), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n822), .A2(KEYINPUT110), .A3(new_n824), .A4(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n826), .A2(new_n828), .ZN(G1339gat));
  AOI21_X1  g628(.A(new_n523), .B1(new_n521), .B2(new_n533), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n539), .A2(new_n540), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n480), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  AND2_X1   g631(.A1(new_n546), .A2(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(new_n660), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n656), .A2(new_n834), .A3(new_n658), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(KEYINPUT111), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT111), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n656), .A2(new_n658), .A3(new_n837), .A4(new_n834), .ZN(new_n838));
  NAND4_X1  g637(.A1(new_n836), .A2(new_n661), .A3(KEYINPUT54), .A4(new_n838), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n834), .B1(new_n656), .B2(new_n658), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT54), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n665), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT55), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  AOI211_X1 g644(.A(new_n844), .B(new_n665), .C1(new_n840), .C2(new_n841), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n666), .B1(new_n846), .B2(new_n839), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n833), .A2(new_n845), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n729), .A2(new_n848), .ZN(new_n849));
  NAND4_X1  g648(.A1(new_n547), .A2(new_n845), .A3(new_n847), .A4(new_n549), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n611), .A2(new_n616), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n833), .A2(new_n671), .ZN(new_n852));
  NAND4_X1  g651(.A1(new_n850), .A2(new_n851), .A3(new_n723), .A4(new_n852), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n849), .A2(new_n650), .A3(new_n853), .ZN(new_n854));
  NAND4_X1  g653(.A1(new_n618), .A2(new_n550), .A3(new_n651), .A4(new_n714), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(KEYINPUT112), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT112), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n854), .A2(new_n858), .A3(new_n855), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n677), .A2(new_n470), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n860), .A2(new_n803), .A3(new_n861), .ZN(new_n862));
  OR3_X1    g661(.A1(new_n862), .A2(G113gat), .A3(new_n550), .ZN(new_n863));
  NOR3_X1   g662(.A1(new_n677), .A2(new_n775), .A3(new_n749), .ZN(new_n864));
  NAND4_X1  g663(.A1(new_n860), .A2(new_n408), .A3(new_n713), .A4(new_n864), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n865), .A2(KEYINPUT113), .A3(G113gat), .ZN(new_n866));
  INV_X1    g665(.A(new_n866), .ZN(new_n867));
  AOI21_X1  g666(.A(KEYINPUT113), .B1(new_n865), .B2(G113gat), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n863), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(KEYINPUT114), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT114), .ZN(new_n871));
  OAI211_X1 g670(.A(new_n871), .B(new_n863), .C1(new_n867), .C2(new_n868), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n870), .A2(new_n872), .ZN(G1340gat));
  AND3_X1   g672(.A1(new_n854), .A2(new_n858), .A3(new_n855), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n858), .B1(new_n854), .B2(new_n855), .ZN(new_n875));
  OAI211_X1 g674(.A(new_n408), .B(new_n864), .C1(new_n874), .C2(new_n875), .ZN(new_n876));
  OAI21_X1  g675(.A(G120gat), .B1(new_n876), .B2(new_n714), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n714), .A2(G120gat), .ZN(new_n878));
  XNOR2_X1  g677(.A(new_n878), .B(KEYINPUT115), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n877), .B1(new_n862), .B2(new_n879), .ZN(new_n880));
  XOR2_X1   g679(.A(new_n880), .B(KEYINPUT116), .Z(G1341gat));
  INV_X1    g680(.A(G127gat), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n650), .A2(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(new_n883), .ZN(new_n884));
  OR3_X1    g683(.A1(new_n876), .A2(KEYINPUT117), .A3(new_n884), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n882), .B1(new_n862), .B2(new_n650), .ZN(new_n886));
  OAI21_X1  g685(.A(KEYINPUT117), .B1(new_n876), .B2(new_n884), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT118), .ZN(new_n889));
  XNOR2_X1  g688(.A(new_n888), .B(new_n889), .ZN(G1342gat));
  OAI21_X1  g689(.A(G134gat), .B1(new_n876), .B2(new_n618), .ZN(new_n891));
  NOR3_X1   g690(.A1(new_n426), .A2(new_n618), .A3(G134gat), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n860), .A2(new_n861), .A3(new_n892), .ZN(new_n893));
  AND3_X1   g692(.A1(new_n893), .A2(KEYINPUT119), .A3(KEYINPUT56), .ZN(new_n894));
  AOI21_X1  g693(.A(KEYINPUT119), .B1(new_n893), .B2(KEYINPUT56), .ZN(new_n895));
  OAI221_X1 g694(.A(new_n891), .B1(KEYINPUT56), .B2(new_n893), .C1(new_n894), .C2(new_n895), .ZN(G1343gat));
  NAND4_X1  g695(.A1(new_n689), .A2(new_n676), .A3(new_n772), .A4(new_n774), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT120), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND4_X1  g698(.A1(new_n803), .A2(KEYINPUT120), .A3(new_n689), .A4(new_n676), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n856), .A2(new_n468), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n901), .B1(KEYINPUT57), .B2(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT57), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n860), .A2(new_n904), .A3(new_n468), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n713), .A2(G141gat), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n874), .A2(new_n875), .ZN(new_n908));
  NOR4_X1   g707(.A1(new_n908), .A2(new_n408), .A3(new_n550), .A4(new_n897), .ZN(new_n909));
  OAI22_X1  g708(.A1(new_n906), .A2(new_n907), .B1(new_n909), .B2(G141gat), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT58), .ZN(new_n911));
  XNOR2_X1  g710(.A(new_n910), .B(new_n911), .ZN(G1344gat));
  INV_X1    g711(.A(G148gat), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n913), .A2(KEYINPUT59), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n914), .B1(new_n906), .B2(new_n714), .ZN(new_n915));
  AOI21_X1  g714(.A(KEYINPUT57), .B1(new_n856), .B2(new_n468), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n408), .A2(new_n904), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n916), .B1(new_n860), .B2(new_n917), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n899), .A2(new_n671), .A3(new_n900), .ZN(new_n919));
  OAI21_X1  g718(.A(G148gat), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  AOI21_X1  g719(.A(KEYINPUT121), .B1(new_n920), .B2(KEYINPUT59), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n917), .B1(new_n874), .B2(new_n875), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n902), .A2(new_n904), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n919), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  OAI211_X1 g723(.A(KEYINPUT121), .B(KEYINPUT59), .C1(new_n924), .C2(new_n913), .ZN(new_n925));
  INV_X1    g724(.A(new_n925), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n915), .B1(new_n921), .B2(new_n926), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n908), .A2(new_n408), .ZN(new_n928));
  INV_X1    g727(.A(new_n897), .ZN(new_n929));
  NAND4_X1  g728(.A1(new_n928), .A2(new_n913), .A3(new_n671), .A4(new_n929), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n927), .A2(new_n930), .ZN(G1345gat));
  OAI21_X1  g730(.A(G155gat), .B1(new_n906), .B2(new_n650), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n650), .A2(G155gat), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n928), .A2(new_n929), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT122), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n932), .A2(KEYINPUT122), .A3(new_n934), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(new_n938), .ZN(G1346gat));
  OAI21_X1  g738(.A(G162gat), .B1(new_n906), .B2(new_n618), .ZN(new_n940));
  NOR3_X1   g739(.A1(new_n426), .A2(new_n618), .A3(G162gat), .ZN(new_n941));
  NAND4_X1  g740(.A1(new_n928), .A2(new_n689), .A3(new_n676), .A4(new_n941), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n940), .A2(new_n942), .ZN(G1347gat));
  OAI21_X1  g742(.A(KEYINPUT123), .B1(new_n908), .B2(new_n676), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT123), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n860), .A2(new_n945), .A3(new_n677), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n803), .A2(new_n470), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n550), .A2(G169gat), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n947), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n677), .A2(new_n426), .A3(new_n472), .ZN(new_n951));
  INV_X1    g750(.A(new_n951), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n860), .A2(new_n408), .A3(new_n952), .ZN(new_n953));
  OAI21_X1  g752(.A(G169gat), .B1(new_n953), .B2(new_n550), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n950), .A2(new_n954), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT124), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n950), .A2(KEYINPUT124), .A3(new_n954), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(G1348gat));
  NAND2_X1  g758(.A1(new_n671), .A2(G176gat), .ZN(new_n960));
  NOR2_X1   g759(.A1(new_n953), .A2(new_n960), .ZN(new_n961));
  XNOR2_X1  g760(.A(new_n961), .B(KEYINPUT125), .ZN(new_n962));
  INV_X1    g761(.A(G176gat), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n947), .A2(new_n671), .A3(new_n948), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n962), .B1(new_n963), .B2(new_n964), .ZN(G1349gat));
  NAND4_X1  g764(.A1(new_n947), .A2(new_n238), .A3(new_n651), .A4(new_n948), .ZN(new_n966));
  OAI21_X1  g765(.A(G183gat), .B1(new_n953), .B2(new_n650), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n968), .A2(KEYINPUT60), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT60), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n966), .A2(new_n970), .A3(new_n967), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n969), .A2(new_n971), .ZN(G1350gat));
  OAI21_X1  g771(.A(G190gat), .B1(new_n953), .B2(new_n618), .ZN(new_n973));
  XNOR2_X1  g772(.A(new_n973), .B(KEYINPUT61), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n947), .A2(new_n948), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n729), .A2(new_n209), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n974), .B1(new_n975), .B2(new_n976), .ZN(G1351gat));
  NAND3_X1  g776(.A1(new_n689), .A2(new_n775), .A3(new_n468), .ZN(new_n978));
  AOI21_X1  g777(.A(new_n978), .B1(new_n944), .B2(new_n946), .ZN(new_n979));
  AOI21_X1  g778(.A(G197gat), .B1(new_n979), .B2(new_n713), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n677), .A2(new_n426), .A3(new_n689), .ZN(new_n981));
  INV_X1    g780(.A(new_n981), .ZN(new_n982));
  INV_X1    g781(.A(new_n922), .ZN(new_n983));
  OAI21_X1  g782(.A(new_n982), .B1(new_n983), .B2(new_n916), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n713), .A2(G197gat), .ZN(new_n985));
  NOR2_X1   g784(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  OAI21_X1  g785(.A(KEYINPUT126), .B1(new_n980), .B2(new_n986), .ZN(new_n987));
  INV_X1    g786(.A(KEYINPUT126), .ZN(new_n988));
  OR3_X1    g787(.A1(new_n918), .A2(new_n981), .A3(new_n985), .ZN(new_n989));
  AOI211_X1 g788(.A(new_n550), .B(new_n978), .C1(new_n944), .C2(new_n946), .ZN(new_n990));
  OAI211_X1 g789(.A(new_n988), .B(new_n989), .C1(new_n990), .C2(G197gat), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n987), .A2(new_n991), .ZN(G1352gat));
  NOR2_X1   g791(.A1(new_n714), .A2(G204gat), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n979), .A2(new_n993), .ZN(new_n994));
  OAI211_X1 g793(.A(new_n671), .B(new_n982), .C1(new_n983), .C2(new_n916), .ZN(new_n995));
  AOI22_X1  g794(.A1(new_n994), .A2(KEYINPUT62), .B1(new_n995), .B2(G204gat), .ZN(new_n996));
  INV_X1    g795(.A(new_n993), .ZN(new_n997));
  AOI211_X1 g796(.A(new_n978), .B(new_n997), .C1(new_n944), .C2(new_n946), .ZN(new_n998));
  INV_X1    g797(.A(KEYINPUT62), .ZN(new_n999));
  AOI21_X1  g798(.A(KEYINPUT127), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  AND4_X1   g799(.A1(KEYINPUT127), .A2(new_n979), .A3(new_n999), .A4(new_n993), .ZN(new_n1001));
  OAI21_X1  g800(.A(new_n996), .B1(new_n1000), .B2(new_n1001), .ZN(G1353gat));
  NAND3_X1  g801(.A1(new_n979), .A2(new_n272), .A3(new_n651), .ZN(new_n1003));
  OAI211_X1 g802(.A(new_n651), .B(new_n982), .C1(new_n983), .C2(new_n916), .ZN(new_n1004));
  AND3_X1   g803(.A1(new_n1004), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1005));
  AOI21_X1  g804(.A(KEYINPUT63), .B1(new_n1004), .B2(G211gat), .ZN(new_n1006));
  OAI21_X1  g805(.A(new_n1003), .B1(new_n1005), .B2(new_n1006), .ZN(G1354gat));
  NAND3_X1  g806(.A1(new_n979), .A2(new_n273), .A3(new_n729), .ZN(new_n1008));
  OAI21_X1  g807(.A(G218gat), .B1(new_n984), .B2(new_n618), .ZN(new_n1009));
  NAND2_X1  g808(.A1(new_n1008), .A2(new_n1009), .ZN(G1355gat));
endmodule


