

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X2 U552 ( .A(n653), .ZN(n638) );
  OR2_X1 U553 ( .A1(n670), .A2(n669), .ZN(n688) );
  INV_X1 U554 ( .A(n695), .ZN(n679) );
  NAND2_X1 U555 ( .A1(n995), .A2(G137), .ZN(n527) );
  NOR2_X1 U556 ( .A1(G651), .A2(n574), .ZN(n791) );
  XOR2_X1 U557 ( .A(KEYINPUT65), .B(n522), .Z(n517) );
  AND2_X1 U558 ( .A1(n531), .A2(n530), .ZN(n518) );
  NOR2_X1 U559 ( .A1(n698), .A2(n697), .ZN(n519) );
  NOR2_X1 U560 ( .A1(n653), .A2(n602), .ZN(n604) );
  NOR2_X1 U561 ( .A1(n965), .A2(n607), .ZN(n618) );
  INV_X1 U562 ( .A(KEYINPUT94), .ZN(n616) );
  NOR2_X1 U563 ( .A1(n801), .A2(n631), .ZN(n633) );
  NOR2_X1 U564 ( .A1(n651), .A2(n650), .ZN(n652) );
  AND2_X1 U565 ( .A1(n688), .A2(n848), .ZN(n671) );
  NAND2_X1 U566 ( .A1(G8), .A2(n653), .ZN(n695) );
  AND2_X1 U567 ( .A1(n601), .A2(G40), .ZN(n701) );
  AND2_X2 U568 ( .A1(n521), .A2(G2105), .ZN(n991) );
  XNOR2_X1 U569 ( .A(KEYINPUT71), .B(KEYINPUT14), .ZN(n595) );
  INV_X1 U570 ( .A(G2104), .ZN(n521) );
  XNOR2_X1 U571 ( .A(n596), .B(n595), .ZN(n597) );
  INV_X1 U572 ( .A(KEYINPUT17), .ZN(n524) );
  NOR2_X2 U573 ( .A1(n521), .A2(G2105), .ZN(n996) );
  XOR2_X1 U574 ( .A(KEYINPUT1), .B(n535), .Z(n790) );
  OR2_X1 U575 ( .A1(n758), .A2(n757), .ZN(n759) );
  BUF_X1 U576 ( .A(n601), .Z(G160) );
  NAND2_X1 U577 ( .A1(G101), .A2(n996), .ZN(n520) );
  XOR2_X1 U578 ( .A(KEYINPUT23), .B(n520), .Z(n523) );
  NAND2_X1 U579 ( .A1(G125), .A2(n991), .ZN(n522) );
  NAND2_X1 U580 ( .A1(n523), .A2(n517), .ZN(n529) );
  NOR2_X1 U581 ( .A1(G2104), .A2(G2105), .ZN(n525) );
  XNOR2_X2 U582 ( .A(n525), .B(n524), .ZN(n995) );
  AND2_X1 U583 ( .A1(G2104), .A2(G2105), .ZN(n992) );
  NAND2_X1 U584 ( .A1(G113), .A2(n992), .ZN(n526) );
  NAND2_X1 U585 ( .A1(n527), .A2(n526), .ZN(n528) );
  NOR2_X1 U586 ( .A1(n529), .A2(n528), .ZN(n601) );
  NAND2_X1 U587 ( .A1(n995), .A2(G138), .ZN(n534) );
  NAND2_X1 U588 ( .A1(G126), .A2(n991), .ZN(n531) );
  NAND2_X1 U589 ( .A1(G114), .A2(n992), .ZN(n530) );
  NAND2_X1 U590 ( .A1(G102), .A2(n996), .ZN(n532) );
  AND2_X1 U591 ( .A1(n518), .A2(n532), .ZN(n533) );
  AND2_X1 U592 ( .A1(n534), .A2(n533), .ZN(G164) );
  INV_X1 U593 ( .A(G651), .ZN(n536) );
  NOR2_X1 U594 ( .A1(G543), .A2(n536), .ZN(n535) );
  NAND2_X1 U595 ( .A1(G65), .A2(n790), .ZN(n538) );
  XOR2_X1 U596 ( .A(G543), .B(KEYINPUT0), .Z(n574) );
  NOR2_X1 U597 ( .A1(n574), .A2(n536), .ZN(n787) );
  NAND2_X1 U598 ( .A1(G78), .A2(n787), .ZN(n537) );
  NAND2_X1 U599 ( .A1(n538), .A2(n537), .ZN(n541) );
  NOR2_X1 U600 ( .A1(G651), .A2(G543), .ZN(n786) );
  NAND2_X1 U601 ( .A1(G91), .A2(n786), .ZN(n539) );
  XNOR2_X1 U602 ( .A(KEYINPUT69), .B(n539), .ZN(n540) );
  NOR2_X1 U603 ( .A1(n541), .A2(n540), .ZN(n543) );
  NAND2_X1 U604 ( .A1(n791), .A2(G53), .ZN(n542) );
  NAND2_X1 U605 ( .A1(n543), .A2(n542), .ZN(G299) );
  XNOR2_X1 U606 ( .A(KEYINPUT68), .B(KEYINPUT9), .ZN(n548) );
  NAND2_X1 U607 ( .A1(G90), .A2(n786), .ZN(n545) );
  NAND2_X1 U608 ( .A1(G77), .A2(n787), .ZN(n544) );
  NAND2_X1 U609 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U610 ( .A(n546), .B(KEYINPUT67), .ZN(n547) );
  XNOR2_X1 U611 ( .A(n548), .B(n547), .ZN(n552) );
  NAND2_X1 U612 ( .A1(G64), .A2(n790), .ZN(n550) );
  NAND2_X1 U613 ( .A1(G52), .A2(n791), .ZN(n549) );
  NAND2_X1 U614 ( .A1(n550), .A2(n549), .ZN(n551) );
  NOR2_X1 U615 ( .A1(n552), .A2(n551), .ZN(G171) );
  INV_X1 U616 ( .A(G171), .ZN(G301) );
  NAND2_X1 U617 ( .A1(G89), .A2(n786), .ZN(n553) );
  XNOR2_X1 U618 ( .A(n553), .B(KEYINPUT74), .ZN(n554) );
  XNOR2_X1 U619 ( .A(n554), .B(KEYINPUT4), .ZN(n556) );
  NAND2_X1 U620 ( .A1(G76), .A2(n787), .ZN(n555) );
  NAND2_X1 U621 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U622 ( .A(n557), .B(KEYINPUT5), .ZN(n562) );
  NAND2_X1 U623 ( .A1(G63), .A2(n790), .ZN(n559) );
  NAND2_X1 U624 ( .A1(G51), .A2(n791), .ZN(n558) );
  NAND2_X1 U625 ( .A1(n559), .A2(n558), .ZN(n560) );
  XOR2_X1 U626 ( .A(KEYINPUT6), .B(n560), .Z(n561) );
  NAND2_X1 U627 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U628 ( .A(n563), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U629 ( .A1(G88), .A2(n786), .ZN(n565) );
  NAND2_X1 U630 ( .A1(G75), .A2(n787), .ZN(n564) );
  NAND2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n568) );
  NAND2_X1 U632 ( .A1(G62), .A2(n790), .ZN(n566) );
  XNOR2_X1 U633 ( .A(KEYINPUT77), .B(n566), .ZN(n567) );
  NOR2_X1 U634 ( .A1(n568), .A2(n567), .ZN(n570) );
  NAND2_X1 U635 ( .A1(n791), .A2(G50), .ZN(n569) );
  NAND2_X1 U636 ( .A1(n570), .A2(n569), .ZN(G303) );
  XOR2_X1 U637 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U638 ( .A1(G49), .A2(n791), .ZN(n572) );
  NAND2_X1 U639 ( .A1(G74), .A2(G651), .ZN(n571) );
  NAND2_X1 U640 ( .A1(n572), .A2(n571), .ZN(n573) );
  NOR2_X1 U641 ( .A1(n790), .A2(n573), .ZN(n576) );
  NAND2_X1 U642 ( .A1(n574), .A2(G87), .ZN(n575) );
  NAND2_X1 U643 ( .A1(n576), .A2(n575), .ZN(G288) );
  NAND2_X1 U644 ( .A1(G61), .A2(n790), .ZN(n578) );
  NAND2_X1 U645 ( .A1(G86), .A2(n786), .ZN(n577) );
  NAND2_X1 U646 ( .A1(n578), .A2(n577), .ZN(n581) );
  NAND2_X1 U647 ( .A1(n787), .A2(G73), .ZN(n579) );
  XOR2_X1 U648 ( .A(KEYINPUT2), .B(n579), .Z(n580) );
  NOR2_X1 U649 ( .A1(n581), .A2(n580), .ZN(n583) );
  NAND2_X1 U650 ( .A1(n791), .A2(G48), .ZN(n582) );
  NAND2_X1 U651 ( .A1(n583), .A2(n582), .ZN(G305) );
  NAND2_X1 U652 ( .A1(G60), .A2(n790), .ZN(n585) );
  NAND2_X1 U653 ( .A1(G47), .A2(n791), .ZN(n584) );
  NAND2_X1 U654 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U655 ( .A(KEYINPUT66), .B(n586), .Z(n590) );
  NAND2_X1 U656 ( .A1(G85), .A2(n786), .ZN(n588) );
  NAND2_X1 U657 ( .A1(G72), .A2(n787), .ZN(n587) );
  AND2_X1 U658 ( .A1(n588), .A2(n587), .ZN(n589) );
  NAND2_X1 U659 ( .A1(n590), .A2(n589), .ZN(G290) );
  NAND2_X1 U660 ( .A1(n786), .A2(G81), .ZN(n591) );
  XNOR2_X1 U661 ( .A(n591), .B(KEYINPUT12), .ZN(n593) );
  NAND2_X1 U662 ( .A1(G68), .A2(n787), .ZN(n592) );
  NAND2_X1 U663 ( .A1(n593), .A2(n592), .ZN(n594) );
  XOR2_X1 U664 ( .A(KEYINPUT13), .B(n594), .Z(n598) );
  NAND2_X1 U665 ( .A1(G56), .A2(n790), .ZN(n596) );
  NOR2_X1 U666 ( .A1(n598), .A2(n597), .ZN(n600) );
  NAND2_X1 U667 ( .A1(n791), .A2(G43), .ZN(n599) );
  NAND2_X1 U668 ( .A1(n600), .A2(n599), .ZN(n965) );
  NOR2_X1 U669 ( .A1(G164), .A2(G1384), .ZN(n703) );
  NAND2_X2 U670 ( .A1(n701), .A2(n703), .ZN(n653) );
  INV_X1 U671 ( .A(G1996), .ZN(n602) );
  XOR2_X1 U672 ( .A(KEYINPUT64), .B(KEYINPUT26), .Z(n603) );
  XNOR2_X1 U673 ( .A(n604), .B(n603), .ZN(n606) );
  NAND2_X1 U674 ( .A1(n653), .A2(G1341), .ZN(n605) );
  NAND2_X1 U675 ( .A1(n606), .A2(n605), .ZN(n607) );
  NAND2_X1 U676 ( .A1(G79), .A2(n787), .ZN(n614) );
  NAND2_X1 U677 ( .A1(G66), .A2(n790), .ZN(n609) );
  NAND2_X1 U678 ( .A1(G54), .A2(n791), .ZN(n608) );
  NAND2_X1 U679 ( .A1(n609), .A2(n608), .ZN(n612) );
  NAND2_X1 U680 ( .A1(n786), .A2(G92), .ZN(n610) );
  XOR2_X1 U681 ( .A(KEYINPUT72), .B(n610), .Z(n611) );
  NOR2_X1 U682 ( .A1(n612), .A2(n611), .ZN(n613) );
  NAND2_X1 U683 ( .A1(n614), .A2(n613), .ZN(n615) );
  XNOR2_X1 U684 ( .A(n615), .B(KEYINPUT15), .ZN(n962) );
  NOR2_X1 U685 ( .A1(n618), .A2(n962), .ZN(n617) );
  XNOR2_X1 U686 ( .A(n617), .B(n616), .ZN(n624) );
  NAND2_X1 U687 ( .A1(n618), .A2(n962), .ZN(n622) );
  NOR2_X1 U688 ( .A1(n638), .A2(G1348), .ZN(n620) );
  NOR2_X1 U689 ( .A1(G2067), .A2(n653), .ZN(n619) );
  NOR2_X1 U690 ( .A1(n620), .A2(n619), .ZN(n621) );
  NAND2_X1 U691 ( .A1(n622), .A2(n621), .ZN(n623) );
  NAND2_X1 U692 ( .A1(n624), .A2(n623), .ZN(n630) );
  INV_X1 U693 ( .A(G299), .ZN(n801) );
  NAND2_X1 U694 ( .A1(G2072), .A2(n638), .ZN(n625) );
  XNOR2_X1 U695 ( .A(n625), .B(KEYINPUT92), .ZN(n626) );
  XNOR2_X1 U696 ( .A(KEYINPUT27), .B(n626), .ZN(n628) );
  INV_X1 U697 ( .A(G1956), .ZN(n894) );
  NOR2_X1 U698 ( .A1(n638), .A2(n894), .ZN(n627) );
  NOR2_X1 U699 ( .A1(n628), .A2(n627), .ZN(n631) );
  NAND2_X1 U700 ( .A1(n801), .A2(n631), .ZN(n629) );
  NAND2_X1 U701 ( .A1(n630), .A2(n629), .ZN(n635) );
  XNOR2_X1 U702 ( .A(KEYINPUT93), .B(KEYINPUT28), .ZN(n632) );
  XNOR2_X1 U703 ( .A(n633), .B(n632), .ZN(n634) );
  NAND2_X1 U704 ( .A1(n635), .A2(n634), .ZN(n636) );
  XNOR2_X1 U705 ( .A(n636), .B(KEYINPUT29), .ZN(n642) );
  NAND2_X1 U706 ( .A1(G1961), .A2(n653), .ZN(n640) );
  XNOR2_X1 U707 ( .A(G2078), .B(KEYINPUT25), .ZN(n637) );
  XNOR2_X1 U708 ( .A(n637), .B(KEYINPUT91), .ZN(n875) );
  NAND2_X1 U709 ( .A1(n638), .A2(n875), .ZN(n639) );
  NAND2_X1 U710 ( .A1(n640), .A2(n639), .ZN(n644) );
  NOR2_X1 U711 ( .A1(G301), .A2(n644), .ZN(n641) );
  NOR2_X1 U712 ( .A1(n642), .A2(n641), .ZN(n643) );
  XNOR2_X1 U713 ( .A(n643), .B(KEYINPUT95), .ZN(n665) );
  NAND2_X1 U714 ( .A1(G301), .A2(n644), .ZN(n645) );
  XNOR2_X1 U715 ( .A(n645), .B(KEYINPUT97), .ZN(n651) );
  NOR2_X1 U716 ( .A1(G1966), .A2(n695), .ZN(n667) );
  NOR2_X1 U717 ( .A1(G2084), .A2(n653), .ZN(n666) );
  NOR2_X1 U718 ( .A1(n667), .A2(n666), .ZN(n646) );
  XNOR2_X1 U719 ( .A(n646), .B(KEYINPUT96), .ZN(n647) );
  NAND2_X1 U720 ( .A1(n647), .A2(G8), .ZN(n648) );
  XNOR2_X1 U721 ( .A(KEYINPUT30), .B(n648), .ZN(n649) );
  NOR2_X1 U722 ( .A1(n649), .A2(G168), .ZN(n650) );
  XOR2_X1 U723 ( .A(KEYINPUT31), .B(n652), .Z(n664) );
  NOR2_X1 U724 ( .A1(G1971), .A2(n695), .ZN(n655) );
  NOR2_X1 U725 ( .A1(G2090), .A2(n653), .ZN(n654) );
  NOR2_X1 U726 ( .A1(n655), .A2(n654), .ZN(n656) );
  NAND2_X1 U727 ( .A1(n656), .A2(G303), .ZN(n658) );
  AND2_X1 U728 ( .A1(n664), .A2(n658), .ZN(n657) );
  NAND2_X1 U729 ( .A1(n665), .A2(n657), .ZN(n662) );
  INV_X1 U730 ( .A(n658), .ZN(n659) );
  OR2_X1 U731 ( .A1(n659), .A2(G286), .ZN(n660) );
  AND2_X1 U732 ( .A1(G8), .A2(n660), .ZN(n661) );
  NAND2_X1 U733 ( .A1(n662), .A2(n661), .ZN(n663) );
  XNOR2_X1 U734 ( .A(n663), .B(KEYINPUT32), .ZN(n687) );
  AND2_X1 U735 ( .A1(n665), .A2(n664), .ZN(n670) );
  AND2_X1 U736 ( .A1(G8), .A2(n666), .ZN(n668) );
  OR2_X1 U737 ( .A1(n668), .A2(n667), .ZN(n669) );
  NAND2_X1 U738 ( .A1(G1976), .A2(G288), .ZN(n848) );
  NAND2_X1 U739 ( .A1(n687), .A2(n671), .ZN(n677) );
  INV_X1 U740 ( .A(n848), .ZN(n675) );
  NOR2_X1 U741 ( .A1(G1971), .A2(G303), .ZN(n673) );
  NOR2_X1 U742 ( .A1(G1976), .A2(G288), .ZN(n672) );
  XOR2_X1 U743 ( .A(KEYINPUT98), .B(n672), .Z(n682) );
  INV_X1 U744 ( .A(n682), .ZN(n851) );
  NOR2_X1 U745 ( .A1(n673), .A2(n851), .ZN(n674) );
  OR2_X1 U746 ( .A1(n675), .A2(n674), .ZN(n676) );
  AND2_X1 U747 ( .A1(n677), .A2(n676), .ZN(n678) );
  XNOR2_X1 U748 ( .A(n678), .B(KEYINPUT99), .ZN(n680) );
  AND2_X1 U749 ( .A1(n680), .A2(n679), .ZN(n681) );
  NOR2_X1 U750 ( .A1(KEYINPUT33), .A2(n681), .ZN(n686) );
  XOR2_X1 U751 ( .A(G1981), .B(G305), .Z(n859) );
  NOR2_X1 U752 ( .A1(n695), .A2(n682), .ZN(n683) );
  NAND2_X1 U753 ( .A1(KEYINPUT33), .A2(n683), .ZN(n684) );
  NAND2_X1 U754 ( .A1(n859), .A2(n684), .ZN(n685) );
  OR2_X1 U755 ( .A1(n686), .A2(n685), .ZN(n699) );
  NAND2_X1 U756 ( .A1(n687), .A2(n688), .ZN(n691) );
  NOR2_X1 U757 ( .A1(G2090), .A2(G303), .ZN(n689) );
  NAND2_X1 U758 ( .A1(G8), .A2(n689), .ZN(n690) );
  NAND2_X1 U759 ( .A1(n691), .A2(n690), .ZN(n692) );
  AND2_X1 U760 ( .A1(n695), .A2(n692), .ZN(n698) );
  NOR2_X1 U761 ( .A1(G1981), .A2(G305), .ZN(n693) );
  XOR2_X1 U762 ( .A(n693), .B(KEYINPUT90), .Z(n694) );
  XNOR2_X1 U763 ( .A(KEYINPUT24), .B(n694), .ZN(n696) );
  NOR2_X1 U764 ( .A1(n696), .A2(n695), .ZN(n697) );
  NAND2_X1 U765 ( .A1(n699), .A2(n519), .ZN(n700) );
  XNOR2_X1 U766 ( .A(n700), .B(KEYINPUT100), .ZN(n705) );
  INV_X1 U767 ( .A(n701), .ZN(n702) );
  NOR2_X1 U768 ( .A1(n703), .A2(n702), .ZN(n754) );
  XNOR2_X1 U769 ( .A(G1986), .B(G290), .ZN(n855) );
  NAND2_X1 U770 ( .A1(n754), .A2(n855), .ZN(n704) );
  NAND2_X1 U771 ( .A1(n705), .A2(n704), .ZN(n742) );
  XNOR2_X1 U772 ( .A(KEYINPUT84), .B(KEYINPUT36), .ZN(n718) );
  NAND2_X1 U773 ( .A1(n991), .A2(G128), .ZN(n706) );
  XOR2_X1 U774 ( .A(KEYINPUT83), .B(n706), .Z(n708) );
  NAND2_X1 U775 ( .A1(n992), .A2(G116), .ZN(n707) );
  NAND2_X1 U776 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U777 ( .A(KEYINPUT35), .B(n709), .ZN(n716) );
  NAND2_X1 U778 ( .A1(G104), .A2(n996), .ZN(n712) );
  NAND2_X1 U779 ( .A1(n995), .A2(G140), .ZN(n710) );
  XOR2_X1 U780 ( .A(KEYINPUT81), .B(n710), .Z(n711) );
  NAND2_X1 U781 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U782 ( .A(n713), .B(KEYINPUT82), .ZN(n714) );
  XOR2_X1 U783 ( .A(KEYINPUT34), .B(n714), .Z(n715) );
  NAND2_X1 U784 ( .A1(n716), .A2(n715), .ZN(n717) );
  XOR2_X1 U785 ( .A(n718), .B(n717), .Z(n1010) );
  XNOR2_X1 U786 ( .A(G2067), .B(KEYINPUT37), .ZN(n752) );
  OR2_X1 U787 ( .A1(n1010), .A2(n752), .ZN(n719) );
  XNOR2_X1 U788 ( .A(n719), .B(KEYINPUT85), .ZN(n927) );
  NAND2_X1 U789 ( .A1(n927), .A2(n754), .ZN(n751) );
  NAND2_X1 U790 ( .A1(G119), .A2(n991), .ZN(n720) );
  XNOR2_X1 U791 ( .A(n720), .B(KEYINPUT86), .ZN(n728) );
  NAND2_X1 U792 ( .A1(G131), .A2(n995), .ZN(n722) );
  NAND2_X1 U793 ( .A1(G95), .A2(n996), .ZN(n721) );
  NAND2_X1 U794 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U795 ( .A(KEYINPUT88), .B(n723), .ZN(n726) );
  NAND2_X1 U796 ( .A1(G107), .A2(n992), .ZN(n724) );
  XNOR2_X1 U797 ( .A(KEYINPUT87), .B(n724), .ZN(n725) );
  NOR2_X1 U798 ( .A1(n726), .A2(n725), .ZN(n727) );
  NAND2_X1 U799 ( .A1(n728), .A2(n727), .ZN(n1002) );
  AND2_X1 U800 ( .A1(n1002), .A2(G1991), .ZN(n738) );
  NAND2_X1 U801 ( .A1(G129), .A2(n991), .ZN(n730) );
  NAND2_X1 U802 ( .A1(G141), .A2(n995), .ZN(n729) );
  NAND2_X1 U803 ( .A1(n730), .A2(n729), .ZN(n734) );
  NAND2_X1 U804 ( .A1(G105), .A2(n996), .ZN(n731) );
  XNOR2_X1 U805 ( .A(n731), .B(KEYINPUT89), .ZN(n732) );
  XNOR2_X1 U806 ( .A(n732), .B(KEYINPUT38), .ZN(n733) );
  NOR2_X1 U807 ( .A1(n734), .A2(n733), .ZN(n736) );
  NAND2_X1 U808 ( .A1(n992), .A2(G117), .ZN(n735) );
  NAND2_X1 U809 ( .A1(n736), .A2(n735), .ZN(n1009) );
  AND2_X1 U810 ( .A1(n1009), .A2(G1996), .ZN(n737) );
  NOR2_X1 U811 ( .A1(n738), .A2(n737), .ZN(n925) );
  INV_X1 U812 ( .A(n754), .ZN(n739) );
  NOR2_X1 U813 ( .A1(n925), .A2(n739), .ZN(n746) );
  INV_X1 U814 ( .A(n746), .ZN(n740) );
  NAND2_X1 U815 ( .A1(n751), .A2(n740), .ZN(n741) );
  NOR2_X1 U816 ( .A1(n742), .A2(n741), .ZN(n758) );
  NOR2_X1 U817 ( .A1(G1996), .A2(n1009), .ZN(n919) );
  NOR2_X1 U818 ( .A1(G1986), .A2(G290), .ZN(n744) );
  NOR2_X1 U819 ( .A1(G1991), .A2(n1002), .ZN(n743) );
  XOR2_X1 U820 ( .A(KEYINPUT101), .B(n743), .Z(n923) );
  NOR2_X1 U821 ( .A1(n744), .A2(n923), .ZN(n745) );
  NOR2_X1 U822 ( .A1(n746), .A2(n745), .ZN(n747) );
  NOR2_X1 U823 ( .A1(n919), .A2(n747), .ZN(n748) );
  XNOR2_X1 U824 ( .A(n748), .B(KEYINPUT102), .ZN(n749) );
  XNOR2_X1 U825 ( .A(n749), .B(KEYINPUT39), .ZN(n750) );
  NAND2_X1 U826 ( .A1(n751), .A2(n750), .ZN(n753) );
  NAND2_X1 U827 ( .A1(n1010), .A2(n752), .ZN(n946) );
  NAND2_X1 U828 ( .A1(n753), .A2(n946), .ZN(n755) );
  NAND2_X1 U829 ( .A1(n755), .A2(n754), .ZN(n756) );
  XNOR2_X1 U830 ( .A(n756), .B(KEYINPUT103), .ZN(n757) );
  XNOR2_X1 U831 ( .A(n759), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U832 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U833 ( .A1(G123), .A2(n991), .ZN(n760) );
  XNOR2_X1 U834 ( .A(n760), .B(KEYINPUT18), .ZN(n767) );
  NAND2_X1 U835 ( .A1(G135), .A2(n995), .ZN(n762) );
  NAND2_X1 U836 ( .A1(G99), .A2(n996), .ZN(n761) );
  NAND2_X1 U837 ( .A1(n762), .A2(n761), .ZN(n765) );
  NAND2_X1 U838 ( .A1(G111), .A2(n992), .ZN(n763) );
  XNOR2_X1 U839 ( .A(KEYINPUT75), .B(n763), .ZN(n764) );
  NOR2_X1 U840 ( .A1(n765), .A2(n764), .ZN(n766) );
  NAND2_X1 U841 ( .A1(n767), .A2(n766), .ZN(n768) );
  XNOR2_X1 U842 ( .A(KEYINPUT76), .B(n768), .ZN(n1008) );
  XNOR2_X1 U843 ( .A(n1008), .B(G2096), .ZN(n769) );
  OR2_X1 U844 ( .A1(G2100), .A2(n769), .ZN(G156) );
  INV_X1 U845 ( .A(G132), .ZN(G219) );
  INV_X1 U846 ( .A(G82), .ZN(G220) );
  INV_X1 U847 ( .A(G57), .ZN(G237) );
  NAND2_X1 U848 ( .A1(G7), .A2(G661), .ZN(n770) );
  XNOR2_X1 U849 ( .A(n770), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U850 ( .A(KEYINPUT70), .B(KEYINPUT11), .Z(n772) );
  INV_X1 U851 ( .A(G223), .ZN(n833) );
  NAND2_X1 U852 ( .A1(G567), .A2(n833), .ZN(n771) );
  XNOR2_X1 U853 ( .A(n772), .B(n771), .ZN(G234) );
  INV_X1 U854 ( .A(G860), .ZN(n779) );
  OR2_X1 U855 ( .A1(n965), .A2(n779), .ZN(G153) );
  NOR2_X1 U856 ( .A1(n962), .A2(G868), .ZN(n773) );
  XNOR2_X1 U857 ( .A(n773), .B(KEYINPUT73), .ZN(n775) );
  NAND2_X1 U858 ( .A1(G868), .A2(G301), .ZN(n774) );
  NAND2_X1 U859 ( .A1(n775), .A2(n774), .ZN(G284) );
  INV_X1 U860 ( .A(G868), .ZN(n776) );
  NOR2_X1 U861 ( .A1(G286), .A2(n776), .ZN(n778) );
  NOR2_X1 U862 ( .A1(G868), .A2(G299), .ZN(n777) );
  NOR2_X1 U863 ( .A1(n778), .A2(n777), .ZN(G297) );
  NAND2_X1 U864 ( .A1(n779), .A2(G559), .ZN(n780) );
  NAND2_X1 U865 ( .A1(n780), .A2(n962), .ZN(n781) );
  XNOR2_X1 U866 ( .A(n781), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U867 ( .A1(G868), .A2(n965), .ZN(n784) );
  NAND2_X1 U868 ( .A1(G868), .A2(n962), .ZN(n782) );
  NOR2_X1 U869 ( .A1(G559), .A2(n782), .ZN(n783) );
  NOR2_X1 U870 ( .A1(n784), .A2(n783), .ZN(G282) );
  NAND2_X1 U871 ( .A1(G559), .A2(n962), .ZN(n785) );
  XNOR2_X1 U872 ( .A(n785), .B(n965), .ZN(n804) );
  NOR2_X1 U873 ( .A1(n804), .A2(G860), .ZN(n796) );
  NAND2_X1 U874 ( .A1(G93), .A2(n786), .ZN(n789) );
  NAND2_X1 U875 ( .A1(G80), .A2(n787), .ZN(n788) );
  NAND2_X1 U876 ( .A1(n789), .A2(n788), .ZN(n795) );
  NAND2_X1 U877 ( .A1(G67), .A2(n790), .ZN(n793) );
  NAND2_X1 U878 ( .A1(G55), .A2(n791), .ZN(n792) );
  NAND2_X1 U879 ( .A1(n793), .A2(n792), .ZN(n794) );
  NOR2_X1 U880 ( .A1(n795), .A2(n794), .ZN(n807) );
  XNOR2_X1 U881 ( .A(n796), .B(n807), .ZN(G145) );
  INV_X1 U882 ( .A(G303), .ZN(G166) );
  XNOR2_X1 U883 ( .A(G166), .B(G305), .ZN(n797) );
  XNOR2_X1 U884 ( .A(n797), .B(G290), .ZN(n800) );
  XOR2_X1 U885 ( .A(KEYINPUT78), .B(KEYINPUT19), .Z(n798) );
  XNOR2_X1 U886 ( .A(G288), .B(n798), .ZN(n799) );
  XOR2_X1 U887 ( .A(n800), .B(n799), .Z(n803) );
  XNOR2_X1 U888 ( .A(n801), .B(n807), .ZN(n802) );
  XNOR2_X1 U889 ( .A(n803), .B(n802), .ZN(n961) );
  XNOR2_X1 U890 ( .A(n961), .B(n804), .ZN(n805) );
  NAND2_X1 U891 ( .A1(n805), .A2(G868), .ZN(n806) );
  XOR2_X1 U892 ( .A(KEYINPUT79), .B(n806), .Z(n809) );
  OR2_X1 U893 ( .A1(n807), .A2(G868), .ZN(n808) );
  NAND2_X1 U894 ( .A1(n809), .A2(n808), .ZN(G295) );
  NAND2_X1 U895 ( .A1(G2078), .A2(G2084), .ZN(n810) );
  XOR2_X1 U896 ( .A(KEYINPUT20), .B(n810), .Z(n811) );
  NAND2_X1 U897 ( .A1(G2090), .A2(n811), .ZN(n812) );
  XNOR2_X1 U898 ( .A(KEYINPUT21), .B(n812), .ZN(n813) );
  NAND2_X1 U899 ( .A1(n813), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U900 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U901 ( .A1(G69), .A2(G120), .ZN(n814) );
  NOR2_X1 U902 ( .A1(G237), .A2(n814), .ZN(n815) );
  NAND2_X1 U903 ( .A1(G108), .A2(n815), .ZN(n959) );
  NAND2_X1 U904 ( .A1(n959), .A2(G567), .ZN(n821) );
  NOR2_X1 U905 ( .A1(G220), .A2(G219), .ZN(n816) );
  XNOR2_X1 U906 ( .A(KEYINPUT22), .B(n816), .ZN(n817) );
  NAND2_X1 U907 ( .A1(n817), .A2(G96), .ZN(n818) );
  NOR2_X1 U908 ( .A1(G218), .A2(n818), .ZN(n819) );
  XOR2_X1 U909 ( .A(KEYINPUT80), .B(n819), .Z(n960) );
  NAND2_X1 U910 ( .A1(G2106), .A2(n960), .ZN(n820) );
  NAND2_X1 U911 ( .A1(n821), .A2(n820), .ZN(n968) );
  NAND2_X1 U912 ( .A1(G661), .A2(G483), .ZN(n822) );
  NOR2_X1 U913 ( .A1(n968), .A2(n822), .ZN(n836) );
  NAND2_X1 U914 ( .A1(n836), .A2(G36), .ZN(G176) );
  XNOR2_X1 U915 ( .A(G2443), .B(G1341), .ZN(n831) );
  XNOR2_X1 U916 ( .A(G2430), .B(G2446), .ZN(n829) );
  XOR2_X1 U917 ( .A(G2454), .B(G2451), .Z(n824) );
  XNOR2_X1 U918 ( .A(G2427), .B(G2435), .ZN(n823) );
  XNOR2_X1 U919 ( .A(n824), .B(n823), .ZN(n825) );
  XOR2_X1 U920 ( .A(n825), .B(G2438), .Z(n827) );
  XNOR2_X1 U921 ( .A(G1348), .B(KEYINPUT104), .ZN(n826) );
  XNOR2_X1 U922 ( .A(n827), .B(n826), .ZN(n828) );
  XNOR2_X1 U923 ( .A(n829), .B(n828), .ZN(n830) );
  XNOR2_X1 U924 ( .A(n831), .B(n830), .ZN(n832) );
  NAND2_X1 U925 ( .A1(n832), .A2(G14), .ZN(n1018) );
  XNOR2_X1 U926 ( .A(KEYINPUT105), .B(n1018), .ZN(G401) );
  NAND2_X1 U927 ( .A1(G2106), .A2(n833), .ZN(G217) );
  AND2_X1 U928 ( .A1(G15), .A2(G2), .ZN(n834) );
  NAND2_X1 U929 ( .A1(G661), .A2(n834), .ZN(G259) );
  NAND2_X1 U930 ( .A1(G3), .A2(G1), .ZN(n835) );
  XNOR2_X1 U931 ( .A(KEYINPUT106), .B(n835), .ZN(n837) );
  NAND2_X1 U932 ( .A1(n837), .A2(n836), .ZN(G188) );
  NAND2_X1 U934 ( .A1(G124), .A2(n991), .ZN(n838) );
  XNOR2_X1 U935 ( .A(n838), .B(KEYINPUT44), .ZN(n839) );
  XNOR2_X1 U936 ( .A(n839), .B(KEYINPUT112), .ZN(n841) );
  NAND2_X1 U937 ( .A1(G100), .A2(n996), .ZN(n840) );
  NAND2_X1 U938 ( .A1(n841), .A2(n840), .ZN(n845) );
  NAND2_X1 U939 ( .A1(G112), .A2(n992), .ZN(n843) );
  NAND2_X1 U940 ( .A1(G136), .A2(n995), .ZN(n842) );
  NAND2_X1 U941 ( .A1(n843), .A2(n842), .ZN(n844) );
  NOR2_X1 U942 ( .A1(n845), .A2(n844), .ZN(G162) );
  XNOR2_X1 U943 ( .A(KEYINPUT56), .B(G16), .ZN(n868) );
  XNOR2_X1 U944 ( .A(n965), .B(G1341), .ZN(n847) );
  XNOR2_X1 U945 ( .A(G299), .B(G1956), .ZN(n846) );
  NOR2_X1 U946 ( .A1(n847), .A2(n846), .ZN(n849) );
  NAND2_X1 U947 ( .A1(n849), .A2(n848), .ZN(n850) );
  NOR2_X1 U948 ( .A1(n851), .A2(n850), .ZN(n857) );
  XNOR2_X1 U949 ( .A(G1348), .B(n962), .ZN(n853) );
  XNOR2_X1 U950 ( .A(G171), .B(G1961), .ZN(n852) );
  NAND2_X1 U951 ( .A1(n853), .A2(n852), .ZN(n854) );
  NOR2_X1 U952 ( .A1(n855), .A2(n854), .ZN(n856) );
  NAND2_X1 U953 ( .A1(n857), .A2(n856), .ZN(n865) );
  XNOR2_X1 U954 ( .A(G1971), .B(G166), .ZN(n858) );
  XNOR2_X1 U955 ( .A(n858), .B(KEYINPUT122), .ZN(n863) );
  XNOR2_X1 U956 ( .A(G1966), .B(G168), .ZN(n860) );
  NAND2_X1 U957 ( .A1(n860), .A2(n859), .ZN(n861) );
  XNOR2_X1 U958 ( .A(n861), .B(KEYINPUT57), .ZN(n862) );
  NAND2_X1 U959 ( .A1(n863), .A2(n862), .ZN(n864) );
  NOR2_X1 U960 ( .A1(n865), .A2(n864), .ZN(n866) );
  XNOR2_X1 U961 ( .A(KEYINPUT123), .B(n866), .ZN(n867) );
  NAND2_X1 U962 ( .A1(n868), .A2(n867), .ZN(n957) );
  XOR2_X1 U963 ( .A(G1991), .B(G25), .Z(n869) );
  NAND2_X1 U964 ( .A1(n869), .A2(G28), .ZN(n870) );
  XNOR2_X1 U965 ( .A(n870), .B(KEYINPUT119), .ZN(n874) );
  XNOR2_X1 U966 ( .A(G2067), .B(G26), .ZN(n872) );
  XNOR2_X1 U967 ( .A(G2072), .B(G33), .ZN(n871) );
  NOR2_X1 U968 ( .A1(n872), .A2(n871), .ZN(n873) );
  NAND2_X1 U969 ( .A1(n874), .A2(n873), .ZN(n880) );
  XOR2_X1 U970 ( .A(n875), .B(G27), .Z(n878) );
  XOR2_X1 U971 ( .A(G32), .B(KEYINPUT120), .Z(n876) );
  XNOR2_X1 U972 ( .A(G1996), .B(n876), .ZN(n877) );
  NAND2_X1 U973 ( .A1(n878), .A2(n877), .ZN(n879) );
  NOR2_X1 U974 ( .A1(n880), .A2(n879), .ZN(n881) );
  XOR2_X1 U975 ( .A(KEYINPUT53), .B(n881), .Z(n885) );
  XNOR2_X1 U976 ( .A(KEYINPUT54), .B(KEYINPUT121), .ZN(n882) );
  XNOR2_X1 U977 ( .A(n882), .B(G34), .ZN(n883) );
  XNOR2_X1 U978 ( .A(G2084), .B(n883), .ZN(n884) );
  NAND2_X1 U979 ( .A1(n885), .A2(n884), .ZN(n887) );
  XNOR2_X1 U980 ( .A(G35), .B(G2090), .ZN(n886) );
  OR2_X1 U981 ( .A1(n887), .A2(n886), .ZN(n914) );
  XOR2_X1 U982 ( .A(KEYINPUT55), .B(KEYINPUT118), .Z(n949) );
  OR2_X1 U983 ( .A1(n914), .A2(n949), .ZN(n888) );
  NAND2_X1 U984 ( .A1(G11), .A2(n888), .ZN(n955) );
  XNOR2_X1 U985 ( .A(G1966), .B(G21), .ZN(n890) );
  XNOR2_X1 U986 ( .A(G5), .B(G1961), .ZN(n889) );
  NOR2_X1 U987 ( .A1(n890), .A2(n889), .ZN(n910) );
  XNOR2_X1 U988 ( .A(G1341), .B(G19), .ZN(n892) );
  XNOR2_X1 U989 ( .A(G1981), .B(G6), .ZN(n891) );
  NOR2_X1 U990 ( .A1(n892), .A2(n891), .ZN(n893) );
  XNOR2_X1 U991 ( .A(KEYINPUT124), .B(n893), .ZN(n896) );
  XNOR2_X1 U992 ( .A(n894), .B(G20), .ZN(n895) );
  NAND2_X1 U993 ( .A1(n896), .A2(n895), .ZN(n899) );
  XOR2_X1 U994 ( .A(KEYINPUT59), .B(G1348), .Z(n897) );
  XNOR2_X1 U995 ( .A(G4), .B(n897), .ZN(n898) );
  NOR2_X1 U996 ( .A1(n899), .A2(n898), .ZN(n900) );
  XNOR2_X1 U997 ( .A(n900), .B(KEYINPUT125), .ZN(n901) );
  XNOR2_X1 U998 ( .A(n901), .B(KEYINPUT60), .ZN(n908) );
  XNOR2_X1 U999 ( .A(G1971), .B(G22), .ZN(n903) );
  XNOR2_X1 U1000 ( .A(G23), .B(G1976), .ZN(n902) );
  NOR2_X1 U1001 ( .A1(n903), .A2(n902), .ZN(n905) );
  XOR2_X1 U1002 ( .A(G1986), .B(G24), .Z(n904) );
  NAND2_X1 U1003 ( .A1(n905), .A2(n904), .ZN(n906) );
  XNOR2_X1 U1004 ( .A(KEYINPUT58), .B(n906), .ZN(n907) );
  NOR2_X1 U1005 ( .A1(n908), .A2(n907), .ZN(n909) );
  NAND2_X1 U1006 ( .A1(n910), .A2(n909), .ZN(n911) );
  XNOR2_X1 U1007 ( .A(n911), .B(KEYINPUT126), .ZN(n912) );
  XNOR2_X1 U1008 ( .A(n912), .B(KEYINPUT61), .ZN(n913) );
  NOR2_X1 U1009 ( .A1(G16), .A2(n913), .ZN(n917) );
  NAND2_X1 U1010 ( .A1(n949), .A2(n914), .ZN(n915) );
  NOR2_X1 U1011 ( .A1(G29), .A2(n915), .ZN(n916) );
  NOR2_X1 U1012 ( .A1(n917), .A2(n916), .ZN(n953) );
  XOR2_X1 U1013 ( .A(G2090), .B(G162), .Z(n918) );
  NOR2_X1 U1014 ( .A1(n919), .A2(n918), .ZN(n920) );
  XOR2_X1 U1015 ( .A(KEYINPUT51), .B(n920), .Z(n930) );
  XNOR2_X1 U1016 ( .A(G160), .B(G2084), .ZN(n921) );
  NAND2_X1 U1017 ( .A1(n921), .A2(n1008), .ZN(n922) );
  NOR2_X1 U1018 ( .A1(n923), .A2(n922), .ZN(n924) );
  NAND2_X1 U1019 ( .A1(n925), .A2(n924), .ZN(n926) );
  NOR2_X1 U1020 ( .A1(n927), .A2(n926), .ZN(n928) );
  XNOR2_X1 U1021 ( .A(n928), .B(KEYINPUT116), .ZN(n929) );
  NAND2_X1 U1022 ( .A1(n930), .A2(n929), .ZN(n944) );
  XOR2_X1 U1023 ( .A(G164), .B(G2078), .Z(n941) );
  NAND2_X1 U1024 ( .A1(G127), .A2(n991), .ZN(n932) );
  NAND2_X1 U1025 ( .A1(G115), .A2(n992), .ZN(n931) );
  NAND2_X1 U1026 ( .A1(n932), .A2(n931), .ZN(n933) );
  XNOR2_X1 U1027 ( .A(n933), .B(KEYINPUT47), .ZN(n935) );
  NAND2_X1 U1028 ( .A1(G139), .A2(n995), .ZN(n934) );
  NAND2_X1 U1029 ( .A1(n935), .A2(n934), .ZN(n938) );
  NAND2_X1 U1030 ( .A1(G103), .A2(n996), .ZN(n936) );
  XNOR2_X1 U1031 ( .A(KEYINPUT113), .B(n936), .ZN(n937) );
  NOR2_X1 U1032 ( .A1(n938), .A2(n937), .ZN(n939) );
  XOR2_X1 U1033 ( .A(KEYINPUT114), .B(n939), .Z(n1004) );
  XNOR2_X1 U1034 ( .A(G2072), .B(n1004), .ZN(n940) );
  NOR2_X1 U1035 ( .A1(n941), .A2(n940), .ZN(n942) );
  XOR2_X1 U1036 ( .A(KEYINPUT50), .B(n942), .Z(n943) );
  NOR2_X1 U1037 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1038 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1039 ( .A(n947), .B(KEYINPUT117), .ZN(n948) );
  XNOR2_X1 U1040 ( .A(KEYINPUT52), .B(n948), .ZN(n950) );
  NAND2_X1 U1041 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1042 ( .A1(n951), .A2(G29), .ZN(n952) );
  NAND2_X1 U1043 ( .A1(n953), .A2(n952), .ZN(n954) );
  NOR2_X1 U1044 ( .A1(n955), .A2(n954), .ZN(n956) );
  NAND2_X1 U1045 ( .A1(n957), .A2(n956), .ZN(n958) );
  XOR2_X1 U1046 ( .A(KEYINPUT62), .B(n958), .Z(G311) );
  XNOR2_X1 U1047 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1048 ( .A(G120), .ZN(G236) );
  INV_X1 U1049 ( .A(G96), .ZN(G221) );
  INV_X1 U1050 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1051 ( .A1(n960), .A2(n959), .ZN(G325) );
  INV_X1 U1052 ( .A(G325), .ZN(G261) );
  XOR2_X1 U1053 ( .A(n961), .B(G286), .Z(n964) );
  XNOR2_X1 U1054 ( .A(G171), .B(n962), .ZN(n963) );
  XNOR2_X1 U1055 ( .A(n964), .B(n963), .ZN(n966) );
  XNOR2_X1 U1056 ( .A(n966), .B(n965), .ZN(n967) );
  NOR2_X1 U1057 ( .A1(G37), .A2(n967), .ZN(G397) );
  INV_X1 U1058 ( .A(n968), .ZN(G319) );
  XNOR2_X1 U1059 ( .A(G2072), .B(G2084), .ZN(n969) );
  XNOR2_X1 U1060 ( .A(n969), .B(G2100), .ZN(n979) );
  XOR2_X1 U1061 ( .A(KEYINPUT108), .B(KEYINPUT107), .Z(n971) );
  XNOR2_X1 U1062 ( .A(G2678), .B(KEYINPUT109), .ZN(n970) );
  XNOR2_X1 U1063 ( .A(n971), .B(n970), .ZN(n975) );
  XOR2_X1 U1064 ( .A(KEYINPUT43), .B(G2096), .Z(n973) );
  XNOR2_X1 U1065 ( .A(G2090), .B(KEYINPUT42), .ZN(n972) );
  XNOR2_X1 U1066 ( .A(n973), .B(n972), .ZN(n974) );
  XOR2_X1 U1067 ( .A(n975), .B(n974), .Z(n977) );
  XNOR2_X1 U1068 ( .A(G2067), .B(G2078), .ZN(n976) );
  XNOR2_X1 U1069 ( .A(n977), .B(n976), .ZN(n978) );
  XNOR2_X1 U1070 ( .A(n979), .B(n978), .ZN(G227) );
  XOR2_X1 U1071 ( .A(KEYINPUT111), .B(G1976), .Z(n981) );
  XNOR2_X1 U1072 ( .A(G1991), .B(G1981), .ZN(n980) );
  XNOR2_X1 U1073 ( .A(n981), .B(n980), .ZN(n982) );
  XOR2_X1 U1074 ( .A(n982), .B(KEYINPUT110), .Z(n984) );
  XNOR2_X1 U1075 ( .A(G1966), .B(G1961), .ZN(n983) );
  XNOR2_X1 U1076 ( .A(n984), .B(n983), .ZN(n988) );
  XOR2_X1 U1077 ( .A(G2474), .B(G1986), .Z(n986) );
  XNOR2_X1 U1078 ( .A(G1956), .B(G1971), .ZN(n985) );
  XNOR2_X1 U1079 ( .A(n986), .B(n985), .ZN(n987) );
  XOR2_X1 U1080 ( .A(n988), .B(n987), .Z(n990) );
  XNOR2_X1 U1081 ( .A(G1996), .B(KEYINPUT41), .ZN(n989) );
  XNOR2_X1 U1082 ( .A(n990), .B(n989), .ZN(G229) );
  NAND2_X1 U1083 ( .A1(G130), .A2(n991), .ZN(n994) );
  NAND2_X1 U1084 ( .A1(G118), .A2(n992), .ZN(n993) );
  NAND2_X1 U1085 ( .A1(n994), .A2(n993), .ZN(n1001) );
  NAND2_X1 U1086 ( .A1(G142), .A2(n995), .ZN(n998) );
  NAND2_X1 U1087 ( .A1(G106), .A2(n996), .ZN(n997) );
  NAND2_X1 U1088 ( .A1(n998), .A2(n997), .ZN(n999) );
  XOR2_X1 U1089 ( .A(n999), .B(KEYINPUT45), .Z(n1000) );
  NOR2_X1 U1090 ( .A1(n1001), .A2(n1000), .ZN(n1003) );
  XNOR2_X1 U1091 ( .A(n1003), .B(n1002), .ZN(n1016) );
  XOR2_X1 U1092 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n1006) );
  XNOR2_X1 U1093 ( .A(G160), .B(n1004), .ZN(n1005) );
  XNOR2_X1 U1094 ( .A(n1006), .B(n1005), .ZN(n1007) );
  XNOR2_X1 U1095 ( .A(G164), .B(n1007), .ZN(n1014) );
  XOR2_X1 U1096 ( .A(n1008), .B(G162), .Z(n1012) );
  XOR2_X1 U1097 ( .A(n1010), .B(n1009), .Z(n1011) );
  XNOR2_X1 U1098 ( .A(n1012), .B(n1011), .ZN(n1013) );
  XNOR2_X1 U1099 ( .A(n1014), .B(n1013), .ZN(n1015) );
  XOR2_X1 U1100 ( .A(n1016), .B(n1015), .Z(n1017) );
  NOR2_X1 U1101 ( .A1(G37), .A2(n1017), .ZN(G395) );
  NAND2_X1 U1102 ( .A1(G319), .A2(n1018), .ZN(n1019) );
  NOR2_X1 U1103 ( .A1(G397), .A2(n1019), .ZN(n1022) );
  NOR2_X1 U1104 ( .A1(G227), .A2(G229), .ZN(n1020) );
  XOR2_X1 U1105 ( .A(KEYINPUT49), .B(n1020), .Z(n1021) );
  NAND2_X1 U1106 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NOR2_X1 U1107 ( .A1(n1023), .A2(G395), .ZN(n1024) );
  XNOR2_X1 U1108 ( .A(n1024), .B(KEYINPUT115), .ZN(G225) );
  INV_X1 U1109 ( .A(G225), .ZN(G308) );
  INV_X1 U1110 ( .A(G108), .ZN(G238) );
endmodule

