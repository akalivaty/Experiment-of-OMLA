

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584;

  XNOR2_X1 U323 ( .A(n342), .B(n341), .ZN(n557) );
  XNOR2_X1 U324 ( .A(n391), .B(n390), .ZN(n520) );
  XOR2_X1 U325 ( .A(n387), .B(n358), .Z(n291) );
  XNOR2_X1 U326 ( .A(KEYINPUT114), .B(KEYINPUT46), .ZN(n324) );
  XNOR2_X1 U327 ( .A(n325), .B(n324), .ZN(n364) );
  XNOR2_X1 U328 ( .A(n372), .B(KEYINPUT48), .ZN(n373) );
  XNOR2_X1 U329 ( .A(n383), .B(n382), .ZN(n384) );
  XNOR2_X1 U330 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U331 ( .A(n374), .B(n373), .ZN(n529) );
  XNOR2_X1 U332 ( .A(n385), .B(n384), .ZN(n386) );
  XNOR2_X1 U333 ( .A(n415), .B(KEYINPUT64), .ZN(n564) );
  XNOR2_X1 U334 ( .A(n330), .B(n329), .ZN(n334) );
  INV_X1 U335 ( .A(n564), .ZN(n566) );
  XOR2_X1 U336 ( .A(n306), .B(n305), .Z(n458) );
  XNOR2_X1 U337 ( .A(n340), .B(n339), .ZN(n341) );
  NOR2_X1 U338 ( .A1(n453), .A2(n530), .ZN(n561) );
  INV_X1 U339 ( .A(G36GAT), .ZN(n476) );
  XOR2_X1 U340 ( .A(KEYINPUT99), .B(n468), .Z(n545) );
  XNOR2_X1 U341 ( .A(n480), .B(G190GAT), .ZN(n481) );
  XNOR2_X1 U342 ( .A(n476), .B(KEYINPUT108), .ZN(n477) );
  XNOR2_X1 U343 ( .A(n482), .B(n481), .ZN(G1351GAT) );
  XNOR2_X1 U344 ( .A(n478), .B(n477), .ZN(G1329GAT) );
  XOR2_X1 U345 ( .A(KEYINPUT73), .B(G92GAT), .Z(n293) );
  XNOR2_X1 U346 ( .A(G204GAT), .B(G85GAT), .ZN(n292) );
  XNOR2_X1 U347 ( .A(n293), .B(n292), .ZN(n306) );
  XOR2_X1 U348 ( .A(G176GAT), .B(G64GAT), .Z(n387) );
  XOR2_X1 U349 ( .A(KEYINPUT70), .B(KEYINPUT13), .Z(n295) );
  XNOR2_X1 U350 ( .A(G71GAT), .B(G78GAT), .ZN(n294) );
  XNOR2_X1 U351 ( .A(n295), .B(n294), .ZN(n358) );
  NAND2_X1 U352 ( .A1(G230GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U353 ( .A(n291), .B(n296), .ZN(n300) );
  XOR2_X1 U354 ( .A(KEYINPUT31), .B(KEYINPUT33), .Z(n298) );
  XNOR2_X1 U355 ( .A(KEYINPUT72), .B(KEYINPUT32), .ZN(n297) );
  XNOR2_X1 U356 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U357 ( .A(n300), .B(n299), .Z(n304) );
  XNOR2_X1 U358 ( .A(G120GAT), .B(G148GAT), .ZN(n301) );
  XNOR2_X1 U359 ( .A(n301), .B(G57GAT), .ZN(n398) );
  XNOR2_X1 U360 ( .A(G99GAT), .B(G106GAT), .ZN(n302) );
  XNOR2_X1 U361 ( .A(n302), .B(KEYINPUT71), .ZN(n335) );
  XNOR2_X1 U362 ( .A(n398), .B(n335), .ZN(n303) );
  XNOR2_X1 U363 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U364 ( .A(n458), .B(KEYINPUT41), .ZN(n507) );
  XOR2_X1 U365 ( .A(KEYINPUT65), .B(KEYINPUT66), .Z(n308) );
  XNOR2_X1 U366 ( .A(G197GAT), .B(KEYINPUT30), .ZN(n307) );
  XNOR2_X1 U367 ( .A(n308), .B(n307), .ZN(n323) );
  XOR2_X1 U368 ( .A(KEYINPUT67), .B(KEYINPUT68), .Z(n310) );
  NAND2_X1 U369 ( .A1(G229GAT), .A2(G233GAT), .ZN(n309) );
  XNOR2_X1 U370 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U371 ( .A(n311), .B(KEYINPUT29), .Z(n315) );
  XNOR2_X1 U372 ( .A(G43GAT), .B(KEYINPUT8), .ZN(n312) );
  XNOR2_X1 U373 ( .A(n312), .B(KEYINPUT7), .ZN(n336) );
  XNOR2_X1 U374 ( .A(G15GAT), .B(G22GAT), .ZN(n313) );
  XNOR2_X1 U375 ( .A(n313), .B(KEYINPUT69), .ZN(n354) );
  XNOR2_X1 U376 ( .A(n336), .B(n354), .ZN(n314) );
  XNOR2_X1 U377 ( .A(n315), .B(n314), .ZN(n319) );
  XOR2_X1 U378 ( .A(G141GAT), .B(G29GAT), .Z(n317) );
  XNOR2_X1 U379 ( .A(G36GAT), .B(G50GAT), .ZN(n316) );
  XNOR2_X1 U380 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U381 ( .A(n319), .B(n318), .Z(n321) );
  XOR2_X1 U382 ( .A(G169GAT), .B(G8GAT), .Z(n383) );
  XOR2_X1 U383 ( .A(G113GAT), .B(G1GAT), .Z(n404) );
  XNOR2_X1 U384 ( .A(n383), .B(n404), .ZN(n320) );
  XNOR2_X1 U385 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U386 ( .A(n323), .B(n322), .Z(n567) );
  NAND2_X1 U387 ( .A1(n507), .A2(n567), .ZN(n325) );
  XNOR2_X1 U388 ( .A(G29GAT), .B(G134GAT), .ZN(n326) );
  XNOR2_X1 U389 ( .A(n326), .B(G85GAT), .ZN(n411) );
  XOR2_X1 U390 ( .A(G50GAT), .B(G162GAT), .Z(n424) );
  XOR2_X1 U391 ( .A(n411), .B(n424), .Z(n330) );
  NAND2_X1 U392 ( .A1(G232GAT), .A2(G233GAT), .ZN(n328) );
  INV_X1 U393 ( .A(KEYINPUT10), .ZN(n327) );
  XOR2_X1 U394 ( .A(G92GAT), .B(G218GAT), .Z(n332) );
  XNOR2_X1 U395 ( .A(G36GAT), .B(G190GAT), .ZN(n331) );
  XNOR2_X1 U396 ( .A(n332), .B(n331), .ZN(n377) );
  XNOR2_X1 U397 ( .A(n377), .B(KEYINPUT74), .ZN(n333) );
  XNOR2_X1 U398 ( .A(n334), .B(n333), .ZN(n342) );
  XNOR2_X1 U399 ( .A(n336), .B(n335), .ZN(n340) );
  XOR2_X1 U400 ( .A(KEYINPUT75), .B(KEYINPUT76), .Z(n338) );
  XNOR2_X1 U401 ( .A(KEYINPUT11), .B(KEYINPUT9), .ZN(n337) );
  XOR2_X1 U402 ( .A(n338), .B(n337), .Z(n339) );
  XOR2_X1 U403 ( .A(KEYINPUT78), .B(KEYINPUT79), .Z(n344) );
  XNOR2_X1 U404 ( .A(KEYINPUT82), .B(KEYINPUT12), .ZN(n343) );
  XNOR2_X1 U405 ( .A(n344), .B(n343), .ZN(n362) );
  XOR2_X1 U406 ( .A(G64GAT), .B(G57GAT), .Z(n346) );
  XNOR2_X1 U407 ( .A(G211GAT), .B(G155GAT), .ZN(n345) );
  XNOR2_X1 U408 ( .A(n346), .B(n345), .ZN(n350) );
  XOR2_X1 U409 ( .A(KEYINPUT81), .B(KEYINPUT80), .Z(n348) );
  XNOR2_X1 U410 ( .A(G8GAT), .B(G1GAT), .ZN(n347) );
  XNOR2_X1 U411 ( .A(n348), .B(n347), .ZN(n349) );
  XOR2_X1 U412 ( .A(n350), .B(n349), .Z(n356) );
  XOR2_X1 U413 ( .A(G183GAT), .B(G127GAT), .Z(n352) );
  NAND2_X1 U414 ( .A1(G231GAT), .A2(G233GAT), .ZN(n351) );
  XNOR2_X1 U415 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U416 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U417 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U418 ( .A(n357), .B(KEYINPUT14), .Z(n360) );
  XNOR2_X1 U419 ( .A(n358), .B(KEYINPUT15), .ZN(n359) );
  XNOR2_X1 U420 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U421 ( .A(n362), .B(n361), .ZN(n555) );
  INV_X1 U422 ( .A(n555), .ZN(n575) );
  NOR2_X1 U423 ( .A1(n557), .A2(n575), .ZN(n363) );
  AND2_X1 U424 ( .A1(n364), .A2(n363), .ZN(n365) );
  XNOR2_X1 U425 ( .A(n365), .B(KEYINPUT47), .ZN(n371) );
  XNOR2_X1 U426 ( .A(KEYINPUT77), .B(n557), .ZN(n479) );
  XNOR2_X1 U427 ( .A(KEYINPUT36), .B(n479), .ZN(n582) );
  NOR2_X1 U428 ( .A1(n582), .A2(n555), .ZN(n366) );
  XNOR2_X1 U429 ( .A(KEYINPUT45), .B(n366), .ZN(n367) );
  NAND2_X1 U430 ( .A1(n367), .A2(n458), .ZN(n368) );
  XNOR2_X1 U431 ( .A(n368), .B(KEYINPUT115), .ZN(n369) );
  INV_X1 U432 ( .A(n567), .ZN(n547) );
  NAND2_X1 U433 ( .A1(n369), .A2(n547), .ZN(n370) );
  NAND2_X1 U434 ( .A1(n371), .A2(n370), .ZN(n374) );
  INV_X1 U435 ( .A(KEYINPUT116), .ZN(n372) );
  XOR2_X1 U436 ( .A(G183GAT), .B(KEYINPUT17), .Z(n376) );
  XNOR2_X1 U437 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n375) );
  XNOR2_X1 U438 ( .A(n376), .B(n375), .ZN(n441) );
  XNOR2_X1 U439 ( .A(n441), .B(n377), .ZN(n391) );
  XOR2_X1 U440 ( .A(KEYINPUT91), .B(G204GAT), .Z(n379) );
  XNOR2_X1 U441 ( .A(G197GAT), .B(G211GAT), .ZN(n378) );
  XNOR2_X1 U442 ( .A(n379), .B(n378), .ZN(n381) );
  XOR2_X1 U443 ( .A(KEYINPUT90), .B(KEYINPUT21), .Z(n380) );
  XNOR2_X1 U444 ( .A(n381), .B(n380), .ZN(n433) );
  INV_X1 U445 ( .A(n433), .ZN(n385) );
  XOR2_X1 U446 ( .A(KEYINPUT100), .B(KEYINPUT101), .Z(n382) );
  XOR2_X1 U447 ( .A(n387), .B(n386), .Z(n389) );
  NAND2_X1 U448 ( .A1(G226GAT), .A2(G233GAT), .ZN(n388) );
  XNOR2_X1 U449 ( .A(n389), .B(n388), .ZN(n390) );
  NOR2_X1 U450 ( .A1(n529), .A2(n520), .ZN(n392) );
  XNOR2_X1 U451 ( .A(KEYINPUT54), .B(n392), .ZN(n414) );
  XOR2_X1 U452 ( .A(KEYINPUT6), .B(KEYINPUT98), .Z(n394) );
  NAND2_X1 U453 ( .A1(G225GAT), .A2(G233GAT), .ZN(n393) );
  XNOR2_X1 U454 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U455 ( .A(n395), .B(KEYINPUT96), .Z(n400) );
  XOR2_X1 U456 ( .A(G155GAT), .B(KEYINPUT2), .Z(n397) );
  XNOR2_X1 U457 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n396) );
  XNOR2_X1 U458 ( .A(n397), .B(n396), .ZN(n425) );
  XNOR2_X1 U459 ( .A(n425), .B(n398), .ZN(n399) );
  XNOR2_X1 U460 ( .A(n400), .B(n399), .ZN(n408) );
  XOR2_X1 U461 ( .A(KEYINPUT1), .B(KEYINPUT97), .Z(n402) );
  XNOR2_X1 U462 ( .A(KEYINPUT4), .B(KEYINPUT95), .ZN(n401) );
  XNOR2_X1 U463 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U464 ( .A(n403), .B(KEYINPUT5), .Z(n406) );
  XNOR2_X1 U465 ( .A(n404), .B(G162GAT), .ZN(n405) );
  XNOR2_X1 U466 ( .A(n406), .B(n405), .ZN(n407) );
  XOR2_X1 U467 ( .A(n408), .B(n407), .Z(n413) );
  XOR2_X1 U468 ( .A(G127GAT), .B(KEYINPUT85), .Z(n410) );
  XNOR2_X1 U469 ( .A(KEYINPUT0), .B(KEYINPUT84), .ZN(n409) );
  XNOR2_X1 U470 ( .A(n410), .B(n409), .ZN(n442) );
  XNOR2_X1 U471 ( .A(n442), .B(n411), .ZN(n412) );
  XNOR2_X1 U472 ( .A(n413), .B(n412), .ZN(n468) );
  NAND2_X1 U473 ( .A1(n414), .A2(n545), .ZN(n415) );
  XOR2_X1 U474 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n417) );
  XNOR2_X1 U475 ( .A(G218GAT), .B(G106GAT), .ZN(n416) );
  XNOR2_X1 U476 ( .A(n417), .B(n416), .ZN(n421) );
  XOR2_X1 U477 ( .A(G78GAT), .B(G148GAT), .Z(n419) );
  XNOR2_X1 U478 ( .A(G22GAT), .B(KEYINPUT22), .ZN(n418) );
  XNOR2_X1 U479 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U480 ( .A(n421), .B(n420), .Z(n431) );
  XOR2_X1 U481 ( .A(KEYINPUT94), .B(KEYINPUT89), .Z(n423) );
  XNOR2_X1 U482 ( .A(KEYINPUT93), .B(KEYINPUT92), .ZN(n422) );
  XNOR2_X1 U483 ( .A(n423), .B(n422), .ZN(n429) );
  XOR2_X1 U484 ( .A(n425), .B(n424), .Z(n427) );
  NAND2_X1 U485 ( .A1(G228GAT), .A2(G233GAT), .ZN(n426) );
  XNOR2_X1 U486 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U487 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U488 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U489 ( .A(n433), .B(n432), .ZN(n464) );
  NOR2_X1 U490 ( .A1(n564), .A2(n464), .ZN(n434) );
  XNOR2_X1 U491 ( .A(n434), .B(KEYINPUT55), .ZN(n453) );
  XOR2_X1 U492 ( .A(KEYINPUT88), .B(G71GAT), .Z(n436) );
  XNOR2_X1 U493 ( .A(G15GAT), .B(KEYINPUT20), .ZN(n435) );
  XNOR2_X1 U494 ( .A(n436), .B(n435), .ZN(n452) );
  XOR2_X1 U495 ( .A(G120GAT), .B(G134GAT), .Z(n438) );
  XNOR2_X1 U496 ( .A(G113GAT), .B(G99GAT), .ZN(n437) );
  XNOR2_X1 U497 ( .A(n438), .B(n437), .ZN(n440) );
  XOR2_X1 U498 ( .A(G43GAT), .B(G190GAT), .Z(n439) );
  XNOR2_X1 U499 ( .A(n440), .B(n439), .ZN(n448) );
  XNOR2_X1 U500 ( .A(n442), .B(n441), .ZN(n446) );
  XOR2_X1 U501 ( .A(KEYINPUT86), .B(KEYINPUT87), .Z(n444) );
  XNOR2_X1 U502 ( .A(G169GAT), .B(G176GAT), .ZN(n443) );
  XNOR2_X1 U503 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U504 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U505 ( .A(n448), .B(n447), .ZN(n450) );
  NAND2_X1 U506 ( .A1(G227GAT), .A2(G233GAT), .ZN(n449) );
  XNOR2_X1 U507 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U508 ( .A(n452), .B(n451), .ZN(n530) );
  NAND2_X1 U509 ( .A1(n561), .A2(n507), .ZN(n457) );
  XOR2_X1 U510 ( .A(KEYINPUT57), .B(KEYINPUT121), .Z(n455) );
  XOR2_X1 U511 ( .A(G176GAT), .B(KEYINPUT56), .Z(n454) );
  XNOR2_X1 U512 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U513 ( .A(n457), .B(n456), .ZN(G1349GAT) );
  INV_X1 U514 ( .A(n458), .ZN(n572) );
  NOR2_X1 U515 ( .A1(n547), .A2(n572), .ZN(n488) );
  XOR2_X1 U516 ( .A(n464), .B(KEYINPUT28), .Z(n525) );
  XOR2_X1 U517 ( .A(n520), .B(KEYINPUT102), .Z(n459) );
  XNOR2_X1 U518 ( .A(KEYINPUT27), .B(n459), .ZN(n466) );
  NAND2_X1 U519 ( .A1(n525), .A2(n466), .ZN(n460) );
  NOR2_X1 U520 ( .A1(n545), .A2(n460), .ZN(n532) );
  AND2_X1 U521 ( .A1(n532), .A2(n530), .ZN(n461) );
  XNOR2_X1 U522 ( .A(n461), .B(KEYINPUT103), .ZN(n471) );
  NOR2_X1 U523 ( .A1(n520), .A2(n530), .ZN(n462) );
  NOR2_X1 U524 ( .A1(n464), .A2(n462), .ZN(n463) );
  XNOR2_X1 U525 ( .A(KEYINPUT25), .B(n463), .ZN(n467) );
  NAND2_X1 U526 ( .A1(n530), .A2(n464), .ZN(n465) );
  XOR2_X1 U527 ( .A(n465), .B(KEYINPUT26), .Z(n565) );
  NAND2_X1 U528 ( .A1(n565), .A2(n466), .ZN(n544) );
  NAND2_X1 U529 ( .A1(n467), .A2(n544), .ZN(n469) );
  NAND2_X1 U530 ( .A1(n469), .A2(n468), .ZN(n470) );
  NAND2_X1 U531 ( .A1(n471), .A2(n470), .ZN(n472) );
  XNOR2_X1 U532 ( .A(n472), .B(KEYINPUT104), .ZN(n486) );
  NOR2_X1 U533 ( .A1(n582), .A2(n575), .ZN(n473) );
  NAND2_X1 U534 ( .A1(n486), .A2(n473), .ZN(n474) );
  XNOR2_X1 U535 ( .A(KEYINPUT37), .B(n474), .ZN(n518) );
  NAND2_X1 U536 ( .A1(n488), .A2(n518), .ZN(n475) );
  XNOR2_X1 U537 ( .A(n475), .B(KEYINPUT38), .ZN(n503) );
  NOR2_X1 U538 ( .A1(n520), .A2(n503), .ZN(n478) );
  INV_X1 U539 ( .A(n479), .ZN(n483) );
  NAND2_X1 U540 ( .A1(n561), .A2(n483), .ZN(n482) );
  XOR2_X1 U541 ( .A(KEYINPUT58), .B(KEYINPUT123), .Z(n480) );
  NAND2_X1 U542 ( .A1(n479), .A2(n575), .ZN(n484) );
  XNOR2_X1 U543 ( .A(n484), .B(KEYINPUT83), .ZN(n485) );
  XNOR2_X1 U544 ( .A(KEYINPUT16), .B(n485), .ZN(n487) );
  AND2_X1 U545 ( .A1(n487), .A2(n486), .ZN(n508) );
  NAND2_X1 U546 ( .A1(n488), .A2(n508), .ZN(n495) );
  NOR2_X1 U547 ( .A1(n545), .A2(n495), .ZN(n489) );
  XOR2_X1 U548 ( .A(G1GAT), .B(n489), .Z(n490) );
  XNOR2_X1 U549 ( .A(KEYINPUT34), .B(n490), .ZN(G1324GAT) );
  NOR2_X1 U550 ( .A1(n520), .A2(n495), .ZN(n492) );
  XNOR2_X1 U551 ( .A(G8GAT), .B(KEYINPUT105), .ZN(n491) );
  XNOR2_X1 U552 ( .A(n492), .B(n491), .ZN(G1325GAT) );
  NOR2_X1 U553 ( .A1(n530), .A2(n495), .ZN(n494) );
  XNOR2_X1 U554 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n493) );
  XNOR2_X1 U555 ( .A(n494), .B(n493), .ZN(G1326GAT) );
  NOR2_X1 U556 ( .A1(n525), .A2(n495), .ZN(n496) );
  XOR2_X1 U557 ( .A(KEYINPUT106), .B(n496), .Z(n497) );
  XNOR2_X1 U558 ( .A(G22GAT), .B(n497), .ZN(G1327GAT) );
  NOR2_X1 U559 ( .A1(n545), .A2(n503), .ZN(n500) );
  XOR2_X1 U560 ( .A(G29GAT), .B(KEYINPUT107), .Z(n498) );
  XNOR2_X1 U561 ( .A(KEYINPUT39), .B(n498), .ZN(n499) );
  XNOR2_X1 U562 ( .A(n500), .B(n499), .ZN(G1328GAT) );
  NOR2_X1 U563 ( .A1(n503), .A2(n530), .ZN(n501) );
  XOR2_X1 U564 ( .A(KEYINPUT40), .B(n501), .Z(n502) );
  XNOR2_X1 U565 ( .A(G43GAT), .B(n502), .ZN(G1330GAT) );
  NOR2_X1 U566 ( .A1(n525), .A2(n503), .ZN(n504) );
  XOR2_X1 U567 ( .A(G50GAT), .B(n504), .Z(G1331GAT) );
  XOR2_X1 U568 ( .A(KEYINPUT110), .B(KEYINPUT42), .Z(n506) );
  XNOR2_X1 U569 ( .A(G57GAT), .B(KEYINPUT109), .ZN(n505) );
  XNOR2_X1 U570 ( .A(n506), .B(n505), .ZN(n510) );
  INV_X1 U571 ( .A(n507), .ZN(n551) );
  NOR2_X1 U572 ( .A1(n567), .A2(n551), .ZN(n517) );
  NAND2_X1 U573 ( .A1(n517), .A2(n508), .ZN(n513) );
  NOR2_X1 U574 ( .A1(n545), .A2(n513), .ZN(n509) );
  XOR2_X1 U575 ( .A(n510), .B(n509), .Z(G1332GAT) );
  NOR2_X1 U576 ( .A1(n520), .A2(n513), .ZN(n511) );
  XOR2_X1 U577 ( .A(G64GAT), .B(n511), .Z(G1333GAT) );
  NOR2_X1 U578 ( .A1(n530), .A2(n513), .ZN(n512) );
  XOR2_X1 U579 ( .A(G71GAT), .B(n512), .Z(G1334GAT) );
  NOR2_X1 U580 ( .A1(n525), .A2(n513), .ZN(n515) );
  XNOR2_X1 U581 ( .A(KEYINPUT43), .B(KEYINPUT111), .ZN(n514) );
  XNOR2_X1 U582 ( .A(n515), .B(n514), .ZN(n516) );
  XOR2_X1 U583 ( .A(G78GAT), .B(n516), .Z(G1335GAT) );
  NAND2_X1 U584 ( .A1(n518), .A2(n517), .ZN(n524) );
  NOR2_X1 U585 ( .A1(n545), .A2(n524), .ZN(n519) );
  XOR2_X1 U586 ( .A(G85GAT), .B(n519), .Z(G1336GAT) );
  NOR2_X1 U587 ( .A1(n520), .A2(n524), .ZN(n521) );
  XOR2_X1 U588 ( .A(KEYINPUT112), .B(n521), .Z(n522) );
  XNOR2_X1 U589 ( .A(G92GAT), .B(n522), .ZN(G1337GAT) );
  NOR2_X1 U590 ( .A1(n530), .A2(n524), .ZN(n523) );
  XOR2_X1 U591 ( .A(G99GAT), .B(n523), .Z(G1338GAT) );
  NOR2_X1 U592 ( .A1(n525), .A2(n524), .ZN(n527) );
  XNOR2_X1 U593 ( .A(KEYINPUT113), .B(KEYINPUT44), .ZN(n526) );
  XNOR2_X1 U594 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U595 ( .A(G106GAT), .B(n528), .ZN(G1339GAT) );
  NOR2_X1 U596 ( .A1(n529), .A2(n530), .ZN(n531) );
  NAND2_X1 U597 ( .A1(n532), .A2(n531), .ZN(n540) );
  NOR2_X1 U598 ( .A1(n547), .A2(n540), .ZN(n533) );
  XOR2_X1 U599 ( .A(G113GAT), .B(n533), .Z(G1340GAT) );
  NOR2_X1 U600 ( .A1(n551), .A2(n540), .ZN(n535) );
  XNOR2_X1 U601 ( .A(KEYINPUT117), .B(KEYINPUT49), .ZN(n534) );
  XNOR2_X1 U602 ( .A(n535), .B(n534), .ZN(n536) );
  XOR2_X1 U603 ( .A(G120GAT), .B(n536), .Z(G1341GAT) );
  NOR2_X1 U604 ( .A1(n555), .A2(n540), .ZN(n538) );
  XNOR2_X1 U605 ( .A(KEYINPUT50), .B(KEYINPUT118), .ZN(n537) );
  XNOR2_X1 U606 ( .A(n538), .B(n537), .ZN(n539) );
  XOR2_X1 U607 ( .A(G127GAT), .B(n539), .Z(G1342GAT) );
  NOR2_X1 U608 ( .A1(n479), .A2(n540), .ZN(n542) );
  XNOR2_X1 U609 ( .A(KEYINPUT119), .B(KEYINPUT51), .ZN(n541) );
  XNOR2_X1 U610 ( .A(n542), .B(n541), .ZN(n543) );
  XOR2_X1 U611 ( .A(G134GAT), .B(n543), .Z(G1343GAT) );
  OR2_X1 U612 ( .A1(n529), .A2(n544), .ZN(n546) );
  NOR2_X1 U613 ( .A1(n546), .A2(n545), .ZN(n558) );
  INV_X1 U614 ( .A(n558), .ZN(n554) );
  NOR2_X1 U615 ( .A1(n547), .A2(n554), .ZN(n548) );
  XOR2_X1 U616 ( .A(G141GAT), .B(n548), .Z(G1344GAT) );
  XOR2_X1 U617 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n550) );
  XNOR2_X1 U618 ( .A(G148GAT), .B(KEYINPUT120), .ZN(n549) );
  XNOR2_X1 U619 ( .A(n550), .B(n549), .ZN(n553) );
  NOR2_X1 U620 ( .A1(n551), .A2(n554), .ZN(n552) );
  XOR2_X1 U621 ( .A(n553), .B(n552), .Z(G1345GAT) );
  NOR2_X1 U622 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U623 ( .A(G155GAT), .B(n556), .Z(G1346GAT) );
  NAND2_X1 U624 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U625 ( .A(n559), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U626 ( .A1(n561), .A2(n567), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n560), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U628 ( .A1(n561), .A2(n575), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n562), .B(KEYINPUT122), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n563), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U631 ( .A1(n566), .A2(n565), .ZN(n581) );
  INV_X1 U632 ( .A(n581), .ZN(n576) );
  NAND2_X1 U633 ( .A1(n576), .A2(n567), .ZN(n571) );
  XOR2_X1 U634 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n569) );
  XNOR2_X1 U635 ( .A(G197GAT), .B(KEYINPUT124), .ZN(n568) );
  XNOR2_X1 U636 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(G1352GAT) );
  XOR2_X1 U638 ( .A(G204GAT), .B(KEYINPUT61), .Z(n574) );
  NAND2_X1 U639 ( .A1(n576), .A2(n572), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(G1353GAT) );
  XOR2_X1 U641 ( .A(G211GAT), .B(KEYINPUT125), .Z(n578) );
  NAND2_X1 U642 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(G1354GAT) );
  XOR2_X1 U644 ( .A(KEYINPUT62), .B(KEYINPUT126), .Z(n580) );
  XNOR2_X1 U645 ( .A(G218GAT), .B(KEYINPUT127), .ZN(n579) );
  XNOR2_X1 U646 ( .A(n580), .B(n579), .ZN(n584) );
  NOR2_X1 U647 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U648 ( .A(n584), .B(n583), .Z(G1355GAT) );
endmodule

