//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 0 1 0 0 1 1 1 1 0 0 0 1 1 1 1 0 0 1 0 0 1 0 0 0 0 1 1 1 0 1 0 0 1 1 0 0 1 0 1 1 0 1 0 1 1 1 0 1 1 1 1 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:44 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n613, new_n614, new_n615,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n651, new_n652, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n667, new_n668, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n890, new_n891, new_n892, new_n893, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  XOR2_X1   g001(.A(KEYINPUT72), .B(G902), .Z(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  AOI21_X1  g003(.A(new_n187), .B1(new_n189), .B2(G234), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT22), .B(G137), .ZN(new_n192));
  INV_X1    g006(.A(G221), .ZN(new_n193));
  INV_X1    g007(.A(G234), .ZN(new_n194));
  NOR3_X1   g008(.A1(new_n193), .A2(new_n194), .A3(G953), .ZN(new_n195));
  XOR2_X1   g009(.A(new_n192), .B(new_n195), .Z(new_n196));
  INV_X1    g010(.A(G119), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G128), .ZN(new_n198));
  INV_X1    g012(.A(G128), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G119), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n198), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(new_n201), .ZN(new_n202));
  XOR2_X1   g016(.A(KEYINPUT24), .B(G110), .Z(new_n203));
  NOR2_X1   g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  XNOR2_X1  g018(.A(new_n200), .B(KEYINPUT23), .ZN(new_n205));
  INV_X1    g019(.A(G110), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n205), .A2(new_n206), .A3(new_n198), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT75), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n204), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n209), .B1(new_n208), .B2(new_n207), .ZN(new_n210));
  INV_X1    g024(.A(G140), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G125), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT16), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT73), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n212), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G125), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G140), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(KEYINPUT73), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n216), .B1(new_n212), .B2(new_n219), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n214), .B1(new_n220), .B2(new_n213), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G146), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n212), .A2(new_n218), .ZN(new_n223));
  OAI211_X1 g037(.A(new_n210), .B(new_n222), .C1(G146), .C2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(G146), .ZN(new_n225));
  OAI211_X1 g039(.A(new_n225), .B(new_n214), .C1(new_n220), .C2(new_n213), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n222), .A2(KEYINPUT74), .A3(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT74), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n221), .A2(new_n228), .A3(G146), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n206), .B1(new_n205), .B2(new_n198), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n230), .B1(new_n202), .B2(new_n203), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n227), .A2(new_n229), .A3(new_n231), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n196), .B1(new_n224), .B2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(new_n233), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n224), .A2(new_n232), .A3(new_n196), .ZN(new_n235));
  AND2_X1   g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n236), .A2(KEYINPUT25), .A3(new_n189), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n234), .A2(new_n189), .A3(new_n235), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT25), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n191), .B1(new_n237), .B2(new_n240), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n190), .A2(G902), .ZN(new_n242));
  AND2_X1   g056(.A1(new_n236), .A2(new_n242), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(G953), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(G227), .ZN(new_n246));
  XNOR2_X1  g060(.A(new_n246), .B(KEYINPUT76), .ZN(new_n247));
  XNOR2_X1  g061(.A(G110), .B(G140), .ZN(new_n248));
  XNOR2_X1  g062(.A(new_n247), .B(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT10), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT78), .ZN(new_n251));
  XNOR2_X1  g065(.A(G104), .B(G107), .ZN(new_n252));
  INV_X1    g066(.A(G101), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n251), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(G104), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G107), .ZN(new_n256));
  INV_X1    g070(.A(G107), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G104), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n259), .A2(KEYINPUT78), .A3(G101), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n257), .A2(G104), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT3), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n262), .B1(new_n255), .B2(G107), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n257), .A2(KEYINPUT3), .A3(G104), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n261), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  AOI22_X1  g079(.A1(new_n254), .A2(new_n260), .B1(new_n265), .B2(new_n253), .ZN(new_n266));
  XNOR2_X1  g080(.A(G143), .B(G146), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n199), .A2(KEYINPUT1), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(G143), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n270), .A2(KEYINPUT1), .A3(G146), .ZN(new_n271));
  OAI211_X1 g085(.A(new_n269), .B(new_n271), .C1(G128), .C2(new_n267), .ZN(new_n272));
  AND3_X1   g086(.A1(new_n266), .A2(KEYINPUT79), .A3(new_n272), .ZN(new_n273));
  AOI21_X1  g087(.A(KEYINPUT79), .B1(new_n266), .B2(new_n272), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n250), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n225), .A2(G143), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n270), .A2(G146), .ZN(new_n277));
  AOI21_X1  g091(.A(G128), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n271), .ZN(new_n279));
  OAI21_X1  g093(.A(KEYINPUT67), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT67), .ZN(new_n281));
  OAI211_X1 g095(.A(new_n271), .B(new_n281), .C1(new_n267), .C2(G128), .ZN(new_n282));
  AOI22_X1  g096(.A1(new_n280), .A2(new_n282), .B1(new_n267), .B2(new_n268), .ZN(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n284), .A2(KEYINPUT10), .A3(new_n266), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT4), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n286), .B1(new_n265), .B2(new_n253), .ZN(new_n287));
  AND3_X1   g101(.A1(new_n257), .A2(KEYINPUT3), .A3(G104), .ZN(new_n288));
  AOI21_X1  g102(.A(KEYINPUT3), .B1(new_n257), .B2(G104), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n256), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(G101), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n287), .A2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT0), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n267), .B1(new_n293), .B2(new_n199), .ZN(new_n294));
  XOR2_X1   g108(.A(KEYINPUT0), .B(G128), .Z(new_n295));
  OAI21_X1  g109(.A(new_n294), .B1(new_n267), .B2(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n290), .A2(new_n286), .A3(G101), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n292), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(KEYINPUT77), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT77), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n292), .A2(new_n300), .A3(new_n296), .A4(new_n297), .ZN(new_n301));
  NAND4_X1  g115(.A1(new_n275), .A2(new_n285), .A3(new_n299), .A4(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT11), .ZN(new_n303));
  XNOR2_X1  g117(.A(KEYINPUT65), .B(G134), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(G137), .ZN(new_n305));
  INV_X1    g119(.A(G137), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(G134), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n303), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n303), .B1(new_n304), .B2(G137), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  OAI21_X1  g124(.A(G131), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(G131), .ZN(new_n312));
  INV_X1    g126(.A(new_n307), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n313), .B1(new_n304), .B2(G137), .ZN(new_n314));
  OAI211_X1 g128(.A(new_n312), .B(new_n309), .C1(new_n314), .C2(new_n303), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n311), .A2(KEYINPUT66), .A3(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT66), .ZN(new_n317));
  OAI211_X1 g131(.A(new_n317), .B(G131), .C1(new_n308), .C2(new_n310), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n249), .B1(new_n302), .B2(new_n320), .ZN(new_n321));
  OAI22_X1  g135(.A1(new_n273), .A2(new_n274), .B1(new_n284), .B2(new_n266), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n320), .A2(KEYINPUT12), .A3(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT12), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n266), .A2(new_n272), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT79), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n266), .A2(new_n272), .A3(KEYINPUT79), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n265), .A2(new_n253), .ZN(new_n329));
  AOI21_X1  g143(.A(KEYINPUT78), .B1(new_n259), .B2(G101), .ZN(new_n330));
  AOI211_X1 g144(.A(new_n251), .B(new_n253), .C1(new_n256), .C2(new_n258), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n329), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  AOI22_X1  g146(.A1(new_n327), .A2(new_n328), .B1(new_n283), .B2(new_n332), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n324), .B1(new_n333), .B2(new_n319), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n321), .B1(new_n323), .B2(new_n334), .ZN(new_n335));
  AND2_X1   g149(.A1(new_n299), .A2(new_n301), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n336), .A2(new_n319), .A3(new_n275), .A4(new_n285), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT81), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n302), .A2(new_n338), .A3(new_n320), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n338), .B1(new_n302), .B2(new_n320), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n337), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(new_n249), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n335), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NOR3_X1   g158(.A1(new_n344), .A2(G469), .A3(new_n188), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n321), .A2(KEYINPUT80), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT80), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n337), .A2(new_n347), .A3(new_n249), .ZN(new_n348));
  OAI211_X1 g162(.A(new_n346), .B(new_n348), .C1(new_n340), .C2(new_n341), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n323), .A2(new_n334), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(new_n337), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(new_n343), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n349), .A2(G469), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(G469), .A2(G902), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n345), .A2(new_n355), .ZN(new_n356));
  OAI21_X1  g170(.A(G214), .B1(G237), .B2(G902), .ZN(new_n357));
  XOR2_X1   g171(.A(new_n357), .B(KEYINPUT82), .Z(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  XOR2_X1   g173(.A(KEYINPUT9), .B(G234), .Z(new_n360));
  INV_X1    g174(.A(G902), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n193), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n359), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n296), .A2(G125), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n365), .B1(new_n283), .B2(G125), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n245), .A2(G224), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(new_n367), .ZN(new_n369));
  OAI211_X1 g183(.A(new_n369), .B(new_n365), .C1(new_n283), .C2(G125), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT6), .ZN(new_n372));
  AND2_X1   g186(.A1(KEYINPUT2), .A2(G113), .ZN(new_n373));
  NOR2_X1   g187(.A1(KEYINPUT2), .A2(G113), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  XNOR2_X1  g190(.A(G116), .B(G119), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n376), .A2(new_n378), .A3(KEYINPUT68), .ZN(new_n379));
  AOI21_X1  g193(.A(KEYINPUT68), .B1(new_n375), .B2(new_n377), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n380), .B1(new_n377), .B2(new_n375), .ZN(new_n381));
  NAND4_X1  g195(.A1(new_n292), .A2(new_n379), .A3(new_n381), .A4(new_n297), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n254), .A2(new_n260), .ZN(new_n383));
  INV_X1    g197(.A(G113), .ZN(new_n384));
  INV_X1    g198(.A(G116), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n385), .A2(G119), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT5), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n384), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n197), .A2(G116), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n385), .A2(G119), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n389), .A2(new_n390), .A3(KEYINPUT5), .ZN(new_n391));
  AOI22_X1  g205(.A1(new_n388), .A2(new_n391), .B1(new_n377), .B2(new_n375), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n383), .A2(new_n392), .A3(new_n329), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT83), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n266), .A2(KEYINPUT83), .A3(new_n392), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n382), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  XNOR2_X1  g211(.A(G110), .B(G122), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n398), .A2(KEYINPUT84), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n382), .A2(new_n395), .A3(new_n398), .A4(new_n396), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n372), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  AOI21_X1  g216(.A(KEYINPUT6), .B1(new_n397), .B2(new_n399), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n371), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  XOR2_X1   g218(.A(new_n398), .B(KEYINPUT8), .Z(new_n405));
  INV_X1    g219(.A(new_n392), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n332), .A2(new_n406), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n405), .B1(new_n407), .B2(new_n393), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT85), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n370), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(new_n405), .ZN(new_n411));
  AND3_X1   g225(.A1(new_n383), .A2(new_n329), .A3(new_n392), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n392), .B1(new_n383), .B2(new_n329), .ZN(new_n413));
  OAI211_X1 g227(.A(new_n409), .B(new_n411), .C1(new_n412), .C2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT7), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n415), .B(new_n365), .C1(new_n283), .C2(G125), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n410), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n366), .A2(KEYINPUT7), .A3(new_n367), .ZN(new_n419));
  AND2_X1   g233(.A1(new_n419), .A2(new_n401), .ZN(new_n420));
  AOI21_X1  g234(.A(G902), .B1(new_n418), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n404), .A2(new_n421), .ZN(new_n422));
  OAI21_X1  g236(.A(G210), .B1(G237), .B2(G902), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n404), .A2(new_n421), .A3(new_n423), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n425), .A2(KEYINPUT86), .A3(new_n426), .ZN(new_n427));
  AND3_X1   g241(.A1(new_n404), .A2(new_n423), .A3(new_n421), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT86), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n427), .A2(new_n430), .ZN(new_n431));
  NOR3_X1   g245(.A1(new_n356), .A2(new_n364), .A3(new_n431), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n304), .A2(G137), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n306), .A2(G134), .ZN(new_n434));
  OAI21_X1  g248(.A(G131), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n284), .A2(new_n315), .A3(new_n435), .ZN(new_n436));
  XNOR2_X1  g250(.A(new_n296), .B(KEYINPUT64), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n436), .B1(new_n319), .B2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT30), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n381), .A2(new_n379), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n296), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n436), .B1(new_n319), .B2(new_n443), .ZN(new_n444));
  OAI211_X1 g258(.A(new_n440), .B(new_n442), .C1(new_n439), .C2(new_n444), .ZN(new_n445));
  XOR2_X1   g259(.A(new_n441), .B(KEYINPUT69), .Z(new_n446));
  OAI211_X1 g260(.A(new_n446), .B(new_n436), .C1(new_n319), .C2(new_n443), .ZN(new_n447));
  XNOR2_X1  g261(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n448));
  INV_X1    g262(.A(G237), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n449), .A2(new_n245), .A3(G210), .ZN(new_n450));
  XNOR2_X1  g264(.A(new_n448), .B(new_n450), .ZN(new_n451));
  XNOR2_X1  g265(.A(KEYINPUT26), .B(G101), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n445), .A2(new_n447), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(KEYINPUT31), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n453), .B(KEYINPUT71), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT28), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n438), .A2(new_n442), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n457), .B1(new_n447), .B2(new_n458), .ZN(new_n459));
  AND2_X1   g273(.A1(new_n447), .A2(new_n457), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n456), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT31), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n445), .A2(new_n462), .A3(new_n447), .A4(new_n453), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n455), .A2(new_n461), .A3(new_n463), .ZN(new_n464));
  NOR2_X1   g278(.A1(G472), .A2(G902), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT32), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n445), .A2(new_n447), .ZN(new_n469));
  INV_X1    g283(.A(new_n453), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT29), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n447), .A2(new_n457), .ZN(new_n473));
  INV_X1    g287(.A(new_n456), .ZN(new_n474));
  AND2_X1   g288(.A1(new_n447), .A2(new_n458), .ZN(new_n475));
  OAI211_X1 g289(.A(new_n473), .B(new_n474), .C1(new_n475), .C2(new_n457), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n471), .A2(new_n472), .A3(new_n476), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n441), .B(KEYINPUT69), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n444), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n447), .A2(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n460), .B1(new_n480), .B2(KEYINPUT28), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n470), .A2(new_n472), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n188), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n477), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(G472), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n464), .A2(KEYINPUT32), .A3(new_n465), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n468), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT20), .ZN(new_n488));
  NOR2_X1   g302(.A1(G475), .A2(G902), .ZN(new_n489));
  INV_X1    g303(.A(G214), .ZN(new_n490));
  NOR3_X1   g304(.A1(new_n490), .A2(G237), .A3(G953), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n491), .B1(KEYINPUT87), .B2(G143), .ZN(new_n492));
  XOR2_X1   g306(.A(KEYINPUT87), .B(G143), .Z(new_n493));
  OAI21_X1  g307(.A(new_n492), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(G131), .ZN(new_n495));
  OAI211_X1 g309(.A(new_n492), .B(new_n312), .C1(new_n491), .C2(new_n493), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  MUX2_X1   g311(.A(new_n497), .B(new_n495), .S(KEYINPUT17), .Z(new_n498));
  NAND2_X1  g312(.A1(new_n227), .A2(new_n229), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n494), .A2(KEYINPUT18), .A3(G131), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT88), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n494), .A2(KEYINPUT88), .A3(KEYINPUT18), .A4(G131), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n223), .A2(G146), .ZN(new_n505));
  INV_X1    g319(.A(new_n220), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n505), .B1(new_n506), .B2(G146), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n496), .B1(new_n494), .B2(KEYINPUT18), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AOI22_X1  g323(.A1(new_n498), .A2(new_n499), .B1(new_n504), .B2(new_n509), .ZN(new_n510));
  XNOR2_X1  g324(.A(G113), .B(G122), .ZN(new_n511));
  XNOR2_X1  g325(.A(KEYINPUT89), .B(G104), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n511), .B(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  AND2_X1   g328(.A1(new_n510), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n504), .A2(new_n509), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n223), .A2(KEYINPUT19), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n517), .B1(new_n506), .B2(KEYINPUT19), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(new_n225), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n519), .A2(new_n222), .A3(new_n497), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n514), .B1(new_n516), .B2(new_n520), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n488), .B(new_n489), .C1(new_n515), .C2(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n521), .B1(new_n510), .B2(new_n514), .ZN(new_n523));
  INV_X1    g337(.A(new_n489), .ZN(new_n524));
  OAI21_X1  g338(.A(KEYINPUT20), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n522), .A2(new_n525), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n510), .A2(new_n514), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n361), .B1(new_n515), .B2(new_n527), .ZN(new_n528));
  XOR2_X1   g342(.A(KEYINPUT90), .B(G475), .Z(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n526), .A2(KEYINPUT91), .A3(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  AOI21_X1  g346(.A(KEYINPUT91), .B1(new_n526), .B2(new_n530), .ZN(new_n533));
  OAI211_X1 g347(.A(G952), .B(new_n245), .C1(new_n194), .C2(new_n449), .ZN(new_n534));
  XNOR2_X1  g348(.A(new_n534), .B(KEYINPUT94), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  OAI211_X1 g350(.A(new_n188), .B(G953), .C1(new_n194), .C2(new_n449), .ZN(new_n537));
  XOR2_X1   g351(.A(new_n537), .B(KEYINPUT95), .Z(new_n538));
  XOR2_X1   g352(.A(KEYINPUT21), .B(G898), .Z(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n536), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n270), .A2(G128), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT13), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n270), .A2(G128), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n542), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n545), .B1(new_n543), .B2(new_n544), .ZN(new_n546));
  AND2_X1   g360(.A1(new_n546), .A2(G134), .ZN(new_n547));
  XOR2_X1   g361(.A(KEYINPUT92), .B(G107), .Z(new_n548));
  XNOR2_X1  g362(.A(G116), .B(G122), .ZN(new_n549));
  OR2_X1    g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  XNOR2_X1  g364(.A(G128), .B(G143), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n304), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n548), .A2(new_n549), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n550), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n547), .A2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(G122), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(G116), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n257), .B1(new_n557), .B2(KEYINPUT14), .ZN(new_n558));
  XNOR2_X1  g372(.A(new_n558), .B(new_n549), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n304), .B(new_n551), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT93), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n559), .A2(KEYINPUT93), .A3(new_n560), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n555), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n360), .ZN(new_n567));
  NOR3_X1   g381(.A1(new_n567), .A2(new_n187), .A3(G953), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n568), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n565), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n569), .A2(new_n189), .A3(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(G478), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n573), .A2(KEYINPUT15), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n572), .B(new_n574), .ZN(new_n575));
  NOR4_X1   g389(.A1(new_n532), .A2(new_n533), .A3(new_n541), .A4(new_n575), .ZN(new_n576));
  AND4_X1   g390(.A1(new_n244), .A2(new_n432), .A3(new_n487), .A4(new_n576), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n577), .B(new_n253), .ZN(G3));
  INV_X1    g392(.A(new_n244), .ZN(new_n579));
  INV_X1    g393(.A(new_n466), .ZN(new_n580));
  INV_X1    g394(.A(G472), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n581), .B1(new_n464), .B2(new_n189), .ZN(new_n582));
  NOR3_X1   g396(.A1(new_n579), .A2(new_n580), .A3(new_n582), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n356), .A2(new_n362), .ZN(new_n584));
  AND2_X1   g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT96), .ZN(new_n586));
  AND2_X1   g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n585), .A2(new_n586), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n358), .B1(new_n425), .B2(new_n426), .ZN(new_n589));
  INV_X1    g403(.A(new_n541), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NOR3_X1   g405(.A1(new_n587), .A2(new_n588), .A3(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT33), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n569), .A2(new_n593), .A3(new_n571), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT97), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n569), .A2(KEYINPUT97), .A3(new_n571), .A4(new_n593), .ZN(new_n597));
  OAI21_X1  g411(.A(KEYINPUT98), .B1(new_n570), .B2(KEYINPUT99), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n566), .A2(new_n598), .ZN(new_n599));
  AOI21_X1  g413(.A(KEYINPUT99), .B1(new_n565), .B2(KEYINPUT98), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n599), .B1(new_n600), .B2(new_n568), .ZN(new_n601));
  AOI22_X1  g415(.A1(new_n596), .A2(new_n597), .B1(KEYINPUT33), .B2(new_n601), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n188), .A2(new_n573), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(KEYINPUT100), .B(G478), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n572), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n607), .B1(new_n532), .B2(new_n533), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n592), .A2(new_n609), .ZN(new_n610));
  XOR2_X1   g424(.A(KEYINPUT34), .B(G104), .Z(new_n611));
  XNOR2_X1  g425(.A(new_n610), .B(new_n611), .ZN(G6));
  AND3_X1   g426(.A1(new_n526), .A2(new_n530), .A3(new_n575), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n592), .A2(new_n613), .ZN(new_n614));
  XOR2_X1   g428(.A(KEYINPUT35), .B(G107), .Z(new_n615));
  XNOR2_X1  g429(.A(new_n614), .B(new_n615), .ZN(G9));
  NOR2_X1   g430(.A1(new_n580), .A2(new_n582), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n224), .A2(new_n232), .ZN(new_n618));
  INV_X1    g432(.A(new_n196), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n619), .A2(KEYINPUT36), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n618), .B(new_n620), .ZN(new_n621));
  AND2_X1   g435(.A1(new_n621), .A2(new_n242), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n241), .A2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n432), .A2(new_n617), .A3(new_n576), .A4(new_n624), .ZN(new_n625));
  XOR2_X1   g439(.A(KEYINPUT37), .B(G110), .Z(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(KEYINPUT101), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n625), .B(new_n627), .ZN(G12));
  INV_X1    g442(.A(G900), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n536), .B1(new_n538), .B2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  AND2_X1   g445(.A1(new_n613), .A2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n589), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n623), .A2(new_n633), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n487), .A2(new_n584), .A3(new_n632), .A4(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(G128), .ZN(G30));
  OAI21_X1  g450(.A(new_n575), .B1(new_n532), .B2(new_n533), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n638), .A2(new_n359), .A3(new_n623), .ZN(new_n639));
  XOR2_X1   g453(.A(new_n639), .B(KEYINPUT102), .Z(new_n640));
  XNOR2_X1  g454(.A(new_n630), .B(KEYINPUT39), .ZN(new_n641));
  OR3_X1    g455(.A1(new_n356), .A2(new_n362), .A3(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(new_n642), .B(KEYINPUT40), .Z(new_n643));
  INV_X1    g457(.A(new_n469), .ZN(new_n644));
  AOI22_X1  g458(.A1(new_n644), .A2(new_n453), .B1(new_n456), .B2(new_n480), .ZN(new_n645));
  OAI21_X1  g459(.A(G472), .B1(new_n645), .B2(G902), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n468), .A2(new_n486), .A3(new_n646), .ZN(new_n647));
  XOR2_X1   g461(.A(new_n431), .B(KEYINPUT38), .Z(new_n648));
  NAND4_X1  g462(.A1(new_n640), .A2(new_n643), .A3(new_n647), .A4(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(G143), .ZN(G45));
  NOR2_X1   g464(.A1(new_n608), .A2(new_n630), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n651), .A2(new_n487), .A3(new_n584), .A4(new_n634), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(G146), .ZN(G48));
  NOR2_X1   g467(.A1(new_n608), .A2(new_n541), .ZN(new_n654));
  OAI21_X1  g468(.A(G469), .B1(new_n344), .B2(new_n188), .ZN(new_n655));
  INV_X1    g469(.A(G469), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n302), .A2(new_n320), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(KEYINPUT81), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(new_n339), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n249), .B1(new_n659), .B2(new_n337), .ZN(new_n660));
  OAI211_X1 g474(.A(new_n656), .B(new_n189), .C1(new_n660), .C2(new_n335), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n655), .A2(new_n661), .ZN(new_n662));
  NOR3_X1   g476(.A1(new_n662), .A2(new_n362), .A3(new_n633), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n654), .A2(new_n487), .A3(new_n244), .A4(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(KEYINPUT41), .B(G113), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G15));
  AND2_X1   g480(.A1(new_n613), .A2(new_n590), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n487), .A2(new_n663), .A3(new_n244), .A4(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(G116), .ZN(G18));
  NOR2_X1   g483(.A1(new_n662), .A2(new_n362), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n487), .A2(new_n576), .A3(new_n634), .A4(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G119), .ZN(G21));
  INV_X1    g486(.A(new_n465), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT103), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n481), .A2(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(new_n480), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n473), .B1(new_n676), .B2(new_n457), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(KEYINPUT103), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n675), .A2(new_n678), .A3(new_n456), .ZN(new_n679));
  AND2_X1   g493(.A1(new_n455), .A2(new_n463), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n673), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NOR3_X1   g495(.A1(new_n681), .A2(new_n579), .A3(new_n582), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n637), .A2(new_n591), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n682), .A2(new_n683), .A3(new_n670), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G122), .ZN(G24));
  NOR3_X1   g499(.A1(new_n681), .A2(new_n582), .A3(new_n623), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n686), .A2(new_n651), .A3(new_n663), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G125), .ZN(G27));
  NAND2_X1  g502(.A1(new_n487), .A2(new_n244), .ZN(new_n689));
  INV_X1    g503(.A(new_n651), .ZN(new_n690));
  OAI21_X1  g504(.A(KEYINPUT104), .B1(new_n345), .B2(new_n355), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT104), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n661), .A2(new_n692), .A3(new_n354), .A4(new_n353), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n691), .A2(new_n363), .A3(new_n693), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n423), .B1(new_n404), .B2(new_n421), .ZN(new_n695));
  NOR3_X1   g509(.A1(new_n428), .A2(new_n695), .A3(new_n429), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n426), .A2(KEYINPUT86), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n359), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(KEYINPUT105), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT105), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n431), .A2(new_n700), .A3(new_n359), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  OAI21_X1  g516(.A(KEYINPUT106), .B1(new_n694), .B2(new_n702), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n700), .B1(new_n431), .B2(new_n359), .ZN(new_n704));
  AOI211_X1 g518(.A(KEYINPUT105), .B(new_n358), .C1(new_n427), .C2(new_n430), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n661), .A2(new_n354), .A3(new_n353), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n362), .B1(new_n707), .B2(KEYINPUT104), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT106), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n706), .A2(new_n708), .A3(new_n709), .A4(new_n693), .ZN(new_n710));
  AOI211_X1 g524(.A(new_n689), .B(new_n690), .C1(new_n703), .C2(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT107), .ZN(new_n712));
  OAI211_X1 g526(.A(KEYINPUT108), .B(KEYINPUT42), .C1(new_n711), .C2(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT108), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n703), .A2(new_n710), .ZN(new_n715));
  INV_X1    g529(.A(new_n689), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n715), .A2(new_n716), .A3(new_n651), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n714), .B1(new_n717), .B2(KEYINPUT107), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT42), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n719), .B1(new_n717), .B2(new_n714), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n713), .B1(new_n718), .B2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G131), .ZN(G33));
  NAND3_X1  g536(.A1(new_n715), .A2(new_n716), .A3(new_n632), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G134), .ZN(G36));
  NOR2_X1   g538(.A1(new_n532), .A2(new_n533), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(new_n607), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT109), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(KEYINPUT43), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(KEYINPUT109), .B(KEYINPUT43), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n729), .B1(new_n726), .B2(new_n730), .ZN(new_n731));
  OAI211_X1 g545(.A(new_n731), .B(new_n624), .C1(new_n580), .C2(new_n582), .ZN(new_n732));
  OR2_X1    g546(.A1(new_n732), .A2(KEYINPUT44), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n732), .A2(KEYINPUT44), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n702), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  AND2_X1   g549(.A1(new_n349), .A2(new_n352), .ZN(new_n736));
  OR2_X1    g550(.A1(new_n736), .A2(KEYINPUT45), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n736), .A2(KEYINPUT45), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n737), .A2(G469), .A3(new_n738), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n739), .A2(KEYINPUT46), .A3(new_n354), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(new_n661), .ZN(new_n741));
  AOI21_X1  g555(.A(KEYINPUT46), .B1(new_n739), .B2(new_n354), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n363), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  OR2_X1    g557(.A1(new_n743), .A2(new_n641), .ZN(new_n744));
  INV_X1    g558(.A(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n735), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G137), .ZN(G39));
  XNOR2_X1  g561(.A(KEYINPUT110), .B(KEYINPUT47), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n743), .B(new_n748), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n651), .A2(new_n579), .A3(new_n706), .ZN(new_n750));
  OR3_X1    g564(.A1(new_n749), .A2(new_n487), .A3(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G140), .ZN(G42));
  NOR3_X1   g566(.A1(new_n648), .A2(new_n364), .A3(new_n726), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n647), .A2(new_n579), .ZN(new_n754));
  XOR2_X1   g568(.A(new_n662), .B(KEYINPUT49), .Z(new_n755));
  NAND3_X1  g569(.A1(new_n753), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT114), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n526), .A2(new_n530), .ZN(new_n758));
  NOR4_X1   g572(.A1(new_n623), .A2(new_n575), .A3(new_n758), .A4(new_n630), .ZN(new_n759));
  AND4_X1   g573(.A1(new_n487), .A2(new_n759), .A3(new_n706), .A4(new_n584), .ZN(new_n760));
  AND2_X1   g574(.A1(new_n686), .A2(new_n651), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n760), .B1(new_n715), .B2(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n762), .A2(KEYINPUT111), .A3(new_n723), .ZN(new_n763));
  INV_X1    g577(.A(new_n533), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n764), .A2(new_n531), .A3(new_n575), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n608), .A2(new_n765), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n583), .A2(new_n432), .A3(new_n766), .A4(new_n590), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n767), .A2(new_n684), .A3(new_n625), .A4(new_n671), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n664), .A2(new_n668), .ZN(new_n769));
  NOR3_X1   g583(.A1(new_n768), .A2(new_n769), .A3(new_n577), .ZN(new_n770));
  AND2_X1   g584(.A1(new_n763), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n762), .A2(new_n723), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT111), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n721), .A2(new_n771), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(KEYINPUT112), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT112), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n721), .A2(new_n771), .A3(new_n777), .A4(new_n774), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n652), .A2(new_n687), .A3(new_n635), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT52), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n624), .A2(new_n630), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n647), .A2(new_n638), .A3(new_n782), .A4(new_n589), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n783), .A2(new_n694), .ZN(new_n784));
  INV_X1    g598(.A(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n780), .A2(new_n781), .A3(new_n785), .ZN(new_n786));
  OAI21_X1  g600(.A(KEYINPUT52), .B1(new_n779), .B2(new_n784), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  AND4_X1   g603(.A1(KEYINPUT53), .A2(new_n776), .A3(new_n778), .A4(new_n789), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n788), .B1(new_n775), .B2(KEYINPUT112), .ZN(new_n791));
  AOI21_X1  g605(.A(KEYINPUT53), .B1(new_n791), .B2(new_n778), .ZN(new_n792));
  OAI21_X1  g606(.A(KEYINPUT54), .B1(new_n790), .B2(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n776), .A2(new_n778), .A3(new_n789), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT53), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT54), .ZN(new_n797));
  AND3_X1   g611(.A1(new_n786), .A2(new_n787), .A3(KEYINPUT53), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n721), .A2(new_n771), .A3(new_n798), .A4(new_n774), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(KEYINPUT113), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n796), .A2(new_n797), .A3(new_n800), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n757), .B1(new_n793), .B2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT113), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n799), .B(new_n803), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n792), .A2(new_n804), .ZN(new_n805));
  AOI21_X1  g619(.A(KEYINPUT114), .B1(new_n805), .B2(new_n797), .ZN(new_n806));
  INV_X1    g620(.A(new_n670), .ZN(new_n807));
  NOR3_X1   g621(.A1(new_n807), .A2(new_n702), .A3(new_n535), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n731), .A2(new_n808), .A3(new_n686), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n754), .ZN(new_n810));
  INV_X1    g624(.A(new_n607), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n725), .A2(new_n811), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n809), .B1(new_n810), .B2(new_n812), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n731), .A2(new_n536), .A3(new_n682), .ZN(new_n814));
  INV_X1    g628(.A(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(new_n706), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(KEYINPUT115), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n749), .B1(new_n363), .B2(new_n662), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n813), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT118), .ZN(new_n820));
  AOI21_X1  g634(.A(KEYINPUT51), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NOR3_X1   g635(.A1(new_n648), .A2(new_n807), .A3(new_n359), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n822), .B(KEYINPUT116), .ZN(new_n823));
  OAI211_X1 g637(.A(new_n823), .B(new_n815), .C1(KEYINPUT117), .C2(KEYINPUT50), .ZN(new_n824));
  NAND2_X1  g638(.A1(KEYINPUT117), .A2(KEYINPUT50), .ZN(new_n825));
  XNOR2_X1  g639(.A(new_n824), .B(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n819), .A2(new_n826), .ZN(new_n827));
  OR2_X1    g641(.A1(new_n821), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n821), .A2(new_n827), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n731), .A2(new_n808), .A3(new_n716), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT48), .ZN(new_n831));
  OAI22_X1  g645(.A1(new_n830), .A2(new_n831), .B1(new_n608), .B2(new_n810), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n815), .A2(new_n663), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n833), .A2(G952), .A3(new_n245), .ZN(new_n834));
  AOI211_X1 g648(.A(new_n832), .B(new_n834), .C1(new_n831), .C2(new_n830), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n828), .A2(new_n829), .A3(new_n835), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n802), .A2(new_n806), .A3(new_n836), .ZN(new_n837));
  NOR2_X1   g651(.A1(G952), .A2(G953), .ZN(new_n838));
  XNOR2_X1  g652(.A(new_n838), .B(KEYINPUT119), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n756), .B1(new_n837), .B2(new_n839), .ZN(G75));
  NOR2_X1   g654(.A1(new_n245), .A2(G952), .ZN(new_n841));
  INV_X1    g655(.A(new_n841), .ZN(new_n842));
  OAI211_X1 g656(.A(new_n188), .B(new_n424), .C1(new_n792), .C2(new_n804), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT56), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n402), .A2(new_n403), .ZN(new_n845));
  XNOR2_X1  g659(.A(new_n845), .B(new_n371), .ZN(new_n846));
  XNOR2_X1  g660(.A(new_n846), .B(KEYINPUT55), .ZN(new_n847));
  AOI22_X1  g661(.A1(new_n843), .A2(new_n844), .B1(KEYINPUT120), .B2(new_n847), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n847), .A2(KEYINPUT120), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n842), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  AOI211_X1 g664(.A(KEYINPUT120), .B(new_n847), .C1(new_n843), .C2(new_n844), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n850), .A2(new_n851), .ZN(G51));
  XOR2_X1   g666(.A(new_n354), .B(KEYINPUT57), .Z(new_n853));
  NOR3_X1   g667(.A1(new_n792), .A2(new_n804), .A3(KEYINPUT54), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n797), .B1(new_n796), .B2(new_n800), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n853), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  XNOR2_X1  g670(.A(new_n344), .B(KEYINPUT121), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  OR3_X1    g672(.A1(new_n805), .A2(new_n189), .A3(new_n739), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n841), .B1(new_n858), .B2(new_n859), .ZN(G54));
  NAND2_X1  g674(.A1(new_n796), .A2(new_n800), .ZN(new_n861));
  AND2_X1   g675(.A1(KEYINPUT58), .A2(G475), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n861), .A2(new_n188), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n863), .A2(new_n523), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n864), .A2(new_n842), .ZN(new_n865));
  OR3_X1    g679(.A1(new_n863), .A2(KEYINPUT122), .A3(new_n523), .ZN(new_n866));
  OAI21_X1  g680(.A(KEYINPUT122), .B1(new_n863), .B2(new_n523), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n865), .B1(new_n866), .B2(new_n867), .ZN(G60));
  INV_X1    g682(.A(new_n602), .ZN(new_n869));
  NAND2_X1  g683(.A1(G478), .A2(G902), .ZN(new_n870));
  XOR2_X1   g684(.A(new_n870), .B(KEYINPUT59), .Z(new_n871));
  NOR2_X1   g685(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n872), .B1(new_n854), .B2(new_n855), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n873), .A2(new_n842), .ZN(new_n874));
  INV_X1    g688(.A(new_n871), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n875), .B1(new_n802), .B2(new_n806), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n874), .B1(new_n876), .B2(new_n869), .ZN(G63));
  INV_X1    g691(.A(new_n236), .ZN(new_n878));
  XNOR2_X1  g692(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n187), .A2(new_n361), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n879), .B(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(new_n881), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n878), .B1(new_n805), .B2(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n861), .A2(new_n621), .A3(new_n881), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n883), .A2(new_n842), .A3(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT61), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n883), .A2(new_n884), .A3(KEYINPUT61), .A4(new_n842), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n887), .A2(new_n888), .ZN(G66));
  AOI21_X1  g703(.A(new_n245), .B1(new_n539), .B2(G224), .ZN(new_n890));
  INV_X1    g704(.A(new_n770), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n890), .B1(new_n891), .B2(new_n245), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n845), .B1(G898), .B2(new_n245), .ZN(new_n893));
  XOR2_X1   g707(.A(new_n892), .B(new_n893), .Z(G69));
  NAND2_X1  g708(.A1(new_n649), .A2(new_n780), .ZN(new_n895));
  XOR2_X1   g709(.A(new_n895), .B(KEYINPUT62), .Z(new_n896));
  INV_X1    g710(.A(new_n766), .ZN(new_n897));
  OR4_X1    g711(.A1(new_n689), .A2(new_n897), .A3(new_n642), .A4(new_n702), .ZN(new_n898));
  AND3_X1   g712(.A1(new_n746), .A2(new_n751), .A3(new_n898), .ZN(new_n899));
  AOI21_X1  g713(.A(G953), .B1(new_n896), .B2(new_n899), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n440), .B1(new_n439), .B2(new_n444), .ZN(new_n901));
  XOR2_X1   g715(.A(new_n901), .B(KEYINPUT124), .Z(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(new_n518), .ZN(new_n903));
  OR3_X1    g717(.A1(new_n900), .A2(KEYINPUT125), .A3(new_n903), .ZN(new_n904));
  NOR3_X1   g718(.A1(new_n689), .A2(new_n633), .A3(new_n637), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n745), .B1(new_n735), .B2(new_n905), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n906), .A2(new_n751), .A3(new_n723), .A4(new_n780), .ZN(new_n907));
  INV_X1    g721(.A(new_n721), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(new_n245), .ZN(new_n910));
  NAND2_X1  g724(.A1(G900), .A2(G953), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n910), .A2(new_n903), .A3(new_n911), .ZN(new_n912));
  OAI21_X1  g726(.A(KEYINPUT125), .B1(new_n900), .B2(new_n903), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n904), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n245), .B1(G227), .B2(G900), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n914), .B(new_n915), .ZN(G72));
  NAND2_X1  g730(.A1(G472), .A2(G902), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n917), .B(KEYINPUT63), .Z(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n919), .B1(new_n909), .B2(new_n770), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n644), .A2(new_n470), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(KEYINPUT126), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n896), .A2(new_n899), .A3(new_n770), .ZN(new_n923));
  AND2_X1   g737(.A1(new_n923), .A2(new_n918), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n469), .A2(new_n453), .ZN(new_n925));
  OAI221_X1 g739(.A(new_n842), .B1(new_n920), .B2(new_n922), .C1(new_n924), .C2(new_n925), .ZN(new_n926));
  OR2_X1    g740(.A1(new_n790), .A2(new_n792), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n919), .B1(new_n471), .B2(new_n454), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n926), .B1(new_n927), .B2(new_n928), .ZN(G57));
endmodule


