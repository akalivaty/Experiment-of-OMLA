//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 0 1 1 0 0 1 0 1 0 1 0 0 1 0 1 0 0 0 0 0 0 0 1 1 0 0 1 1 1 1 1 0 0 1 1 1 1 0 0 1 1 1 1 1 0 1 0 0 0 0 0 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n717,
    new_n718, new_n719, new_n720, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n728, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n762, new_n763, new_n764, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n803,
    new_n804, new_n805, new_n806, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n860, new_n861, new_n863,
    new_n864, new_n865, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n967, new_n968, new_n969, new_n970, new_n971, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n981,
    new_n982;
  XOR2_X1   g000(.A(G8gat), .B(G36gat), .Z(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT71), .ZN(new_n203));
  XNOR2_X1  g002(.A(G64gat), .B(G92gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n205), .B(KEYINPUT72), .ZN(new_n206));
  INV_X1    g005(.A(G226gat), .ZN(new_n207));
  INV_X1    g006(.A(G233gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT24), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n211), .A2(G183gat), .A3(G190gat), .ZN(new_n212));
  XNOR2_X1  g011(.A(G183gat), .B(G190gat), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n212), .B1(new_n213), .B2(new_n211), .ZN(new_n214));
  NAND2_X1  g013(.A1(G169gat), .A2(G176gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(KEYINPUT23), .ZN(new_n216));
  INV_X1    g015(.A(G169gat), .ZN(new_n217));
  INV_X1    g016(.A(G176gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n216), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT25), .ZN(new_n221));
  NOR2_X1   g020(.A1(G169gat), .A2(G176gat), .ZN(new_n222));
  AOI21_X1  g021(.A(new_n221), .B1(new_n222), .B2(KEYINPUT23), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n220), .A2(new_n223), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n214), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT65), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n218), .A2(KEYINPUT23), .ZN(new_n227));
  AND2_X1   g026(.A1(KEYINPUT64), .A2(G169gat), .ZN(new_n228));
  NOR2_X1   g027(.A1(KEYINPUT64), .A2(G169gat), .ZN(new_n229));
  NOR3_X1   g028(.A1(new_n227), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n222), .B1(KEYINPUT23), .B2(new_n215), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n226), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT23), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n233), .A2(G176gat), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT64), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(new_n217), .ZN(new_n236));
  NAND2_X1  g035(.A1(KEYINPUT64), .A2(G169gat), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n234), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n238), .A2(new_n220), .A3(KEYINPUT65), .ZN(new_n239));
  INV_X1    g038(.A(new_n212), .ZN(new_n240));
  XOR2_X1   g039(.A(G183gat), .B(G190gat), .Z(new_n241));
  AOI21_X1  g040(.A(new_n240), .B1(new_n241), .B2(KEYINPUT24), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n232), .A2(new_n239), .A3(new_n242), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n225), .B1(new_n243), .B2(new_n221), .ZN(new_n244));
  AOI21_X1  g043(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT66), .ZN(new_n246));
  OR3_X1    g045(.A1(new_n245), .A2(new_n222), .A3(new_n246), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n246), .B1(new_n245), .B2(new_n222), .ZN(new_n248));
  OAI211_X1 g047(.A(new_n247), .B(new_n248), .C1(KEYINPUT26), .C2(new_n219), .ZN(new_n249));
  XNOR2_X1  g048(.A(KEYINPUT27), .B(G183gat), .ZN(new_n250));
  INV_X1    g049(.A(G190gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  OR2_X1    g051(.A1(new_n252), .A2(KEYINPUT28), .ZN(new_n253));
  AOI22_X1  g052(.A1(new_n252), .A2(KEYINPUT28), .B1(G183gat), .B2(G190gat), .ZN(new_n254));
  AND3_X1   g053(.A1(new_n249), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n244), .A2(new_n255), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n210), .B1(new_n256), .B2(KEYINPUT29), .ZN(new_n257));
  XNOR2_X1  g056(.A(G197gat), .B(G204gat), .ZN(new_n258));
  INV_X1    g057(.A(G211gat), .ZN(new_n259));
  INV_X1    g058(.A(G218gat), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n258), .B1(KEYINPUT22), .B2(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(G211gat), .B(G218gat), .ZN(new_n263));
  XNOR2_X1  g062(.A(new_n262), .B(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(new_n225), .ZN(new_n266));
  AND3_X1   g065(.A1(new_n238), .A2(KEYINPUT65), .A3(new_n220), .ZN(new_n267));
  AOI21_X1  g066(.A(KEYINPUT65), .B1(new_n238), .B2(new_n220), .ZN(new_n268));
  NOR3_X1   g067(.A1(new_n267), .A2(new_n268), .A3(new_n214), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n266), .B1(new_n269), .B2(KEYINPUT25), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n249), .A2(new_n253), .A3(new_n254), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(new_n209), .ZN(new_n273));
  AND3_X1   g072(.A1(new_n257), .A2(new_n265), .A3(new_n273), .ZN(new_n274));
  XOR2_X1   g073(.A(KEYINPUT70), .B(KEYINPUT29), .Z(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n210), .B1(new_n256), .B2(new_n276), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n265), .B1(new_n277), .B2(new_n273), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n206), .B1(new_n274), .B2(new_n278), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n209), .B1(new_n272), .B2(new_n275), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n256), .A2(new_n210), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n264), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n257), .A2(new_n265), .A3(new_n273), .ZN(new_n283));
  NAND4_X1  g082(.A1(new_n282), .A2(new_n283), .A3(KEYINPUT30), .A4(new_n205), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n279), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT30), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n282), .A2(new_n283), .A3(new_n205), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n285), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(G228gat), .A2(G233gat), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT3), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n291), .B1(new_n264), .B2(new_n276), .ZN(new_n292));
  INV_X1    g091(.A(G141gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(G148gat), .ZN(new_n294));
  INV_X1    g093(.A(G148gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(G141gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT74), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(G141gat), .B(G148gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(KEYINPUT74), .ZN(new_n301));
  NAND2_X1  g100(.A1(G155gat), .A2(G162gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(KEYINPUT2), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n299), .A2(new_n301), .A3(new_n303), .ZN(new_n304));
  OR2_X1    g103(.A1(G155gat), .A2(G162gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(new_n302), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT75), .ZN(new_n308));
  AND3_X1   g107(.A1(new_n294), .A2(new_n296), .A3(new_n308), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n295), .A2(KEYINPUT75), .A3(G141gat), .ZN(new_n310));
  INV_X1    g109(.A(new_n302), .ZN(new_n311));
  NOR2_X1   g110(.A1(G155gat), .A2(G162gat), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n310), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n309), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT76), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n303), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n302), .A2(KEYINPUT76), .A3(KEYINPUT2), .ZN(new_n317));
  AND2_X1   g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  AOI22_X1  g117(.A1(new_n304), .A2(new_n307), .B1(new_n314), .B2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  AND2_X1   g119(.A1(new_n292), .A2(new_n320), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n303), .B1(new_n300), .B2(KEYINPUT74), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n297), .A2(new_n298), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n307), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n313), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n294), .A2(new_n296), .A3(new_n308), .ZN(new_n326));
  NAND4_X1  g125(.A1(new_n325), .A2(new_n326), .A3(new_n316), .A4(new_n317), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n324), .A2(new_n291), .A3(new_n327), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n265), .B1(new_n328), .B2(new_n275), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n290), .B1(new_n321), .B2(new_n329), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n291), .B1(new_n264), .B2(KEYINPUT29), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(new_n320), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n332), .A2(G228gat), .A3(G233gat), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n330), .B1(new_n329), .B2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT80), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(G22gat), .ZN(new_n336));
  XNOR2_X1  g135(.A(G78gat), .B(G106gat), .ZN(new_n337));
  XNOR2_X1  g136(.A(KEYINPUT31), .B(G50gat), .ZN(new_n338));
  XNOR2_X1  g137(.A(new_n337), .B(new_n338), .ZN(new_n339));
  MUX2_X1   g138(.A(G22gat), .B(new_n336), .S(new_n339), .Z(new_n340));
  XOR2_X1   g139(.A(new_n334), .B(new_n340), .Z(new_n341));
  NOR3_X1   g140(.A1(new_n289), .A2(KEYINPUT35), .A3(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT67), .ZN(new_n343));
  INV_X1    g142(.A(G120gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(G113gat), .ZN(new_n345));
  INV_X1    g144(.A(G113gat), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(G120gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  XNOR2_X1  g147(.A(G127gat), .B(G134gat), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT1), .ZN(new_n350));
  AND3_X1   g149(.A1(new_n348), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n349), .B1(new_n350), .B2(new_n348), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  NAND4_X1  g153(.A1(new_n270), .A2(new_n343), .A3(new_n354), .A4(new_n271), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n343), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n353), .A2(KEYINPUT67), .ZN(new_n357));
  OAI211_X1 g156(.A(new_n356), .B(new_n357), .C1(new_n244), .C2(new_n255), .ZN(new_n358));
  NAND2_X1  g157(.A1(G227gat), .A2(G233gat), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n355), .A2(new_n358), .A3(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(KEYINPUT32), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT33), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  XOR2_X1   g163(.A(G15gat), .B(G43gat), .Z(new_n365));
  XNOR2_X1  g164(.A(G71gat), .B(G99gat), .ZN(new_n366));
  XNOR2_X1  g165(.A(new_n365), .B(new_n366), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n362), .A2(new_n364), .A3(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n367), .ZN(new_n369));
  OAI211_X1 g168(.A(new_n361), .B(KEYINPUT32), .C1(new_n363), .C2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n358), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(new_n359), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT69), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n373), .A2(new_n374), .A3(KEYINPUT34), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT34), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n360), .B1(new_n355), .B2(new_n358), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n376), .B1(new_n377), .B2(KEYINPUT69), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n375), .A2(new_n378), .ZN(new_n379));
  OR2_X1    g178(.A1(new_n371), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n371), .A2(new_n379), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT5), .ZN(new_n384));
  XNOR2_X1  g183(.A(G113gat), .B(G120gat), .ZN(new_n385));
  INV_X1    g184(.A(G127gat), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n386), .A2(G134gat), .ZN(new_n387));
  INV_X1    g186(.A(G134gat), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n388), .A2(G127gat), .ZN(new_n389));
  OAI22_X1  g188(.A1(new_n385), .A2(KEYINPUT1), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n348), .A2(new_n349), .A3(new_n350), .ZN(new_n391));
  AND3_X1   g190(.A1(new_n390), .A2(new_n391), .A3(KEYINPUT77), .ZN(new_n392));
  AOI21_X1  g191(.A(KEYINPUT77), .B1(new_n390), .B2(new_n391), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT2), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n394), .B1(G155gat), .B2(G162gat), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n395), .B1(new_n297), .B2(new_n298), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n306), .B1(new_n396), .B2(new_n301), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n326), .A2(new_n306), .A3(new_n310), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n316), .A2(new_n317), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  OAI22_X1  g199(.A1(new_n392), .A2(new_n393), .B1(new_n397), .B2(new_n400), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n353), .A2(new_n324), .A3(new_n327), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(G225gat), .A2(G233gat), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n384), .B1(new_n403), .B2(new_n405), .ZN(new_n406));
  OAI21_X1  g205(.A(KEYINPUT3), .B1(new_n397), .B2(new_n400), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT77), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n408), .B1(new_n351), .B2(new_n352), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n390), .A2(new_n391), .A3(KEYINPUT77), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n407), .A2(new_n411), .A3(new_n328), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT4), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n402), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n319), .A2(KEYINPUT4), .A3(new_n353), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n412), .A2(new_n404), .A3(new_n414), .A4(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n406), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(KEYINPUT4), .B1(new_n319), .B2(new_n353), .ZN(new_n418));
  AND4_X1   g217(.A1(KEYINPUT4), .A2(new_n353), .A3(new_n324), .A4(new_n327), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n420), .A2(new_n384), .A3(new_n404), .A4(new_n412), .ZN(new_n421));
  XNOR2_X1  g220(.A(G1gat), .B(G29gat), .ZN(new_n422));
  XNOR2_X1  g221(.A(new_n422), .B(KEYINPUT0), .ZN(new_n423));
  XOR2_X1   g222(.A(G57gat), .B(G85gat), .Z(new_n424));
  XNOR2_X1  g223(.A(new_n423), .B(new_n424), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n417), .A2(new_n421), .A3(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT78), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT6), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n417), .A2(new_n421), .A3(KEYINPUT78), .A4(new_n425), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n428), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  AND2_X1   g230(.A1(new_n417), .A2(new_n421), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n432), .A2(new_n425), .ZN(new_n433));
  OR2_X1    g232(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(KEYINPUT6), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n342), .A2(new_n383), .A3(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT79), .ZN(new_n438));
  AND2_X1   g237(.A1(new_n426), .A2(new_n427), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n430), .A2(new_n429), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n438), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(new_n433), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n428), .A2(KEYINPUT79), .A3(new_n429), .A4(new_n430), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n441), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(new_n435), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT73), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n285), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n279), .A2(new_n284), .A3(KEYINPUT73), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n287), .A2(new_n286), .ZN(new_n449));
  AND3_X1   g248(.A1(new_n447), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT68), .ZN(new_n451));
  AOI21_X1  g250(.A(KEYINPUT34), .B1(new_n373), .B2(new_n374), .ZN(new_n452));
  NOR3_X1   g251(.A1(new_n377), .A2(KEYINPUT69), .A3(new_n376), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n451), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(new_n371), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n379), .A2(new_n451), .A3(new_n368), .A4(new_n370), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n341), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n445), .A2(new_n450), .A3(new_n457), .ZN(new_n458));
  AND3_X1   g257(.A1(new_n458), .A2(KEYINPUT86), .A3(KEYINPUT35), .ZN(new_n459));
  AOI21_X1  g258(.A(KEYINPUT86), .B1(new_n458), .B2(KEYINPUT35), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n437), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  XNOR2_X1  g260(.A(new_n334), .B(new_n340), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n462), .B1(new_n445), .B2(new_n450), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT36), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n380), .A2(new_n464), .A3(new_n381), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n455), .A2(KEYINPUT36), .A3(new_n456), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  OAI21_X1  g266(.A(KEYINPUT81), .B1(new_n463), .B2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n467), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT81), .ZN(new_n470));
  INV_X1    g269(.A(new_n435), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n433), .B1(new_n431), .B2(new_n438), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n471), .B1(new_n472), .B2(new_n443), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n447), .A2(new_n448), .A3(new_n449), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n469), .B(new_n470), .C1(new_n475), .C2(new_n462), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n401), .A2(new_n404), .A3(new_n402), .ZN(new_n477));
  XNOR2_X1  g276(.A(new_n477), .B(KEYINPUT83), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n412), .A2(new_n414), .A3(new_n415), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(new_n405), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n478), .A2(KEYINPUT39), .A3(new_n480), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n425), .B1(new_n480), .B2(KEYINPUT39), .ZN(new_n482));
  AND2_X1   g281(.A1(new_n482), .A2(KEYINPUT82), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n482), .A2(KEYINPUT82), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n481), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT40), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n433), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  OAI211_X1 g286(.A(KEYINPUT40), .B(new_n481), .C1(new_n483), .C2(new_n484), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT84), .ZN(new_n489));
  AND2_X1   g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n488), .A2(new_n489), .ZN(new_n491));
  OAI211_X1 g290(.A(new_n289), .B(new_n487), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT38), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT37), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n282), .A2(new_n283), .A3(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT85), .ZN(new_n496));
  XNOR2_X1  g295(.A(new_n495), .B(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n282), .A2(new_n283), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n205), .B1(new_n498), .B2(KEYINPUT37), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n493), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n206), .A2(new_n493), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n277), .A2(new_n273), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n494), .B1(new_n502), .B2(new_n265), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n257), .A2(new_n264), .A3(new_n273), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n501), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n497), .A2(new_n505), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n506), .A2(new_n435), .A3(new_n287), .A4(new_n434), .ZN(new_n507));
  OAI211_X1 g306(.A(new_n492), .B(new_n462), .C1(new_n500), .C2(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n468), .A2(new_n476), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n461), .A2(new_n509), .ZN(new_n510));
  XNOR2_X1  g309(.A(G15gat), .B(G22gat), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT16), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n511), .B1(new_n512), .B2(G1gat), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n513), .B1(G1gat), .B2(new_n511), .ZN(new_n514));
  INV_X1    g313(.A(G8gat), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n514), .B(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(new_n516), .ZN(new_n517));
  XNOR2_X1  g316(.A(G43gat), .B(G50gat), .ZN(new_n518));
  INV_X1    g317(.A(G29gat), .ZN(new_n519));
  INV_X1    g318(.A(G36gat), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n519), .A2(new_n520), .A3(KEYINPUT14), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT14), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n522), .B1(G29gat), .B2(G36gat), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT87), .ZN(new_n525));
  OAI22_X1  g324(.A1(new_n524), .A2(new_n525), .B1(new_n519), .B2(new_n520), .ZN(new_n526));
  AOI21_X1  g325(.A(KEYINPUT87), .B1(new_n521), .B2(new_n523), .ZN(new_n527));
  OAI211_X1 g326(.A(KEYINPUT15), .B(new_n518), .C1(new_n526), .C2(new_n527), .ZN(new_n528));
  AOI22_X1  g327(.A1(new_n518), .A2(KEYINPUT15), .B1(G29gat), .B2(G36gat), .ZN(new_n529));
  INV_X1    g328(.A(new_n524), .ZN(new_n530));
  OAI211_X1 g329(.A(new_n529), .B(new_n530), .C1(KEYINPUT15), .C2(new_n518), .ZN(new_n531));
  AND2_X1   g330(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT88), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT17), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n528), .A2(new_n531), .ZN(new_n536));
  NAND2_X1  g335(.A1(KEYINPUT88), .A2(KEYINPUT17), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n533), .A2(new_n534), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n517), .B1(new_n535), .B2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT89), .ZN(new_n541));
  AOI22_X1  g340(.A1(new_n540), .A2(new_n541), .B1(new_n517), .B2(new_n536), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n535), .A2(new_n539), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(new_n516), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n544), .A2(KEYINPUT89), .ZN(new_n545));
  NAND2_X1  g344(.A1(G229gat), .A2(G233gat), .ZN(new_n546));
  NAND4_X1  g345(.A1(new_n542), .A2(new_n545), .A3(KEYINPUT18), .A4(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT92), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n532), .B(new_n516), .ZN(new_n550));
  XOR2_X1   g349(.A(new_n546), .B(KEYINPUT13), .Z(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  AND2_X1   g351(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  AND2_X1   g352(.A1(new_n542), .A2(new_n545), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT90), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n554), .A2(new_n555), .A3(new_n546), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n542), .A2(new_n545), .A3(new_n546), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(KEYINPUT90), .ZN(new_n558));
  XOR2_X1   g357(.A(KEYINPUT91), .B(KEYINPUT18), .Z(new_n559));
  NAND3_X1  g358(.A1(new_n556), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  OR2_X1    g359(.A1(new_n547), .A2(new_n548), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n553), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(G113gat), .B(G141gat), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n563), .B(G197gat), .ZN(new_n564));
  XOR2_X1   g363(.A(KEYINPUT11), .B(G169gat), .Z(new_n565));
  XNOR2_X1  g364(.A(new_n564), .B(new_n565), .ZN(new_n566));
  XOR2_X1   g365(.A(new_n566), .B(KEYINPUT12), .Z(new_n567));
  NAND2_X1  g366(.A1(new_n562), .A2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n567), .ZN(new_n569));
  NAND4_X1  g368(.A1(new_n553), .A2(new_n560), .A3(new_n569), .A4(new_n561), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(G230gat), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n572), .A2(new_n208), .ZN(new_n573));
  XOR2_X1   g372(.A(G57gat), .B(G64gat), .Z(new_n574));
  INV_X1    g373(.A(KEYINPUT9), .ZN(new_n575));
  INV_X1    g374(.A(G71gat), .ZN(new_n576));
  INV_X1    g375(.A(G78gat), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n575), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n574), .A2(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(G71gat), .B(G78gat), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n574), .A2(new_n580), .A3(new_n578), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT99), .ZN(new_n585));
  XNOR2_X1  g384(.A(G99gat), .B(G106gat), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n584), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  XOR2_X1   g386(.A(KEYINPUT96), .B(G92gat), .Z(new_n588));
  INV_X1    g387(.A(G85gat), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(G85gat), .A2(G92gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n591), .B(KEYINPUT7), .ZN(new_n592));
  INV_X1    g391(.A(G99gat), .ZN(new_n593));
  INV_X1    g392(.A(G106gat), .ZN(new_n594));
  OAI21_X1  g393(.A(KEYINPUT8), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND4_X1  g394(.A1(new_n590), .A2(new_n586), .A3(new_n592), .A4(new_n595), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n590), .A2(new_n592), .A3(new_n595), .ZN(new_n597));
  INV_X1    g396(.A(new_n586), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n597), .A2(KEYINPUT99), .A3(new_n598), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n587), .A2(new_n596), .A3(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT100), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND4_X1  g401(.A1(new_n587), .A2(KEYINPUT100), .A3(new_n596), .A4(new_n599), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT10), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n597), .A2(new_n598), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n606), .A2(new_n596), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n607), .A2(new_n584), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n604), .A2(new_n605), .A3(new_n608), .ZN(new_n609));
  NOR3_X1   g408(.A1(new_n607), .A2(new_n605), .A3(new_n584), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(KEYINPUT101), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n573), .B1(new_n609), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n604), .A2(new_n608), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n612), .B1(new_n573), .B2(new_n613), .ZN(new_n614));
  XOR2_X1   g413(.A(G120gat), .B(G148gat), .Z(new_n615));
  XNOR2_X1  g414(.A(G176gat), .B(G204gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n615), .B(new_n616), .ZN(new_n617));
  OR2_X1    g416(.A1(new_n614), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n614), .A2(new_n617), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  XOR2_X1   g420(.A(G134gat), .B(G162gat), .Z(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT95), .ZN(new_n624));
  NAND3_X1  g423(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n625), .B1(new_n532), .B2(new_n607), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT97), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  OAI211_X1 g427(.A(KEYINPUT97), .B(new_n625), .C1(new_n532), .C2(new_n607), .ZN(new_n629));
  AOI22_X1  g428(.A1(new_n628), .A2(new_n629), .B1(new_n543), .B2(new_n607), .ZN(new_n630));
  XNOR2_X1  g429(.A(G190gat), .B(G218gat), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT98), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n624), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  AND2_X1   g434(.A1(new_n628), .A2(new_n629), .ZN(new_n636));
  AND2_X1   g435(.A1(new_n543), .A2(new_n607), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n631), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n630), .A2(new_n632), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n638), .A2(new_n639), .A3(KEYINPUT98), .ZN(new_n640));
  AOI21_X1  g439(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n635), .A2(new_n640), .A3(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n642), .B1(new_n635), .B2(new_n640), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n623), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n635), .A2(new_n640), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n647), .A2(new_n641), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n648), .A2(new_n622), .A3(new_n643), .ZN(new_n649));
  XNOR2_X1  g448(.A(KEYINPUT93), .B(KEYINPUT21), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n584), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(G127gat), .B(G155gat), .ZN(new_n652));
  XOR2_X1   g451(.A(new_n651), .B(new_n652), .Z(new_n653));
  INV_X1    g452(.A(KEYINPUT21), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n516), .B1(new_n654), .B2(new_n584), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n653), .B(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(G231gat), .A2(G233gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(KEYINPUT94), .ZN(new_n658));
  XOR2_X1   g457(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n659));
  XNOR2_X1  g458(.A(new_n658), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g459(.A(G183gat), .B(G211gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n656), .B(new_n662), .ZN(new_n663));
  AND3_X1   g462(.A1(new_n646), .A2(new_n649), .A3(new_n663), .ZN(new_n664));
  AND4_X1   g463(.A1(new_n510), .A2(new_n571), .A3(new_n621), .A4(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n665), .A2(new_n473), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g466(.A1(new_n665), .A2(new_n289), .ZN(new_n668));
  XOR2_X1   g467(.A(KEYINPUT16), .B(G8gat), .Z(new_n669));
  AND2_X1   g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n668), .A2(new_n515), .ZN(new_n671));
  OAI21_X1  g470(.A(KEYINPUT42), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n672), .B1(KEYINPUT42), .B2(new_n670), .ZN(G1325gat));
  INV_X1    g472(.A(G15gat), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n665), .A2(new_n674), .A3(new_n383), .ZN(new_n675));
  AND2_X1   g474(.A1(new_n665), .A2(new_n467), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n675), .B1(new_n676), .B2(new_n674), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(KEYINPUT102), .ZN(G1326gat));
  NAND2_X1  g477(.A1(new_n665), .A2(new_n341), .ZN(new_n679));
  XNOR2_X1  g478(.A(KEYINPUT43), .B(G22gat), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(G1327gat));
  NAND2_X1  g480(.A1(new_n646), .A2(new_n649), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n510), .A2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  AND2_X1   g483(.A1(new_n568), .A2(new_n570), .ZN(new_n685));
  NOR3_X1   g484(.A1(new_n685), .A2(new_n620), .A3(new_n663), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  NOR3_X1   g486(.A1(new_n687), .A2(G29gat), .A3(new_n445), .ZN(new_n688));
  XOR2_X1   g487(.A(new_n688), .B(KEYINPUT45), .Z(new_n689));
  INV_X1    g488(.A(new_n682), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n690), .A2(KEYINPUT44), .ZN(new_n691));
  OAI211_X1 g490(.A(KEYINPUT104), .B(new_n437), .C1(new_n459), .C2(new_n460), .ZN(new_n692));
  OAI211_X1 g491(.A(new_n508), .B(new_n469), .C1(new_n462), .C2(new_n475), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT86), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n454), .A2(new_n371), .ZN(new_n696));
  AOI22_X1  g495(.A1(new_n379), .A2(new_n451), .B1(new_n368), .B2(new_n370), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n462), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  NOR3_X1   g497(.A1(new_n473), .A2(new_n698), .A3(new_n474), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT35), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n695), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n458), .A2(KEYINPUT86), .A3(KEYINPUT35), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  AOI21_X1  g502(.A(KEYINPUT104), .B1(new_n703), .B2(new_n437), .ZN(new_n704));
  OAI211_X1 g503(.A(KEYINPUT105), .B(new_n691), .C1(new_n694), .C2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n683), .A2(KEYINPUT44), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT104), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n461), .A2(new_n708), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n709), .A2(new_n692), .A3(new_n693), .ZN(new_n710));
  AOI21_X1  g509(.A(KEYINPUT105), .B1(new_n710), .B2(new_n691), .ZN(new_n711));
  OR2_X1    g510(.A1(new_n707), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n686), .B(KEYINPUT103), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n712), .A2(new_n473), .A3(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n689), .B1(new_n715), .B2(new_n519), .ZN(G1328gat));
  NOR3_X1   g515(.A1(new_n687), .A2(G36gat), .A3(new_n288), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(KEYINPUT46), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n712), .A2(new_n289), .A3(new_n713), .ZN(new_n719));
  INV_X1    g518(.A(new_n719), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n718), .B1(new_n720), .B2(new_n520), .ZN(G1329gat));
  NOR3_X1   g520(.A1(new_n687), .A2(G43gat), .A3(new_n382), .ZN(new_n722));
  OAI211_X1 g521(.A(new_n467), .B(new_n713), .C1(new_n707), .C2(new_n711), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n722), .B1(new_n723), .B2(G43gat), .ZN(new_n724));
  XOR2_X1   g523(.A(KEYINPUT106), .B(KEYINPUT47), .Z(new_n725));
  XNOR2_X1  g524(.A(new_n724), .B(new_n725), .ZN(G1330gat));
  NOR3_X1   g525(.A1(new_n687), .A2(G50gat), .A3(new_n462), .ZN(new_n727));
  OAI211_X1 g526(.A(new_n341), .B(new_n713), .C1(new_n707), .C2(new_n711), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n727), .B1(new_n728), .B2(G50gat), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(KEYINPUT48), .ZN(G1331gat));
  NAND3_X1  g529(.A1(new_n685), .A2(new_n664), .A3(new_n620), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(KEYINPUT107), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT107), .ZN(new_n733));
  NAND4_X1  g532(.A1(new_n685), .A2(new_n664), .A3(new_n733), .A4(new_n620), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n735), .B1(new_n694), .B2(new_n704), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(KEYINPUT108), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT108), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n710), .A2(new_n738), .A3(new_n735), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n737), .A2(new_n473), .A3(new_n739), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(G57gat), .ZN(G1332gat));
  AND3_X1   g540(.A1(new_n737), .A2(KEYINPUT109), .A3(new_n739), .ZN(new_n742));
  AOI21_X1  g541(.A(KEYINPUT109), .B1(new_n737), .B2(new_n739), .ZN(new_n743));
  OR2_X1    g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT49), .ZN(new_n745));
  INV_X1    g544(.A(G64gat), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n288), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(KEYINPUT110), .ZN(new_n749));
  AND3_X1   g548(.A1(new_n744), .A2(new_n747), .A3(new_n749), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n747), .B1(new_n744), .B2(new_n749), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n750), .A2(new_n751), .ZN(G1333gat));
  INV_X1    g551(.A(KEYINPUT50), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n467), .B1(new_n742), .B2(new_n743), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(G71gat), .ZN(new_n755));
  XOR2_X1   g554(.A(new_n382), .B(KEYINPUT111), .Z(new_n756));
  NAND4_X1  g555(.A1(new_n737), .A2(new_n739), .A3(new_n576), .A4(new_n756), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n753), .B1(new_n755), .B2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(new_n757), .ZN(new_n759));
  AOI211_X1 g558(.A(KEYINPUT50), .B(new_n759), .C1(new_n754), .C2(G71gat), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n758), .A2(new_n760), .ZN(G1334gat));
  NAND2_X1  g560(.A1(new_n744), .A2(new_n341), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(G78gat), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n744), .A2(new_n577), .A3(new_n341), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(G1335gat));
  NOR2_X1   g564(.A1(new_n445), .A2(G85gat), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n571), .A2(new_n663), .ZN(new_n767));
  INV_X1    g566(.A(new_n767), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n768), .A2(new_n690), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n769), .B1(new_n694), .B2(new_n704), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(KEYINPUT51), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT51), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n710), .A2(new_n772), .A3(new_n769), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n771), .A2(new_n773), .ZN(new_n774));
  AND2_X1   g573(.A1(new_n774), .A2(KEYINPUT113), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n774), .A2(KEYINPUT113), .ZN(new_n776));
  OAI211_X1 g575(.A(new_n620), .B(new_n766), .C1(new_n775), .C2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT112), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n768), .A2(new_n621), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n712), .A2(new_n779), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n778), .B1(new_n780), .B2(new_n445), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(G85gat), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n780), .A2(new_n778), .A3(new_n445), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n777), .B1(new_n782), .B2(new_n783), .ZN(G1336gat));
  OAI211_X1 g583(.A(new_n289), .B(new_n779), .C1(new_n707), .C2(new_n711), .ZN(new_n785));
  INV_X1    g584(.A(new_n588), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT52), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n621), .A2(G92gat), .A3(new_n288), .ZN(new_n789));
  INV_X1    g588(.A(new_n789), .ZN(new_n790));
  OAI211_X1 g589(.A(new_n787), .B(new_n788), .C1(new_n774), .C2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT115), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n770), .A2(new_n792), .A3(new_n772), .ZN(new_n793));
  OAI211_X1 g592(.A(new_n710), .B(new_n769), .C1(KEYINPUT115), .C2(KEYINPUT51), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  XNOR2_X1  g594(.A(new_n789), .B(KEYINPUT114), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(KEYINPUT116), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT116), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n795), .A2(new_n799), .A3(new_n796), .ZN(new_n800));
  AND3_X1   g599(.A1(new_n798), .A2(new_n787), .A3(new_n800), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n791), .B1(new_n801), .B2(new_n788), .ZN(G1337gat));
  NOR2_X1   g601(.A1(new_n382), .A2(G99gat), .ZN(new_n803));
  OAI211_X1 g602(.A(new_n620), .B(new_n803), .C1(new_n775), .C2(new_n776), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n712), .A2(new_n467), .A3(new_n779), .ZN(new_n805));
  INV_X1    g604(.A(new_n805), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n804), .B1(new_n806), .B2(new_n593), .ZN(G1338gat));
  INV_X1    g606(.A(KEYINPUT118), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT53), .ZN(new_n809));
  OAI211_X1 g608(.A(new_n341), .B(new_n779), .C1(new_n707), .C2(new_n711), .ZN(new_n810));
  XOR2_X1   g609(.A(KEYINPUT117), .B(G106gat), .Z(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NOR3_X1   g611(.A1(new_n621), .A2(G106gat), .A3(new_n462), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n795), .A2(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n809), .B1(new_n812), .B2(new_n814), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n771), .A2(new_n773), .A3(new_n813), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(new_n809), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n817), .B1(new_n810), .B2(new_n811), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n808), .B1(new_n815), .B2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(new_n817), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n812), .A2(new_n820), .ZN(new_n821));
  AOI22_X1  g620(.A1(new_n810), .A2(new_n811), .B1(new_n795), .B2(new_n813), .ZN(new_n822));
  OAI211_X1 g621(.A(new_n821), .B(KEYINPUT118), .C1(new_n809), .C2(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n819), .A2(new_n823), .ZN(G1339gat));
  INV_X1    g623(.A(KEYINPUT54), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n617), .B1(new_n612), .B2(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(new_n608), .ZN(new_n827));
  AOI211_X1 g626(.A(KEYINPUT10), .B(new_n827), .C1(new_n602), .C2(new_n603), .ZN(new_n828));
  XOR2_X1   g627(.A(new_n610), .B(KEYINPUT101), .Z(new_n829));
  OAI22_X1  g628(.A1(new_n828), .A2(new_n829), .B1(new_n572), .B2(new_n208), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n609), .A2(new_n573), .A3(new_n611), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n830), .A2(new_n831), .A3(KEYINPUT54), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n826), .A2(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT55), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n826), .A2(new_n832), .A3(KEYINPUT55), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n835), .A2(new_n619), .A3(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n837), .B1(new_n568), .B2(new_n570), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n554), .A2(new_n546), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n550), .A2(new_n551), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n566), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  AND3_X1   g640(.A1(new_n620), .A2(new_n570), .A3(new_n841), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n690), .B1(new_n838), .B2(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(new_n837), .ZN(new_n844));
  NAND4_X1  g643(.A1(new_n682), .A2(new_n844), .A3(new_n570), .A4(new_n841), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n663), .B1(new_n846), .B2(KEYINPUT119), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT119), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n843), .A2(new_n848), .A3(new_n845), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n685), .A2(new_n664), .A3(new_n621), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n445), .A2(new_n289), .ZN(new_n853));
  NAND4_X1  g652(.A1(new_n852), .A2(new_n462), .A3(new_n383), .A4(new_n853), .ZN(new_n854));
  NOR3_X1   g653(.A1(new_n854), .A2(new_n346), .A3(new_n685), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n852), .A2(new_n473), .A3(new_n457), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n856), .A2(new_n289), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(new_n571), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n855), .B1(new_n858), .B2(new_n346), .ZN(G1340gat));
  NOR3_X1   g658(.A1(new_n854), .A2(new_n344), .A3(new_n621), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n857), .A2(new_n620), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n860), .B1(new_n861), .B2(new_n344), .ZN(G1341gat));
  NAND3_X1  g661(.A1(new_n857), .A2(new_n386), .A3(new_n663), .ZN(new_n863));
  INV_X1    g662(.A(new_n663), .ZN(new_n864));
  OAI21_X1  g663(.A(G127gat), .B1(new_n854), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n863), .A2(new_n865), .ZN(G1342gat));
  NAND2_X1  g665(.A1(new_n682), .A2(new_n288), .ZN(new_n867));
  XOR2_X1   g666(.A(new_n867), .B(KEYINPUT120), .Z(new_n868));
  OR2_X1    g667(.A1(new_n868), .A2(G134gat), .ZN(new_n869));
  OR3_X1    g668(.A1(new_n856), .A2(KEYINPUT56), .A3(new_n869), .ZN(new_n870));
  OAI21_X1  g669(.A(KEYINPUT56), .B1(new_n856), .B2(new_n869), .ZN(new_n871));
  OAI21_X1  g670(.A(G134gat), .B1(new_n854), .B2(new_n690), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n870), .A2(new_n871), .A3(new_n872), .ZN(G1343gat));
  INV_X1    g672(.A(KEYINPUT57), .ZN(new_n874));
  INV_X1    g673(.A(new_n851), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n875), .B1(new_n847), .B2(new_n849), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n874), .B1(new_n876), .B2(new_n462), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n875), .B1(new_n846), .B2(new_n864), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n462), .A2(new_n874), .ZN(new_n879));
  INV_X1    g678(.A(new_n879), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n877), .A2(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(new_n853), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n884), .A2(new_n467), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n883), .A2(new_n571), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(G141gat), .ZN(new_n887));
  OAI21_X1  g686(.A(KEYINPUT121), .B1(new_n876), .B2(new_n445), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT121), .ZN(new_n889));
  AND3_X1   g688(.A1(new_n843), .A2(new_n848), .A3(new_n845), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n848), .B1(new_n843), .B2(new_n845), .ZN(new_n891));
  NOR3_X1   g690(.A1(new_n890), .A2(new_n891), .A3(new_n663), .ZN(new_n892));
  OAI211_X1 g691(.A(new_n889), .B(new_n473), .C1(new_n892), .C2(new_n875), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n467), .A2(new_n462), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n888), .A2(new_n893), .A3(new_n288), .A4(new_n894), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n685), .A2(G141gat), .ZN(new_n896));
  INV_X1    g695(.A(new_n896), .ZN(new_n897));
  OR2_X1    g696(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT58), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n887), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(new_n885), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n901), .B1(new_n877), .B2(new_n882), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n293), .B1(new_n902), .B2(new_n571), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n895), .A2(new_n897), .ZN(new_n904));
  OAI21_X1  g703(.A(KEYINPUT58), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n900), .A2(new_n905), .ZN(G1344gat));
  OAI21_X1  g705(.A(KEYINPUT59), .B1(new_n895), .B2(new_n621), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(new_n295), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n879), .B1(new_n892), .B2(new_n875), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n874), .B1(new_n878), .B2(new_n462), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT122), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  OAI211_X1 g711(.A(KEYINPUT122), .B(new_n874), .C1(new_n878), .C2(new_n462), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n909), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n914), .A2(new_n620), .A3(new_n885), .ZN(new_n915));
  AND2_X1   g714(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n621), .A2(KEYINPUT59), .ZN(new_n917));
  AOI22_X1  g716(.A1(new_n915), .A2(new_n916), .B1(new_n902), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n908), .A2(new_n918), .ZN(G1345gat));
  AND3_X1   g718(.A1(new_n902), .A2(G155gat), .A3(new_n663), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n895), .A2(new_n864), .ZN(new_n921));
  AOI21_X1  g720(.A(G155gat), .B1(new_n921), .B2(KEYINPUT123), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT123), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n923), .B1(new_n895), .B2(new_n864), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n920), .B1(new_n922), .B2(new_n924), .ZN(G1346gat));
  INV_X1    g724(.A(new_n902), .ZN(new_n926));
  OAI21_X1  g725(.A(G162gat), .B1(new_n926), .B2(new_n690), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n868), .A2(G162gat), .ZN(new_n928));
  NAND4_X1  g727(.A1(new_n888), .A2(new_n893), .A3(new_n894), .A4(new_n928), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT124), .ZN(new_n930));
  AND2_X1   g729(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n929), .A2(new_n930), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n927), .B1(new_n931), .B2(new_n932), .ZN(G1347gat));
  NOR2_X1   g732(.A1(new_n473), .A2(new_n288), .ZN(new_n934));
  INV_X1    g733(.A(new_n934), .ZN(new_n935));
  NOR3_X1   g734(.A1(new_n876), .A2(new_n341), .A3(new_n935), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n936), .A2(new_n756), .ZN(new_n937));
  OAI21_X1  g736(.A(G169gat), .B1(new_n937), .B2(new_n685), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n455), .A2(new_n456), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n936), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n571), .A2(new_n236), .A3(new_n237), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n938), .B1(new_n940), .B2(new_n941), .ZN(G1348gat));
  OAI21_X1  g741(.A(G176gat), .B1(new_n937), .B2(new_n621), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n620), .A2(new_n218), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n943), .B1(new_n940), .B2(new_n944), .ZN(G1349gat));
  NAND3_X1  g744(.A1(new_n936), .A2(new_n663), .A3(new_n756), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n946), .A2(G183gat), .ZN(new_n947));
  INV_X1    g746(.A(new_n947), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n663), .A2(new_n250), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n940), .A2(new_n949), .ZN(new_n950));
  OAI21_X1  g749(.A(KEYINPUT60), .B1(new_n948), .B2(new_n950), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT60), .ZN(new_n952));
  OAI211_X1 g751(.A(new_n947), .B(new_n952), .C1(new_n940), .C2(new_n949), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n951), .A2(new_n953), .ZN(G1350gat));
  NAND3_X1  g753(.A1(new_n936), .A2(new_n682), .A3(new_n756), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT61), .ZN(new_n956));
  AND3_X1   g755(.A1(new_n955), .A2(new_n956), .A3(G190gat), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n956), .B1(new_n955), .B2(G190gat), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n682), .A2(new_n251), .ZN(new_n959));
  OAI22_X1  g758(.A1(new_n957), .A2(new_n958), .B1(new_n940), .B2(new_n959), .ZN(G1351gat));
  NOR4_X1   g759(.A1(new_n876), .A2(new_n462), .A3(new_n467), .A4(new_n935), .ZN(new_n961));
  XNOR2_X1  g760(.A(KEYINPUT125), .B(G197gat), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n961), .A2(new_n571), .A3(new_n962), .ZN(new_n963));
  NOR2_X1   g762(.A1(new_n935), .A2(new_n467), .ZN(new_n964));
  AND3_X1   g763(.A1(new_n914), .A2(new_n571), .A3(new_n964), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n963), .B1(new_n965), .B2(new_n962), .ZN(G1352gat));
  INV_X1    g765(.A(G204gat), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n961), .A2(new_n967), .A3(new_n620), .ZN(new_n968));
  OR2_X1    g767(.A1(new_n968), .A2(KEYINPUT62), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n968), .A2(KEYINPUT62), .ZN(new_n970));
  AND3_X1   g769(.A1(new_n914), .A2(new_n620), .A3(new_n964), .ZN(new_n971));
  OAI211_X1 g770(.A(new_n969), .B(new_n970), .C1(new_n967), .C2(new_n971), .ZN(G1353gat));
  NAND3_X1  g771(.A1(new_n961), .A2(new_n259), .A3(new_n663), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n914), .A2(new_n663), .A3(new_n964), .ZN(new_n974));
  AND2_X1   g773(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n975));
  OAI21_X1  g774(.A(G211gat), .B1(KEYINPUT126), .B2(KEYINPUT63), .ZN(new_n976));
  INV_X1    g775(.A(new_n976), .ZN(new_n977));
  AND3_X1   g776(.A1(new_n974), .A2(new_n975), .A3(new_n977), .ZN(new_n978));
  AOI21_X1  g777(.A(new_n975), .B1(new_n974), .B2(new_n977), .ZN(new_n979));
  OAI21_X1  g778(.A(new_n973), .B1(new_n978), .B2(new_n979), .ZN(G1354gat));
  NAND3_X1  g779(.A1(new_n961), .A2(new_n260), .A3(new_n682), .ZN(new_n981));
  AND3_X1   g780(.A1(new_n914), .A2(new_n682), .A3(new_n964), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n981), .B1(new_n982), .B2(new_n260), .ZN(G1355gat));
endmodule


