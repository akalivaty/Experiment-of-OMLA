//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 0 0 0 1 0 1 1 0 1 1 0 1 0 0 1 0 1 1 1 1 0 1 0 0 1 1 0 0 1 1 0 0 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 0 0 1 1 1 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:40 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n644, new_n645,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n727, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n821, new_n822, new_n823, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n889, new_n890, new_n891, new_n892, new_n894, new_n895, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n909, new_n910, new_n911, new_n913, new_n914,
    new_n915, new_n916, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n925, new_n926, new_n927, new_n928, new_n930, new_n931,
    new_n932, new_n933, new_n935, new_n936, new_n937;
  XNOR2_X1  g000(.A(G1gat), .B(G29gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT0), .ZN(new_n203));
  XNOR2_X1  g002(.A(G57gat), .B(G85gat), .ZN(new_n204));
  XOR2_X1   g003(.A(new_n203), .B(new_n204), .Z(new_n205));
  XOR2_X1   g004(.A(G127gat), .B(G134gat), .Z(new_n206));
  XNOR2_X1  g005(.A(G113gat), .B(G120gat), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n206), .B1(KEYINPUT1), .B2(new_n207), .ZN(new_n208));
  XOR2_X1   g007(.A(G113gat), .B(G120gat), .Z(new_n209));
  INV_X1    g008(.A(KEYINPUT1), .ZN(new_n210));
  XNOR2_X1  g009(.A(G127gat), .B(G134gat), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n209), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n208), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT73), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n208), .A2(new_n212), .A3(KEYINPUT73), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT72), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT2), .ZN(new_n219));
  INV_X1    g018(.A(G155gat), .ZN(new_n220));
  INV_X1    g019(.A(G162gat), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n219), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(G155gat), .A2(G162gat), .ZN(new_n223));
  INV_X1    g022(.A(G148gat), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n224), .A2(G141gat), .ZN(new_n225));
  AOI22_X1  g024(.A1(new_n222), .A2(new_n223), .B1(new_n225), .B2(KEYINPUT71), .ZN(new_n226));
  XNOR2_X1  g025(.A(G141gat), .B(G148gat), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT71), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(G141gat), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n230), .A2(G148gat), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n219), .B1(new_n225), .B2(new_n231), .ZN(new_n232));
  XOR2_X1   g031(.A(G155gat), .B(G162gat), .Z(new_n233));
  AOI22_X1  g032(.A1(new_n226), .A2(new_n229), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT3), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n218), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n226), .A2(new_n229), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n232), .A2(new_n233), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n239), .A2(KEYINPUT72), .A3(KEYINPUT3), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n234), .A2(new_n235), .ZN(new_n241));
  NAND4_X1  g040(.A1(new_n217), .A2(new_n236), .A3(new_n240), .A4(new_n241), .ZN(new_n242));
  NAND4_X1  g041(.A1(new_n237), .A2(new_n238), .A3(new_n212), .A4(new_n208), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n243), .B(KEYINPUT4), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT5), .ZN(new_n245));
  NAND2_X1  g044(.A1(G225gat), .A2(G233gat), .ZN(new_n246));
  NAND4_X1  g045(.A1(new_n242), .A2(new_n244), .A3(new_n245), .A4(new_n246), .ZN(new_n247));
  AND3_X1   g046(.A1(new_n242), .A2(new_n244), .A3(new_n246), .ZN(new_n248));
  INV_X1    g047(.A(new_n243), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n249), .B1(new_n217), .B2(new_n239), .ZN(new_n250));
  OAI21_X1  g049(.A(KEYINPUT5), .B1(new_n250), .B2(new_n246), .ZN(new_n251));
  OAI211_X1 g050(.A(new_n205), .B(new_n247), .C1(new_n248), .C2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT6), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n247), .B1(new_n248), .B2(new_n251), .ZN(new_n256));
  INV_X1    g055(.A(new_n205), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n258), .A2(KEYINPUT79), .ZN(new_n259));
  AND3_X1   g058(.A1(new_n208), .A2(new_n212), .A3(KEYINPUT73), .ZN(new_n260));
  AOI21_X1  g059(.A(KEYINPUT73), .B1(new_n208), .B2(new_n212), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n239), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(new_n243), .ZN(new_n263));
  INV_X1    g062(.A(new_n246), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n245), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n242), .A2(new_n244), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n265), .B1(new_n266), .B2(new_n264), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n205), .B1(new_n267), .B2(new_n247), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT79), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND4_X1  g069(.A1(new_n255), .A2(new_n259), .A3(KEYINPUT80), .A4(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n268), .A2(KEYINPUT6), .ZN(new_n272));
  AND2_X1   g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT82), .ZN(new_n274));
  AND2_X1   g073(.A1(G226gat), .A2(G233gat), .ZN(new_n275));
  XNOR2_X1  g074(.A(KEYINPUT27), .B(G183gat), .ZN(new_n276));
  INV_X1    g075(.A(G190gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT66), .ZN(new_n279));
  OR2_X1    g078(.A1(new_n279), .A2(KEYINPUT28), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n278), .B(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(G169gat), .ZN(new_n283));
  INV_X1    g082(.A(G176gat), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n283), .A2(new_n284), .A3(KEYINPUT26), .ZN(new_n285));
  NAND2_X1  g084(.A1(G183gat), .A2(G190gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(G169gat), .A2(G176gat), .ZN(new_n288));
  AOI21_X1  g087(.A(KEYINPUT26), .B1(new_n283), .B2(new_n284), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n287), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n282), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT64), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT24), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n293), .A2(G183gat), .A3(G190gat), .ZN(new_n294));
  XNOR2_X1  g093(.A(G183gat), .B(G190gat), .ZN(new_n295));
  OAI211_X1 g094(.A(new_n292), .B(new_n294), .C1(new_n295), .C2(new_n293), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT25), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n294), .B1(new_n295), .B2(new_n293), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n283), .A2(new_n284), .A3(KEYINPUT23), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT23), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n300), .B1(G169gat), .B2(G176gat), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n299), .A2(new_n301), .A3(new_n288), .ZN(new_n302));
  OAI211_X1 g101(.A(new_n296), .B(new_n297), .C1(new_n298), .C2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT65), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n286), .A2(KEYINPUT24), .ZN(new_n305));
  INV_X1    g104(.A(G183gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(G190gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n277), .A2(G183gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n305), .B1(new_n309), .B2(KEYINPUT24), .ZN(new_n310));
  INV_X1    g109(.A(new_n302), .ZN(new_n311));
  OAI211_X1 g110(.A(new_n310), .B(new_n311), .C1(new_n292), .C2(KEYINPUT25), .ZN(new_n312));
  AND3_X1   g111(.A1(new_n303), .A2(new_n304), .A3(new_n312), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n304), .B1(new_n303), .B2(new_n312), .ZN(new_n314));
  OAI211_X1 g113(.A(new_n275), .B(new_n291), .C1(new_n313), .C2(new_n314), .ZN(new_n315));
  XOR2_X1   g114(.A(G211gat), .B(G218gat), .Z(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  OR2_X1    g116(.A1(new_n317), .A2(KEYINPUT69), .ZN(new_n318));
  XNOR2_X1  g117(.A(G197gat), .B(G204gat), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT22), .ZN(new_n320));
  INV_X1    g119(.A(G211gat), .ZN(new_n321));
  INV_X1    g120(.A(G218gat), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n320), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n319), .A2(new_n323), .ZN(new_n324));
  XNOR2_X1  g123(.A(new_n318), .B(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n303), .A2(new_n312), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n291), .A2(new_n326), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n275), .A2(KEYINPUT29), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n315), .A2(new_n325), .A3(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT81), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n291), .B1(new_n313), .B2(new_n314), .ZN(new_n332));
  INV_X1    g131(.A(new_n327), .ZN(new_n333));
  AOI22_X1  g132(.A1(new_n332), .A2(new_n328), .B1(new_n333), .B2(new_n275), .ZN(new_n334));
  OAI211_X1 g133(.A(new_n330), .B(new_n331), .C1(new_n334), .C2(new_n325), .ZN(new_n335));
  OR2_X1    g134(.A1(new_n330), .A2(new_n331), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n335), .A2(new_n336), .A3(KEYINPUT37), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT38), .ZN(new_n339));
  XNOR2_X1  g138(.A(G8gat), .B(G36gat), .ZN(new_n340));
  XNOR2_X1  g139(.A(G64gat), .B(G92gat), .ZN(new_n341));
  XOR2_X1   g140(.A(new_n340), .B(new_n341), .Z(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n334), .A2(new_n325), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n325), .B1(new_n315), .B2(new_n329), .ZN(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  OAI211_X1 g146(.A(new_n339), .B(new_n343), .C1(new_n347), .C2(KEYINPUT37), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n274), .B1(new_n338), .B2(new_n348), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n345), .B1(new_n325), .B2(new_n334), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT37), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n342), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n352), .A2(KEYINPUT82), .A3(new_n337), .A4(new_n339), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n349), .A2(new_n353), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n352), .B1(new_n351), .B2(new_n350), .ZN(new_n355));
  AOI22_X1  g154(.A1(new_n355), .A2(KEYINPUT38), .B1(new_n342), .B2(new_n350), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n255), .A2(new_n259), .A3(new_n270), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT80), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND4_X1  g158(.A1(new_n273), .A2(new_n354), .A3(new_n356), .A4(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(G228gat), .A2(G233gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n361), .B(KEYINPUT75), .ZN(new_n362));
  INV_X1    g161(.A(new_n325), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT29), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n363), .B1(new_n364), .B2(new_n241), .ZN(new_n365));
  AOI21_X1  g164(.A(KEYINPUT29), .B1(new_n317), .B2(new_n324), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n366), .B1(new_n324), .B2(new_n317), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n234), .B1(new_n367), .B2(new_n235), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n362), .B1(new_n365), .B2(new_n368), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n235), .B1(new_n325), .B2(KEYINPUT29), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(new_n239), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n371), .A2(G228gat), .A3(G233gat), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n369), .B1(new_n372), .B2(new_n365), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT76), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(G22gat), .ZN(new_n375));
  XNOR2_X1  g174(.A(G78gat), .B(G106gat), .ZN(new_n376));
  XNOR2_X1  g175(.A(KEYINPUT31), .B(G50gat), .ZN(new_n377));
  XNOR2_X1  g176(.A(new_n376), .B(new_n377), .ZN(new_n378));
  MUX2_X1   g177(.A(G22gat), .B(new_n375), .S(new_n378), .Z(new_n379));
  XOR2_X1   g178(.A(new_n373), .B(new_n379), .Z(new_n380));
  NAND3_X1  g179(.A1(new_n344), .A2(new_n346), .A3(new_n342), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT30), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n347), .A2(new_n343), .ZN(new_n384));
  NAND4_X1  g183(.A1(new_n344), .A2(new_n346), .A3(KEYINPUT30), .A4(new_n342), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n383), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  AND3_X1   g185(.A1(new_n386), .A2(new_n259), .A3(new_n270), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n266), .A2(new_n264), .ZN(new_n388));
  OAI211_X1 g187(.A(new_n388), .B(KEYINPUT39), .C1(new_n264), .C2(new_n263), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT39), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n266), .A2(new_n390), .A3(new_n264), .ZN(new_n391));
  AND3_X1   g190(.A1(new_n391), .A2(KEYINPUT77), .A3(new_n205), .ZN(new_n392));
  AOI21_X1  g191(.A(KEYINPUT77), .B1(new_n391), .B2(new_n205), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n389), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT78), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n395), .A2(KEYINPUT40), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  XNOR2_X1  g196(.A(new_n394), .B(new_n397), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n380), .B1(new_n387), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n360), .A2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT74), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n401), .B1(new_n254), .B2(new_n268), .ZN(new_n402));
  NAND4_X1  g201(.A1(new_n258), .A2(KEYINPUT74), .A3(new_n253), .A4(new_n252), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n402), .A2(new_n403), .A3(new_n272), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n384), .A2(new_n385), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT70), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n384), .A2(KEYINPUT70), .A3(new_n385), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n404), .A2(new_n383), .A3(new_n407), .A4(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(new_n380), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT36), .ZN(new_n411));
  NAND2_X1  g210(.A1(G227gat), .A2(G233gat), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n213), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n326), .A2(KEYINPUT65), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n303), .A2(new_n312), .A3(new_n304), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n414), .B1(new_n417), .B2(new_n291), .ZN(new_n418));
  OAI211_X1 g217(.A(new_n414), .B(new_n291), .C1(new_n313), .C2(new_n314), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n413), .B1(new_n418), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(KEYINPUT32), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT33), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  XNOR2_X1  g223(.A(G15gat), .B(G43gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(new_n425), .B(KEYINPUT67), .ZN(new_n426));
  INV_X1    g225(.A(G71gat), .ZN(new_n427));
  XNOR2_X1  g226(.A(new_n426), .B(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(G99gat), .ZN(new_n429));
  XNOR2_X1  g228(.A(new_n428), .B(new_n429), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n422), .A2(new_n424), .A3(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n430), .ZN(new_n432));
  OAI211_X1 g231(.A(new_n421), .B(KEYINPUT32), .C1(new_n423), .C2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n332), .A2(new_n213), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(new_n419), .ZN(new_n436));
  OAI21_X1  g235(.A(KEYINPUT34), .B1(new_n436), .B2(new_n413), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT34), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n435), .A2(new_n438), .A3(new_n412), .A4(new_n419), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n434), .A2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n431), .A2(new_n440), .A3(new_n433), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n411), .B1(new_n443), .B2(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n412), .B1(new_n435), .B2(new_n419), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n430), .B1(new_n447), .B2(KEYINPUT33), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT32), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  AOI221_X4 g250(.A(new_n449), .B1(new_n430), .B2(KEYINPUT33), .C1(new_n436), .C2(new_n413), .ZN(new_n452));
  OAI21_X1  g251(.A(KEYINPUT68), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(new_n440), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n434), .A2(KEYINPUT68), .A3(new_n441), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n454), .A2(KEYINPUT36), .A3(new_n455), .ZN(new_n456));
  NAND4_X1  g255(.A1(new_n400), .A2(new_n410), .A3(new_n446), .A4(new_n456), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n380), .B1(new_n444), .B2(new_n442), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT35), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n359), .A2(new_n272), .A3(new_n271), .ZN(new_n460));
  INV_X1    g259(.A(new_n386), .ZN(new_n461));
  NAND4_X1  g260(.A1(new_n458), .A2(new_n459), .A3(new_n460), .A4(new_n461), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n380), .B1(new_n454), .B2(new_n455), .ZN(new_n463));
  AND4_X1   g262(.A1(new_n404), .A2(new_n383), .A3(new_n407), .A4(new_n408), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n459), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n462), .B1(new_n465), .B2(KEYINPUT83), .ZN(new_n466));
  XNOR2_X1  g265(.A(new_n373), .B(new_n379), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n441), .B1(new_n434), .B2(KEYINPUT68), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT68), .ZN(new_n469));
  AOI211_X1 g268(.A(new_n469), .B(new_n440), .C1(new_n431), .C2(new_n433), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n467), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  OAI211_X1 g270(.A(KEYINPUT83), .B(KEYINPUT35), .C1(new_n471), .C2(new_n409), .ZN(new_n472));
  INV_X1    g271(.A(new_n472), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n457), .B1(new_n466), .B2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT84), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  OAI211_X1 g275(.A(new_n457), .B(KEYINPUT84), .C1(new_n466), .C2(new_n473), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT87), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT15), .ZN(new_n480));
  XNOR2_X1  g279(.A(KEYINPUT14), .B(G29gat), .ZN(new_n481));
  INV_X1    g280(.A(G36gat), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(G29gat), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n484), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT85), .ZN(new_n487));
  XNOR2_X1  g286(.A(G43gat), .B(G50gat), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n486), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(new_n488), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n483), .A2(new_n490), .A3(new_n485), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n480), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  AOI22_X1  g291(.A1(new_n483), .A2(new_n485), .B1(new_n490), .B2(KEYINPUT85), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n493), .A2(KEYINPUT15), .ZN(new_n494));
  OAI21_X1  g293(.A(KEYINPUT86), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(new_n491), .ZN(new_n496));
  OAI21_X1  g295(.A(KEYINPUT15), .B1(new_n496), .B2(new_n493), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n489), .A2(new_n480), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT86), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n497), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n495), .A2(new_n500), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n479), .B1(new_n501), .B2(KEYINPUT17), .ZN(new_n502));
  XNOR2_X1  g301(.A(G15gat), .B(G22gat), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT16), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n503), .B1(new_n504), .B2(G1gat), .ZN(new_n505));
  OAI211_X1 g304(.A(new_n505), .B(KEYINPUT88), .C1(G1gat), .C2(new_n503), .ZN(new_n506));
  INV_X1    g305(.A(G8gat), .ZN(new_n507));
  XNOR2_X1  g306(.A(new_n506), .B(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT17), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n495), .A2(KEYINPUT87), .A3(new_n500), .A4(new_n509), .ZN(new_n510));
  OAI21_X1  g309(.A(KEYINPUT17), .B1(new_n492), .B2(new_n494), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n502), .A2(new_n508), .A3(new_n510), .A4(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(G229gat), .A2(G233gat), .ZN(new_n513));
  INV_X1    g312(.A(new_n501), .ZN(new_n514));
  INV_X1    g313(.A(new_n508), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n512), .A2(new_n513), .A3(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT18), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n512), .A2(KEYINPUT18), .A3(new_n513), .A4(new_n516), .ZN(new_n520));
  AOI21_X1  g319(.A(KEYINPUT89), .B1(new_n501), .B2(new_n508), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n516), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n514), .A2(KEYINPUT89), .A3(new_n515), .ZN(new_n523));
  XOR2_X1   g322(.A(new_n513), .B(KEYINPUT13), .Z(new_n524));
  NAND3_X1  g323(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n519), .A2(new_n520), .A3(new_n525), .ZN(new_n526));
  XNOR2_X1  g325(.A(G113gat), .B(G141gat), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n527), .B(G197gat), .ZN(new_n528));
  XOR2_X1   g327(.A(KEYINPUT11), .B(G169gat), .Z(new_n529));
  XNOR2_X1  g328(.A(new_n528), .B(new_n529), .ZN(new_n530));
  XOR2_X1   g329(.A(new_n530), .B(KEYINPUT12), .Z(new_n531));
  NAND2_X1  g330(.A1(new_n526), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(new_n531), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n519), .A2(new_n533), .A3(new_n520), .A4(new_n525), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT90), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n532), .A2(KEYINPUT90), .A3(new_n534), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT102), .ZN(new_n541));
  INV_X1    g340(.A(G230gat), .ZN(new_n542));
  INV_X1    g341(.A(G233gat), .ZN(new_n543));
  NOR2_X1   g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  XOR2_X1   g343(.A(G99gat), .B(G106gat), .Z(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(G85gat), .A2(G92gat), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n547), .B(KEYINPUT7), .ZN(new_n548));
  XNOR2_X1  g347(.A(KEYINPUT95), .B(G92gat), .ZN(new_n549));
  INV_X1    g348(.A(G85gat), .ZN(new_n550));
  NAND2_X1  g349(.A1(G99gat), .A2(G106gat), .ZN(new_n551));
  AOI22_X1  g350(.A1(new_n549), .A2(new_n550), .B1(KEYINPUT8), .B2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT96), .ZN(new_n553));
  AND2_X1   g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n552), .A2(new_n553), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n548), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n546), .B1(new_n556), .B2(KEYINPUT99), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n557), .B1(KEYINPUT99), .B2(new_n556), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n558), .A2(KEYINPUT100), .ZN(new_n559));
  XNOR2_X1  g358(.A(G57gat), .B(G64gat), .ZN(new_n560));
  AOI21_X1  g359(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n561));
  OR2_X1    g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(G71gat), .B(G78gat), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n562), .B(new_n563), .ZN(new_n564));
  OR2_X1    g363(.A1(new_n556), .A2(new_n545), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT100), .ZN(new_n566));
  OAI211_X1 g365(.A(new_n557), .B(new_n566), .C1(KEYINPUT99), .C2(new_n556), .ZN(new_n567));
  NAND4_X1  g366(.A1(new_n559), .A2(new_n564), .A3(new_n565), .A4(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT10), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n556), .B(new_n546), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n570), .A2(new_n564), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n568), .A2(new_n569), .A3(new_n572), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n570), .A2(KEYINPUT10), .A3(new_n564), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n544), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  AOI211_X1 g374(.A(new_n542), .B(new_n543), .C1(new_n568), .C2(new_n572), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n541), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  XOR2_X1   g376(.A(G120gat), .B(G148gat), .Z(new_n578));
  XNOR2_X1  g377(.A(new_n578), .B(KEYINPUT101), .ZN(new_n579));
  XNOR2_X1  g378(.A(G176gat), .B(G204gat), .ZN(new_n580));
  XOR2_X1   g379(.A(new_n579), .B(new_n580), .Z(new_n581));
  XNOR2_X1  g380(.A(new_n577), .B(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n570), .ZN(new_n584));
  NAND4_X1  g383(.A1(new_n502), .A2(new_n510), .A3(new_n511), .A4(new_n584), .ZN(new_n585));
  AND3_X1   g384(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n586), .B1(new_n514), .B2(new_n570), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(G190gat), .B(G218gat), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n588), .A2(new_n589), .ZN(new_n592));
  XOR2_X1   g391(.A(G134gat), .B(G162gat), .Z(new_n593));
  AOI21_X1  g392(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n593), .B(new_n594), .ZN(new_n595));
  NOR3_X1   g394(.A1(new_n591), .A2(new_n592), .A3(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT97), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n597), .B1(new_n588), .B2(new_n589), .ZN(new_n598));
  INV_X1    g397(.A(new_n589), .ZN(new_n599));
  NAND4_X1  g398(.A1(new_n585), .A2(KEYINPUT97), .A3(new_n587), .A4(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n598), .A2(new_n600), .A3(new_n590), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n595), .B(KEYINPUT94), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n603), .A2(KEYINPUT98), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT98), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n601), .A2(new_n605), .A3(new_n602), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n596), .B1(new_n604), .B2(new_n606), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n515), .B1(KEYINPUT21), .B2(new_n564), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(KEYINPUT93), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n564), .A2(KEYINPUT21), .ZN(new_n610));
  XNOR2_X1  g409(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n610), .B(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n609), .B(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(G127gat), .B(G155gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(KEYINPUT92), .ZN(new_n615));
  NAND2_X1  g414(.A1(G231gat), .A2(G233gat), .ZN(new_n616));
  XOR2_X1   g415(.A(new_n616), .B(KEYINPUT91), .Z(new_n617));
  XNOR2_X1  g416(.A(new_n615), .B(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(G183gat), .B(G211gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n613), .B(new_n620), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n583), .A2(new_n607), .A3(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n478), .A2(new_n540), .A3(new_n623), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n624), .A2(new_n404), .ZN(new_n625));
  XOR2_X1   g424(.A(new_n625), .B(G1gat), .Z(G1324gat));
  NOR2_X1   g425(.A1(new_n624), .A2(new_n461), .ZN(new_n627));
  XOR2_X1   g426(.A(KEYINPUT16), .B(G8gat), .Z(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT103), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT42), .ZN(new_n631));
  NOR3_X1   g430(.A1(new_n629), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n629), .A2(new_n631), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n633), .A2(KEYINPUT103), .ZN(new_n634));
  OAI21_X1  g433(.A(KEYINPUT42), .B1(new_n627), .B2(new_n507), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n635), .A2(new_n629), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n632), .B1(new_n634), .B2(new_n636), .ZN(G1325gat));
  NAND2_X1  g436(.A1(new_n446), .A2(new_n456), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  OAI21_X1  g438(.A(G15gat), .B1(new_n624), .B2(new_n639), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n443), .A2(new_n445), .ZN(new_n641));
  OR2_X1    g440(.A1(new_n641), .A2(G15gat), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n640), .B1(new_n624), .B2(new_n642), .ZN(G1326gat));
  NOR2_X1   g442(.A1(new_n624), .A2(new_n467), .ZN(new_n644));
  XOR2_X1   g443(.A(KEYINPUT43), .B(G22gat), .Z(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(G1327gat));
  NOR2_X1   g445(.A1(new_n582), .A2(new_n621), .ZN(new_n647));
  INV_X1    g446(.A(new_n596), .ZN(new_n648));
  INV_X1    g447(.A(new_n606), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n605), .B1(new_n601), .B2(new_n602), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n648), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n647), .A2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n477), .ZN(new_n654));
  OAI21_X1  g453(.A(KEYINPUT35), .B1(new_n471), .B2(new_n409), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT83), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n657), .A2(new_n472), .A3(new_n462), .ZN(new_n658));
  AOI21_X1  g457(.A(KEYINPUT84), .B1(new_n658), .B2(new_n457), .ZN(new_n659));
  OAI211_X1 g458(.A(new_n540), .B(new_n653), .C1(new_n654), .C2(new_n659), .ZN(new_n660));
  NOR3_X1   g459(.A1(new_n660), .A2(G29gat), .A3(new_n404), .ZN(new_n661));
  XOR2_X1   g460(.A(new_n661), .B(KEYINPUT45), .Z(new_n662));
  INV_X1    g461(.A(KEYINPUT44), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n607), .A2(new_n663), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n664), .B1(new_n654), .B2(new_n659), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n474), .A2(new_n651), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n666), .A2(new_n663), .ZN(new_n667));
  AND2_X1   g466(.A1(new_n647), .A2(new_n535), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n665), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT104), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n404), .ZN(new_n672));
  NAND4_X1  g471(.A1(new_n665), .A2(KEYINPUT104), .A3(new_n667), .A4(new_n668), .ZN(new_n673));
  AND3_X1   g472(.A1(new_n671), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n662), .B1(new_n484), .B2(new_n674), .ZN(G1328gat));
  NOR3_X1   g474(.A1(new_n660), .A2(G36gat), .A3(new_n461), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(KEYINPUT46), .ZN(new_n677));
  AND3_X1   g476(.A1(new_n671), .A2(new_n386), .A3(new_n673), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n677), .B1(new_n482), .B2(new_n678), .ZN(G1329gat));
  OAI21_X1  g478(.A(G43gat), .B1(new_n669), .B2(new_n639), .ZN(new_n680));
  OR3_X1    g479(.A1(new_n660), .A2(G43gat), .A3(new_n641), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n680), .A2(KEYINPUT47), .A3(new_n681), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n671), .A2(new_n638), .A3(new_n673), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT105), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n683), .A2(new_n684), .A3(G43gat), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT47), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n681), .A2(KEYINPUT105), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n688), .B1(new_n683), .B2(G43gat), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n682), .B1(new_n687), .B2(new_n689), .ZN(G1330gat));
  INV_X1    g489(.A(KEYINPUT107), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT106), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n660), .A2(new_n692), .ZN(new_n693));
  NAND4_X1  g492(.A1(new_n478), .A2(KEYINPUT106), .A3(new_n540), .A4(new_n653), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n467), .A2(G50gat), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n693), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  AND2_X1   g495(.A1(new_n696), .A2(KEYINPUT48), .ZN(new_n697));
  OAI21_X1  g496(.A(G50gat), .B1(new_n669), .B2(new_n467), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n691), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  AND4_X1   g498(.A1(new_n691), .A2(new_n698), .A3(KEYINPUT48), .A4(new_n696), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n671), .A2(new_n380), .A3(new_n673), .ZN(new_n701));
  AND2_X1   g500(.A1(new_n694), .A2(new_n695), .ZN(new_n702));
  AOI22_X1  g501(.A1(new_n701), .A2(G50gat), .B1(new_n693), .B2(new_n702), .ZN(new_n703));
  OAI22_X1  g502(.A1(new_n699), .A2(new_n700), .B1(new_n703), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g503(.A1(new_n607), .A2(new_n621), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n705), .A2(new_n535), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(new_n582), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n707), .B(KEYINPUT108), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(new_n474), .ZN(new_n709));
  INV_X1    g508(.A(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(new_n672), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n711), .B(G57gat), .ZN(G1332gat));
  XNOR2_X1  g511(.A(new_n386), .B(KEYINPUT109), .ZN(new_n713));
  INV_X1    g512(.A(new_n713), .ZN(new_n714));
  XNOR2_X1  g513(.A(KEYINPUT49), .B(G64gat), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n710), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  OAI22_X1  g515(.A1(new_n709), .A2(new_n713), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT110), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n718), .B(new_n719), .ZN(G1333gat));
  OAI21_X1  g519(.A(G71gat), .B1(new_n709), .B2(new_n639), .ZN(new_n721));
  INV_X1    g520(.A(new_n641), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(new_n427), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n721), .B1(new_n709), .B2(new_n723), .ZN(new_n724));
  XNOR2_X1  g523(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n724), .B(new_n725), .ZN(G1334gat));
  NAND2_X1  g525(.A1(new_n710), .A2(new_n380), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g527(.A1(new_n621), .A2(new_n535), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n474), .A2(new_n651), .A3(new_n729), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(KEYINPUT51), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(KEYINPUT112), .ZN(new_n732));
  NAND4_X1  g531(.A1(new_n732), .A2(new_n550), .A3(new_n672), .A4(new_n582), .ZN(new_n733));
  AND2_X1   g532(.A1(new_n665), .A2(new_n667), .ZN(new_n734));
  AND2_X1   g533(.A1(new_n729), .A2(new_n582), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  OAI21_X1  g535(.A(G85gat), .B1(new_n736), .B2(new_n404), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n733), .A2(new_n737), .ZN(G1336gat));
  INV_X1    g537(.A(KEYINPUT52), .ZN(new_n739));
  NOR3_X1   g538(.A1(new_n583), .A2(G92gat), .A3(new_n713), .ZN(new_n740));
  INV_X1    g539(.A(new_n740), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n665), .A2(new_n667), .A3(new_n714), .A4(new_n735), .ZN(new_n742));
  AND2_X1   g541(.A1(new_n742), .A2(KEYINPUT116), .ZN(new_n743));
  INV_X1    g542(.A(new_n549), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n744), .B1(new_n742), .B2(KEYINPUT116), .ZN(new_n745));
  OAI221_X1 g544(.A(new_n739), .B1(new_n731), .B2(new_n741), .C1(new_n743), .C2(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT51), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT113), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n730), .A2(new_n748), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n747), .B1(new_n749), .B2(KEYINPUT114), .ZN(new_n750));
  OAI21_X1  g549(.A(KEYINPUT113), .B1(new_n747), .B2(KEYINPUT114), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n730), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n750), .A2(new_n740), .A3(new_n752), .ZN(new_n753));
  NAND4_X1  g552(.A1(new_n665), .A2(new_n386), .A3(new_n667), .A4(new_n735), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(new_n744), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  AND3_X1   g555(.A1(new_n756), .A2(KEYINPUT115), .A3(KEYINPUT52), .ZN(new_n757));
  AOI21_X1  g556(.A(KEYINPUT115), .B1(new_n756), .B2(KEYINPUT52), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n746), .B1(new_n757), .B2(new_n758), .ZN(G1337gat));
  NAND4_X1  g558(.A1(new_n732), .A2(new_n429), .A3(new_n722), .A4(new_n582), .ZN(new_n760));
  OAI21_X1  g559(.A(G99gat), .B1(new_n736), .B2(new_n639), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(G1338gat));
  AND2_X1   g561(.A1(new_n750), .A2(new_n752), .ZN(new_n763));
  NOR3_X1   g562(.A1(new_n583), .A2(G106gat), .A3(new_n467), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n734), .A2(new_n380), .A3(new_n735), .ZN(new_n765));
  AOI22_X1  g564(.A1(new_n763), .A2(new_n764), .B1(new_n765), .B2(G106gat), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT53), .ZN(new_n767));
  AND2_X1   g566(.A1(new_n765), .A2(G106gat), .ZN(new_n768));
  INV_X1    g567(.A(new_n764), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n767), .B1(new_n731), .B2(new_n769), .ZN(new_n770));
  OAI22_X1  g569(.A1(new_n766), .A2(new_n767), .B1(new_n768), .B2(new_n770), .ZN(G1339gat));
  INV_X1    g570(.A(KEYINPUT118), .ZN(new_n772));
  INV_X1    g571(.A(new_n621), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n565), .A2(new_n564), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n774), .B1(KEYINPUT100), .B2(new_n558), .ZN(new_n775));
  AOI211_X1 g574(.A(KEYINPUT10), .B(new_n571), .C1(new_n775), .C2(new_n567), .ZN(new_n776));
  INV_X1    g575(.A(new_n574), .ZN(new_n777));
  OAI22_X1  g576(.A1(new_n776), .A2(new_n777), .B1(new_n542), .B2(new_n543), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n573), .A2(new_n544), .A3(new_n574), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n778), .A2(KEYINPUT54), .A3(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT54), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n581), .B1(new_n575), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT55), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n575), .A2(new_n576), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(new_n581), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n780), .A2(new_n782), .A3(KEYINPUT55), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n785), .A2(new_n535), .A3(new_n787), .A4(new_n788), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n513), .B1(new_n512), .B2(new_n516), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n524), .B1(new_n522), .B2(new_n523), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n530), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(KEYINPUT117), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT117), .ZN(new_n794));
  OAI211_X1 g593(.A(new_n794), .B(new_n530), .C1(new_n790), .C2(new_n791), .ZN(new_n795));
  AND3_X1   g594(.A1(new_n793), .A2(new_n534), .A3(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n582), .A2(new_n796), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n651), .B1(new_n789), .B2(new_n797), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n785), .A2(new_n796), .A3(new_n787), .A4(new_n788), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n799), .A2(new_n607), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n773), .B1(new_n798), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n706), .A2(new_n583), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  AND2_X1   g602(.A1(new_n803), .A2(new_n458), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n714), .A2(new_n404), .ZN(new_n805));
  AND2_X1   g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(new_n540), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n772), .B1(new_n807), .B2(G113gat), .ZN(new_n808));
  INV_X1    g607(.A(G113gat), .ZN(new_n809));
  AOI211_X1 g608(.A(KEYINPUT118), .B(new_n809), .C1(new_n806), .C2(new_n540), .ZN(new_n810));
  NOR3_X1   g609(.A1(new_n705), .A2(new_n535), .A3(new_n582), .ZN(new_n811));
  AND2_X1   g610(.A1(new_n788), .A2(new_n787), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n651), .A2(new_n796), .A3(new_n812), .A4(new_n785), .ZN(new_n813));
  AND2_X1   g612(.A1(new_n789), .A2(new_n797), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n813), .B1(new_n814), .B2(new_n651), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n811), .B1(new_n815), .B2(new_n773), .ZN(new_n816));
  NOR3_X1   g615(.A1(new_n816), .A2(new_n404), .A3(new_n471), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(new_n713), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n535), .A2(new_n809), .ZN(new_n819));
  OAI22_X1  g618(.A1(new_n808), .A2(new_n810), .B1(new_n818), .B2(new_n819), .ZN(G1340gat));
  NAND3_X1  g619(.A1(new_n817), .A2(new_n582), .A3(new_n713), .ZN(new_n821));
  INV_X1    g620(.A(G120gat), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n583), .A2(new_n822), .ZN(new_n823));
  AOI22_X1  g622(.A1(new_n821), .A2(new_n822), .B1(new_n806), .B2(new_n823), .ZN(G1341gat));
  INV_X1    g623(.A(G127gat), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n825), .B1(new_n818), .B2(new_n773), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n773), .A2(new_n825), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n804), .A2(new_n805), .A3(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT119), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n806), .A2(KEYINPUT119), .A3(new_n827), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n826), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT120), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n826), .A2(new_n831), .A3(KEYINPUT120), .A4(new_n830), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(G1342gat));
  NOR3_X1   g635(.A1(new_n607), .A2(G134gat), .A3(new_n386), .ZN(new_n837));
  AND2_X1   g636(.A1(new_n817), .A2(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT56), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT121), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n838), .A2(KEYINPUT121), .A3(new_n839), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n806), .A2(new_n651), .ZN(new_n844));
  AOI21_X1  g643(.A(KEYINPUT56), .B1(new_n844), .B2(G134gat), .ZN(new_n845));
  OAI211_X1 g644(.A(new_n842), .B(new_n843), .C1(new_n845), .C2(new_n838), .ZN(G1343gat));
  NOR2_X1   g645(.A1(new_n816), .A2(new_n404), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n638), .A2(new_n467), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n539), .A2(G141gat), .ZN(new_n849));
  NAND4_X1  g648(.A1(new_n847), .A2(new_n713), .A3(new_n848), .A4(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n850), .B1(KEYINPUT123), .B2(KEYINPUT58), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT122), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT57), .ZN(new_n853));
  OAI211_X1 g652(.A(new_n852), .B(new_n853), .C1(new_n816), .C2(new_n467), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n467), .B1(new_n801), .B2(new_n802), .ZN(new_n855));
  OAI21_X1  g654(.A(KEYINPUT122), .B1(new_n855), .B2(KEYINPUT57), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n785), .A2(new_n787), .A3(new_n788), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n797), .B1(new_n539), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n800), .B1(new_n858), .B2(new_n607), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n802), .B1(new_n859), .B2(new_n621), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n467), .A2(new_n853), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n854), .A2(new_n856), .A3(new_n862), .ZN(new_n863));
  NOR3_X1   g662(.A1(new_n638), .A2(new_n404), .A3(new_n714), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n863), .A2(new_n535), .A3(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT58), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n866), .A2(new_n230), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n851), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n863), .A2(new_n540), .A3(new_n864), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(G141gat), .ZN(new_n870));
  OR2_X1    g669(.A1(new_n850), .A2(KEYINPUT123), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n868), .B1(new_n872), .B2(new_n866), .ZN(G1344gat));
  NOR2_X1   g672(.A1(new_n224), .A2(KEYINPUT59), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n863), .A2(new_n864), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n874), .B1(new_n875), .B2(new_n583), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n864), .A2(new_n582), .ZN(new_n877));
  OAI22_X1  g676(.A1(new_n859), .A2(new_n621), .B1(new_n540), .B2(new_n622), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(new_n380), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(new_n853), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n803), .A2(new_n861), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n877), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  OAI21_X1  g681(.A(KEYINPUT59), .B1(new_n882), .B2(new_n224), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n876), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n847), .A2(new_n848), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n885), .A2(new_n714), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n886), .A2(new_n224), .A3(new_n582), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n884), .A2(new_n887), .ZN(G1345gat));
  AOI21_X1  g687(.A(G155gat), .B1(new_n886), .B2(new_n621), .ZN(new_n889));
  INV_X1    g688(.A(new_n875), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n621), .A2(G155gat), .ZN(new_n891));
  XNOR2_X1  g690(.A(new_n891), .B(KEYINPUT124), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n889), .B1(new_n890), .B2(new_n892), .ZN(G1346gat));
  OAI21_X1  g692(.A(G162gat), .B1(new_n875), .B2(new_n607), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n651), .A2(new_n221), .A3(new_n461), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n894), .B1(new_n885), .B2(new_n895), .ZN(G1347gat));
  NOR2_X1   g695(.A1(new_n816), .A2(new_n672), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n714), .A2(new_n463), .ZN(new_n898));
  XOR2_X1   g697(.A(new_n898), .B(KEYINPUT125), .Z(new_n899));
  AND2_X1   g698(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g699(.A(G169gat), .B1(new_n900), .B2(new_n535), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n672), .A2(new_n461), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n804), .A2(new_n902), .ZN(new_n903));
  NOR3_X1   g702(.A1(new_n903), .A2(new_n283), .A3(new_n539), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n901), .A2(new_n904), .ZN(G1348gat));
  NAND3_X1  g704(.A1(new_n900), .A2(new_n284), .A3(new_n582), .ZN(new_n906));
  OAI21_X1  g705(.A(G176gat), .B1(new_n903), .B2(new_n583), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(G1349gat));
  NAND3_X1  g707(.A1(new_n900), .A2(new_n276), .A3(new_n621), .ZN(new_n909));
  OAI21_X1  g708(.A(G183gat), .B1(new_n903), .B2(new_n773), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  XNOR2_X1  g710(.A(new_n911), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g711(.A1(new_n900), .A2(new_n277), .A3(new_n651), .ZN(new_n913));
  OAI21_X1  g712(.A(G190gat), .B1(new_n903), .B2(new_n607), .ZN(new_n914));
  AND2_X1   g713(.A1(new_n914), .A2(KEYINPUT61), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n914), .A2(KEYINPUT61), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n913), .B1(new_n915), .B2(new_n916), .ZN(G1351gat));
  AND4_X1   g716(.A1(new_n404), .A2(new_n803), .A3(new_n714), .A4(new_n848), .ZN(new_n918));
  AOI21_X1  g717(.A(G197gat), .B1(new_n918), .B2(new_n535), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n880), .A2(new_n881), .ZN(new_n920));
  NOR3_X1   g719(.A1(new_n638), .A2(new_n672), .A3(new_n461), .ZN(new_n921));
  AND2_X1   g720(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  AND2_X1   g721(.A1(new_n540), .A2(G197gat), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n919), .B1(new_n922), .B2(new_n923), .ZN(G1352gat));
  INV_X1    g723(.A(G204gat), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n918), .A2(new_n925), .A3(new_n582), .ZN(new_n926));
  XOR2_X1   g725(.A(new_n926), .B(KEYINPUT62), .Z(new_n927));
  AND2_X1   g726(.A1(new_n922), .A2(new_n582), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n927), .B1(new_n928), .B2(new_n925), .ZN(G1353gat));
  NAND3_X1  g728(.A1(new_n918), .A2(new_n321), .A3(new_n621), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n920), .A2(new_n621), .A3(new_n921), .ZN(new_n931));
  AND3_X1   g730(.A1(new_n931), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n932));
  AOI21_X1  g731(.A(KEYINPUT63), .B1(new_n931), .B2(G211gat), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n930), .B1(new_n932), .B2(new_n933), .ZN(G1354gat));
  AOI21_X1  g733(.A(G218gat), .B1(new_n918), .B2(new_n651), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n607), .A2(new_n322), .ZN(new_n936));
  XNOR2_X1  g735(.A(new_n936), .B(KEYINPUT126), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n935), .B1(new_n922), .B2(new_n937), .ZN(G1355gat));
endmodule


