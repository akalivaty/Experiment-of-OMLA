//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 0 1 1 1 0 0 0 1 1 0 0 0 0 0 1 0 0 1 0 0 1 1 0 0 1 0 1 1 0 1 1 1 1 1 1 0 1 1 1 0 0 0 0 0 1 0 0 1 1 1 1 1 0 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:05 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n632, new_n633, new_n634, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n680, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n791, new_n792,
    new_n793, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n802, new_n803, new_n804, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n842, new_n843, new_n845, new_n846, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n861, new_n862, new_n863,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n894, new_n895,
    new_n896, new_n897, new_n899, new_n900, new_n901, new_n902, new_n904,
    new_n905;
  INV_X1    g000(.A(KEYINPUT76), .ZN(new_n202));
  INV_X1    g001(.A(G113gat), .ZN(new_n203));
  INV_X1    g002(.A(G120gat), .ZN(new_n204));
  AOI21_X1  g003(.A(KEYINPUT1), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n205), .B1(new_n203), .B2(new_n204), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT73), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  XOR2_X1   g007(.A(G127gat), .B(G134gat), .Z(new_n209));
  XNOR2_X1  g008(.A(new_n208), .B(new_n209), .ZN(new_n210));
  NOR2_X1   g009(.A1(G169gat), .A2(G176gat), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n211), .B(KEYINPUT26), .ZN(new_n212));
  NAND2_X1  g011(.A1(G169gat), .A2(G176gat), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT69), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND3_X1  g014(.A1(KEYINPUT69), .A2(G169gat), .A3(G176gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n212), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(G183gat), .A2(G190gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT28), .ZN(new_n221));
  NOR2_X1   g020(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n222));
  XNOR2_X1  g021(.A(KEYINPUT71), .B(G183gat), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n222), .B1(new_n223), .B2(KEYINPUT27), .ZN(new_n224));
  XNOR2_X1  g023(.A(KEYINPUT72), .B(G190gat), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n221), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(new_n225), .ZN(new_n227));
  XNOR2_X1  g026(.A(KEYINPUT27), .B(G183gat), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n227), .A2(KEYINPUT28), .A3(new_n228), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n220), .B1(new_n226), .B2(new_n229), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n225), .A2(new_n223), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n219), .A2(KEYINPUT24), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT24), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n233), .A2(G183gat), .A3(G190gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n231), .A2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT68), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n238), .B1(new_n211), .B2(KEYINPUT23), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT23), .ZN(new_n240));
  OAI211_X1 g039(.A(new_n240), .B(KEYINPUT68), .C1(G169gat), .C2(G176gat), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n217), .A2(new_n239), .A3(new_n241), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n240), .A2(G176gat), .ZN(new_n243));
  INV_X1    g042(.A(G169gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(KEYINPUT25), .ZN(new_n246));
  NOR3_X1   g045(.A1(new_n237), .A2(new_n242), .A3(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT25), .ZN(new_n248));
  OAI21_X1  g047(.A(KEYINPUT65), .B1(G183gat), .B2(G190gat), .ZN(new_n249));
  OR3_X1    g048(.A1(KEYINPUT65), .A2(G183gat), .A3(G190gat), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n235), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n211), .A2(KEYINPUT23), .ZN(new_n252));
  AOI22_X1  g051(.A1(new_n252), .A2(KEYINPUT68), .B1(new_n215), .B2(new_n216), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n251), .A2(new_n253), .A3(new_n239), .ZN(new_n254));
  XNOR2_X1  g053(.A(KEYINPUT66), .B(G169gat), .ZN(new_n255));
  AOI21_X1  g054(.A(KEYINPUT67), .B1(new_n255), .B2(new_n243), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n244), .A2(KEYINPUT66), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT66), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n258), .A2(G169gat), .ZN(new_n259));
  AND4_X1   g058(.A1(KEYINPUT67), .A2(new_n243), .A3(new_n257), .A4(new_n259), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n256), .A2(new_n260), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n248), .B1(new_n254), .B2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT70), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n247), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n243), .A2(new_n257), .A3(new_n259), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT67), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n255), .A2(KEYINPUT67), .A3(new_n243), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  AND3_X1   g068(.A1(new_n217), .A2(new_n239), .A3(new_n241), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n269), .A2(new_n270), .A3(new_n251), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n271), .A2(KEYINPUT70), .A3(new_n248), .ZN(new_n272));
  AOI211_X1 g071(.A(new_n210), .B(new_n230), .C1(new_n264), .C2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(new_n210), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n262), .A2(new_n263), .ZN(new_n275));
  INV_X1    g074(.A(new_n247), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n275), .A2(new_n272), .A3(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(new_n230), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n274), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n273), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(G227gat), .A2(G233gat), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n281), .B(KEYINPUT64), .ZN(new_n282));
  AOI21_X1  g081(.A(KEYINPUT74), .B1(new_n280), .B2(new_n282), .ZN(new_n283));
  AND3_X1   g082(.A1(new_n271), .A2(KEYINPUT70), .A3(new_n248), .ZN(new_n284));
  AOI21_X1  g083(.A(KEYINPUT70), .B1(new_n271), .B2(new_n248), .ZN(new_n285));
  NOR3_X1   g084(.A1(new_n284), .A2(new_n285), .A3(new_n247), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n210), .B1(new_n286), .B2(new_n230), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n277), .A2(new_n274), .A3(new_n278), .ZN(new_n288));
  NAND4_X1  g087(.A1(new_n287), .A2(KEYINPUT74), .A3(new_n282), .A4(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  OAI21_X1  g089(.A(KEYINPUT32), .B1(new_n283), .B2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT33), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n292), .B1(new_n283), .B2(new_n290), .ZN(new_n293));
  XOR2_X1   g092(.A(G15gat), .B(G43gat), .Z(new_n294));
  XNOR2_X1  g093(.A(G71gat), .B(G99gat), .ZN(new_n295));
  XNOR2_X1  g094(.A(new_n294), .B(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n291), .A2(new_n293), .A3(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT32), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n287), .A2(new_n282), .A3(new_n288), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT74), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n298), .B1(new_n301), .B2(new_n289), .ZN(new_n302));
  AOI21_X1  g101(.A(KEYINPUT33), .B1(new_n301), .B2(new_n289), .ZN(new_n303));
  INV_X1    g102(.A(new_n296), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n302), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n297), .A2(new_n305), .ZN(new_n306));
  OR3_X1    g105(.A1(new_n280), .A2(KEYINPUT34), .A3(new_n282), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n287), .A2(new_n288), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(new_n281), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(KEYINPUT34), .ZN(new_n310));
  AND2_X1   g109(.A1(new_n307), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n202), .B1(new_n306), .B2(new_n312), .ZN(new_n313));
  AOI211_X1 g112(.A(KEYINPUT76), .B(new_n311), .C1(new_n297), .C2(new_n305), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n297), .A2(new_n305), .A3(new_n311), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(KEYINPUT75), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT75), .ZN(new_n318));
  NAND4_X1  g117(.A1(new_n297), .A2(new_n305), .A3(new_n318), .A4(new_n311), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  OAI21_X1  g119(.A(KEYINPUT86), .B1(new_n315), .B2(new_n320), .ZN(new_n321));
  NOR3_X1   g120(.A1(new_n302), .A2(new_n303), .A3(new_n304), .ZN(new_n322));
  AOI221_X4 g121(.A(new_n298), .B1(KEYINPUT33), .B2(new_n296), .C1(new_n301), .C2(new_n289), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n312), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(KEYINPUT76), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n306), .A2(new_n202), .A3(new_n312), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  AND2_X1   g126(.A1(new_n317), .A2(new_n319), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT86), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n327), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT35), .ZN(new_n331));
  NAND2_X1  g130(.A1(G228gat), .A2(G233gat), .ZN(new_n332));
  XNOR2_X1  g131(.A(G197gat), .B(G204gat), .ZN(new_n333));
  INV_X1    g132(.A(G211gat), .ZN(new_n334));
  INV_X1    g133(.A(G218gat), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n333), .B1(KEYINPUT22), .B2(new_n336), .ZN(new_n337));
  XNOR2_X1  g136(.A(G211gat), .B(G218gat), .ZN(new_n338));
  XNOR2_X1  g137(.A(new_n337), .B(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  XOR2_X1   g139(.A(G155gat), .B(G162gat), .Z(new_n341));
  XNOR2_X1  g140(.A(G141gat), .B(G148gat), .ZN(new_n342));
  XNOR2_X1  g141(.A(KEYINPUT77), .B(KEYINPUT2), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n341), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT78), .ZN(new_n345));
  XNOR2_X1  g144(.A(new_n344), .B(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT3), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n341), .A2(new_n342), .ZN(new_n348));
  INV_X1    g147(.A(G155gat), .ZN(new_n349));
  INV_X1    g148(.A(G162gat), .ZN(new_n350));
  OAI21_X1  g149(.A(KEYINPUT2), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n348), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n346), .A2(new_n347), .A3(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT29), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n340), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT82), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n332), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n346), .A2(new_n352), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n347), .B1(new_n339), .B2(KEYINPUT29), .ZN(new_n359));
  AND2_X1   g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n355), .A2(new_n360), .ZN(new_n361));
  OR2_X1    g160(.A1(new_n357), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n357), .A2(new_n361), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  OR2_X1    g163(.A1(new_n364), .A2(G22gat), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(G22gat), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  XNOR2_X1  g166(.A(G78gat), .B(G106gat), .ZN(new_n368));
  XNOR2_X1  g167(.A(KEYINPUT31), .B(G50gat), .ZN(new_n369));
  XNOR2_X1  g168(.A(new_n368), .B(new_n369), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n364), .A2(G22gat), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n370), .B1(new_n371), .B2(KEYINPUT83), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n367), .A2(new_n372), .ZN(new_n373));
  NAND4_X1  g172(.A1(new_n365), .A2(KEYINPUT83), .A3(new_n366), .A4(new_n370), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n277), .A2(new_n278), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(new_n354), .ZN(new_n377));
  NAND2_X1  g176(.A1(G226gat), .A2(G233gat), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n376), .A2(G226gat), .A3(G233gat), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n379), .A2(new_n340), .A3(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  XNOR2_X1  g181(.A(G8gat), .B(G36gat), .ZN(new_n383));
  XNOR2_X1  g182(.A(G64gat), .B(G92gat), .ZN(new_n384));
  XOR2_X1   g183(.A(new_n383), .B(new_n384), .Z(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n340), .B1(new_n379), .B2(new_n380), .ZN(new_n387));
  OR4_X1    g186(.A1(KEYINPUT30), .A2(new_n382), .A3(new_n386), .A4(new_n387), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n386), .B1(new_n382), .B2(new_n387), .ZN(new_n389));
  INV_X1    g188(.A(new_n387), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n390), .A2(new_n385), .A3(new_n381), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n389), .A2(new_n391), .A3(KEYINPUT30), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n388), .A2(new_n392), .ZN(new_n393));
  XOR2_X1   g192(.A(G1gat), .B(G29gat), .Z(new_n394));
  XNOR2_X1  g193(.A(new_n394), .B(KEYINPUT0), .ZN(new_n395));
  XNOR2_X1  g194(.A(G57gat), .B(G85gat), .ZN(new_n396));
  XNOR2_X1  g195(.A(new_n395), .B(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n210), .A2(new_n346), .A3(new_n352), .ZN(new_n398));
  OR2_X1    g197(.A1(new_n398), .A2(KEYINPUT4), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(KEYINPUT4), .ZN(new_n400));
  AOI21_X1  g199(.A(KEYINPUT5), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT81), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n210), .B1(new_n358), .B2(KEYINPUT3), .ZN(new_n403));
  AOI22_X1  g202(.A1(new_n403), .A2(new_n353), .B1(G225gat), .B2(G233gat), .ZN(new_n404));
  AND3_X1   g203(.A1(new_n401), .A2(new_n402), .A3(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n402), .B1(new_n401), .B2(new_n404), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n399), .A2(KEYINPUT79), .ZN(new_n408));
  OR3_X1    g207(.A1(new_n398), .A2(KEYINPUT79), .A3(KEYINPUT4), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n408), .A2(new_n409), .A3(new_n400), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(new_n404), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT80), .ZN(new_n412));
  NAND2_X1  g211(.A1(G225gat), .A2(G233gat), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n358), .A2(new_n274), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n413), .B1(new_n414), .B2(new_n398), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT5), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n412), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  OR3_X1    g216(.A1(new_n415), .A2(new_n412), .A3(new_n416), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n411), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n397), .B1(new_n407), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(KEYINPUT6), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n407), .A2(new_n419), .A3(new_n397), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT6), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  XNOR2_X1  g223(.A(new_n397), .B(KEYINPUT84), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n426), .B1(new_n407), .B2(new_n419), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n421), .B1(new_n424), .B2(new_n427), .ZN(new_n428));
  AND4_X1   g227(.A1(new_n331), .A2(new_n375), .A3(new_n393), .A4(new_n428), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n321), .A2(new_n330), .A3(new_n429), .ZN(new_n430));
  AND2_X1   g229(.A1(new_n324), .A2(new_n316), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n421), .B1(new_n424), .B2(new_n420), .ZN(new_n432));
  NAND4_X1  g231(.A1(new_n431), .A2(new_n432), .A3(new_n393), .A4(new_n375), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(KEYINPUT35), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n430), .A2(new_n434), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n375), .B1(new_n432), .B2(new_n393), .ZN(new_n436));
  OAI211_X1 g235(.A(new_n421), .B(new_n391), .C1(new_n424), .C2(new_n427), .ZN(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT85), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n390), .A2(new_n439), .A3(new_n381), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(KEYINPUT37), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT38), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT37), .ZN(new_n443));
  NAND4_X1  g242(.A1(new_n390), .A2(new_n439), .A3(new_n443), .A4(new_n381), .ZN(new_n444));
  NAND4_X1  g243(.A1(new_n441), .A2(new_n442), .A3(new_n386), .A4(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n441), .A2(new_n386), .A3(new_n444), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(KEYINPUT38), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n438), .A2(new_n445), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n399), .A2(new_n400), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n403), .A2(new_n353), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n413), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT39), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n425), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n414), .A2(new_n398), .A3(new_n413), .ZN(new_n454));
  AOI22_X1  g253(.A1(new_n399), .A2(new_n400), .B1(new_n353), .B2(new_n403), .ZN(new_n455));
  OAI211_X1 g254(.A(KEYINPUT39), .B(new_n454), .C1(new_n455), .C2(new_n413), .ZN(new_n456));
  AND3_X1   g255(.A1(new_n453), .A2(KEYINPUT40), .A3(new_n456), .ZN(new_n457));
  AOI21_X1  g256(.A(KEYINPUT40), .B1(new_n453), .B2(new_n456), .ZN(new_n458));
  NOR3_X1   g257(.A1(new_n427), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n459), .A2(new_n392), .A3(new_n388), .ZN(new_n460));
  AND2_X1   g259(.A1(new_n460), .A2(new_n375), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n436), .B1(new_n448), .B2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT36), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n431), .A2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n327), .A2(new_n328), .ZN(new_n466));
  OAI211_X1 g265(.A(new_n462), .B(new_n465), .C1(KEYINPUT36), .C2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n435), .A2(new_n467), .ZN(new_n468));
  XNOR2_X1  g267(.A(G15gat), .B(G22gat), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT16), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n469), .B1(new_n470), .B2(G1gat), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n471), .B1(G1gat), .B2(new_n469), .ZN(new_n472));
  INV_X1    g271(.A(G8gat), .ZN(new_n473));
  XNOR2_X1  g272(.A(new_n472), .B(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  AND2_X1   g274(.A1(G71gat), .A2(G78gat), .ZN(new_n476));
  NOR2_X1   g275(.A1(G71gat), .A2(G78gat), .ZN(new_n477));
  XOR2_X1   g276(.A(G57gat), .B(G64gat), .Z(new_n478));
  AOI211_X1 g277(.A(new_n476), .B(new_n477), .C1(new_n478), .C2(KEYINPUT9), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n476), .B1(KEYINPUT9), .B2(new_n477), .ZN(new_n480));
  XNOR2_X1  g279(.A(KEYINPUT92), .B(G57gat), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(G64gat), .ZN(new_n482));
  INV_X1    g281(.A(G64gat), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(G57gat), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n480), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n479), .A2(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n475), .B1(KEYINPUT21), .B2(new_n486), .ZN(new_n487));
  XOR2_X1   g286(.A(KEYINPUT95), .B(KEYINPUT96), .Z(new_n488));
  XNOR2_X1  g287(.A(new_n487), .B(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(G231gat), .A2(G233gat), .ZN(new_n490));
  XNOR2_X1  g289(.A(new_n490), .B(KEYINPUT94), .ZN(new_n491));
  XOR2_X1   g290(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n492));
  XNOR2_X1  g291(.A(new_n491), .B(new_n492), .ZN(new_n493));
  XNOR2_X1  g292(.A(new_n489), .B(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(new_n486), .ZN(new_n495));
  XOR2_X1   g294(.A(KEYINPUT93), .B(KEYINPUT21), .Z(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  XOR2_X1   g296(.A(G127gat), .B(G155gat), .Z(new_n498));
  XNOR2_X1  g297(.A(new_n497), .B(new_n498), .ZN(new_n499));
  XNOR2_X1  g298(.A(G183gat), .B(G211gat), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n499), .B(new_n500), .ZN(new_n501));
  OR2_X1    g300(.A1(new_n494), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n494), .A2(new_n501), .ZN(new_n503));
  AND2_X1   g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(G232gat), .A2(G233gat), .ZN(new_n505));
  XOR2_X1   g304(.A(new_n505), .B(KEYINPUT97), .Z(new_n506));
  INV_X1    g305(.A(new_n506), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n507), .A2(KEYINPUT41), .ZN(new_n508));
  XNOR2_X1  g307(.A(G134gat), .B(G162gat), .ZN(new_n509));
  XOR2_X1   g308(.A(new_n508), .B(new_n509), .Z(new_n510));
  NAND2_X1  g309(.A1(G85gat), .A2(G92gat), .ZN(new_n511));
  NAND2_X1  g310(.A1(KEYINPUT98), .A2(KEYINPUT7), .ZN(new_n512));
  XOR2_X1   g311(.A(new_n511), .B(new_n512), .Z(new_n513));
  XOR2_X1   g312(.A(G99gat), .B(G106gat), .Z(new_n514));
  INV_X1    g313(.A(KEYINPUT99), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(G99gat), .A2(G106gat), .ZN(new_n517));
  INV_X1    g316(.A(G85gat), .ZN(new_n518));
  INV_X1    g317(.A(G92gat), .ZN(new_n519));
  AOI22_X1  g318(.A1(KEYINPUT8), .A2(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n513), .A2(new_n516), .A3(new_n520), .ZN(new_n521));
  OR2_X1    g320(.A1(new_n514), .A2(new_n515), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n521), .B(new_n522), .ZN(new_n523));
  XOR2_X1   g322(.A(G43gat), .B(G50gat), .Z(new_n524));
  INV_X1    g323(.A(KEYINPUT15), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT88), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n526), .B(new_n527), .ZN(new_n528));
  NOR2_X1   g327(.A1(G29gat), .A2(G36gat), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n529), .B(KEYINPUT14), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n524), .A2(new_n525), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n532), .B1(G29gat), .B2(G36gat), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n528), .A2(new_n531), .A3(new_n533), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n531), .A2(KEYINPUT87), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT87), .ZN(new_n536));
  INV_X1    g335(.A(G29gat), .ZN(new_n537));
  INV_X1    g336(.A(G36gat), .ZN(new_n538));
  OAI22_X1  g337(.A1(new_n530), .A2(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n532), .B1(new_n535), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n534), .A2(new_n540), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n541), .A2(KEYINPUT17), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT17), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n543), .B1(new_n534), .B2(new_n540), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n523), .B1(new_n542), .B2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(new_n523), .ZN(new_n546));
  AOI22_X1  g345(.A1(new_n541), .A2(new_n546), .B1(KEYINPUT41), .B2(new_n507), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(G190gat), .B(G218gat), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n548), .A2(new_n550), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n510), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT100), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  OAI211_X1 g355(.A(KEYINPUT100), .B(new_n510), .C1(new_n552), .C2(new_n553), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n552), .A2(KEYINPUT101), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT101), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n559), .B1(new_n549), .B2(new_n551), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n553), .A2(new_n510), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n558), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n556), .A2(new_n557), .A3(new_n562), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n504), .A2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n541), .B(new_n474), .ZN(new_n566));
  NAND2_X1  g365(.A1(G229gat), .A2(G233gat), .ZN(new_n567));
  XOR2_X1   g366(.A(new_n567), .B(KEYINPUT89), .Z(new_n568));
  XOR2_X1   g367(.A(new_n568), .B(KEYINPUT13), .Z(new_n569));
  OR2_X1    g368(.A1(new_n566), .A2(new_n569), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n474), .B1(new_n542), .B2(new_n544), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n541), .A2(new_n475), .ZN(new_n572));
  INV_X1    g371(.A(new_n568), .ZN(new_n573));
  NAND4_X1  g372(.A1(new_n571), .A2(KEYINPUT18), .A3(new_n572), .A4(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n570), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT90), .ZN(new_n577));
  AOI21_X1  g376(.A(KEYINPUT18), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n571), .A2(KEYINPUT90), .A3(new_n572), .A4(new_n573), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n575), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(G113gat), .B(G141gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(G197gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(KEYINPUT11), .B(G169gat), .ZN(new_n583));
  XOR2_X1   g382(.A(new_n582), .B(new_n583), .Z(new_n584));
  XOR2_X1   g383(.A(new_n584), .B(KEYINPUT12), .Z(new_n585));
  INV_X1    g384(.A(KEYINPUT91), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n585), .B1(new_n575), .B2(new_n586), .ZN(new_n587));
  AND2_X1   g386(.A1(new_n580), .A2(new_n587), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n580), .A2(new_n587), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n546), .A2(new_n486), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT10), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n523), .A2(new_n495), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n546), .A2(KEYINPUT10), .A3(new_n486), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(G230gat), .A2(G233gat), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n591), .A2(new_n593), .ZN(new_n599));
  INV_X1    g398(.A(new_n597), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(G120gat), .B(G148gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(G176gat), .B(G204gat), .ZN(new_n604));
  XOR2_X1   g403(.A(new_n603), .B(new_n604), .Z(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n602), .A2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n602), .A2(new_n606), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NOR3_X1   g409(.A1(new_n565), .A2(new_n590), .A3(new_n610), .ZN(new_n611));
  AND2_X1   g410(.A1(new_n468), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n432), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(G1gat), .ZN(G1324gat));
  INV_X1    g414(.A(new_n612), .ZN(new_n616));
  XNOR2_X1  g415(.A(KEYINPUT16), .B(G8gat), .ZN(new_n617));
  NOR3_X1   g416(.A1(new_n616), .A2(new_n393), .A3(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n393), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n473), .B1(new_n612), .B2(new_n619), .ZN(new_n620));
  OAI21_X1  g419(.A(KEYINPUT42), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n621), .B1(KEYINPUT42), .B2(new_n618), .ZN(G1325gat));
  NAND2_X1  g421(.A1(new_n321), .A2(new_n330), .ZN(new_n623));
  OR3_X1    g422(.A1(new_n616), .A2(G15gat), .A3(new_n623), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n465), .B1(new_n466), .B2(KEYINPUT36), .ZN(new_n625));
  OR2_X1    g424(.A1(new_n625), .A2(KEYINPUT102), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(KEYINPUT102), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  OAI21_X1  g428(.A(G15gat), .B1(new_n616), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n624), .A2(new_n630), .ZN(G1326gat));
  INV_X1    g430(.A(new_n375), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n612), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(KEYINPUT43), .B(G22gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n633), .B(new_n634), .ZN(G1327gat));
  INV_X1    g434(.A(new_n563), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n636), .B1(new_n435), .B2(new_n467), .ZN(new_n637));
  INV_X1    g436(.A(new_n504), .ZN(new_n638));
  NOR3_X1   g437(.A1(new_n638), .A2(new_n590), .A3(new_n610), .ZN(new_n639));
  AND2_X1   g438(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n640), .A2(new_n537), .A3(new_n613), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(KEYINPUT45), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n468), .A2(KEYINPUT103), .A3(new_n563), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT44), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n644), .A2(KEYINPUT103), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n645), .A2(KEYINPUT44), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n643), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n637), .A2(KEYINPUT103), .A3(KEYINPUT44), .ZN(new_n648));
  AND2_X1   g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  AND3_X1   g448(.A1(new_n649), .A2(new_n613), .A3(new_n639), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n642), .B1(new_n650), .B2(new_n537), .ZN(G1328gat));
  NAND3_X1  g450(.A1(new_n649), .A2(new_n619), .A3(new_n639), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n538), .B1(new_n652), .B2(KEYINPUT104), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n653), .B1(KEYINPUT104), .B2(new_n652), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n640), .A2(new_n538), .A3(new_n619), .ZN(new_n655));
  XOR2_X1   g454(.A(new_n655), .B(KEYINPUT46), .Z(new_n656));
  NAND2_X1  g455(.A1(new_n654), .A2(new_n656), .ZN(G1329gat));
  NAND3_X1  g456(.A1(new_n649), .A2(new_n625), .A3(new_n639), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n658), .A2(G43gat), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n623), .A2(G43gat), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n640), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n659), .A2(KEYINPUT47), .A3(new_n661), .ZN(new_n662));
  NAND4_X1  g461(.A1(new_n647), .A2(new_n628), .A3(new_n639), .A4(new_n648), .ZN(new_n663));
  AND3_X1   g462(.A1(new_n663), .A2(KEYINPUT105), .A3(G43gat), .ZN(new_n664));
  AOI21_X1  g463(.A(KEYINPUT105), .B1(new_n663), .B2(G43gat), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT106), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n661), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n640), .A2(KEYINPUT106), .A3(new_n660), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NOR3_X1   g468(.A1(new_n664), .A2(new_n665), .A3(new_n669), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n662), .B1(new_n670), .B2(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g470(.A1(new_n647), .A2(new_n632), .A3(new_n639), .A4(new_n648), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n672), .A2(G50gat), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n375), .A2(G50gat), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(KEYINPUT107), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n640), .A2(new_n675), .ZN(new_n676));
  AOI22_X1  g475(.A1(new_n673), .A2(new_n676), .B1(KEYINPUT108), .B2(KEYINPUT48), .ZN(new_n677));
  NOR2_X1   g476(.A1(KEYINPUT108), .A2(KEYINPUT48), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n677), .B(new_n678), .ZN(G1331gat));
  INV_X1    g478(.A(new_n590), .ZN(new_n680));
  INV_X1    g479(.A(new_n610), .ZN(new_n681));
  NOR3_X1   g480(.A1(new_n565), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n468), .A2(new_n682), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n683), .A2(new_n432), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(new_n481), .ZN(G1332gat));
  NOR2_X1   g484(.A1(new_n683), .A2(new_n393), .ZN(new_n686));
  NOR2_X1   g485(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n687));
  AND2_X1   g486(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n686), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n689), .B1(new_n686), .B2(new_n687), .ZN(G1333gat));
  INV_X1    g489(.A(new_n683), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n691), .A2(G71gat), .A3(new_n628), .ZN(new_n692));
  OAI21_X1  g491(.A(KEYINPUT109), .B1(new_n683), .B2(new_n623), .ZN(new_n693));
  INV_X1    g492(.A(G71gat), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NOR3_X1   g494(.A1(new_n683), .A2(KEYINPUT109), .A3(new_n623), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n692), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n697), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g497(.A1(new_n691), .A2(new_n632), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g499(.A1(new_n638), .A2(new_n680), .ZN(new_n701));
  INV_X1    g500(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n702), .A2(new_n681), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n647), .A2(new_n648), .A3(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT110), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND4_X1  g505(.A1(new_n647), .A2(KEYINPUT110), .A3(new_n648), .A4(new_n703), .ZN(new_n707));
  AND3_X1   g506(.A1(new_n706), .A2(new_n613), .A3(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT111), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n315), .A2(new_n320), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n464), .B1(new_n710), .B2(new_n463), .ZN(new_n711));
  AOI22_X1  g510(.A1(new_n434), .A2(new_n430), .B1(new_n711), .B2(new_n462), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n709), .B1(new_n712), .B2(new_n636), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n468), .A2(KEYINPUT111), .A3(new_n563), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n713), .A2(new_n714), .A3(new_n701), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT51), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n702), .B1(new_n637), .B2(KEYINPUT111), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n718), .A2(KEYINPUT51), .A3(new_n713), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n613), .A2(new_n518), .A3(new_n610), .ZN(new_n722));
  OAI22_X1  g521(.A1(new_n708), .A2(new_n518), .B1(new_n721), .B2(new_n722), .ZN(G1336gat));
  INV_X1    g522(.A(KEYINPUT52), .ZN(new_n724));
  OAI211_X1 g523(.A(new_n724), .B(G92gat), .C1(new_n704), .C2(new_n393), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n619), .A2(new_n519), .A3(new_n610), .ZN(new_n726));
  OAI221_X1 g525(.A(new_n725), .B1(KEYINPUT112), .B2(new_n724), .C1(new_n721), .C2(new_n726), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n706), .A2(new_n619), .A3(new_n707), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT112), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n726), .B1(new_n717), .B2(new_n719), .ZN(new_n730));
  AOI22_X1  g529(.A1(new_n728), .A2(G92gat), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n727), .B1(new_n731), .B2(new_n724), .ZN(G1337gat));
  NAND3_X1  g531(.A1(new_n706), .A2(new_n628), .A3(new_n707), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(G99gat), .ZN(new_n734));
  OR3_X1    g533(.A1(new_n623), .A2(G99gat), .A3(new_n681), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n734), .B1(new_n721), .B2(new_n735), .ZN(G1338gat));
  INV_X1    g535(.A(KEYINPUT113), .ZN(new_n737));
  NOR3_X1   g536(.A1(new_n375), .A2(G106gat), .A3(new_n681), .ZN(new_n738));
  AOI21_X1  g537(.A(KEYINPUT53), .B1(new_n720), .B2(new_n738), .ZN(new_n739));
  OAI21_X1  g538(.A(G106gat), .B1(new_n704), .B2(new_n375), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n737), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  AND4_X1   g540(.A1(KEYINPUT51), .A2(new_n713), .A3(new_n714), .A4(new_n701), .ZN(new_n742));
  AOI21_X1  g541(.A(KEYINPUT51), .B1(new_n718), .B2(new_n713), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n738), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT53), .ZN(new_n745));
  AND4_X1   g544(.A1(new_n737), .A2(new_n744), .A3(new_n745), .A4(new_n740), .ZN(new_n746));
  INV_X1    g545(.A(new_n738), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n747), .B1(new_n717), .B2(new_n719), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n706), .A2(new_n632), .A3(new_n707), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n748), .B1(new_n749), .B2(G106gat), .ZN(new_n750));
  OAI22_X1  g549(.A1(new_n741), .A2(new_n746), .B1(new_n750), .B2(new_n745), .ZN(G1339gat));
  INV_X1    g550(.A(KEYINPUT114), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n594), .A2(new_n595), .A3(new_n600), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n598), .A2(KEYINPUT54), .A3(new_n753), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n600), .B1(new_n594), .B2(new_n595), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT54), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n605), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n754), .A2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT55), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n752), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n754), .A2(new_n757), .A3(KEYINPUT114), .A4(KEYINPUT55), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n607), .B1(new_n759), .B2(new_n758), .ZN(new_n763));
  OAI211_X1 g562(.A(new_n762), .B(new_n763), .C1(new_n588), .C2(new_n589), .ZN(new_n764));
  INV_X1    g563(.A(new_n585), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n566), .A2(new_n569), .ZN(new_n766));
  AND2_X1   g565(.A1(new_n571), .A2(new_n572), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n766), .B1(new_n767), .B2(new_n573), .ZN(new_n768));
  AOI22_X1  g567(.A1(new_n580), .A2(new_n765), .B1(new_n584), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(new_n610), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n563), .B1(new_n764), .B2(new_n770), .ZN(new_n771));
  AND4_X1   g570(.A1(new_n563), .A2(new_n769), .A3(new_n762), .A4(new_n763), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n504), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n564), .A2(new_n590), .A3(new_n681), .ZN(new_n774));
  AND3_X1   g573(.A1(new_n773), .A2(KEYINPUT115), .A3(new_n774), .ZN(new_n775));
  AOI21_X1  g574(.A(KEYINPUT115), .B1(new_n773), .B2(new_n774), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n375), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n623), .B1(new_n777), .B2(KEYINPUT116), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n619), .A2(new_n432), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT116), .ZN(new_n780));
  OAI211_X1 g579(.A(new_n780), .B(new_n375), .C1(new_n775), .C2(new_n776), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n778), .A2(new_n779), .A3(new_n781), .ZN(new_n782));
  OAI21_X1  g581(.A(G113gat), .B1(new_n782), .B2(new_n590), .ZN(new_n783));
  OR2_X1    g582(.A1(new_n775), .A2(new_n776), .ZN(new_n784));
  AND2_X1   g583(.A1(new_n784), .A2(new_n779), .ZN(new_n785));
  AND2_X1   g584(.A1(new_n431), .A2(new_n375), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n680), .A2(new_n203), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n788), .B(KEYINPUT117), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n783), .B1(new_n787), .B2(new_n789), .ZN(G1340gat));
  OAI21_X1  g589(.A(G120gat), .B1(new_n782), .B2(new_n681), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n610), .A2(new_n204), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n791), .B1(new_n787), .B2(new_n792), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n793), .B(KEYINPUT118), .ZN(G1341gat));
  INV_X1    g593(.A(KEYINPUT119), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n638), .A2(G127gat), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n795), .B1(new_n782), .B2(new_n796), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n787), .A2(new_n504), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n797), .B1(new_n798), .B2(G127gat), .ZN(new_n799));
  NOR3_X1   g598(.A1(new_n782), .A2(new_n795), .A3(new_n796), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n799), .A2(new_n800), .ZN(G1342gat));
  NOR3_X1   g600(.A1(new_n787), .A2(G134gat), .A3(new_n636), .ZN(new_n802));
  XNOR2_X1  g601(.A(new_n802), .B(KEYINPUT56), .ZN(new_n803));
  OAI21_X1  g602(.A(G134gat), .B1(new_n782), .B2(new_n636), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(G1343gat));
  NOR2_X1   g604(.A1(new_n628), .A2(new_n375), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n785), .A2(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(G141gat), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n808), .A2(new_n809), .A3(new_n680), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n711), .A2(new_n779), .ZN(new_n811));
  INV_X1    g610(.A(new_n811), .ZN(new_n812));
  XOR2_X1   g611(.A(KEYINPUT120), .B(KEYINPUT57), .Z(new_n813));
  INV_X1    g612(.A(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n814), .B1(new_n784), .B2(new_n632), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n773), .A2(new_n774), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(new_n632), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT57), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n812), .B1(new_n815), .B2(new_n819), .ZN(new_n820));
  OAI21_X1  g619(.A(G141gat), .B1(new_n820), .B2(new_n590), .ZN(new_n821));
  NAND2_X1  g620(.A1(KEYINPUT121), .A2(KEYINPUT58), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n810), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  NOR2_X1   g622(.A1(KEYINPUT121), .A2(KEYINPUT58), .ZN(new_n824));
  INV_X1    g623(.A(new_n824), .ZN(new_n825));
  XNOR2_X1  g624(.A(new_n823), .B(new_n825), .ZN(G1344gat));
  INV_X1    g625(.A(G148gat), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n808), .A2(new_n827), .A3(new_n610), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n827), .A2(KEYINPUT59), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n829), .B1(new_n820), .B2(new_n681), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT122), .ZN(new_n831));
  XNOR2_X1  g630(.A(new_n830), .B(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT59), .ZN(new_n833));
  OAI211_X1 g632(.A(new_n632), .B(new_n814), .C1(new_n775), .C2(new_n776), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n817), .A2(new_n818), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n811), .A2(new_n681), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n833), .B1(new_n838), .B2(G148gat), .ZN(new_n839));
  XNOR2_X1  g638(.A(new_n839), .B(KEYINPUT123), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n828), .B1(new_n832), .B2(new_n840), .ZN(G1345gat));
  NAND3_X1  g640(.A1(new_n808), .A2(new_n349), .A3(new_n638), .ZN(new_n842));
  OAI21_X1  g641(.A(G155gat), .B1(new_n820), .B2(new_n504), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(G1346gat));
  AOI21_X1  g643(.A(G162gat), .B1(new_n808), .B2(new_n563), .ZN(new_n845));
  NOR3_X1   g644(.A1(new_n820), .A2(new_n350), .A3(new_n636), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n845), .A2(new_n846), .ZN(G1347gat));
  NOR2_X1   g646(.A1(new_n613), .A2(new_n393), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n784), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(new_n786), .ZN(new_n850));
  INV_X1    g649(.A(new_n850), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n851), .A2(new_n255), .A3(new_n680), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n777), .A2(KEYINPUT116), .ZN(new_n853));
  INV_X1    g652(.A(new_n623), .ZN(new_n854));
  NAND4_X1  g653(.A1(new_n853), .A2(new_n854), .A3(new_n781), .A4(new_n848), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(KEYINPUT124), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT124), .ZN(new_n857));
  NAND4_X1  g656(.A1(new_n778), .A2(new_n857), .A3(new_n781), .A4(new_n848), .ZN(new_n858));
  AND3_X1   g657(.A1(new_n856), .A2(new_n680), .A3(new_n858), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n852), .B1(new_n859), .B2(new_n244), .ZN(G1348gat));
  NAND3_X1  g659(.A1(new_n856), .A2(new_n610), .A3(new_n858), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(G176gat), .ZN(new_n862));
  OR2_X1    g661(.A1(new_n681), .A2(G176gat), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n862), .B1(new_n850), .B2(new_n863), .ZN(G1349gat));
  NAND3_X1  g663(.A1(new_n856), .A2(new_n638), .A3(new_n858), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(new_n223), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n638), .A2(new_n228), .ZN(new_n867));
  OAI21_X1  g666(.A(KEYINPUT125), .B1(new_n850), .B2(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT125), .ZN(new_n869));
  INV_X1    g668(.A(new_n867), .ZN(new_n870));
  NAND4_X1  g669(.A1(new_n849), .A2(new_n869), .A3(new_n786), .A4(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n868), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n866), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(KEYINPUT60), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT60), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n866), .A2(new_n875), .A3(new_n872), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n874), .A2(new_n876), .ZN(G1350gat));
  NAND3_X1  g676(.A1(new_n851), .A2(new_n227), .A3(new_n563), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n856), .A2(new_n563), .A3(new_n858), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT61), .ZN(new_n880));
  AND4_X1   g679(.A1(KEYINPUT126), .A2(new_n879), .A3(new_n880), .A4(G190gat), .ZN(new_n881));
  INV_X1    g680(.A(G190gat), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT126), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n882), .B1(new_n883), .B2(KEYINPUT61), .ZN(new_n884));
  AOI22_X1  g683(.A1(new_n879), .A2(new_n884), .B1(KEYINPUT126), .B2(new_n880), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n878), .B1(new_n881), .B2(new_n885), .ZN(G1351gat));
  NAND2_X1  g685(.A1(new_n849), .A2(new_n806), .ZN(new_n887));
  OR3_X1    g686(.A1(new_n887), .A2(G197gat), .A3(new_n590), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n836), .A2(new_n629), .A3(new_n848), .ZN(new_n889));
  OAI21_X1  g688(.A(KEYINPUT127), .B1(new_n889), .B2(new_n590), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(G197gat), .ZN(new_n891));
  NOR3_X1   g690(.A1(new_n889), .A2(KEYINPUT127), .A3(new_n590), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n888), .B1(new_n891), .B2(new_n892), .ZN(G1352gat));
  OR3_X1    g692(.A1(new_n887), .A2(G204gat), .A3(new_n681), .ZN(new_n894));
  OR2_X1    g693(.A1(new_n894), .A2(KEYINPUT62), .ZN(new_n895));
  OAI21_X1  g694(.A(G204gat), .B1(new_n889), .B2(new_n681), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n894), .A2(KEYINPUT62), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(G1353gat));
  OR2_X1    g697(.A1(new_n889), .A2(new_n504), .ZN(new_n899));
  AND3_X1   g698(.A1(new_n899), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n900));
  AOI21_X1  g699(.A(KEYINPUT63), .B1(new_n899), .B2(G211gat), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n638), .A2(new_n334), .ZN(new_n902));
  OAI22_X1  g701(.A1(new_n900), .A2(new_n901), .B1(new_n887), .B2(new_n902), .ZN(G1354gat));
  OAI21_X1  g702(.A(G218gat), .B1(new_n889), .B2(new_n636), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n563), .A2(new_n335), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n904), .B1(new_n887), .B2(new_n905), .ZN(G1355gat));
endmodule


