//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 0 1 1 0 0 0 0 1 1 1 0 0 1 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 1 1 0 1 0 0 1 1 1 1 0 0 1 0 1 0 0 1 0 1 0 0 0 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:35 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n536, new_n537, new_n538, new_n539, new_n540, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n550, new_n551,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n584, new_n585,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n602,
    new_n603, new_n606, new_n608, new_n609, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT64), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT65), .B(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT66), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(KEYINPUT67), .B(KEYINPUT2), .Z(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n455), .A2(G567), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT68), .ZN(new_n459));
  AOI21_X1  g034(.A(new_n459), .B1(G2106), .B2(new_n453), .ZN(G319));
  OR2_X1    g035(.A1(KEYINPUT70), .A2(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(KEYINPUT70), .A2(G2104), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n461), .A2(KEYINPUT3), .A3(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n463), .A2(KEYINPUT71), .A3(new_n465), .ZN(new_n466));
  AND2_X1   g041(.A1(KEYINPUT70), .A2(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(KEYINPUT70), .A2(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT71), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n469), .A2(new_n470), .A3(KEYINPUT3), .ZN(new_n471));
  AOI21_X1  g046(.A(G2105), .B1(new_n466), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G137), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n469), .A2(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G101), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(G125), .ZN(new_n477));
  INV_X1    g052(.A(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(KEYINPUT3), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n465), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(KEYINPUT69), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT69), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n465), .A2(new_n479), .A3(new_n482), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n477), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(G113), .A2(G2104), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(new_n486));
  OAI21_X1  g061(.A(G2105), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n476), .A2(new_n488), .ZN(G160));
  OAI21_X1  g064(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(G112), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n490), .B1(new_n491), .B2(G2105), .ZN(new_n492));
  INV_X1    g067(.A(G2105), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n493), .B1(new_n466), .B2(new_n471), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G124), .ZN(new_n495));
  XNOR2_X1  g070(.A(new_n495), .B(KEYINPUT72), .ZN(new_n496));
  AOI211_X1 g071(.A(new_n492), .B(new_n496), .C1(G136), .C2(new_n472), .ZN(G162));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n498), .A2(new_n493), .A3(G138), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n499), .B1(new_n481), .B2(new_n483), .ZN(new_n500));
  OAI21_X1  g075(.A(KEYINPUT71), .B1(new_n478), .B2(KEYINPUT3), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n501), .B1(new_n469), .B2(KEYINPUT3), .ZN(new_n502));
  NOR4_X1   g077(.A1(new_n467), .A2(new_n468), .A3(KEYINPUT71), .A4(new_n464), .ZN(new_n503));
  OAI211_X1 g078(.A(G138), .B(new_n493), .C1(new_n502), .C2(new_n503), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n500), .B1(new_n504), .B2(KEYINPUT4), .ZN(new_n505));
  OAI211_X1 g080(.A(G126), .B(G2105), .C1(new_n502), .C2(new_n503), .ZN(new_n506));
  OAI21_X1  g081(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n507));
  INV_X1    g082(.A(G114), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n507), .B1(new_n508), .B2(G2105), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n506), .A2(new_n510), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n505), .A2(new_n511), .ZN(G164));
  INV_X1    g087(.A(G50), .ZN(new_n513));
  AND2_X1   g088(.A1(KEYINPUT6), .A2(G651), .ZN(new_n514));
  NOR2_X1   g089(.A1(KEYINPUT6), .A2(G651), .ZN(new_n515));
  OR2_X1    g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G543), .ZN(new_n517));
  XNOR2_X1  g092(.A(KEYINPUT5), .B(G543), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(G88), .ZN(new_n520));
  OAI22_X1  g095(.A1(new_n513), .A2(new_n517), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n518), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n522));
  INV_X1    g097(.A(G651), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n521), .A2(new_n524), .ZN(G166));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  XNOR2_X1  g101(.A(new_n526), .B(KEYINPUT7), .ZN(new_n527));
  INV_X1    g102(.A(G51), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n527), .B1(new_n517), .B2(new_n528), .ZN(new_n529));
  XOR2_X1   g104(.A(KEYINPUT5), .B(G543), .Z(new_n530));
  NAND2_X1  g105(.A1(new_n516), .A2(G89), .ZN(new_n531));
  NAND2_X1  g106(.A1(G63), .A2(G651), .ZN(new_n532));
  AOI21_X1  g107(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  OR2_X1    g108(.A1(new_n529), .A2(new_n533), .ZN(G286));
  INV_X1    g109(.A(G286), .ZN(G168));
  INV_X1    g110(.A(G52), .ZN(new_n536));
  INV_X1    g111(.A(G90), .ZN(new_n537));
  OAI22_X1  g112(.A1(new_n536), .A2(new_n517), .B1(new_n519), .B2(new_n537), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n518), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n539), .A2(new_n523), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n538), .A2(new_n540), .ZN(G171));
  INV_X1    g116(.A(G43), .ZN(new_n542));
  INV_X1    g117(.A(G81), .ZN(new_n543));
  OAI22_X1  g118(.A1(new_n542), .A2(new_n517), .B1(new_n519), .B2(new_n543), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n518), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n545), .A2(new_n523), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(G153));
  NAND4_X1  g123(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g124(.A1(G1), .A2(G3), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT8), .ZN(new_n551));
  NAND4_X1  g126(.A1(G319), .A2(G483), .A3(G661), .A4(new_n551), .ZN(G188));
  NOR2_X1   g127(.A1(new_n514), .A2(new_n515), .ZN(new_n553));
  INV_X1    g128(.A(G543), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  AOI21_X1  g130(.A(KEYINPUT73), .B1(new_n555), .B2(G53), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT9), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n530), .A2(new_n553), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G91), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n518), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n561));
  OAI211_X1 g136(.A(new_n558), .B(new_n560), .C1(new_n523), .C2(new_n561), .ZN(new_n562));
  AND3_X1   g137(.A1(new_n555), .A2(KEYINPUT73), .A3(G53), .ZN(new_n563));
  NOR3_X1   g138(.A1(new_n563), .A2(new_n556), .A3(new_n557), .ZN(new_n564));
  NOR2_X1   g139(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(new_n565), .ZN(G299));
  INV_X1    g141(.A(G171), .ZN(G301));
  INV_X1    g142(.A(G166), .ZN(G303));
  NAND2_X1  g143(.A1(new_n559), .A2(G87), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n555), .A2(G49), .ZN(new_n570));
  INV_X1    g145(.A(G74), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n530), .A2(new_n571), .ZN(new_n572));
  AOI21_X1  g147(.A(KEYINPUT74), .B1(new_n572), .B2(G651), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT74), .ZN(new_n574));
  AOI211_X1 g149(.A(new_n574), .B(new_n523), .C1(new_n530), .C2(new_n571), .ZN(new_n575));
  OAI211_X1 g150(.A(new_n569), .B(new_n570), .C1(new_n573), .C2(new_n575), .ZN(G288));
  NAND2_X1  g151(.A1(new_n559), .A2(G86), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n555), .A2(G48), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n518), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n580), .A2(new_n523), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  XNOR2_X1  g157(.A(new_n582), .B(KEYINPUT75), .ZN(G305));
  AOI22_X1  g158(.A1(new_n559), .A2(G85), .B1(new_n555), .B2(G47), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n518), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n523), .B2(new_n585), .ZN(G290));
  INV_X1    g161(.A(G868), .ZN(new_n587));
  NOR2_X1   g162(.A1(G301), .A2(new_n587), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n518), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n589));
  INV_X1    g164(.A(G54), .ZN(new_n590));
  OAI22_X1  g165(.A1(new_n523), .A2(new_n589), .B1(new_n517), .B2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT76), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n591), .B(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n559), .A2(G92), .ZN(new_n594));
  XOR2_X1   g169(.A(new_n594), .B(KEYINPUT10), .Z(new_n595));
  AND2_X1   g170(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n596), .A2(KEYINPUT77), .ZN(new_n597));
  AND3_X1   g172(.A1(new_n593), .A2(KEYINPUT77), .A3(new_n595), .ZN(new_n598));
  OR2_X1    g173(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n588), .B1(new_n599), .B2(new_n587), .ZN(G284));
  AOI21_X1  g175(.A(new_n588), .B1(new_n599), .B2(new_n587), .ZN(G321));
  NAND2_X1  g176(.A1(G286), .A2(G868), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n602), .B(KEYINPUT78), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n603), .B1(G868), .B2(new_n565), .ZN(G297));
  OAI21_X1  g179(.A(new_n603), .B1(G868), .B2(new_n565), .ZN(G280));
  XNOR2_X1  g180(.A(KEYINPUT79), .B(G559), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n599), .B1(G860), .B2(new_n606), .ZN(G148));
  NAND2_X1  g182(.A1(new_n599), .A2(new_n606), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(G868), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(G868), .B2(new_n547), .ZN(G323));
  XNOR2_X1  g185(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g186(.A1(new_n481), .A2(new_n483), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(new_n474), .ZN(new_n613));
  XOR2_X1   g188(.A(new_n613), .B(KEYINPUT12), .Z(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT13), .ZN(new_n615));
  XOR2_X1   g190(.A(new_n615), .B(G2100), .Z(new_n616));
  NAND2_X1  g191(.A1(new_n472), .A2(G135), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n494), .A2(G123), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n493), .A2(G111), .ZN(new_n619));
  OAI21_X1  g194(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n620));
  OAI211_X1 g195(.A(new_n617), .B(new_n618), .C1(new_n619), .C2(new_n620), .ZN(new_n621));
  INV_X1    g196(.A(G2096), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n621), .B(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n616), .A2(new_n623), .ZN(G156));
  XOR2_X1   g199(.A(G2451), .B(G2454), .Z(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT16), .ZN(new_n626));
  XNOR2_X1  g201(.A(G1341), .B(G1348), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  INV_X1    g203(.A(KEYINPUT14), .ZN(new_n629));
  XNOR2_X1  g204(.A(G2427), .B(G2438), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2430), .ZN(new_n631));
  XNOR2_X1  g206(.A(KEYINPUT15), .B(G2435), .ZN(new_n632));
  AOI21_X1  g207(.A(new_n629), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n633), .B1(new_n632), .B2(new_n631), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n628), .B(new_n634), .Z(new_n635));
  XNOR2_X1  g210(.A(G2443), .B(G2446), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n637), .A2(G14), .ZN(new_n638));
  NOR2_X1   g213(.A1(new_n635), .A2(new_n636), .ZN(new_n639));
  NOR2_X1   g214(.A1(new_n638), .A2(new_n639), .ZN(G401));
  XNOR2_X1  g215(.A(G2067), .B(G2678), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT80), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT81), .ZN(new_n643));
  XOR2_X1   g218(.A(G2072), .B(G2078), .Z(new_n644));
  NAND2_X1  g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2084), .B(G2090), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n644), .B(KEYINPUT17), .ZN(new_n647));
  OAI211_X1 g222(.A(new_n645), .B(new_n646), .C1(new_n643), .C2(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(KEYINPUT82), .Z(new_n649));
  NOR3_X1   g224(.A1(new_n642), .A2(new_n644), .A3(new_n646), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n650), .B(KEYINPUT18), .Z(new_n651));
  INV_X1    g226(.A(new_n647), .ZN(new_n652));
  NOR2_X1   g227(.A1(new_n652), .A2(new_n646), .ZN(new_n653));
  AOI21_X1  g228(.A(new_n651), .B1(new_n643), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n649), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(new_n622), .ZN(new_n656));
  XNOR2_X1  g231(.A(KEYINPUT83), .B(G2100), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(G227));
  XNOR2_X1  g234(.A(G1956), .B(G2474), .ZN(new_n660));
  XNOR2_X1  g235(.A(G1961), .B(G1966), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G1971), .B(G1976), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT19), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n660), .A2(new_n661), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(new_n666));
  OAI21_X1  g241(.A(new_n662), .B1(new_n664), .B2(new_n666), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n664), .A2(KEYINPUT84), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n664), .A2(new_n665), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT20), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1991), .B(G1996), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1981), .B(G1986), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(G229));
  NOR2_X1   g253(.A1(G6), .A2(G16), .ZN(new_n679));
  INV_X1    g254(.A(G305), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n679), .B1(new_n680), .B2(G16), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT32), .B(G1981), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(G288), .ZN(new_n684));
  INV_X1    g259(.A(G16), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n686), .B1(new_n685), .B2(G23), .ZN(new_n687));
  XOR2_X1   g262(.A(KEYINPUT33), .B(G1976), .Z(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(new_n689));
  OR2_X1    g264(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n687), .A2(new_n689), .ZN(new_n691));
  NOR2_X1   g266(.A1(G166), .A2(new_n685), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n692), .B1(new_n685), .B2(G22), .ZN(new_n693));
  INV_X1    g268(.A(G1971), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  OR2_X1    g270(.A1(new_n693), .A2(new_n694), .ZN(new_n696));
  NAND4_X1  g271(.A1(new_n690), .A2(new_n691), .A3(new_n695), .A4(new_n696), .ZN(new_n697));
  OR3_X1    g272(.A1(new_n683), .A2(KEYINPUT34), .A3(new_n697), .ZN(new_n698));
  OAI21_X1  g273(.A(KEYINPUT34), .B1(new_n683), .B2(new_n697), .ZN(new_n699));
  NOR2_X1   g274(.A1(G25), .A2(G29), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n472), .A2(G131), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n494), .A2(G119), .ZN(new_n702));
  OR2_X1    g277(.A1(G95), .A2(G2105), .ZN(new_n703));
  OAI211_X1 g278(.A(new_n703), .B(G2104), .C1(G107), .C2(new_n493), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n701), .A2(new_n702), .A3(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n700), .B1(new_n706), .B2(G29), .ZN(new_n707));
  XOR2_X1   g282(.A(KEYINPUT35), .B(G1991), .Z(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT85), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n707), .A2(new_n709), .ZN(new_n711));
  MUX2_X1   g286(.A(G24), .B(G290), .S(G16), .Z(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(G1986), .ZN(new_n713));
  INV_X1    g288(.A(KEYINPUT86), .ZN(new_n714));
  AOI211_X1 g289(.A(new_n711), .B(new_n713), .C1(new_n714), .C2(KEYINPUT36), .ZN(new_n715));
  NAND4_X1  g290(.A1(new_n698), .A2(new_n699), .A3(new_n710), .A4(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(KEYINPUT36), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(KEYINPUT86), .ZN(new_n718));
  XOR2_X1   g293(.A(new_n716), .B(new_n718), .Z(new_n719));
  NAND2_X1  g294(.A1(new_n472), .A2(G141), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT91), .ZN(new_n721));
  AND2_X1   g296(.A1(new_n494), .A2(G129), .ZN(new_n722));
  NAND3_X1  g297(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT26), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n474), .A2(G105), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT92), .ZN(new_n726));
  NOR4_X1   g301(.A1(new_n721), .A2(new_n722), .A3(new_n724), .A4(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n727), .A2(G29), .ZN(new_n728));
  OAI211_X1 g303(.A(new_n728), .B(KEYINPUT93), .C1(G29), .C2(G32), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(KEYINPUT93), .B2(new_n728), .ZN(new_n730));
  XOR2_X1   g305(.A(KEYINPUT27), .B(G1996), .Z(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(KEYINPUT94), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n730), .B(new_n732), .ZN(new_n733));
  AOI22_X1  g308(.A1(new_n612), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n734), .A2(new_n493), .ZN(new_n735));
  OR2_X1    g310(.A1(new_n735), .A2(KEYINPUT90), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n735), .A2(KEYINPUT90), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n493), .A2(G103), .A3(G2104), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT25), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(new_n472), .B2(G139), .ZN(new_n740));
  NAND3_X1  g315(.A1(new_n736), .A2(new_n737), .A3(new_n740), .ZN(new_n741));
  MUX2_X1   g316(.A(G33), .B(new_n741), .S(G29), .Z(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(G2072), .Z(new_n743));
  INV_X1    g318(.A(G29), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n744), .A2(G27), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(G164), .B2(new_n744), .ZN(new_n746));
  INV_X1    g321(.A(G2078), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n746), .B(new_n747), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n733), .A2(new_n743), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n744), .A2(G35), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G162), .B2(new_n744), .ZN(new_n751));
  XOR2_X1   g326(.A(KEYINPUT29), .B(G2090), .Z(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n685), .A2(G20), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(KEYINPUT23), .Z(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(G299), .B2(G16), .ZN(new_n756));
  INV_X1    g331(.A(G1956), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n685), .A2(G19), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT88), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(new_n547), .B2(new_n685), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(G1341), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n685), .A2(G5), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(G171), .B2(new_n685), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(G1961), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n685), .A2(G21), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(G168), .B2(new_n685), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(G1966), .ZN(new_n768));
  NOR4_X1   g343(.A1(new_n758), .A2(new_n762), .A3(new_n765), .A4(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(G160), .A2(G29), .ZN(new_n770));
  INV_X1    g345(.A(G34), .ZN(new_n771));
  AOI21_X1  g346(.A(G29), .B1(new_n771), .B2(KEYINPUT24), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(KEYINPUT24), .B2(new_n771), .ZN(new_n773));
  AOI21_X1  g348(.A(G2084), .B1(new_n770), .B2(new_n773), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n770), .A2(G2084), .A3(new_n773), .ZN(new_n775));
  INV_X1    g350(.A(KEYINPUT95), .ZN(new_n776));
  XNOR2_X1  g351(.A(KEYINPUT30), .B(G28), .ZN(new_n777));
  OR2_X1    g352(.A1(KEYINPUT31), .A2(G11), .ZN(new_n778));
  NAND2_X1  g353(.A1(KEYINPUT31), .A2(G11), .ZN(new_n779));
  AOI22_X1  g354(.A1(new_n777), .A2(new_n744), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(new_n621), .B2(new_n744), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n775), .B1(new_n776), .B2(new_n781), .ZN(new_n782));
  AOI211_X1 g357(.A(new_n774), .B(new_n782), .C1(new_n776), .C2(new_n781), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n744), .A2(G26), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n784), .B(KEYINPUT28), .Z(new_n785));
  NAND2_X1  g360(.A1(new_n494), .A2(G128), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n472), .A2(G140), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n493), .A2(G116), .ZN(new_n788));
  OAI21_X1  g363(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n789));
  OAI211_X1 g364(.A(new_n786), .B(new_n787), .C1(new_n788), .C2(new_n789), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n785), .B1(new_n790), .B2(G29), .ZN(new_n791));
  XNOR2_X1  g366(.A(KEYINPUT89), .B(G2067), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  NAND4_X1  g368(.A1(new_n753), .A2(new_n769), .A3(new_n783), .A4(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(G4), .A2(G16), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT87), .ZN(new_n796));
  INV_X1    g371(.A(new_n599), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n796), .B1(new_n797), .B2(new_n685), .ZN(new_n798));
  INV_X1    g373(.A(G1348), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  OR3_X1    g375(.A1(new_n749), .A2(new_n794), .A3(new_n800), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n719), .A2(new_n801), .ZN(G311));
  INV_X1    g377(.A(G311), .ZN(G150));
  NAND2_X1  g378(.A1(new_n599), .A2(G559), .ZN(new_n804));
  XNOR2_X1  g379(.A(KEYINPUT96), .B(KEYINPUT38), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  AOI22_X1  g381(.A1(new_n559), .A2(G93), .B1(new_n555), .B2(G55), .ZN(new_n807));
  AOI22_X1  g382(.A1(new_n518), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n807), .B1(new_n523), .B2(new_n808), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n547), .B(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(new_n810), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n806), .B(new_n811), .ZN(new_n812));
  AND2_X1   g387(.A1(new_n812), .A2(KEYINPUT39), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n812), .A2(KEYINPUT39), .ZN(new_n814));
  NOR3_X1   g389(.A1(new_n813), .A2(new_n814), .A3(G860), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n809), .A2(G860), .ZN(new_n816));
  XOR2_X1   g391(.A(KEYINPUT97), .B(KEYINPUT37), .Z(new_n817));
  XOR2_X1   g392(.A(new_n816), .B(new_n817), .Z(new_n818));
  OR2_X1    g393(.A1(new_n815), .A2(new_n818), .ZN(G145));
  XNOR2_X1  g394(.A(G164), .B(new_n790), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(new_n741), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(new_n727), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n494), .A2(G130), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n493), .A2(G118), .ZN(new_n824));
  OAI21_X1  g399(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n823), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n826), .B1(G142), .B2(new_n472), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(new_n614), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(new_n705), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n822), .B(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(G160), .B(new_n621), .ZN(new_n831));
  XNOR2_X1  g406(.A(G162), .B(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  OR2_X1    g408(.A1(new_n822), .A2(KEYINPUT98), .ZN(new_n834));
  OR2_X1    g409(.A1(new_n822), .A2(new_n829), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n832), .B(KEYINPUT99), .Z(new_n836));
  NAND3_X1  g411(.A1(new_n822), .A2(KEYINPUT98), .A3(new_n829), .ZN(new_n837));
  NAND4_X1  g412(.A1(new_n834), .A2(new_n835), .A3(new_n836), .A4(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(G37), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n833), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT40), .ZN(G395));
  AOI21_X1  g416(.A(KEYINPUT103), .B1(new_n809), .B2(new_n587), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n608), .B(new_n810), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n596), .A2(new_n565), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n593), .A2(new_n595), .ZN(new_n845));
  NAND2_X1  g420(.A1(G299), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n847), .A2(KEYINPUT41), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT41), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n844), .A2(new_n846), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n843), .A2(new_n851), .ZN(new_n852));
  OR2_X1    g427(.A1(new_n852), .A2(KEYINPUT101), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(KEYINPUT101), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT100), .ZN(new_n855));
  OR3_X1    g430(.A1(new_n843), .A2(new_n855), .A3(new_n847), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n855), .B1(new_n843), .B2(new_n847), .ZN(new_n857));
  AOI22_X1  g432(.A1(new_n853), .A2(new_n854), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n680), .A2(new_n684), .ZN(new_n859));
  XOR2_X1   g434(.A(G166), .B(G290), .Z(new_n860));
  NAND2_X1  g435(.A1(G305), .A2(G288), .ZN(new_n861));
  AND3_X1   g436(.A1(new_n859), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n860), .B1(new_n859), .B2(new_n861), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  XOR2_X1   g439(.A(KEYINPUT102), .B(KEYINPUT42), .Z(new_n865));
  XOR2_X1   g440(.A(new_n864), .B(new_n865), .Z(new_n866));
  NAND2_X1  g441(.A1(new_n858), .A2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  OAI21_X1  g443(.A(G868), .B1(new_n858), .B2(new_n866), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n842), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n853), .A2(new_n854), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n856), .A2(new_n857), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n866), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n587), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n875), .A2(KEYINPUT103), .A3(new_n867), .ZN(new_n876));
  AND2_X1   g451(.A1(new_n870), .A2(new_n876), .ZN(G295));
  AND2_X1   g452(.A1(new_n870), .A2(new_n876), .ZN(G331));
  INV_X1    g453(.A(KEYINPUT44), .ZN(new_n879));
  XNOR2_X1  g454(.A(G286), .B(G171), .ZN(new_n880));
  OR2_X1    g455(.A1(new_n880), .A2(new_n810), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n810), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n851), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n881), .A2(new_n882), .A3(KEYINPUT104), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT104), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n880), .A2(new_n810), .A3(new_n886), .ZN(new_n887));
  AND2_X1   g462(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n884), .B1(new_n888), .B2(new_n847), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n864), .A2(KEYINPUT105), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT105), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n891), .B1(new_n862), .B2(new_n863), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n889), .A2(new_n890), .A3(new_n892), .ZN(new_n893));
  OAI211_X1 g468(.A(new_n884), .B(new_n864), .C1(new_n847), .C2(new_n888), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n893), .A2(new_n839), .A3(new_n894), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n895), .A2(KEYINPUT43), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n890), .A2(new_n892), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n883), .A2(new_n847), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT106), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n850), .A2(new_n899), .ZN(new_n900));
  NAND4_X1  g475(.A1(new_n844), .A2(new_n846), .A3(KEYINPUT106), .A4(new_n849), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n900), .A2(new_n848), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n888), .A2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT107), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n898), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n888), .A2(new_n902), .A3(KEYINPUT107), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n897), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n894), .A2(new_n839), .ZN(new_n908));
  OAI21_X1  g483(.A(KEYINPUT43), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n896), .B1(new_n909), .B2(KEYINPUT108), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT108), .ZN(new_n911));
  OAI211_X1 g486(.A(new_n911), .B(KEYINPUT43), .C1(new_n907), .C2(new_n908), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n879), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  OR3_X1    g488(.A1(new_n907), .A2(KEYINPUT43), .A3(new_n908), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n895), .A2(KEYINPUT43), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n914), .A2(new_n879), .A3(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  OAI21_X1  g492(.A(KEYINPUT109), .B1(new_n913), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n909), .A2(KEYINPUT108), .ZN(new_n919));
  INV_X1    g494(.A(new_n896), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n919), .A2(new_n912), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(KEYINPUT44), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT109), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n922), .A2(new_n923), .A3(new_n916), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n918), .A2(new_n924), .ZN(G397));
  XNOR2_X1  g500(.A(new_n565), .B(KEYINPUT57), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n509), .B1(new_n494), .B2(G126), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n498), .B1(new_n472), .B2(G138), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n927), .B1(new_n928), .B2(new_n500), .ZN(new_n929));
  INV_X1    g504(.A(G1384), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n929), .A2(KEYINPUT45), .A3(new_n930), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n930), .B1(new_n505), .B2(new_n511), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT45), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND4_X1  g509(.A1(new_n473), .A2(new_n487), .A3(G40), .A4(new_n475), .ZN(new_n935));
  INV_X1    g510(.A(new_n935), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n931), .A2(new_n934), .A3(new_n936), .ZN(new_n937));
  XOR2_X1   g512(.A(KEYINPUT56), .B(G2072), .Z(new_n938));
  OR2_X1    g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g514(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n940), .B1(new_n505), .B2(new_n511), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT114), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  OAI211_X1 g518(.A(KEYINPUT114), .B(new_n940), .C1(new_n505), .C2(new_n511), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n935), .B1(new_n932), .B2(KEYINPUT50), .ZN(new_n946));
  AOI211_X1 g521(.A(KEYINPUT117), .B(G1956), .C1(new_n945), .C2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT117), .ZN(new_n948));
  AOI21_X1  g523(.A(KEYINPUT114), .B1(new_n929), .B2(new_n940), .ZN(new_n949));
  INV_X1    g524(.A(new_n944), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n946), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n948), .B1(new_n951), .B2(new_n757), .ZN(new_n952));
  OAI211_X1 g527(.A(new_n926), .B(new_n939), .C1(new_n947), .C2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n951), .A2(new_n757), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(KEYINPUT117), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n951), .A2(new_n948), .A3(new_n757), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n926), .B1(new_n957), .B2(new_n939), .ZN(new_n958));
  AOI21_X1  g533(.A(KEYINPUT111), .B1(new_n929), .B2(new_n940), .ZN(new_n959));
  OAI211_X1 g534(.A(KEYINPUT111), .B(new_n940), .C1(new_n505), .C2(new_n511), .ZN(new_n960));
  INV_X1    g535(.A(new_n960), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n946), .B1(new_n959), .B2(new_n961), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n932), .A2(new_n935), .ZN(new_n963));
  INV_X1    g538(.A(G2067), .ZN(new_n964));
  AOI22_X1  g539(.A1(new_n962), .A2(new_n799), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n797), .A2(new_n965), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n953), .B1(new_n958), .B2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT61), .ZN(new_n968));
  INV_X1    g543(.A(new_n953), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n968), .B1(new_n958), .B2(new_n969), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n939), .B1(new_n947), .B2(new_n952), .ZN(new_n971));
  INV_X1    g546(.A(new_n926), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n973), .A2(KEYINPUT61), .A3(new_n953), .ZN(new_n974));
  XNOR2_X1  g549(.A(KEYINPUT58), .B(G1341), .ZN(new_n975));
  OAI22_X1  g550(.A1(new_n937), .A2(G1996), .B1(new_n963), .B2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT59), .ZN(new_n977));
  AND3_X1   g552(.A1(new_n976), .A2(new_n977), .A3(new_n547), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n977), .B1(new_n976), .B2(new_n547), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(new_n980), .ZN(new_n981));
  NAND4_X1  g556(.A1(new_n970), .A2(KEYINPUT118), .A3(new_n974), .A4(new_n981), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n965), .B1(new_n599), .B2(KEYINPUT60), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n599), .A2(KEYINPUT60), .ZN(new_n984));
  XNOR2_X1  g559(.A(new_n983), .B(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n982), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n973), .A2(new_n953), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n980), .B1(new_n987), .B2(new_n968), .ZN(new_n988));
  AOI21_X1  g563(.A(KEYINPUT118), .B1(new_n988), .B2(new_n974), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n967), .B1(new_n986), .B2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT53), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n991), .B1(new_n937), .B2(G2078), .ZN(new_n992));
  INV_X1    g567(.A(G1961), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n962), .A2(new_n993), .ZN(new_n994));
  AND2_X1   g569(.A1(new_n992), .A2(new_n994), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n931), .A2(KEYINPUT53), .A3(new_n747), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n934), .A2(new_n936), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n996), .B1(KEYINPUT122), .B2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT122), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n934), .A2(new_n999), .A3(new_n936), .ZN(new_n1000));
  AOI21_X1  g575(.A(KEYINPUT123), .B1(new_n998), .B2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n997), .A2(KEYINPUT122), .ZN(new_n1002));
  AND3_X1   g577(.A1(new_n931), .A2(KEYINPUT53), .A3(new_n747), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1002), .A2(new_n1003), .A3(new_n1000), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT123), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  OAI211_X1 g581(.A(G301), .B(new_n995), .C1(new_n1001), .C2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(KEYINPUT124), .ZN(new_n1008));
  XNOR2_X1  g583(.A(new_n1004), .B(new_n1005), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT124), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n1009), .A2(new_n1010), .A3(G301), .A4(new_n995), .ZN(new_n1011));
  OR3_X1    g586(.A1(new_n937), .A2(new_n991), .A3(G2078), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n995), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(G171), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1008), .A2(new_n1011), .A3(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT54), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(G286), .A2(G8), .ZN(new_n1018));
  XNOR2_X1  g593(.A(new_n1018), .B(KEYINPUT119), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(G1966), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n937), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(G2084), .ZN(new_n1023));
  OAI211_X1 g598(.A(new_n946), .B(new_n1023), .C1(new_n959), .C2(new_n961), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1020), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1025));
  XNOR2_X1  g600(.A(new_n1025), .B(KEYINPUT120), .ZN(new_n1026));
  INV_X1    g601(.A(G8), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1027), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT51), .ZN(new_n1029));
  OR3_X1    g604(.A1(new_n1028), .A2(new_n1029), .A3(new_n1019), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1029), .B1(new_n1028), .B2(new_n1019), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1026), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT121), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1026), .A2(KEYINPUT121), .A3(new_n1030), .A4(new_n1031), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n1012), .A2(G301), .A3(new_n992), .A4(new_n994), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(KEYINPUT54), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1009), .A2(new_n995), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1038), .B1(new_n1039), .B2(G171), .ZN(new_n1040));
  INV_X1    g615(.A(G1976), .ZN(new_n1041));
  OAI221_X1 g616(.A(G8), .B1(new_n1041), .B2(G288), .C1(new_n932), .C2(new_n935), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1042), .ZN(new_n1043));
  AOI21_X1  g618(.A(KEYINPUT52), .B1(G288), .B2(new_n1041), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT113), .ZN(new_n1045));
  XNOR2_X1  g620(.A(new_n1044), .B(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1043), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1042), .A2(KEYINPUT52), .ZN(new_n1048));
  OAI21_X1  g623(.A(G1981), .B1(new_n579), .B2(new_n581), .ZN(new_n1049));
  INV_X1    g624(.A(new_n581), .ZN(new_n1050));
  INV_X1    g625(.A(G1981), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1050), .A2(new_n1051), .A3(new_n577), .A4(new_n578), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1049), .A2(new_n1052), .ZN(new_n1053));
  XNOR2_X1  g628(.A(new_n1053), .B(KEYINPUT49), .ZN(new_n1054));
  INV_X1    g629(.A(new_n963), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1054), .A2(new_n1055), .A3(G8), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1047), .A2(new_n1048), .A3(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n937), .A2(new_n694), .ZN(new_n1058));
  INV_X1    g633(.A(G2090), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n945), .A2(new_n1059), .A3(new_n946), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(G8), .ZN(new_n1062));
  NAND2_X1  g637(.A1(G303), .A2(G8), .ZN(new_n1063));
  XNOR2_X1  g638(.A(new_n1063), .B(KEYINPUT55), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1057), .B1(new_n1062), .B2(new_n1064), .ZN(new_n1065));
  OAI211_X1 g640(.A(new_n946), .B(new_n1059), .C1(new_n959), .C2(new_n961), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1058), .A2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT112), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1058), .A2(KEYINPUT112), .A3(new_n1066), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1064), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1069), .A2(G8), .A3(new_n1070), .A4(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1065), .A2(new_n1072), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1040), .A2(new_n1073), .ZN(new_n1074));
  AND3_X1   g649(.A1(new_n1017), .A2(new_n1036), .A3(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n990), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1036), .A2(KEYINPUT62), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT62), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1034), .A2(new_n1078), .A3(new_n1035), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1073), .A2(new_n1014), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1077), .A2(new_n1079), .A3(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT116), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1028), .A2(G168), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1065), .A2(new_n1072), .A3(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT63), .ZN(new_n1086));
  AND3_X1   g661(.A1(new_n1085), .A2(KEYINPUT115), .A3(new_n1086), .ZN(new_n1087));
  AOI21_X1  g662(.A(KEYINPUT115), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1069), .A2(G8), .A3(new_n1070), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(new_n1064), .ZN(new_n1090));
  NOR3_X1   g665(.A1(new_n1083), .A2(new_n1086), .A3(new_n1057), .ZN(new_n1091));
  AND3_X1   g666(.A1(new_n1090), .A2(new_n1091), .A3(new_n1072), .ZN(new_n1092));
  NOR3_X1   g667(.A1(new_n1087), .A2(new_n1088), .A3(new_n1092), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1072), .A2(new_n1057), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1056), .A2(new_n1041), .A3(new_n684), .ZN(new_n1095));
  AOI211_X1 g670(.A(new_n1027), .B(new_n963), .C1(new_n1095), .C2(new_n1052), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1097), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1082), .B1(new_n1093), .B2(new_n1098), .ZN(new_n1099));
  OR2_X1    g674(.A1(new_n1088), .A2(new_n1092), .ZN(new_n1100));
  OAI211_X1 g675(.A(KEYINPUT116), .B(new_n1097), .C1(new_n1100), .C2(new_n1087), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1076), .A2(new_n1081), .A3(new_n1099), .A4(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(G1996), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n934), .A2(new_n935), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n727), .A2(new_n1103), .A3(new_n1104), .ZN(new_n1105));
  XNOR2_X1  g680(.A(new_n1105), .B(KEYINPUT110), .ZN(new_n1106));
  XNOR2_X1  g681(.A(new_n790), .B(new_n964), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1107), .B1(new_n727), .B2(new_n1103), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(new_n1104), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1106), .A2(new_n1109), .ZN(new_n1110));
  XNOR2_X1  g685(.A(new_n705), .B(new_n709), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1110), .B1(new_n1104), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1112), .ZN(new_n1113));
  XNOR2_X1  g688(.A(G290), .B(G1986), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1113), .B1(new_n1104), .B2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1102), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1104), .A2(new_n1103), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT46), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  XNOR2_X1  g694(.A(new_n1119), .B(KEYINPUT125), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n727), .A2(new_n1107), .ZN(new_n1121));
  AOI22_X1  g696(.A1(new_n1121), .A2(new_n1104), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1123));
  XNOR2_X1  g698(.A(new_n1123), .B(KEYINPUT47), .ZN(new_n1124));
  NOR3_X1   g699(.A1(new_n1110), .A2(new_n709), .A3(new_n705), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n790), .A2(G2067), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1104), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  NOR2_X1   g702(.A1(G290), .A2(G1986), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1104), .A2(new_n1128), .ZN(new_n1129));
  XOR2_X1   g704(.A(new_n1129), .B(KEYINPUT48), .Z(new_n1130));
  OAI211_X1 g705(.A(new_n1124), .B(new_n1127), .C1(new_n1113), .C2(new_n1130), .ZN(new_n1131));
  XOR2_X1   g706(.A(new_n1131), .B(KEYINPUT126), .Z(new_n1132));
  NAND2_X1  g707(.A1(new_n1116), .A2(new_n1132), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g708(.A(G319), .B1(new_n638), .B2(new_n639), .ZN(new_n1135));
  NOR2_X1   g709(.A1(G229), .A2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g710(.A1(new_n658), .A2(new_n1136), .ZN(new_n1137));
  XOR2_X1   g711(.A(new_n1137), .B(KEYINPUT127), .Z(new_n1138));
  NAND2_X1  g712(.A1(new_n914), .A2(new_n915), .ZN(new_n1139));
  NAND3_X1  g713(.A1(new_n1138), .A2(new_n840), .A3(new_n1139), .ZN(G225));
  INV_X1    g714(.A(G225), .ZN(G308));
endmodule


