//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 1 1 1 0 0 1 1 0 0 0 1 1 1 1 1 0 1 0 1 1 0 0 1 0 1 0 0 1 1 1 0 1 0 1 0 0 0 0 1 1 1 0 0 0 0 0 0 1 0 1 1 0 0 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n682, new_n683, new_n684, new_n685,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n724, new_n725, new_n726,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n781, new_n782, new_n783, new_n785, new_n786,
    new_n787, new_n788, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n846,
    new_n847, new_n848, new_n850, new_n851, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n861, new_n862, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n901, new_n902;
  XNOR2_X1  g000(.A(G197gat), .B(G204gat), .ZN(new_n202));
  INV_X1    g001(.A(G211gat), .ZN(new_n203));
  INV_X1    g002(.A(G218gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n202), .B1(KEYINPUT22), .B2(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(G211gat), .B(G218gat), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  OR2_X1    g008(.A1(new_n209), .A2(KEYINPUT74), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT29), .ZN(new_n211));
  OAI211_X1 g010(.A(new_n207), .B(new_n202), .C1(KEYINPUT22), .C2(new_n205), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n209), .A2(KEYINPUT74), .A3(new_n212), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n210), .A2(new_n211), .A3(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT3), .ZN(new_n215));
  XOR2_X1   g014(.A(G155gat), .B(G162gat), .Z(new_n216));
  XNOR2_X1  g015(.A(G141gat), .B(G148gat), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n216), .B1(KEYINPUT2), .B2(new_n217), .ZN(new_n218));
  XOR2_X1   g017(.A(G141gat), .B(G148gat), .Z(new_n219));
  XNOR2_X1  g018(.A(G155gat), .B(G162gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT2), .ZN(new_n222));
  XNOR2_X1  g021(.A(KEYINPUT80), .B(G162gat), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n222), .B1(new_n223), .B2(G155gat), .ZN(new_n224));
  OR2_X1    g023(.A1(new_n221), .A2(new_n224), .ZN(new_n225));
  AOI22_X1  g024(.A1(new_n214), .A2(new_n215), .B1(new_n218), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n213), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n218), .B1(new_n221), .B2(new_n224), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n211), .B1(new_n228), .B2(KEYINPUT3), .ZN(new_n229));
  AND2_X1   g028(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  OAI211_X1 g029(.A(G228gat), .B(G233gat), .C1(new_n226), .C2(new_n230), .ZN(new_n231));
  AOI21_X1  g030(.A(KEYINPUT29), .B1(new_n209), .B2(new_n212), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(new_n228), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT86), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n228), .A2(KEYINPUT3), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n233), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n227), .A2(new_n229), .ZN(new_n237));
  NAND2_X1  g036(.A1(G228gat), .A2(G233gat), .ZN(new_n238));
  OAI211_X1 g037(.A(KEYINPUT86), .B(new_n228), .C1(new_n232), .C2(KEYINPUT3), .ZN(new_n239));
  NAND4_X1  g038(.A1(new_n236), .A2(new_n237), .A3(new_n238), .A4(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n231), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(G22gat), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT85), .ZN(new_n243));
  INV_X1    g042(.A(G22gat), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n231), .A2(new_n244), .A3(new_n240), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n242), .A2(new_n243), .A3(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(G78gat), .ZN(new_n247));
  INV_X1    g046(.A(G78gat), .ZN(new_n248));
  NAND4_X1  g047(.A1(new_n242), .A2(new_n243), .A3(new_n248), .A4(new_n245), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(KEYINPUT31), .B(G50gat), .ZN(new_n251));
  INV_X1    g050(.A(G106gat), .ZN(new_n252));
  XNOR2_X1  g051(.A(new_n251), .B(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n250), .A2(new_n254), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n247), .A2(new_n249), .A3(new_n253), .ZN(new_n256));
  AND2_X1   g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  XOR2_X1   g056(.A(G113gat), .B(G120gat), .Z(new_n258));
  INV_X1    g057(.A(KEYINPUT1), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(G134gat), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(G127gat), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT70), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  OAI21_X1  g063(.A(KEYINPUT71), .B1(new_n261), .B2(G127gat), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT71), .ZN(new_n266));
  INV_X1    g065(.A(G127gat), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n266), .A2(new_n267), .A3(G134gat), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n261), .A2(KEYINPUT70), .A3(G127gat), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n264), .A2(new_n265), .A3(new_n268), .A4(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n260), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n267), .A2(G134gat), .ZN(new_n272));
  NAND4_X1  g071(.A1(new_n258), .A2(new_n259), .A3(new_n262), .A4(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n274), .B(new_n228), .ZN(new_n275));
  NAND2_X1  g074(.A1(G225gat), .A2(G233gat), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT81), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n225), .A2(new_n215), .A3(new_n218), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n281), .A2(new_n274), .A3(new_n235), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT4), .ZN(new_n283));
  OR3_X1    g082(.A1(new_n274), .A2(new_n228), .A3(new_n283), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n283), .B1(new_n274), .B2(new_n228), .ZN(new_n285));
  NAND4_X1  g084(.A1(new_n282), .A2(new_n284), .A3(new_n276), .A4(new_n285), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n275), .A2(KEYINPUT81), .A3(new_n277), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n280), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(KEYINPUT82), .B(KEYINPUT5), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  XNOR2_X1  g089(.A(G57gat), .B(G85gat), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n291), .B(KEYINPUT84), .ZN(new_n292));
  XOR2_X1   g091(.A(KEYINPUT83), .B(KEYINPUT0), .Z(new_n293));
  XNOR2_X1  g092(.A(new_n292), .B(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(G1gat), .B(G29gat), .ZN(new_n295));
  XNOR2_X1  g094(.A(new_n294), .B(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n286), .ZN(new_n297));
  OR2_X1    g096(.A1(new_n297), .A2(new_n289), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n290), .A2(new_n296), .A3(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT88), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n299), .B(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n290), .A2(new_n298), .ZN(new_n302));
  INV_X1    g101(.A(new_n296), .ZN(new_n303));
  AOI21_X1  g102(.A(KEYINPUT6), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(new_n299), .ZN(new_n305));
  AOI22_X1  g104(.A1(new_n301), .A2(new_n304), .B1(KEYINPUT6), .B2(new_n305), .ZN(new_n306));
  NOR3_X1   g105(.A1(new_n257), .A2(KEYINPUT35), .A3(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT75), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT69), .ZN(new_n309));
  NOR2_X1   g108(.A1(G169gat), .A2(G176gat), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT68), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT26), .ZN(new_n313));
  OAI21_X1  g112(.A(KEYINPUT68), .B1(G169gat), .B2(G176gat), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n312), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(G169gat), .A2(G176gat), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(new_n310), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n317), .B1(new_n318), .B2(KEYINPUT26), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n315), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(G183gat), .A2(G190gat), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n309), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n321), .ZN(new_n323));
  AOI211_X1 g122(.A(KEYINPUT69), .B(new_n323), .C1(new_n315), .C2(new_n319), .ZN(new_n324));
  XNOR2_X1  g123(.A(KEYINPUT27), .B(G183gat), .ZN(new_n325));
  INV_X1    g124(.A(new_n325), .ZN(new_n326));
  OAI21_X1  g125(.A(KEYINPUT28), .B1(new_n326), .B2(G190gat), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT28), .ZN(new_n328));
  INV_X1    g127(.A(G190gat), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n325), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n327), .A2(new_n330), .ZN(new_n331));
  NOR3_X1   g130(.A1(new_n322), .A2(new_n324), .A3(new_n331), .ZN(new_n332));
  OR2_X1    g131(.A1(KEYINPUT66), .A2(KEYINPUT23), .ZN(new_n333));
  NAND2_X1  g132(.A1(KEYINPUT66), .A2(KEYINPUT23), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n310), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT25), .ZN(new_n336));
  NOR3_X1   g135(.A1(new_n335), .A2(new_n336), .A3(new_n317), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n312), .A2(KEYINPUT23), .A3(new_n314), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT24), .ZN(new_n339));
  INV_X1    g138(.A(G183gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(G190gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n329), .A2(G183gat), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n339), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n321), .A2(KEYINPUT24), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AND3_X1   g144(.A1(new_n337), .A2(new_n338), .A3(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT65), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n347), .B1(new_n343), .B2(new_n344), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n323), .A2(new_n339), .ZN(new_n349));
  XNOR2_X1  g148(.A(G183gat), .B(G190gat), .ZN(new_n350));
  OAI211_X1 g149(.A(new_n349), .B(KEYINPUT65), .C1(new_n350), .C2(new_n339), .ZN(new_n351));
  INV_X1    g150(.A(G169gat), .ZN(new_n352));
  INV_X1    g151(.A(G176gat), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n352), .A2(new_n353), .A3(KEYINPUT23), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(new_n316), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n335), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n348), .A2(new_n351), .A3(new_n356), .ZN(new_n357));
  XOR2_X1   g156(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n346), .B1(new_n359), .B2(KEYINPUT67), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT67), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n357), .A2(new_n361), .A3(new_n358), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n332), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(G226gat), .A2(G233gat), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n308), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(new_n364), .ZN(new_n366));
  INV_X1    g165(.A(new_n362), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n361), .B1(new_n357), .B2(new_n358), .ZN(new_n368));
  NOR3_X1   g167(.A1(new_n367), .A2(new_n368), .A3(new_n346), .ZN(new_n369));
  OAI211_X1 g168(.A(KEYINPUT75), .B(new_n366), .C1(new_n369), .C2(new_n332), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n211), .B1(new_n369), .B2(new_n332), .ZN(new_n371));
  AOI22_X1  g170(.A1(new_n365), .A2(new_n370), .B1(new_n371), .B2(new_n364), .ZN(new_n372));
  INV_X1    g171(.A(new_n227), .ZN(new_n373));
  OAI21_X1  g172(.A(KEYINPUT76), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n364), .B1(new_n363), .B2(KEYINPUT29), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n359), .A2(KEYINPUT67), .ZN(new_n376));
  INV_X1    g175(.A(new_n346), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n376), .A2(new_n362), .A3(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n332), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  AOI21_X1  g179(.A(KEYINPUT75), .B1(new_n380), .B2(new_n366), .ZN(new_n381));
  AOI211_X1 g180(.A(new_n308), .B(new_n364), .C1(new_n378), .C2(new_n379), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n375), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT76), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n383), .A2(new_n384), .A3(new_n227), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n363), .A2(new_n364), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n386), .B1(new_n364), .B2(new_n371), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(new_n373), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n374), .A2(new_n385), .A3(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(KEYINPUT77), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT77), .ZN(new_n391));
  NAND4_X1  g190(.A1(new_n374), .A2(new_n385), .A3(new_n388), .A4(new_n391), .ZN(new_n392));
  XNOR2_X1  g191(.A(G8gat), .B(G36gat), .ZN(new_n393));
  XNOR2_X1  g192(.A(G64gat), .B(G92gat), .ZN(new_n394));
  XOR2_X1   g193(.A(new_n393), .B(new_n394), .Z(new_n395));
  XOR2_X1   g194(.A(new_n395), .B(KEYINPUT78), .Z(new_n396));
  NAND3_X1  g195(.A1(new_n390), .A2(new_n392), .A3(new_n396), .ZN(new_n397));
  NAND4_X1  g196(.A1(new_n374), .A2(new_n385), .A3(new_n388), .A4(new_n395), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT30), .ZN(new_n399));
  OR2_X1    g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n398), .A2(new_n399), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n397), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  XNOR2_X1  g202(.A(G15gat), .B(G43gat), .ZN(new_n404));
  XNOR2_X1  g203(.A(new_n404), .B(KEYINPUT72), .ZN(new_n405));
  INV_X1    g204(.A(G71gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(new_n405), .B(new_n406), .ZN(new_n407));
  XNOR2_X1  g206(.A(new_n407), .B(G99gat), .ZN(new_n408));
  INV_X1    g207(.A(new_n274), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n380), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n363), .A2(new_n274), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n410), .A2(new_n411), .A3(G227gat), .A4(G233gat), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT33), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n408), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n412), .A2(KEYINPUT32), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  OAI211_X1 g215(.A(new_n412), .B(KEYINPUT32), .C1(new_n413), .C2(new_n408), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n410), .A2(new_n411), .ZN(new_n419));
  NAND2_X1  g218(.A1(G227gat), .A2(G233gat), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  OR2_X1    g220(.A1(new_n421), .A2(KEYINPUT34), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(KEYINPUT34), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n418), .A2(new_n424), .ZN(new_n425));
  OR2_X1    g224(.A1(new_n425), .A2(KEYINPUT73), .ZN(new_n426));
  NAND4_X1  g225(.A1(new_n416), .A2(new_n422), .A3(new_n423), .A4(new_n417), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n425), .A2(KEYINPUT73), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n307), .A2(new_n403), .A3(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT79), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n397), .A2(new_n431), .A3(new_n400), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n304), .A2(new_n299), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n305), .A2(KEYINPUT6), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  AND2_X1   g234(.A1(new_n435), .A2(new_n401), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n432), .A2(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n431), .B1(new_n397), .B2(new_n400), .ZN(new_n438));
  AND2_X1   g237(.A1(new_n425), .A2(new_n427), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n255), .A2(new_n256), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NOR3_X1   g240(.A1(new_n437), .A2(new_n438), .A3(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT35), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n430), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n257), .B1(new_n437), .B2(new_n438), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT36), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n439), .A2(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n448), .B1(new_n447), .B2(new_n429), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n389), .A2(KEYINPUT37), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n387), .A2(new_n227), .ZN(new_n452));
  OAI211_X1 g251(.A(new_n452), .B(KEYINPUT37), .C1(new_n227), .C2(new_n372), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT38), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n453), .A2(new_n454), .A3(new_n396), .ZN(new_n455));
  OAI211_X1 g254(.A(new_n306), .B(new_n398), .C1(new_n451), .C2(new_n455), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n451), .A2(new_n395), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n390), .A2(KEYINPUT37), .A3(new_n392), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n454), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  OR2_X1    g258(.A1(new_n456), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n282), .A2(new_n284), .A3(new_n285), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(new_n277), .ZN(new_n462));
  OAI211_X1 g261(.A(new_n462), .B(KEYINPUT39), .C1(new_n277), .C2(new_n275), .ZN(new_n463));
  OAI211_X1 g262(.A(new_n463), .B(new_n303), .C1(KEYINPUT39), .C2(new_n462), .ZN(new_n464));
  XNOR2_X1  g263(.A(new_n464), .B(KEYINPUT40), .ZN(new_n465));
  AND2_X1   g264(.A1(new_n301), .A2(new_n465), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n257), .B1(new_n402), .B2(new_n466), .ZN(new_n467));
  AOI22_X1  g266(.A1(new_n450), .A2(KEYINPUT87), .B1(new_n460), .B2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT87), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n446), .A2(new_n449), .A3(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n445), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT14), .ZN(new_n472));
  INV_X1    g271(.A(G29gat), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n475));
  AOI21_X1  g274(.A(G36gat), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(G36gat), .ZN(new_n477));
  NOR3_X1   g276(.A1(new_n472), .A2(new_n477), .A3(G29gat), .ZN(new_n478));
  OR3_X1    g277(.A1(new_n476), .A2(KEYINPUT15), .A3(new_n478), .ZN(new_n479));
  OAI21_X1  g278(.A(KEYINPUT15), .B1(new_n476), .B2(new_n478), .ZN(new_n480));
  XNOR2_X1  g279(.A(G43gat), .B(G50gat), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n479), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n482), .B1(new_n480), .B2(new_n481), .ZN(new_n483));
  XNOR2_X1  g282(.A(new_n483), .B(KEYINPUT17), .ZN(new_n484));
  XNOR2_X1  g283(.A(G15gat), .B(G22gat), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT16), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n485), .B1(new_n486), .B2(G1gat), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n487), .B1(G1gat), .B2(new_n485), .ZN(new_n488));
  INV_X1    g287(.A(G8gat), .ZN(new_n489));
  XNOR2_X1  g288(.A(new_n488), .B(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n484), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(G229gat), .A2(G233gat), .ZN(new_n492));
  XOR2_X1   g291(.A(new_n492), .B(KEYINPUT89), .Z(new_n493));
  INV_X1    g292(.A(new_n490), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(new_n483), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n491), .A2(new_n493), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(KEYINPUT90), .ZN(new_n497));
  OR2_X1    g296(.A1(new_n497), .A2(KEYINPUT18), .ZN(new_n498));
  XNOR2_X1  g297(.A(new_n483), .B(new_n490), .ZN(new_n499));
  XNOR2_X1  g298(.A(new_n493), .B(KEYINPUT13), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n501), .B1(new_n497), .B2(KEYINPUT18), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n498), .A2(new_n502), .ZN(new_n503));
  XNOR2_X1  g302(.A(G113gat), .B(G141gat), .ZN(new_n504));
  XNOR2_X1  g303(.A(new_n504), .B(G197gat), .ZN(new_n505));
  XOR2_X1   g304(.A(KEYINPUT11), .B(G169gat), .Z(new_n506));
  XNOR2_X1  g305(.A(new_n505), .B(new_n506), .ZN(new_n507));
  XOR2_X1   g306(.A(new_n507), .B(KEYINPUT12), .Z(new_n508));
  NAND2_X1  g307(.A1(new_n503), .A2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(new_n508), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n498), .A2(new_n510), .A3(new_n502), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(G71gat), .A2(G78gat), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n406), .A2(new_n248), .ZN(new_n515));
  XNOR2_X1  g314(.A(G57gat), .B(G64gat), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT9), .ZN(new_n517));
  OAI211_X1 g316(.A(new_n514), .B(new_n515), .C1(new_n516), .C2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT91), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n518), .B(new_n519), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n406), .A2(new_n248), .A3(KEYINPUT9), .ZN(new_n521));
  AOI22_X1  g320(.A1(new_n516), .A2(KEYINPUT92), .B1(new_n514), .B2(new_n521), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n522), .B1(KEYINPUT92), .B2(new_n516), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n520), .A2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT21), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n490), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  XOR2_X1   g325(.A(KEYINPUT94), .B(KEYINPUT20), .Z(new_n527));
  XNOR2_X1  g326(.A(new_n526), .B(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n524), .A2(new_n525), .ZN(new_n530));
  NAND2_X1  g329(.A1(G231gat), .A2(G233gat), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n530), .B(new_n531), .ZN(new_n532));
  XNOR2_X1  g331(.A(KEYINPUT93), .B(KEYINPUT19), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n532), .B(new_n533), .ZN(new_n534));
  XOR2_X1   g333(.A(G127gat), .B(G155gat), .Z(new_n535));
  XNOR2_X1  g334(.A(new_n534), .B(new_n535), .ZN(new_n536));
  XOR2_X1   g335(.A(G183gat), .B(G211gat), .Z(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n536), .A2(new_n538), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n529), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(new_n541), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n543), .A2(new_n539), .A3(new_n528), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  XOR2_X1   g344(.A(G134gat), .B(G162gat), .Z(new_n546));
  INV_X1    g345(.A(KEYINPUT8), .ZN(new_n547));
  NAND2_X1  g346(.A1(G99gat), .A2(G106gat), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n547), .B1(new_n548), .B2(KEYINPUT98), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT98), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n550), .A2(G99gat), .A3(G106gat), .ZN(new_n551));
  INV_X1    g350(.A(G85gat), .ZN(new_n552));
  INV_X1    g351(.A(G92gat), .ZN(new_n553));
  AOI22_X1  g352(.A1(new_n549), .A2(new_n551), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT7), .ZN(new_n555));
  OAI211_X1 g354(.A(KEYINPUT97), .B(new_n555), .C1(new_n552), .C2(new_n553), .ZN(new_n556));
  OAI21_X1  g355(.A(KEYINPUT97), .B1(new_n552), .B2(new_n553), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT97), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n558), .A2(G85gat), .A3(G92gat), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n557), .A2(new_n559), .A3(KEYINPUT7), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n554), .A2(new_n556), .A3(new_n560), .ZN(new_n561));
  XOR2_X1   g360(.A(G99gat), .B(G106gat), .Z(new_n562));
  XNOR2_X1  g361(.A(new_n561), .B(new_n562), .ZN(new_n563));
  XOR2_X1   g362(.A(new_n563), .B(KEYINPUT99), .Z(new_n564));
  NAND2_X1  g363(.A1(new_n564), .A2(new_n483), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n563), .B(KEYINPUT99), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n484), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(G232gat), .A2(G233gat), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n568), .B(KEYINPUT95), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n570), .A2(KEYINPUT41), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n565), .A2(new_n567), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(G190gat), .ZN(new_n573));
  NAND4_X1  g372(.A1(new_n565), .A2(new_n329), .A3(new_n567), .A4(new_n571), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(new_n204), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n573), .A2(G218gat), .A3(new_n574), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n576), .A2(KEYINPUT96), .A3(new_n577), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n570), .A2(KEYINPUT41), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n579), .ZN(new_n581));
  NAND4_X1  g380(.A1(new_n576), .A2(KEYINPUT96), .A3(new_n581), .A4(new_n577), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n546), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n580), .A2(new_n546), .A3(new_n582), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n524), .B(new_n563), .ZN(new_n586));
  OR2_X1    g385(.A1(new_n586), .A2(KEYINPUT10), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT100), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n520), .A2(KEYINPUT10), .A3(new_n523), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n564), .A2(new_n588), .A3(new_n590), .ZN(new_n591));
  OAI21_X1  g390(.A(KEYINPUT100), .B1(new_n566), .B2(new_n589), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n587), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(G230gat), .A2(G233gat), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n594), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n586), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(G120gat), .B(G148gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(G176gat), .B(G204gat), .ZN(new_n600));
  XOR2_X1   g399(.A(new_n599), .B(new_n600), .Z(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n598), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n595), .A2(new_n597), .A3(new_n601), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  NAND4_X1  g405(.A1(new_n545), .A2(new_n584), .A3(new_n585), .A4(new_n606), .ZN(new_n607));
  NOR3_X1   g406(.A1(new_n471), .A2(new_n513), .A3(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n435), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(KEYINPUT101), .B(G1gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n610), .B(new_n611), .ZN(G1324gat));
  NOR4_X1   g411(.A1(new_n471), .A2(new_n513), .A3(new_n403), .A4(new_n607), .ZN(new_n613));
  XOR2_X1   g412(.A(KEYINPUT16), .B(G8gat), .Z(new_n614));
  NAND3_X1  g413(.A1(new_n613), .A2(KEYINPUT42), .A3(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT103), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n615), .B(new_n616), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n613), .A2(new_n489), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n618), .B(KEYINPUT102), .ZN(new_n619));
  AND2_X1   g418(.A1(new_n613), .A2(new_n614), .ZN(new_n620));
  OR2_X1    g419(.A1(new_n620), .A2(KEYINPUT42), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n617), .A2(new_n619), .A3(new_n621), .ZN(G1325gat));
  INV_X1    g421(.A(new_n608), .ZN(new_n623));
  OAI21_X1  g422(.A(G15gat), .B1(new_n623), .B2(new_n449), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n471), .A2(new_n513), .ZN(new_n625));
  INV_X1    g424(.A(new_n429), .ZN(new_n626));
  NOR3_X1   g425(.A1(new_n607), .A2(G15gat), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n624), .A2(new_n628), .ZN(G1326gat));
  INV_X1    g428(.A(KEYINPUT104), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n630), .B1(new_n623), .B2(new_n440), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n608), .A2(KEYINPUT104), .A3(new_n257), .ZN(new_n632));
  XNOR2_X1  g431(.A(KEYINPUT43), .B(G22gat), .ZN(new_n633));
  AND3_X1   g432(.A1(new_n631), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n633), .B1(new_n631), .B2(new_n632), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n634), .A2(new_n635), .ZN(G1327gat));
  INV_X1    g435(.A(new_n585), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n637), .A2(new_n583), .ZN(new_n638));
  NOR3_X1   g437(.A1(new_n638), .A2(new_n545), .A3(new_n605), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n625), .A2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT45), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n609), .A2(new_n473), .ZN(new_n642));
  OR3_X1    g441(.A1(new_n640), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n402), .A2(new_n466), .ZN(new_n644));
  OAI211_X1 g443(.A(new_n644), .B(new_n440), .C1(new_n459), .C2(new_n456), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n645), .A2(new_n446), .A3(new_n449), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n444), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n584), .A2(new_n585), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT44), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n545), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n652), .A2(new_n512), .A3(new_n606), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(KEYINPUT105), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n648), .A2(KEYINPUT44), .ZN(new_n655));
  OAI211_X1 g454(.A(new_n651), .B(new_n654), .C1(new_n471), .C2(new_n655), .ZN(new_n656));
  OAI21_X1  g455(.A(G29gat), .B1(new_n656), .B2(new_n435), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n641), .B1(new_n640), .B2(new_n642), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n643), .A2(new_n657), .A3(new_n658), .ZN(G1328gat));
  NAND4_X1  g458(.A1(new_n625), .A2(new_n477), .A3(new_n402), .A4(new_n639), .ZN(new_n660));
  AND2_X1   g459(.A1(KEYINPUT106), .A2(KEYINPUT46), .ZN(new_n661));
  NOR2_X1   g460(.A1(KEYINPUT106), .A2(KEYINPUT46), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n660), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  OAI21_X1  g462(.A(G36gat), .B1(new_n656), .B2(new_n403), .ZN(new_n664));
  OAI211_X1 g463(.A(new_n663), .B(new_n664), .C1(new_n661), .C2(new_n660), .ZN(G1329gat));
  INV_X1    g464(.A(G43gat), .ZN(new_n666));
  NAND4_X1  g465(.A1(new_n625), .A2(new_n666), .A3(new_n429), .A4(new_n639), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n656), .A2(new_n449), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n667), .B1(new_n668), .B2(new_n666), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT47), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  OAI211_X1 g470(.A(KEYINPUT47), .B(new_n667), .C1(new_n668), .C2(new_n666), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(G1330gat));
  INV_X1    g472(.A(G50gat), .ZN(new_n674));
  NAND4_X1  g473(.A1(new_n625), .A2(new_n674), .A3(new_n257), .A4(new_n639), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n656), .A2(new_n440), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n675), .B1(new_n676), .B2(new_n674), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT48), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  OAI211_X1 g478(.A(KEYINPUT48), .B(new_n675), .C1(new_n676), .C2(new_n674), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(G1331gat));
  AND3_X1   g480(.A1(new_n545), .A2(new_n585), .A3(new_n584), .ZN(new_n682));
  AND4_X1   g481(.A1(new_n513), .A2(new_n647), .A3(new_n682), .A4(new_n605), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(new_n609), .ZN(new_n684));
  XNOR2_X1  g483(.A(KEYINPUT107), .B(G57gat), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n684), .B(new_n685), .ZN(G1332gat));
  NAND2_X1  g485(.A1(new_n683), .A2(new_n402), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n687), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n688));
  XOR2_X1   g487(.A(KEYINPUT49), .B(G64gat), .Z(new_n689));
  OAI21_X1  g488(.A(new_n688), .B1(new_n687), .B2(new_n689), .ZN(G1333gat));
  NAND3_X1  g489(.A1(new_n683), .A2(new_n406), .A3(new_n429), .ZN(new_n691));
  INV_X1    g490(.A(new_n449), .ZN(new_n692));
  AND2_X1   g491(.A1(new_n683), .A2(new_n692), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n691), .B1(new_n693), .B2(new_n406), .ZN(new_n694));
  XOR2_X1   g493(.A(new_n694), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g494(.A1(new_n683), .A2(new_n257), .ZN(new_n696));
  XNOR2_X1  g495(.A(KEYINPUT108), .B(G78gat), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n696), .B(new_n697), .ZN(G1335gat));
  INV_X1    g497(.A(KEYINPUT51), .ZN(new_n699));
  AOI211_X1 g498(.A(new_n512), .B(new_n545), .C1(KEYINPUT111), .C2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT110), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n701), .B1(new_n647), .B2(new_n648), .ZN(new_n702));
  AOI211_X1 g501(.A(KEYINPUT110), .B(new_n638), .C1(new_n444), .C2(new_n646), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n700), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n699), .A2(KEYINPUT111), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(new_n705), .ZN(new_n707));
  OAI211_X1 g506(.A(new_n707), .B(new_n700), .C1(new_n702), .C2(new_n703), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n609), .A2(new_n552), .A3(new_n605), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(KEYINPUT112), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n706), .A2(new_n708), .A3(new_n710), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n652), .A2(new_n513), .A3(new_n605), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  OAI211_X1 g512(.A(new_n651), .B(new_n713), .C1(new_n471), .C2(new_n655), .ZN(new_n714));
  OAI21_X1  g513(.A(KEYINPUT109), .B1(new_n714), .B2(new_n435), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(G85gat), .ZN(new_n716));
  NOR3_X1   g515(.A1(new_n714), .A2(KEYINPUT109), .A3(new_n435), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n711), .B1(new_n716), .B2(new_n717), .ZN(G1336gat));
  NOR3_X1   g517(.A1(new_n403), .A2(G92gat), .A3(new_n606), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n706), .A2(new_n708), .A3(new_n719), .ZN(new_n720));
  OAI21_X1  g519(.A(G92gat), .B1(new_n714), .B2(new_n403), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(KEYINPUT52), .ZN(G1337gat));
  NOR3_X1   g522(.A1(new_n626), .A2(G99gat), .A3(new_n606), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n706), .A2(new_n708), .A3(new_n724), .ZN(new_n725));
  OAI21_X1  g524(.A(G99gat), .B1(new_n714), .B2(new_n449), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(G1338gat));
  NAND2_X1  g526(.A1(new_n450), .A2(KEYINPUT87), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n728), .A2(new_n470), .A3(new_n645), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n655), .B1(new_n729), .B2(new_n444), .ZN(new_n730));
  AOI21_X1  g529(.A(KEYINPUT44), .B1(new_n647), .B2(new_n648), .ZN(new_n731));
  NOR4_X1   g530(.A1(new_n730), .A2(new_n731), .A3(new_n440), .A4(new_n712), .ZN(new_n732));
  XNOR2_X1  g531(.A(KEYINPUT113), .B(G106gat), .ZN(new_n733));
  OAI21_X1  g532(.A(KEYINPUT114), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NOR3_X1   g533(.A1(new_n440), .A2(new_n606), .A3(G106gat), .ZN(new_n735));
  NAND4_X1  g534(.A1(new_n706), .A2(KEYINPUT115), .A3(new_n708), .A4(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT114), .ZN(new_n737));
  INV_X1    g536(.A(new_n733), .ZN(new_n738));
  OAI211_X1 g537(.A(new_n737), .B(new_n738), .C1(new_n714), .C2(new_n440), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n734), .A2(new_n736), .A3(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(KEYINPUT53), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n706), .A2(new_n708), .A3(new_n735), .ZN(new_n742));
  NAND2_X1  g541(.A1(KEYINPUT115), .A2(KEYINPUT53), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n738), .B1(new_n714), .B2(new_n440), .ZN(new_n744));
  OAI211_X1 g543(.A(new_n742), .B(new_n743), .C1(new_n744), .C2(KEYINPUT53), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n741), .A2(new_n745), .ZN(G1339gat));
  AOI21_X1  g545(.A(new_n493), .B1(new_n491), .B2(new_n495), .ZN(new_n747));
  AND2_X1   g546(.A1(new_n499), .A2(new_n500), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n507), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  AND2_X1   g548(.A1(new_n511), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(new_n605), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT54), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n752), .B1(new_n593), .B2(new_n594), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n753), .B1(new_n594), .B2(new_n593), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n593), .A2(new_n752), .A3(new_n594), .ZN(new_n755));
  AND2_X1   g554(.A1(new_n755), .A2(new_n602), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT55), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(new_n512), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n754), .A2(new_n756), .A3(KEYINPUT55), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(new_n604), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n751), .B1(new_n760), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n638), .A2(new_n763), .ZN(new_n764));
  AND4_X1   g563(.A1(new_n604), .A2(new_n759), .A3(new_n750), .A4(new_n761), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n648), .A2(new_n765), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n545), .B1(new_n764), .B2(new_n766), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n607), .A2(new_n512), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n402), .A2(new_n435), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n626), .A2(new_n257), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n770), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  OAI21_X1  g572(.A(G113gat), .B1(new_n773), .B2(new_n513), .ZN(new_n774));
  NOR3_X1   g573(.A1(new_n769), .A2(new_n435), .A3(new_n402), .ZN(new_n775));
  INV_X1    g574(.A(new_n441), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n513), .A2(G113gat), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n778), .B(KEYINPUT116), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n774), .B1(new_n777), .B2(new_n779), .ZN(G1340gat));
  INV_X1    g579(.A(G120gat), .ZN(new_n781));
  NOR3_X1   g580(.A1(new_n773), .A2(new_n781), .A3(new_n606), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n775), .A2(new_n776), .A3(new_n605), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n782), .B1(new_n781), .B2(new_n783), .ZN(G1341gat));
  NOR3_X1   g583(.A1(new_n773), .A2(new_n267), .A3(new_n652), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n777), .A2(new_n652), .ZN(new_n786));
  OR2_X1    g585(.A1(new_n786), .A2(KEYINPUT117), .ZN(new_n787));
  AOI21_X1  g586(.A(G127gat), .B1(new_n786), .B2(KEYINPUT117), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n785), .B1(new_n787), .B2(new_n788), .ZN(G1342gat));
  NOR2_X1   g588(.A1(new_n638), .A2(G134gat), .ZN(new_n790));
  INV_X1    g589(.A(new_n790), .ZN(new_n791));
  OAI21_X1  g590(.A(KEYINPUT56), .B1(new_n777), .B2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT56), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n775), .A2(new_n793), .A3(new_n776), .A4(new_n790), .ZN(new_n794));
  OAI21_X1  g593(.A(G134gat), .B1(new_n773), .B2(new_n638), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n792), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(KEYINPUT118), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT118), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n792), .A2(new_n798), .A3(new_n794), .A4(new_n795), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n797), .A2(new_n799), .ZN(G1343gat));
  INV_X1    g599(.A(G141gat), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n449), .A2(new_n771), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT57), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n440), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n763), .A2(KEYINPUT119), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT119), .ZN(new_n806));
  OAI211_X1 g605(.A(new_n751), .B(new_n806), .C1(new_n760), .C2(new_n762), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n805), .A2(new_n638), .A3(new_n807), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n545), .B1(new_n808), .B2(new_n766), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT120), .ZN(new_n810));
  OAI22_X1  g609(.A1(new_n809), .A2(new_n810), .B1(new_n512), .B2(new_n607), .ZN(new_n811));
  AOI211_X1 g610(.A(KEYINPUT120), .B(new_n545), .C1(new_n808), .C2(new_n766), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n804), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n803), .B1(new_n769), .B2(new_n440), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n802), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n801), .B1(new_n815), .B2(new_n512), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n449), .A2(new_n257), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n817), .A2(KEYINPUT121), .ZN(new_n818));
  INV_X1    g617(.A(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n817), .A2(KEYINPUT121), .ZN(new_n820));
  AND3_X1   g619(.A1(new_n775), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n513), .A2(G141gat), .ZN(new_n822));
  AND2_X1   g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  OAI21_X1  g622(.A(KEYINPUT58), .B1(new_n816), .B2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT58), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n821), .A2(new_n822), .ZN(new_n826));
  AOI211_X1 g625(.A(new_n513), .B(new_n802), .C1(new_n813), .C2(new_n814), .ZN(new_n827));
  OAI211_X1 g626(.A(new_n825), .B(new_n826), .C1(new_n827), .C2(new_n801), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n824), .A2(new_n828), .ZN(G1344gat));
  INV_X1    g628(.A(G148gat), .ZN(new_n830));
  AND2_X1   g629(.A1(new_n821), .A2(new_n605), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT59), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n830), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT122), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n682), .A2(new_n834), .A3(new_n513), .A4(new_n606), .ZN(new_n835));
  OAI21_X1  g634(.A(KEYINPUT122), .B1(new_n607), .B2(new_n512), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n257), .B1(new_n837), .B2(new_n809), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(new_n803), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n770), .A2(new_n804), .ZN(new_n840));
  AND2_X1   g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n449), .A2(new_n605), .A3(new_n771), .ZN(new_n842));
  OAI211_X1 g641(.A(KEYINPUT59), .B(G148gat), .C1(new_n841), .C2(new_n842), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n815), .A2(new_n832), .A3(new_n605), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n833), .A2(new_n843), .A3(new_n844), .ZN(G1345gat));
  INV_X1    g644(.A(G155gat), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n821), .A2(new_n846), .A3(new_n545), .ZN(new_n847));
  AND2_X1   g646(.A1(new_n815), .A2(new_n545), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n847), .B1(new_n848), .B2(new_n846), .ZN(G1346gat));
  AOI21_X1  g648(.A(new_n223), .B1(new_n821), .B2(new_n648), .ZN(new_n850));
  AND2_X1   g649(.A1(new_n648), .A2(new_n223), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n850), .B1(new_n815), .B2(new_n851), .ZN(G1347gat));
  NOR2_X1   g651(.A1(new_n403), .A2(new_n609), .ZN(new_n853));
  OAI211_X1 g652(.A(new_n772), .B(new_n853), .C1(new_n767), .C2(new_n768), .ZN(new_n854));
  OAI21_X1  g653(.A(G169gat), .B1(new_n854), .B2(new_n513), .ZN(new_n855));
  XNOR2_X1  g654(.A(new_n855), .B(KEYINPUT123), .ZN(new_n856));
  OAI211_X1 g655(.A(new_n776), .B(new_n853), .C1(new_n767), .C2(new_n768), .ZN(new_n857));
  INV_X1    g656(.A(new_n857), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n858), .A2(new_n352), .A3(new_n512), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n856), .A2(new_n859), .ZN(G1348gat));
  OAI21_X1  g659(.A(G176gat), .B1(new_n854), .B2(new_n606), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n605), .A2(new_n353), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n861), .B1(new_n857), .B2(new_n862), .ZN(G1349gat));
  OAI21_X1  g662(.A(G183gat), .B1(new_n854), .B2(new_n652), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT124), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n545), .A2(new_n325), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n865), .B1(new_n857), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n864), .A2(new_n867), .ZN(new_n868));
  NOR3_X1   g667(.A1(new_n857), .A2(new_n865), .A3(new_n866), .ZN(new_n869));
  OAI22_X1  g668(.A1(new_n868), .A2(new_n869), .B1(KEYINPUT125), .B2(KEYINPUT60), .ZN(new_n870));
  NAND2_X1  g669(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n871));
  XNOR2_X1  g670(.A(new_n870), .B(new_n871), .ZN(G1350gat));
  NAND3_X1  g671(.A1(new_n858), .A2(new_n329), .A3(new_n648), .ZN(new_n873));
  OAI21_X1  g672(.A(G190gat), .B1(new_n854), .B2(new_n638), .ZN(new_n874));
  OR2_X1    g673(.A1(new_n874), .A2(KEYINPUT126), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT61), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n874), .A2(KEYINPUT126), .ZN(new_n877));
  AND3_X1   g676(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n876), .B1(new_n875), .B2(new_n877), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n873), .B1(new_n878), .B2(new_n879), .ZN(G1351gat));
  NAND2_X1  g679(.A1(new_n449), .A2(new_n853), .ZN(new_n881));
  NOR3_X1   g680(.A1(new_n769), .A2(new_n440), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(G197gat), .B1(new_n882), .B2(new_n512), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n881), .B1(new_n839), .B2(new_n840), .ZN(new_n884));
  AND2_X1   g683(.A1(new_n512), .A2(G197gat), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n883), .B1(new_n884), .B2(new_n885), .ZN(G1352gat));
  INV_X1    g685(.A(KEYINPUT127), .ZN(new_n887));
  AOI21_X1  g686(.A(G204gat), .B1(new_n887), .B2(KEYINPUT62), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n882), .A2(new_n605), .A3(new_n888), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n887), .A2(KEYINPUT62), .ZN(new_n890));
  XNOR2_X1  g689(.A(new_n889), .B(new_n890), .ZN(new_n891));
  AND2_X1   g690(.A1(new_n884), .A2(new_n605), .ZN(new_n892));
  INV_X1    g691(.A(G204gat), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n891), .B1(new_n892), .B2(new_n893), .ZN(G1353gat));
  NAND3_X1  g693(.A1(new_n882), .A2(new_n203), .A3(new_n545), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n884), .A2(new_n545), .ZN(new_n896));
  AOI21_X1  g695(.A(KEYINPUT63), .B1(new_n896), .B2(G211gat), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT63), .ZN(new_n898));
  AOI211_X1 g697(.A(new_n898), .B(new_n203), .C1(new_n884), .C2(new_n545), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n895), .B1(new_n897), .B2(new_n899), .ZN(G1354gat));
  NAND3_X1  g699(.A1(new_n882), .A2(new_n204), .A3(new_n648), .ZN(new_n901));
  AND2_X1   g700(.A1(new_n884), .A2(new_n648), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n901), .B1(new_n902), .B2(new_n204), .ZN(G1355gat));
endmodule


