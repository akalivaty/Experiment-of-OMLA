

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U557 ( .A(G2104), .ZN(n537) );
  NOR2_X1 U558 ( .A1(n702), .A2(G168), .ZN(n703) );
  BUF_X1 U559 ( .A(n577), .Z(n578) );
  AND2_X2 U560 ( .A1(n537), .A2(G2105), .ZN(n904) );
  AND2_X2 U561 ( .A1(G2105), .A2(G2104), .ZN(n905) );
  OR2_X2 U562 ( .A1(n605), .A2(n604), .ZN(n1018) );
  NOR2_X1 U563 ( .A1(n757), .A2(n762), .ZN(n699) );
  INV_X1 U564 ( .A(KEYINPUT14), .ZN(n599) );
  XNOR2_X1 U565 ( .A(n701), .B(KEYINPUT30), .ZN(n702) );
  XNOR2_X1 U566 ( .A(n542), .B(n541), .ZN(n577) );
  INV_X1 U567 ( .A(KEYINPUT66), .ZN(n540) );
  NAND2_X1 U568 ( .A1(n530), .A2(n603), .ZN(n604) );
  NOR2_X1 U569 ( .A1(G543), .A2(G651), .ZN(n652) );
  XOR2_X1 U570 ( .A(KEYINPUT68), .B(G651), .Z(n524) );
  AND2_X1 U571 ( .A1(n764), .A2(n533), .ZN(n525) );
  AND2_X1 U572 ( .A1(n529), .A2(n768), .ZN(n526) );
  NOR2_X1 U573 ( .A1(n838), .A2(n843), .ZN(n527) );
  OR2_X1 U574 ( .A1(n835), .A2(n826), .ZN(n528) );
  NOR2_X1 U575 ( .A1(n835), .A2(n767), .ZN(n529) );
  XOR2_X1 U576 ( .A(n602), .B(n601), .Z(n530) );
  AND2_X1 U577 ( .A1(n727), .A2(n726), .ZN(n531) );
  OR2_X1 U578 ( .A1(n834), .A2(n833), .ZN(n532) );
  XOR2_X1 U579 ( .A(n763), .B(KEYINPUT106), .Z(n533) );
  INV_X1 U580 ( .A(KEYINPUT109), .ZN(n768) );
  NOR2_X1 U581 ( .A1(n531), .A2(n733), .ZN(n734) );
  INV_X1 U582 ( .A(KEYINPUT107), .ZN(n746) );
  XNOR2_X1 U583 ( .A(n698), .B(n697), .ZN(n748) );
  BUF_X1 U584 ( .A(n748), .Z(n835) );
  NAND2_X1 U585 ( .A1(n666), .A2(G66), .ZN(n616) );
  XNOR2_X1 U586 ( .A(n600), .B(n599), .ZN(n601) );
  XNOR2_X1 U587 ( .A(n540), .B(KEYINPUT17), .ZN(n542) );
  AND2_X1 U588 ( .A1(n827), .A2(n528), .ZN(n828) );
  INV_X1 U589 ( .A(KEYINPUT1), .ZN(n550) );
  NOR2_X1 U590 ( .A1(n662), .A2(n524), .ZN(n653) );
  AND2_X1 U591 ( .A1(n845), .A2(n844), .ZN(n846) );
  XOR2_X1 U592 ( .A(n621), .B(KEYINPUT15), .Z(n917) );
  NOR2_X1 U593 ( .A1(G651), .A2(n662), .ZN(n667) );
  XNOR2_X1 U594 ( .A(n536), .B(KEYINPUT85), .ZN(n539) );
  NOR2_X1 U595 ( .A1(n545), .A2(n544), .ZN(G164) );
  NAND2_X1 U596 ( .A1(G126), .A2(n904), .ZN(n535) );
  NAND2_X1 U597 ( .A1(G114), .A2(n905), .ZN(n534) );
  NAND2_X1 U598 ( .A1(n535), .A2(n534), .ZN(n536) );
  NOR2_X4 U599 ( .A1(G2105), .A2(n537), .ZN(n901) );
  NAND2_X1 U600 ( .A1(G102), .A2(n901), .ZN(n538) );
  NAND2_X1 U601 ( .A1(n539), .A2(n538), .ZN(n545) );
  NOR2_X1 U602 ( .A1(G2105), .A2(G2104), .ZN(n541) );
  NAND2_X1 U603 ( .A1(n577), .A2(G138), .ZN(n543) );
  XOR2_X1 U604 ( .A(n543), .B(KEYINPUT86), .Z(n544) );
  NAND2_X1 U605 ( .A1(n652), .A2(G89), .ZN(n546) );
  XNOR2_X1 U606 ( .A(n546), .B(KEYINPUT4), .ZN(n548) );
  XOR2_X1 U607 ( .A(G543), .B(KEYINPUT0), .Z(n662) );
  NAND2_X1 U608 ( .A1(G76), .A2(n653), .ZN(n547) );
  NAND2_X1 U609 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U610 ( .A(n549), .B(KEYINPUT5), .ZN(n556) );
  NAND2_X1 U611 ( .A1(G51), .A2(n667), .ZN(n553) );
  NOR2_X1 U612 ( .A1(G543), .A2(n524), .ZN(n551) );
  XNOR2_X2 U613 ( .A(n551), .B(n550), .ZN(n666) );
  NAND2_X1 U614 ( .A1(G63), .A2(n666), .ZN(n552) );
  NAND2_X1 U615 ( .A1(n553), .A2(n552), .ZN(n554) );
  XOR2_X1 U616 ( .A(KEYINPUT6), .B(n554), .Z(n555) );
  NAND2_X1 U617 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U618 ( .A(n557), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U619 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U620 ( .A1(G137), .A2(n577), .ZN(n558) );
  XNOR2_X1 U621 ( .A(n558), .B(KEYINPUT67), .ZN(n566) );
  AND2_X1 U622 ( .A1(n904), .A2(G125), .ZN(n561) );
  NAND2_X1 U623 ( .A1(G113), .A2(n905), .ZN(n559) );
  XNOR2_X1 U624 ( .A(n559), .B(KEYINPUT65), .ZN(n560) );
  NOR2_X1 U625 ( .A1(n561), .A2(n560), .ZN(n564) );
  NAND2_X1 U626 ( .A1(G101), .A2(n901), .ZN(n562) );
  XOR2_X1 U627 ( .A(KEYINPUT23), .B(n562), .Z(n563) );
  NAND2_X1 U628 ( .A1(n564), .A2(n563), .ZN(n565) );
  NOR2_X2 U629 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X2 U630 ( .A(n567), .B(KEYINPUT64), .ZN(G160) );
  NAND2_X1 U631 ( .A1(n652), .A2(G91), .ZN(n569) );
  NAND2_X1 U632 ( .A1(G78), .A2(n653), .ZN(n568) );
  NAND2_X1 U633 ( .A1(n569), .A2(n568), .ZN(n573) );
  NAND2_X1 U634 ( .A1(G53), .A2(n667), .ZN(n571) );
  NAND2_X1 U635 ( .A1(G65), .A2(n666), .ZN(n570) );
  NAND2_X1 U636 ( .A1(n571), .A2(n570), .ZN(n572) );
  OR2_X1 U637 ( .A1(n573), .A2(n572), .ZN(G299) );
  AND2_X1 U638 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U639 ( .A1(n904), .A2(G123), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n574), .B(KEYINPUT18), .ZN(n576) );
  NAND2_X1 U641 ( .A1(G99), .A2(n901), .ZN(n575) );
  NAND2_X1 U642 ( .A1(n576), .A2(n575), .ZN(n582) );
  NAND2_X1 U643 ( .A1(G111), .A2(n905), .ZN(n580) );
  NAND2_X1 U644 ( .A1(G135), .A2(n578), .ZN(n579) );
  NAND2_X1 U645 ( .A1(n580), .A2(n579), .ZN(n581) );
  NOR2_X1 U646 ( .A1(n582), .A2(n581), .ZN(n992) );
  XNOR2_X1 U647 ( .A(n992), .B(G2096), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n583), .B(KEYINPUT79), .ZN(n584) );
  OR2_X1 U649 ( .A1(G2100), .A2(n584), .ZN(G156) );
  INV_X1 U650 ( .A(G57), .ZN(G237) );
  INV_X1 U651 ( .A(G132), .ZN(G219) );
  NAND2_X1 U652 ( .A1(n652), .A2(G88), .ZN(n586) );
  NAND2_X1 U653 ( .A1(G75), .A2(n653), .ZN(n585) );
  NAND2_X1 U654 ( .A1(n586), .A2(n585), .ZN(n591) );
  NAND2_X1 U655 ( .A1(G50), .A2(n667), .ZN(n588) );
  NAND2_X1 U656 ( .A1(G62), .A2(n666), .ZN(n587) );
  NAND2_X1 U657 ( .A1(n588), .A2(n587), .ZN(n589) );
  XOR2_X1 U658 ( .A(KEYINPUT83), .B(n589), .Z(n590) );
  NOR2_X1 U659 ( .A1(n591), .A2(n590), .ZN(G166) );
  NAND2_X1 U660 ( .A1(G7), .A2(G661), .ZN(n592) );
  XOR2_X1 U661 ( .A(n592), .B(KEYINPUT10), .Z(n850) );
  NAND2_X1 U662 ( .A1(n850), .A2(G567), .ZN(n593) );
  XOR2_X1 U663 ( .A(KEYINPUT11), .B(n593), .Z(G234) );
  NAND2_X1 U664 ( .A1(G68), .A2(n653), .ZN(n594) );
  XNOR2_X1 U665 ( .A(KEYINPUT75), .B(n594), .ZN(n597) );
  NAND2_X1 U666 ( .A1(n652), .A2(G81), .ZN(n595) );
  XOR2_X1 U667 ( .A(KEYINPUT12), .B(n595), .Z(n596) );
  NOR2_X1 U668 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X1 U669 ( .A(KEYINPUT13), .B(n598), .ZN(n605) );
  NAND2_X1 U670 ( .A1(G56), .A2(n666), .ZN(n602) );
  XOR2_X1 U671 ( .A(KEYINPUT74), .B(KEYINPUT73), .Z(n600) );
  NAND2_X1 U672 ( .A1(n667), .A2(G43), .ZN(n603) );
  INV_X1 U673 ( .A(G860), .ZN(n634) );
  OR2_X1 U674 ( .A1(n1018), .A2(n634), .ZN(G153) );
  NAND2_X1 U675 ( .A1(n666), .A2(G64), .ZN(n606) );
  XNOR2_X1 U676 ( .A(n606), .B(KEYINPUT71), .ZN(n613) );
  NAND2_X1 U677 ( .A1(n652), .A2(G90), .ZN(n608) );
  NAND2_X1 U678 ( .A1(G77), .A2(n653), .ZN(n607) );
  NAND2_X1 U679 ( .A1(n608), .A2(n607), .ZN(n609) );
  XNOR2_X1 U680 ( .A(n609), .B(KEYINPUT9), .ZN(n611) );
  NAND2_X1 U681 ( .A1(G52), .A2(n667), .ZN(n610) );
  NAND2_X1 U682 ( .A1(n611), .A2(n610), .ZN(n612) );
  NOR2_X1 U683 ( .A1(n613), .A2(n612), .ZN(G171) );
  INV_X1 U684 ( .A(G171), .ZN(G301) );
  NAND2_X1 U685 ( .A1(G868), .A2(G301), .ZN(n623) );
  NAND2_X1 U686 ( .A1(n667), .A2(G54), .ZN(n615) );
  NAND2_X1 U687 ( .A1(G79), .A2(n653), .ZN(n614) );
  NAND2_X1 U688 ( .A1(n615), .A2(n614), .ZN(n620) );
  NAND2_X1 U689 ( .A1(n652), .A2(G92), .ZN(n617) );
  NAND2_X1 U690 ( .A1(n617), .A2(n616), .ZN(n618) );
  XNOR2_X1 U691 ( .A(KEYINPUT76), .B(n618), .ZN(n619) );
  NOR2_X1 U692 ( .A1(n620), .A2(n619), .ZN(n621) );
  INV_X1 U693 ( .A(n917), .ZN(n1017) );
  INV_X1 U694 ( .A(G868), .ZN(n678) );
  NAND2_X1 U695 ( .A1(n1017), .A2(n678), .ZN(n622) );
  NAND2_X1 U696 ( .A1(n623), .A2(n622), .ZN(G284) );
  NOR2_X1 U697 ( .A1(G286), .A2(n678), .ZN(n625) );
  NOR2_X1 U698 ( .A1(G868), .A2(G299), .ZN(n624) );
  NOR2_X1 U699 ( .A1(n625), .A2(n624), .ZN(G297) );
  NAND2_X1 U700 ( .A1(G559), .A2(n634), .ZN(n626) );
  XOR2_X1 U701 ( .A(KEYINPUT77), .B(n626), .Z(n627) );
  NAND2_X1 U702 ( .A1(n627), .A2(n917), .ZN(n628) );
  XNOR2_X1 U703 ( .A(n628), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U704 ( .A1(G868), .A2(n1018), .ZN(n631) );
  NAND2_X1 U705 ( .A1(G868), .A2(n917), .ZN(n629) );
  NOR2_X1 U706 ( .A1(G559), .A2(n629), .ZN(n630) );
  NOR2_X1 U707 ( .A1(n631), .A2(n630), .ZN(n632) );
  XNOR2_X1 U708 ( .A(KEYINPUT78), .B(n632), .ZN(G282) );
  NAND2_X1 U709 ( .A1(G559), .A2(n917), .ZN(n633) );
  XOR2_X1 U710 ( .A(n1018), .B(n633), .Z(n675) );
  NAND2_X1 U711 ( .A1(n634), .A2(n675), .ZN(n642) );
  NAND2_X1 U712 ( .A1(G55), .A2(n667), .ZN(n636) );
  NAND2_X1 U713 ( .A1(G67), .A2(n666), .ZN(n635) );
  NAND2_X1 U714 ( .A1(n636), .A2(n635), .ZN(n637) );
  XNOR2_X1 U715 ( .A(KEYINPUT80), .B(n637), .ZN(n641) );
  NAND2_X1 U716 ( .A1(n652), .A2(G93), .ZN(n639) );
  NAND2_X1 U717 ( .A1(G80), .A2(n653), .ZN(n638) );
  NAND2_X1 U718 ( .A1(n639), .A2(n638), .ZN(n640) );
  NOR2_X1 U719 ( .A1(n641), .A2(n640), .ZN(n677) );
  XOR2_X1 U720 ( .A(n642), .B(n677), .Z(G145) );
  NAND2_X1 U721 ( .A1(G73), .A2(n653), .ZN(n644) );
  XNOR2_X1 U722 ( .A(KEYINPUT2), .B(KEYINPUT82), .ZN(n643) );
  XNOR2_X1 U723 ( .A(n644), .B(n643), .ZN(n651) );
  NAND2_X1 U724 ( .A1(G48), .A2(n667), .ZN(n646) );
  NAND2_X1 U725 ( .A1(G86), .A2(n652), .ZN(n645) );
  NAND2_X1 U726 ( .A1(n646), .A2(n645), .ZN(n649) );
  NAND2_X1 U727 ( .A1(G61), .A2(n666), .ZN(n647) );
  XNOR2_X1 U728 ( .A(KEYINPUT81), .B(n647), .ZN(n648) );
  NOR2_X1 U729 ( .A1(n649), .A2(n648), .ZN(n650) );
  NAND2_X1 U730 ( .A1(n651), .A2(n650), .ZN(G305) );
  NAND2_X1 U731 ( .A1(n652), .A2(G85), .ZN(n660) );
  NAND2_X1 U732 ( .A1(G72), .A2(n653), .ZN(n655) );
  NAND2_X1 U733 ( .A1(G60), .A2(n666), .ZN(n654) );
  NAND2_X1 U734 ( .A1(n655), .A2(n654), .ZN(n658) );
  NAND2_X1 U735 ( .A1(G47), .A2(n667), .ZN(n656) );
  XNOR2_X1 U736 ( .A(KEYINPUT69), .B(n656), .ZN(n657) );
  NOR2_X1 U737 ( .A1(n658), .A2(n657), .ZN(n659) );
  NAND2_X1 U738 ( .A1(n660), .A2(n659), .ZN(n661) );
  XNOR2_X1 U739 ( .A(n661), .B(KEYINPUT70), .ZN(G290) );
  INV_X1 U740 ( .A(G166), .ZN(G303) );
  NAND2_X1 U741 ( .A1(G87), .A2(n662), .ZN(n664) );
  NAND2_X1 U742 ( .A1(G74), .A2(G651), .ZN(n663) );
  NAND2_X1 U743 ( .A1(n664), .A2(n663), .ZN(n665) );
  NOR2_X1 U744 ( .A1(n666), .A2(n665), .ZN(n669) );
  NAND2_X1 U745 ( .A1(n667), .A2(G49), .ZN(n668) );
  NAND2_X1 U746 ( .A1(n669), .A2(n668), .ZN(G288) );
  XNOR2_X1 U747 ( .A(G305), .B(n677), .ZN(n671) );
  XOR2_X1 U748 ( .A(G290), .B(G303), .Z(n670) );
  XNOR2_X1 U749 ( .A(n671), .B(n670), .ZN(n674) );
  XOR2_X1 U750 ( .A(KEYINPUT19), .B(G299), .Z(n672) );
  XNOR2_X1 U751 ( .A(G288), .B(n672), .ZN(n673) );
  XNOR2_X1 U752 ( .A(n674), .B(n673), .ZN(n916) );
  XOR2_X1 U753 ( .A(n916), .B(n675), .Z(n676) );
  NOR2_X1 U754 ( .A1(n678), .A2(n676), .ZN(n680) );
  AND2_X1 U755 ( .A1(n678), .A2(n677), .ZN(n679) );
  NOR2_X1 U756 ( .A1(n680), .A2(n679), .ZN(G295) );
  NAND2_X1 U757 ( .A1(G2078), .A2(G2084), .ZN(n681) );
  XOR2_X1 U758 ( .A(KEYINPUT20), .B(n681), .Z(n682) );
  NAND2_X1 U759 ( .A1(G2090), .A2(n682), .ZN(n683) );
  XNOR2_X1 U760 ( .A(KEYINPUT21), .B(n683), .ZN(n684) );
  NAND2_X1 U761 ( .A1(n684), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U762 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U763 ( .A(KEYINPUT72), .B(G82), .Z(G220) );
  NOR2_X1 U764 ( .A1(G220), .A2(G219), .ZN(n685) );
  XOR2_X1 U765 ( .A(KEYINPUT22), .B(n685), .Z(n686) );
  NOR2_X1 U766 ( .A1(G218), .A2(n686), .ZN(n687) );
  NAND2_X1 U767 ( .A1(G96), .A2(n687), .ZN(n855) );
  NAND2_X1 U768 ( .A1(G2106), .A2(n855), .ZN(n691) );
  NAND2_X1 U769 ( .A1(G69), .A2(G120), .ZN(n688) );
  NOR2_X1 U770 ( .A1(G237), .A2(n688), .ZN(n689) );
  NAND2_X1 U771 ( .A1(G108), .A2(n689), .ZN(n856) );
  NAND2_X1 U772 ( .A1(G567), .A2(n856), .ZN(n690) );
  NAND2_X1 U773 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U774 ( .A(KEYINPUT84), .B(n692), .ZN(n854) );
  NAND2_X1 U775 ( .A1(G661), .A2(G483), .ZN(n693) );
  NOR2_X1 U776 ( .A1(n854), .A2(n693), .ZN(n853) );
  NAND2_X1 U777 ( .A1(n853), .A2(G36), .ZN(G176) );
  NOR2_X1 U778 ( .A1(G164), .A2(G1384), .ZN(n803) );
  INV_X1 U779 ( .A(n803), .ZN(n694) );
  NAND2_X1 U780 ( .A1(G40), .A2(G160), .ZN(n802) );
  NOR2_X1 U781 ( .A1(n694), .A2(n802), .ZN(n710) );
  INV_X1 U782 ( .A(n710), .ZN(n714) );
  INV_X1 U783 ( .A(n714), .ZN(n695) );
  INV_X1 U784 ( .A(n695), .ZN(n749) );
  NOR2_X1 U785 ( .A1(n749), .A2(G2084), .ZN(n696) );
  XNOR2_X1 U786 ( .A(n696), .B(KEYINPUT94), .ZN(n757) );
  NAND2_X1 U787 ( .A1(n714), .A2(G8), .ZN(n698) );
  INV_X1 U788 ( .A(KEYINPUT93), .ZN(n697) );
  NOR2_X1 U789 ( .A1(G1966), .A2(n748), .ZN(n762) );
  XNOR2_X1 U790 ( .A(n699), .B(KEYINPUT104), .ZN(n700) );
  NAND2_X1 U791 ( .A1(n700), .A2(G8), .ZN(n701) );
  XNOR2_X1 U792 ( .A(n703), .B(KEYINPUT105), .ZN(n708) );
  XOR2_X1 U793 ( .A(G1961), .B(KEYINPUT96), .Z(n958) );
  NAND2_X1 U794 ( .A1(n958), .A2(n749), .ZN(n704) );
  XNOR2_X1 U795 ( .A(n704), .B(KEYINPUT97), .ZN(n706) );
  XOR2_X1 U796 ( .A(KEYINPUT25), .B(G2078), .Z(n940) );
  NOR2_X1 U797 ( .A1(n749), .A2(n940), .ZN(n705) );
  NOR2_X1 U798 ( .A1(n706), .A2(n705), .ZN(n741) );
  NAND2_X1 U799 ( .A1(n741), .A2(G301), .ZN(n707) );
  NAND2_X1 U800 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U801 ( .A(n709), .B(KEYINPUT31), .ZN(n745) );
  NAND2_X1 U802 ( .A1(G1348), .A2(n714), .ZN(n712) );
  BUF_X1 U803 ( .A(n710), .Z(n729) );
  NAND2_X1 U804 ( .A1(G2067), .A2(n729), .ZN(n711) );
  NAND2_X1 U805 ( .A1(n712), .A2(n711), .ZN(n713) );
  XOR2_X1 U806 ( .A(KEYINPUT100), .B(n713), .Z(n721) );
  NAND2_X1 U807 ( .A1(G1341), .A2(n714), .ZN(n715) );
  XNOR2_X1 U808 ( .A(n715), .B(KEYINPUT99), .ZN(n716) );
  NOR2_X1 U809 ( .A1(n716), .A2(n1018), .ZN(n719) );
  NAND2_X1 U810 ( .A1(G1996), .A2(n729), .ZN(n717) );
  XNOR2_X1 U811 ( .A(KEYINPUT26), .B(n717), .ZN(n718) );
  NAND2_X1 U812 ( .A1(n719), .A2(n718), .ZN(n723) );
  NOR2_X1 U813 ( .A1(n723), .A2(n1017), .ZN(n720) );
  NOR2_X1 U814 ( .A1(n721), .A2(n720), .ZN(n722) );
  XNOR2_X1 U815 ( .A(n722), .B(KEYINPUT101), .ZN(n727) );
  AND2_X1 U816 ( .A1(n1017), .A2(n723), .ZN(n724) );
  XNOR2_X1 U817 ( .A(KEYINPUT102), .B(n724), .ZN(n725) );
  INV_X1 U818 ( .A(n725), .ZN(n726) );
  NAND2_X1 U819 ( .A1(G1956), .A2(n749), .ZN(n728) );
  XNOR2_X1 U820 ( .A(KEYINPUT98), .B(n728), .ZN(n732) );
  NAND2_X1 U821 ( .A1(n729), .A2(G2072), .ZN(n730) );
  XOR2_X1 U822 ( .A(KEYINPUT27), .B(n730), .Z(n731) );
  NAND2_X1 U823 ( .A1(n732), .A2(n731), .ZN(n735) );
  NOR2_X1 U824 ( .A1(G299), .A2(n735), .ZN(n733) );
  XNOR2_X1 U825 ( .A(n734), .B(KEYINPUT103), .ZN(n738) );
  NAND2_X1 U826 ( .A1(G299), .A2(n735), .ZN(n736) );
  XNOR2_X1 U827 ( .A(KEYINPUT28), .B(n736), .ZN(n737) );
  NAND2_X1 U828 ( .A1(n738), .A2(n737), .ZN(n740) );
  INV_X1 U829 ( .A(KEYINPUT29), .ZN(n739) );
  XNOR2_X1 U830 ( .A(n740), .B(n739), .ZN(n743) );
  OR2_X1 U831 ( .A1(n741), .A2(G301), .ZN(n742) );
  NAND2_X1 U832 ( .A1(n743), .A2(n742), .ZN(n744) );
  NAND2_X1 U833 ( .A1(n745), .A2(n744), .ZN(n759) );
  NAND2_X1 U834 ( .A1(n759), .A2(G286), .ZN(n747) );
  XNOR2_X1 U835 ( .A(n747), .B(n746), .ZN(n754) );
  NOR2_X1 U836 ( .A1(G1971), .A2(n835), .ZN(n751) );
  NOR2_X1 U837 ( .A1(G2090), .A2(n749), .ZN(n750) );
  NOR2_X1 U838 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U839 ( .A1(G303), .A2(n752), .ZN(n753) );
  NAND2_X1 U840 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U841 ( .A1(n755), .A2(G8), .ZN(n756) );
  XNOR2_X1 U842 ( .A(n756), .B(KEYINPUT32), .ZN(n764) );
  NAND2_X1 U843 ( .A1(G8), .A2(n757), .ZN(n758) );
  XOR2_X1 U844 ( .A(KEYINPUT95), .B(n758), .Z(n760) );
  NAND2_X1 U845 ( .A1(n760), .A2(n759), .ZN(n761) );
  NOR2_X1 U846 ( .A1(n762), .A2(n761), .ZN(n763) );
  XNOR2_X1 U847 ( .A(n525), .B(KEYINPUT108), .ZN(n834) );
  INV_X1 U848 ( .A(G1971), .ZN(n1028) );
  NAND2_X1 U849 ( .A1(G166), .A2(n1028), .ZN(n766) );
  NOR2_X1 U850 ( .A1(G1976), .A2(G288), .ZN(n823) );
  INV_X1 U851 ( .A(n823), .ZN(n765) );
  NAND2_X1 U852 ( .A1(n766), .A2(n765), .ZN(n1030) );
  OR2_X1 U853 ( .A1(n834), .A2(n1030), .ZN(n769) );
  NAND2_X1 U854 ( .A1(G1976), .A2(G288), .ZN(n1032) );
  INV_X1 U855 ( .A(n1032), .ZN(n767) );
  NAND2_X1 U856 ( .A1(n769), .A2(n526), .ZN(n771) );
  INV_X1 U857 ( .A(KEYINPUT33), .ZN(n770) );
  NAND2_X1 U858 ( .A1(n771), .A2(n770), .ZN(n829) );
  XOR2_X1 U859 ( .A(G1981), .B(G305), .Z(n1021) );
  XOR2_X1 U860 ( .A(KEYINPUT89), .B(KEYINPUT36), .Z(n783) );
  NAND2_X1 U861 ( .A1(G128), .A2(n904), .ZN(n773) );
  NAND2_X1 U862 ( .A1(G116), .A2(n905), .ZN(n772) );
  NAND2_X1 U863 ( .A1(n773), .A2(n772), .ZN(n774) );
  XOR2_X1 U864 ( .A(KEYINPUT35), .B(n774), .Z(n781) );
  XNOR2_X1 U865 ( .A(KEYINPUT87), .B(KEYINPUT88), .ZN(n778) );
  NAND2_X1 U866 ( .A1(n901), .A2(G104), .ZN(n776) );
  NAND2_X1 U867 ( .A1(G140), .A2(n578), .ZN(n775) );
  NAND2_X1 U868 ( .A1(n776), .A2(n775), .ZN(n777) );
  XNOR2_X1 U869 ( .A(n778), .B(n777), .ZN(n779) );
  XOR2_X1 U870 ( .A(n779), .B(KEYINPUT34), .Z(n780) );
  NOR2_X1 U871 ( .A1(n781), .A2(n780), .ZN(n782) );
  XNOR2_X1 U872 ( .A(n783), .B(n782), .ZN(n898) );
  XNOR2_X1 U873 ( .A(G2067), .B(KEYINPUT37), .ZN(n811) );
  AND2_X1 U874 ( .A1(n898), .A2(n811), .ZN(n784) );
  XNOR2_X1 U875 ( .A(KEYINPUT111), .B(n784), .ZN(n1000) );
  NAND2_X1 U876 ( .A1(n901), .A2(G105), .ZN(n785) );
  XNOR2_X1 U877 ( .A(n785), .B(KEYINPUT38), .ZN(n787) );
  NAND2_X1 U878 ( .A1(G117), .A2(n905), .ZN(n786) );
  NAND2_X1 U879 ( .A1(n787), .A2(n786), .ZN(n790) );
  NAND2_X1 U880 ( .A1(G129), .A2(n904), .ZN(n788) );
  XNOR2_X1 U881 ( .A(KEYINPUT91), .B(n788), .ZN(n789) );
  NOR2_X1 U882 ( .A1(n790), .A2(n789), .ZN(n791) );
  XNOR2_X1 U883 ( .A(n791), .B(KEYINPUT92), .ZN(n793) );
  NAND2_X1 U884 ( .A1(G141), .A2(n578), .ZN(n792) );
  NAND2_X1 U885 ( .A1(n793), .A2(n792), .ZN(n895) );
  NOR2_X1 U886 ( .A1(G1996), .A2(n895), .ZN(n987) );
  NAND2_X1 U887 ( .A1(n901), .A2(G95), .ZN(n795) );
  NAND2_X1 U888 ( .A1(G131), .A2(n578), .ZN(n794) );
  NAND2_X1 U889 ( .A1(n795), .A2(n794), .ZN(n799) );
  NAND2_X1 U890 ( .A1(G119), .A2(n904), .ZN(n797) );
  NAND2_X1 U891 ( .A1(G107), .A2(n905), .ZN(n796) );
  NAND2_X1 U892 ( .A1(n797), .A2(n796), .ZN(n798) );
  OR2_X1 U893 ( .A1(n799), .A2(n798), .ZN(n882) );
  AND2_X1 U894 ( .A1(n882), .A2(G1991), .ZN(n801) );
  AND2_X1 U895 ( .A1(G1996), .A2(n895), .ZN(n800) );
  NOR2_X1 U896 ( .A1(n801), .A2(n800), .ZN(n990) );
  INV_X1 U897 ( .A(n990), .ZN(n804) );
  NOR2_X1 U898 ( .A1(n803), .A2(n802), .ZN(n816) );
  NAND2_X1 U899 ( .A1(n804), .A2(n816), .ZN(n817) );
  INV_X1 U900 ( .A(n817), .ZN(n807) );
  NOR2_X1 U901 ( .A1(G290), .A2(G1986), .ZN(n805) );
  NOR2_X1 U902 ( .A1(G1991), .A2(n882), .ZN(n993) );
  NOR2_X1 U903 ( .A1(n805), .A2(n993), .ZN(n806) );
  NOR2_X1 U904 ( .A1(n807), .A2(n806), .ZN(n808) );
  NOR2_X1 U905 ( .A1(n987), .A2(n808), .ZN(n809) );
  XNOR2_X1 U906 ( .A(KEYINPUT110), .B(n809), .ZN(n810) );
  XNOR2_X1 U907 ( .A(n810), .B(KEYINPUT39), .ZN(n813) );
  NOR2_X1 U908 ( .A1(n811), .A2(n898), .ZN(n812) );
  XNOR2_X1 U909 ( .A(n812), .B(KEYINPUT90), .ZN(n1003) );
  NAND2_X1 U910 ( .A1(n816), .A2(n1003), .ZN(n818) );
  NAND2_X1 U911 ( .A1(n813), .A2(n818), .ZN(n814) );
  NAND2_X1 U912 ( .A1(n1000), .A2(n814), .ZN(n815) );
  NAND2_X1 U913 ( .A1(n815), .A2(n816), .ZN(n836) );
  INV_X1 U914 ( .A(n836), .ZN(n831) );
  XNOR2_X1 U915 ( .A(G290), .B(G1986), .ZN(n1025) );
  AND2_X1 U916 ( .A1(n1025), .A2(n816), .ZN(n820) );
  NAND2_X1 U917 ( .A1(n818), .A2(n817), .ZN(n819) );
  NOR2_X1 U918 ( .A1(n820), .A2(n819), .ZN(n821) );
  OR2_X1 U919 ( .A1(n831), .A2(n821), .ZN(n837) );
  AND2_X1 U920 ( .A1(n1021), .A2(n837), .ZN(n827) );
  NAND2_X1 U921 ( .A1(n823), .A2(KEYINPUT33), .ZN(n822) );
  NAND2_X1 U922 ( .A1(n768), .A2(n822), .ZN(n825) );
  NAND2_X1 U923 ( .A1(n823), .A2(KEYINPUT109), .ZN(n824) );
  NAND2_X1 U924 ( .A1(n825), .A2(n824), .ZN(n826) );
  NAND2_X1 U925 ( .A1(n829), .A2(n828), .ZN(n847) );
  NAND2_X1 U926 ( .A1(G166), .A2(G8), .ZN(n830) );
  NOR2_X1 U927 ( .A1(G2090), .A2(n830), .ZN(n832) );
  OR2_X1 U928 ( .A1(n832), .A2(n831), .ZN(n833) );
  INV_X1 U929 ( .A(n835), .ZN(n840) );
  AND2_X1 U930 ( .A1(n836), .A2(n840), .ZN(n838) );
  INV_X1 U931 ( .A(n837), .ZN(n843) );
  NAND2_X1 U932 ( .A1(n532), .A2(n527), .ZN(n845) );
  NOR2_X1 U933 ( .A1(G1981), .A2(G305), .ZN(n839) );
  XNOR2_X1 U934 ( .A(n839), .B(KEYINPUT24), .ZN(n841) );
  NAND2_X1 U935 ( .A1(n841), .A2(n840), .ZN(n842) );
  OR2_X1 U936 ( .A1(n843), .A2(n842), .ZN(n844) );
  NAND2_X1 U937 ( .A1(n847), .A2(n846), .ZN(n849) );
  XNOR2_X1 U938 ( .A(KEYINPUT40), .B(KEYINPUT112), .ZN(n848) );
  XNOR2_X1 U939 ( .A(n849), .B(n848), .ZN(G329) );
  NAND2_X1 U940 ( .A1(G2106), .A2(n850), .ZN(G217) );
  INV_X1 U941 ( .A(n850), .ZN(G223) );
  AND2_X1 U942 ( .A1(G15), .A2(G2), .ZN(n851) );
  NAND2_X1 U943 ( .A1(G661), .A2(n851), .ZN(G259) );
  NAND2_X1 U944 ( .A1(G3), .A2(G1), .ZN(n852) );
  NAND2_X1 U945 ( .A1(n853), .A2(n852), .ZN(G188) );
  INV_X1 U946 ( .A(n854), .ZN(G319) );
  INV_X1 U948 ( .A(G120), .ZN(G236) );
  INV_X1 U949 ( .A(G96), .ZN(G221) );
  INV_X1 U950 ( .A(G69), .ZN(G235) );
  NOR2_X1 U951 ( .A1(n856), .A2(n855), .ZN(G325) );
  INV_X1 U952 ( .A(G325), .ZN(G261) );
  XOR2_X1 U953 ( .A(G2100), .B(G2096), .Z(n858) );
  XNOR2_X1 U954 ( .A(KEYINPUT42), .B(G2678), .ZN(n857) );
  XNOR2_X1 U955 ( .A(n858), .B(n857), .ZN(n862) );
  XOR2_X1 U956 ( .A(KEYINPUT43), .B(G2072), .Z(n860) );
  XNOR2_X1 U957 ( .A(G2067), .B(G2090), .ZN(n859) );
  XNOR2_X1 U958 ( .A(n860), .B(n859), .ZN(n861) );
  XOR2_X1 U959 ( .A(n862), .B(n861), .Z(n864) );
  XNOR2_X1 U960 ( .A(G2078), .B(G2084), .ZN(n863) );
  XNOR2_X1 U961 ( .A(n864), .B(n863), .ZN(G227) );
  XOR2_X1 U962 ( .A(G1976), .B(G1956), .Z(n866) );
  XNOR2_X1 U963 ( .A(G1991), .B(G1961), .ZN(n865) );
  XNOR2_X1 U964 ( .A(n866), .B(n865), .ZN(n870) );
  XNOR2_X1 U965 ( .A(G1981), .B(n1028), .ZN(n868) );
  XNOR2_X1 U966 ( .A(G1986), .B(G1966), .ZN(n867) );
  XNOR2_X1 U967 ( .A(n868), .B(n867), .ZN(n869) );
  XOR2_X1 U968 ( .A(n870), .B(n869), .Z(n872) );
  XNOR2_X1 U969 ( .A(G2474), .B(KEYINPUT113), .ZN(n871) );
  XNOR2_X1 U970 ( .A(n872), .B(n871), .ZN(n873) );
  XNOR2_X1 U971 ( .A(KEYINPUT41), .B(n873), .ZN(n874) );
  XOR2_X1 U972 ( .A(n874), .B(G1996), .Z(G229) );
  NAND2_X1 U973 ( .A1(n904), .A2(G124), .ZN(n875) );
  XNOR2_X1 U974 ( .A(n875), .B(KEYINPUT44), .ZN(n877) );
  NAND2_X1 U975 ( .A1(G100), .A2(n901), .ZN(n876) );
  NAND2_X1 U976 ( .A1(n877), .A2(n876), .ZN(n881) );
  NAND2_X1 U977 ( .A1(G112), .A2(n905), .ZN(n879) );
  NAND2_X1 U978 ( .A1(G136), .A2(n578), .ZN(n878) );
  NAND2_X1 U979 ( .A1(n879), .A2(n878), .ZN(n880) );
  NOR2_X1 U980 ( .A1(n881), .A2(n880), .ZN(G162) );
  XNOR2_X1 U981 ( .A(G164), .B(G160), .ZN(n883) );
  XNOR2_X1 U982 ( .A(n883), .B(n882), .ZN(n887) );
  XOR2_X1 U983 ( .A(KEYINPUT116), .B(KEYINPUT46), .Z(n885) );
  XNOR2_X1 U984 ( .A(KEYINPUT115), .B(KEYINPUT48), .ZN(n884) );
  XNOR2_X1 U985 ( .A(n885), .B(n884), .ZN(n886) );
  XOR2_X1 U986 ( .A(n887), .B(n886), .Z(n900) );
  NAND2_X1 U987 ( .A1(G130), .A2(n904), .ZN(n889) );
  NAND2_X1 U988 ( .A1(G118), .A2(n905), .ZN(n888) );
  NAND2_X1 U989 ( .A1(n889), .A2(n888), .ZN(n894) );
  NAND2_X1 U990 ( .A1(n901), .A2(G106), .ZN(n891) );
  NAND2_X1 U991 ( .A1(G142), .A2(n578), .ZN(n890) );
  NAND2_X1 U992 ( .A1(n891), .A2(n890), .ZN(n892) );
  XOR2_X1 U993 ( .A(n892), .B(KEYINPUT45), .Z(n893) );
  NOR2_X1 U994 ( .A1(n894), .A2(n893), .ZN(n896) );
  XNOR2_X1 U995 ( .A(n896), .B(n895), .ZN(n897) );
  XOR2_X1 U996 ( .A(n898), .B(n897), .Z(n899) );
  XNOR2_X1 U997 ( .A(n900), .B(n899), .ZN(n912) );
  NAND2_X1 U998 ( .A1(n901), .A2(G103), .ZN(n903) );
  NAND2_X1 U999 ( .A1(G139), .A2(n578), .ZN(n902) );
  NAND2_X1 U1000 ( .A1(n903), .A2(n902), .ZN(n910) );
  NAND2_X1 U1001 ( .A1(G127), .A2(n904), .ZN(n907) );
  NAND2_X1 U1002 ( .A1(G115), .A2(n905), .ZN(n906) );
  NAND2_X1 U1003 ( .A1(n907), .A2(n906), .ZN(n908) );
  XOR2_X1 U1004 ( .A(KEYINPUT47), .B(n908), .Z(n909) );
  NOR2_X1 U1005 ( .A1(n910), .A2(n909), .ZN(n911) );
  XOR2_X1 U1006 ( .A(KEYINPUT114), .B(n911), .Z(n982) );
  XOR2_X1 U1007 ( .A(n912), .B(n982), .Z(n914) );
  XNOR2_X1 U1008 ( .A(n992), .B(G162), .ZN(n913) );
  XNOR2_X1 U1009 ( .A(n914), .B(n913), .ZN(n915) );
  NOR2_X1 U1010 ( .A1(G37), .A2(n915), .ZN(G395) );
  XOR2_X1 U1011 ( .A(n916), .B(G286), .Z(n919) );
  XOR2_X1 U1012 ( .A(G301), .B(n917), .Z(n918) );
  XNOR2_X1 U1013 ( .A(n919), .B(n918), .ZN(n920) );
  XNOR2_X1 U1014 ( .A(n920), .B(n1018), .ZN(n921) );
  NOR2_X1 U1015 ( .A1(G37), .A2(n921), .ZN(G397) );
  XOR2_X1 U1016 ( .A(G2451), .B(G2430), .Z(n923) );
  XNOR2_X1 U1017 ( .A(G2438), .B(G2443), .ZN(n922) );
  XNOR2_X1 U1018 ( .A(n923), .B(n922), .ZN(n929) );
  XOR2_X1 U1019 ( .A(G2435), .B(G2454), .Z(n925) );
  XNOR2_X1 U1020 ( .A(G1341), .B(G1348), .ZN(n924) );
  XNOR2_X1 U1021 ( .A(n925), .B(n924), .ZN(n927) );
  XOR2_X1 U1022 ( .A(G2446), .B(G2427), .Z(n926) );
  XNOR2_X1 U1023 ( .A(n927), .B(n926), .ZN(n928) );
  XOR2_X1 U1024 ( .A(n929), .B(n928), .Z(n930) );
  NAND2_X1 U1025 ( .A1(G14), .A2(n930), .ZN(n936) );
  NAND2_X1 U1026 ( .A1(n936), .A2(G319), .ZN(n933) );
  NOR2_X1 U1027 ( .A1(G227), .A2(G229), .ZN(n931) );
  XNOR2_X1 U1028 ( .A(KEYINPUT49), .B(n931), .ZN(n932) );
  NOR2_X1 U1029 ( .A1(n933), .A2(n932), .ZN(n935) );
  NOR2_X1 U1030 ( .A1(G395), .A2(G397), .ZN(n934) );
  NAND2_X1 U1031 ( .A1(n935), .A2(n934), .ZN(G225) );
  INV_X1 U1032 ( .A(G225), .ZN(G308) );
  INV_X1 U1033 ( .A(G108), .ZN(G238) );
  INV_X1 U1034 ( .A(n936), .ZN(G401) );
  INV_X1 U1035 ( .A(KEYINPUT55), .ZN(n1008) );
  XOR2_X1 U1036 ( .A(G25), .B(G1991), .Z(n937) );
  NAND2_X1 U1037 ( .A1(n937), .A2(G28), .ZN(n946) );
  XNOR2_X1 U1038 ( .A(G1996), .B(G32), .ZN(n939) );
  XNOR2_X1 U1039 ( .A(G33), .B(G2072), .ZN(n938) );
  NOR2_X1 U1040 ( .A1(n939), .A2(n938), .ZN(n944) );
  XNOR2_X1 U1041 ( .A(G2067), .B(G26), .ZN(n942) );
  XNOR2_X1 U1042 ( .A(G27), .B(n940), .ZN(n941) );
  NOR2_X1 U1043 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1044 ( .A1(n944), .A2(n943), .ZN(n945) );
  NOR2_X1 U1045 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1046 ( .A(n947), .B(KEYINPUT53), .ZN(n948) );
  XNOR2_X1 U1047 ( .A(n948), .B(KEYINPUT123), .ZN(n951) );
  XOR2_X1 U1048 ( .A(G2084), .B(KEYINPUT54), .Z(n949) );
  XNOR2_X1 U1049 ( .A(G34), .B(n949), .ZN(n950) );
  NAND2_X1 U1050 ( .A1(n951), .A2(n950), .ZN(n954) );
  XNOR2_X1 U1051 ( .A(KEYINPUT122), .B(G2090), .ZN(n952) );
  XNOR2_X1 U1052 ( .A(G35), .B(n952), .ZN(n953) );
  NOR2_X1 U1053 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1054 ( .A(n1008), .B(n955), .ZN(n956) );
  NOR2_X1 U1055 ( .A1(G29), .A2(n956), .ZN(n957) );
  XOR2_X1 U1056 ( .A(KEYINPUT124), .B(n957), .Z(n1015) );
  XOR2_X1 U1057 ( .A(G1966), .B(G21), .Z(n960) );
  XNOR2_X1 U1058 ( .A(n958), .B(G5), .ZN(n959) );
  NAND2_X1 U1059 ( .A1(n960), .A2(n959), .ZN(n978) );
  XOR2_X1 U1060 ( .A(G22), .B(G1971), .Z(n964) );
  XNOR2_X1 U1061 ( .A(G1986), .B(G24), .ZN(n962) );
  XNOR2_X1 U1062 ( .A(G1976), .B(G23), .ZN(n961) );
  NOR2_X1 U1063 ( .A1(n962), .A2(n961), .ZN(n963) );
  NAND2_X1 U1064 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1065 ( .A(n965), .B(KEYINPUT127), .ZN(n966) );
  XNOR2_X1 U1066 ( .A(n966), .B(KEYINPUT58), .ZN(n976) );
  XOR2_X1 U1067 ( .A(G1348), .B(KEYINPUT59), .Z(n967) );
  XNOR2_X1 U1068 ( .A(G4), .B(n967), .ZN(n969) );
  XNOR2_X1 U1069 ( .A(G20), .B(G1956), .ZN(n968) );
  NOR2_X1 U1070 ( .A1(n969), .A2(n968), .ZN(n973) );
  XNOR2_X1 U1071 ( .A(G1341), .B(G19), .ZN(n971) );
  XNOR2_X1 U1072 ( .A(G6), .B(G1981), .ZN(n970) );
  NOR2_X1 U1073 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1074 ( .A1(n973), .A2(n972), .ZN(n974) );
  XOR2_X1 U1075 ( .A(KEYINPUT60), .B(n974), .Z(n975) );
  NAND2_X1 U1076 ( .A1(n976), .A2(n975), .ZN(n977) );
  NOR2_X1 U1077 ( .A1(n978), .A2(n977), .ZN(n979) );
  XNOR2_X1 U1078 ( .A(KEYINPUT61), .B(n979), .ZN(n980) );
  INV_X1 U1079 ( .A(G16), .ZN(n1016) );
  NAND2_X1 U1080 ( .A1(n980), .A2(n1016), .ZN(n981) );
  NAND2_X1 U1081 ( .A1(n981), .A2(G11), .ZN(n1013) );
  XOR2_X1 U1082 ( .A(G164), .B(G2078), .Z(n984) );
  XNOR2_X1 U1083 ( .A(G2072), .B(n982), .ZN(n983) );
  NOR2_X1 U1084 ( .A1(n984), .A2(n983), .ZN(n985) );
  XOR2_X1 U1085 ( .A(KEYINPUT50), .B(n985), .Z(n1006) );
  XOR2_X1 U1086 ( .A(G2090), .B(G162), .Z(n986) );
  NOR2_X1 U1087 ( .A1(n987), .A2(n986), .ZN(n988) );
  XNOR2_X1 U1088 ( .A(n988), .B(KEYINPUT119), .ZN(n989) );
  XNOR2_X1 U1089 ( .A(n989), .B(KEYINPUT51), .ZN(n991) );
  NAND2_X1 U1090 ( .A1(n991), .A2(n990), .ZN(n999) );
  XOR2_X1 U1091 ( .A(G160), .B(G2084), .Z(n996) );
  NOR2_X1 U1092 ( .A1(n993), .A2(n992), .ZN(n994) );
  XNOR2_X1 U1093 ( .A(KEYINPUT117), .B(n994), .ZN(n995) );
  NOR2_X1 U1094 ( .A1(n996), .A2(n995), .ZN(n997) );
  XOR2_X1 U1095 ( .A(KEYINPUT118), .B(n997), .Z(n998) );
  NOR2_X1 U1096 ( .A1(n999), .A2(n998), .ZN(n1001) );
  NAND2_X1 U1097 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NOR2_X1 U1098 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XOR2_X1 U1099 ( .A(KEYINPUT120), .B(n1004), .Z(n1005) );
  NOR2_X1 U1100 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1101 ( .A(n1007), .B(KEYINPUT52), .ZN(n1009) );
  NAND2_X1 U1102 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1103 ( .A1(G29), .A2(n1010), .ZN(n1011) );
  XNOR2_X1 U1104 ( .A(KEYINPUT121), .B(n1011), .ZN(n1012) );
  NOR2_X1 U1105 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1106 ( .A1(n1015), .A2(n1014), .ZN(n1044) );
  XNOR2_X1 U1107 ( .A(n1016), .B(KEYINPUT56), .ZN(n1042) );
  XOR2_X1 U1108 ( .A(n1017), .B(G1348), .Z(n1020) );
  XOR2_X1 U1109 ( .A(G1341), .B(n1018), .Z(n1019) );
  NAND2_X1 U1110 ( .A1(n1020), .A2(n1019), .ZN(n1039) );
  XNOR2_X1 U1111 ( .A(G1966), .B(G168), .ZN(n1022) );
  NAND2_X1 U1112 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XNOR2_X1 U1113 ( .A(n1023), .B(KEYINPUT57), .ZN(n1037) );
  XOR2_X1 U1114 ( .A(G301), .B(G1961), .Z(n1027) );
  XNOR2_X1 U1115 ( .A(G1956), .B(G299), .ZN(n1024) );
  NOR2_X1 U1116 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NAND2_X1 U1117 ( .A1(n1027), .A2(n1026), .ZN(n1035) );
  NOR2_X1 U1118 ( .A1(G166), .A2(n1028), .ZN(n1029) );
  NOR2_X1 U1119 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NAND2_X1 U1120 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  XOR2_X1 U1121 ( .A(KEYINPUT125), .B(n1033), .Z(n1034) );
  NOR2_X1 U1122 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  NAND2_X1 U1123 ( .A1(n1037), .A2(n1036), .ZN(n1038) );
  NOR2_X1 U1124 ( .A1(n1039), .A2(n1038), .ZN(n1040) );
  XNOR2_X1 U1125 ( .A(KEYINPUT126), .B(n1040), .ZN(n1041) );
  NOR2_X1 U1126 ( .A1(n1042), .A2(n1041), .ZN(n1043) );
  NOR2_X1 U1127 ( .A1(n1044), .A2(n1043), .ZN(n1045) );
  XOR2_X1 U1128 ( .A(n1045), .B(KEYINPUT62), .Z(G150) );
  INV_X1 U1129 ( .A(G150), .ZN(G311) );
endmodule

