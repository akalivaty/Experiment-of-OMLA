//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 1 0 1 1 1 0 0 1 0 1 1 0 1 0 1 0 0 0 1 0 1 0 0 1 1 1 0 1 0 0 1 1 1 0 0 1 0 0 1 1 0 0 1 0 1 1 0 0 1 0 1 0 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:53 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n241, new_n242, new_n243, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n251, new_n252,
    new_n254, new_n255, new_n256, new_n257, new_n258, new_n259, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1259, new_n1260, new_n1261, new_n1262, new_n1263,
    new_n1264, new_n1265, new_n1266;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  AOI22_X1  g0005(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n206));
  INV_X1    g0006(.A(G87), .ZN(new_n207));
  INV_X1    g0007(.A(G250), .ZN(new_n208));
  INV_X1    g0008(.A(G107), .ZN(new_n209));
  INV_X1    g0009(.A(G264), .ZN(new_n210));
  OAI221_X1 g0010(.A(new_n206), .B1(new_n207), .B2(new_n208), .C1(new_n209), .C2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(KEYINPUT65), .ZN(new_n212));
  OR2_X1    g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G116), .A2(G270), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n211), .A2(new_n212), .ZN(new_n215));
  INV_X1    g0015(.A(G226), .ZN(new_n216));
  INV_X1    g0016(.A(G68), .ZN(new_n217));
  INV_X1    g0017(.A(G238), .ZN(new_n218));
  OAI22_X1  g0018(.A1(new_n202), .A2(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  AOI21_X1  g0019(.A(new_n219), .B1(G77), .B2(G244), .ZN(new_n220));
  NAND4_X1  g0020(.A1(new_n213), .A2(new_n214), .A3(new_n215), .A4(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(G1), .ZN(new_n222));
  INV_X1    g0022(.A(G20), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g0024(.A(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n221), .A2(new_n225), .ZN(new_n226));
  XOR2_X1   g0026(.A(new_n226), .B(KEYINPUT1), .Z(new_n227));
  NOR2_X1   g0027(.A1(new_n225), .A2(G13), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  INV_X1    g0029(.A(G257), .ZN(new_n230));
  AOI211_X1 g0030(.A(new_n208), .B(new_n229), .C1(new_n230), .C2(new_n210), .ZN(new_n231));
  NAND2_X1  g0031(.A1(G1), .A2(G13), .ZN(new_n232));
  INV_X1    g0032(.A(KEYINPUT64), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g0034(.A1(KEYINPUT64), .A2(G1), .A3(G13), .ZN(new_n235));
  NAND2_X1  g0035(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  INV_X1    g0036(.A(new_n236), .ZN(new_n237));
  NOR2_X1   g0037(.A1(new_n237), .A2(new_n223), .ZN(new_n238));
  INV_X1    g0038(.A(new_n201), .ZN(new_n239));
  NAND2_X1  g0039(.A1(new_n239), .A2(G50), .ZN(new_n240));
  INV_X1    g0040(.A(new_n240), .ZN(new_n241));
  AOI22_X1  g0041(.A1(new_n231), .A2(KEYINPUT0), .B1(new_n238), .B2(new_n241), .ZN(new_n242));
  OAI211_X1 g0042(.A(new_n227), .B(new_n242), .C1(KEYINPUT0), .C2(new_n231), .ZN(new_n243));
  INV_X1    g0043(.A(new_n243), .ZN(G361));
  XNOR2_X1  g0044(.A(G238), .B(G244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(G232), .ZN(new_n246));
  XNOR2_X1  g0046(.A(KEYINPUT2), .B(G226), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n246), .B(new_n247), .Z(new_n248));
  XOR2_X1   g0048(.A(new_n248), .B(KEYINPUT66), .Z(new_n249));
  XNOR2_X1  g0049(.A(G250), .B(G257), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G264), .B(G270), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n249), .B(new_n252), .ZN(G358));
  XOR2_X1   g0053(.A(G68), .B(G77), .Z(new_n254));
  XNOR2_X1  g0054(.A(G50), .B(G58), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n254), .B(new_n255), .ZN(new_n256));
  XOR2_X1   g0056(.A(G87), .B(G97), .Z(new_n257));
  XNOR2_X1  g0057(.A(G107), .B(G116), .ZN(new_n258));
  XNOR2_X1  g0058(.A(new_n257), .B(new_n258), .ZN(new_n259));
  XNOR2_X1  g0059(.A(new_n256), .B(new_n259), .ZN(G351));
  NAND3_X1  g0060(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n234), .A2(new_n235), .A3(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT16), .ZN(new_n263));
  NAND2_X1  g0063(.A1(G58), .A2(G68), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n223), .B1(new_n239), .B2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT3), .ZN(new_n266));
  INV_X1    g0066(.A(G33), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(KEYINPUT3), .A2(G33), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n268), .A2(new_n223), .A3(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT7), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND4_X1  g0072(.A1(new_n268), .A2(KEYINPUT7), .A3(new_n223), .A4(new_n269), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n265), .B1(new_n274), .B2(G68), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n223), .A2(new_n267), .ZN(new_n276));
  INV_X1    g0076(.A(G159), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n263), .B1(new_n275), .B2(new_n279), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n217), .B1(new_n272), .B2(new_n273), .ZN(new_n281));
  NOR4_X1   g0081(.A1(new_n281), .A2(KEYINPUT16), .A3(new_n278), .A4(new_n265), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n262), .B1(new_n280), .B2(new_n282), .ZN(new_n283));
  XNOR2_X1  g0083(.A(KEYINPUT8), .B(G58), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n222), .A2(G13), .A3(G20), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n262), .B1(new_n222), .B2(G20), .ZN(new_n288));
  INV_X1    g0088(.A(new_n284), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n283), .A2(new_n287), .A3(new_n290), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n222), .B1(G41), .B2(G45), .ZN(new_n292));
  INV_X1    g0092(.A(G274), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(G33), .A2(G41), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n295), .A2(G1), .A3(G13), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(new_n292), .ZN(new_n297));
  INV_X1    g0097(.A(G232), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n216), .A2(G1698), .ZN(new_n300));
  AND2_X1   g0100(.A1(KEYINPUT3), .A2(G33), .ZN(new_n301));
  NOR2_X1   g0101(.A1(KEYINPUT3), .A2(G33), .ZN(new_n302));
  OAI221_X1 g0102(.A(new_n300), .B1(G223), .B2(G1698), .C1(new_n301), .C2(new_n302), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n303), .B1(new_n267), .B2(new_n207), .ZN(new_n304));
  AOI22_X1  g0104(.A1(new_n234), .A2(new_n235), .B1(G33), .B2(G41), .ZN(new_n305));
  AOI211_X1 g0105(.A(new_n294), .B(new_n299), .C1(new_n304), .C2(new_n305), .ZN(new_n306));
  OR2_X1    g0106(.A1(new_n306), .A2(G169), .ZN(new_n307));
  INV_X1    g0107(.A(G179), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n291), .A2(new_n307), .A3(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT18), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n291), .A2(KEYINPUT18), .A3(new_n307), .A4(new_n309), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT17), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n301), .A2(new_n302), .ZN(new_n316));
  AOI21_X1  g0116(.A(KEYINPUT7), .B1(new_n316), .B2(new_n223), .ZN(new_n317));
  INV_X1    g0117(.A(new_n273), .ZN(new_n318));
  OAI21_X1  g0118(.A(G68), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n265), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n319), .A2(new_n279), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(KEYINPUT16), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n275), .A2(new_n263), .A3(new_n279), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  AOI22_X1  g0124(.A1(new_n324), .A2(new_n262), .B1(new_n284), .B2(new_n286), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n304), .A2(new_n305), .ZN(new_n326));
  INV_X1    g0126(.A(G190), .ZN(new_n327));
  INV_X1    g0127(.A(new_n294), .ZN(new_n328));
  INV_X1    g0128(.A(new_n299), .ZN(new_n329));
  NAND4_X1  g0129(.A1(new_n326), .A2(new_n327), .A3(new_n328), .A4(new_n329), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n330), .B1(new_n306), .B2(G200), .ZN(new_n331));
  NAND4_X1  g0131(.A1(new_n325), .A2(KEYINPUT70), .A3(new_n290), .A4(new_n331), .ZN(new_n332));
  NAND4_X1  g0132(.A1(new_n283), .A2(new_n287), .A3(new_n290), .A4(new_n331), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT70), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n315), .B1(new_n332), .B2(new_n335), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n333), .A2(KEYINPUT17), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n314), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT69), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT14), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT13), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n236), .A2(new_n295), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n268), .A2(new_n269), .ZN(new_n345));
  INV_X1    g0145(.A(G1698), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n216), .A2(new_n346), .ZN(new_n347));
  OAI211_X1 g0147(.A(new_n345), .B(new_n347), .C1(G232), .C2(new_n346), .ZN(new_n348));
  NAND2_X1  g0148(.A1(G33), .A2(G97), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n344), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n350), .A2(new_n294), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n297), .A2(new_n218), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n343), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  NOR4_X1   g0154(.A1(new_n350), .A2(KEYINPUT13), .A3(new_n352), .A4(new_n294), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(G169), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n342), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  OAI221_X1 g0158(.A(G169), .B1(new_n340), .B2(new_n341), .C1(new_n354), .C2(new_n355), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n356), .A2(G179), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n358), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n223), .A2(G33), .ZN(new_n362));
  INV_X1    g0162(.A(G77), .ZN(new_n363));
  OAI22_X1  g0163(.A1(new_n276), .A2(new_n202), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n223), .A2(G68), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n262), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT11), .ZN(new_n367));
  OR2_X1    g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n288), .A2(G68), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n366), .A2(new_n367), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n365), .A2(new_n222), .A3(G13), .ZN(new_n371));
  XNOR2_X1  g0171(.A(new_n371), .B(KEYINPUT12), .ZN(new_n372));
  AND4_X1   g0172(.A1(new_n368), .A2(new_n369), .A3(new_n370), .A4(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n361), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n356), .A2(G190), .ZN(new_n376));
  OAI21_X1  g0176(.A(G200), .B1(new_n354), .B2(new_n355), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n376), .A2(new_n373), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(G238), .A2(G1698), .ZN(new_n379));
  OAI221_X1 g0179(.A(new_n379), .B1(new_n298), .B2(G1698), .C1(new_n301), .C2(new_n302), .ZN(new_n380));
  OAI211_X1 g0180(.A(new_n380), .B(new_n305), .C1(G107), .C2(new_n345), .ZN(new_n381));
  INV_X1    g0181(.A(new_n297), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(G244), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n381), .A2(new_n328), .A3(new_n383), .ZN(new_n384));
  OR2_X1    g0184(.A1(new_n384), .A2(G179), .ZN(new_n385));
  XNOR2_X1  g0185(.A(KEYINPUT15), .B(G87), .ZN(new_n386));
  OAI22_X1  g0186(.A1(new_n284), .A2(new_n276), .B1(new_n386), .B2(new_n362), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n223), .A2(new_n363), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n262), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n288), .A2(G77), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n286), .A2(new_n363), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n389), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n384), .A2(new_n357), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n385), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT68), .ZN(new_n395));
  XNOR2_X1  g0195(.A(KEYINPUT67), .B(G200), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n384), .A2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n395), .B1(new_n398), .B2(new_n392), .ZN(new_n399));
  OR2_X1    g0199(.A1(new_n384), .A2(new_n327), .ZN(new_n400));
  INV_X1    g0200(.A(new_n392), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n401), .A2(new_n397), .A3(KEYINPUT68), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n399), .A2(new_n400), .A3(new_n402), .ZN(new_n403));
  AND4_X1   g0203(.A1(new_n375), .A2(new_n378), .A3(new_n394), .A4(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n203), .A2(G20), .ZN(new_n405));
  INV_X1    g0205(.A(G150), .ZN(new_n406));
  OAI221_X1 g0206(.A(new_n405), .B1(new_n406), .B2(new_n276), .C1(new_n284), .C2(new_n362), .ZN(new_n407));
  AOI22_X1  g0207(.A1(new_n407), .A2(new_n262), .B1(new_n202), .B2(new_n286), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n288), .A2(G50), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT9), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n346), .A2(G222), .ZN(new_n413));
  NAND2_X1  g0213(.A1(G223), .A2(G1698), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n345), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  OAI211_X1 g0215(.A(new_n415), .B(new_n305), .C1(G77), .C2(new_n345), .ZN(new_n416));
  OAI211_X1 g0216(.A(new_n416), .B(new_n328), .C1(new_n216), .C2(new_n297), .ZN(new_n417));
  OR2_X1    g0217(.A1(new_n417), .A2(new_n327), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n408), .A2(KEYINPUT9), .A3(new_n409), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n417), .A2(new_n396), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n412), .A2(new_n418), .A3(new_n419), .A4(new_n420), .ZN(new_n421));
  XNOR2_X1  g0221(.A(new_n421), .B(KEYINPUT10), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n417), .A2(new_n357), .ZN(new_n423));
  OAI211_X1 g0223(.A(new_n423), .B(new_n410), .C1(G179), .C2(new_n417), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n339), .A2(new_n404), .A3(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(G20), .B1(G33), .B2(G283), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n267), .A2(G97), .ZN(new_n430));
  INV_X1    g0230(.A(G116), .ZN(new_n431));
  AOI22_X1  g0231(.A1(new_n429), .A2(new_n430), .B1(G20), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(new_n262), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT20), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n432), .A2(new_n262), .A3(KEYINPUT20), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n285), .A2(new_n431), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n285), .B1(G1), .B2(new_n267), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n262), .A2(new_n439), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n438), .B1(new_n440), .B2(new_n431), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n437), .A2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT5), .ZN(new_n443));
  OR3_X1    g0243(.A1(new_n443), .A2(KEYINPUT74), .A3(G41), .ZN(new_n444));
  OAI21_X1  g0244(.A(KEYINPUT74), .B1(new_n443), .B2(G41), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n444), .A2(G274), .A3(new_n296), .A4(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(G41), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n448), .A2(KEYINPUT5), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n222), .A2(G45), .ZN(new_n450));
  OAI21_X1  g0250(.A(KEYINPUT72), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(G45), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n452), .A2(G1), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT72), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n443), .A2(G41), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n453), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  AND3_X1   g0256(.A1(new_n451), .A2(KEYINPUT73), .A3(new_n456), .ZN(new_n457));
  AOI21_X1  g0257(.A(KEYINPUT73), .B1(new_n451), .B2(new_n456), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n447), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(G264), .A2(G1698), .ZN(new_n460));
  OAI211_X1 g0260(.A(new_n345), .B(new_n460), .C1(new_n230), .C2(G1698), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n461), .B(new_n305), .C1(G303), .C2(new_n345), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n451), .A2(new_n456), .A3(new_n444), .A4(new_n445), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n463), .A2(G270), .A3(new_n296), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n459), .A2(new_n462), .A3(new_n464), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n442), .B1(new_n465), .B2(G200), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n466), .B1(new_n327), .B2(new_n465), .ZN(new_n467));
  AND3_X1   g0267(.A1(new_n459), .A2(new_n462), .A3(new_n464), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n468), .A2(KEYINPUT78), .A3(G179), .A4(new_n442), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT78), .ZN(new_n470));
  INV_X1    g0270(.A(new_n442), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n459), .A2(G179), .A3(new_n462), .A4(new_n464), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n357), .B1(new_n437), .B2(new_n441), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT21), .ZN(new_n475));
  AND3_X1   g0275(.A1(new_n465), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n475), .B1(new_n465), .B2(new_n474), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n469), .B(new_n473), .C1(new_n476), .C2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n230), .A2(G1698), .ZN(new_n479));
  OAI221_X1 g0279(.A(new_n479), .B1(G250), .B2(G1698), .C1(new_n301), .C2(new_n302), .ZN(new_n480));
  INV_X1    g0280(.A(G294), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n480), .B1(new_n267), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(new_n305), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n463), .A2(G264), .A3(new_n296), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT73), .ZN(new_n486));
  NOR3_X1   g0286(.A1(new_n449), .A2(new_n450), .A3(KEYINPUT72), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n454), .B1(new_n453), .B2(new_n455), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n486), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n451), .A2(KEYINPUT73), .A3(new_n456), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n446), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n357), .B1(new_n485), .B2(new_n491), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n459), .A2(new_n308), .A3(new_n483), .A4(new_n484), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  OAI21_X1  g0294(.A(KEYINPUT23), .B1(new_n223), .B2(G107), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT23), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n496), .A2(new_n209), .A3(G20), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n223), .A2(G33), .A3(G116), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n495), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT79), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n495), .A2(new_n497), .A3(new_n498), .A4(KEYINPUT79), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n223), .B(G87), .C1(new_n301), .C2(new_n302), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(KEYINPUT22), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT22), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n345), .A2(new_n506), .A3(new_n223), .A4(G87), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n503), .A2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT80), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n503), .A2(new_n508), .A3(KEYINPUT80), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n511), .A2(KEYINPUT24), .A3(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT24), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n509), .A2(new_n510), .A3(new_n514), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n513), .A2(new_n262), .A3(new_n515), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n286), .B(new_n209), .C1(KEYINPUT81), .C2(KEYINPUT25), .ZN(new_n517));
  NAND2_X1  g0317(.A1(KEYINPUT81), .A2(KEYINPUT25), .ZN(new_n518));
  OR2_X1    g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n517), .A2(new_n518), .ZN(new_n520));
  AOI22_X1  g0320(.A1(new_n519), .A2(new_n520), .B1(G107), .B2(new_n440), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n494), .B1(new_n516), .B2(new_n521), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n478), .A2(new_n522), .ZN(new_n523));
  OAI21_X1  g0323(.A(G244), .B1(new_n301), .B2(new_n302), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT4), .ZN(new_n525));
  AOI22_X1  g0325(.A1(new_n524), .A2(new_n525), .B1(G33), .B2(G283), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n345), .A2(KEYINPUT4), .A3(G244), .A4(new_n346), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n525), .B1(new_n345), .B2(G250), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n526), .B(new_n527), .C1(new_n346), .C2(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n491), .B1(new_n305), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n463), .A2(G257), .A3(new_n296), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n530), .A2(new_n308), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n529), .A2(new_n305), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n533), .A2(new_n459), .A3(new_n531), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(new_n357), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n223), .A2(new_n267), .A3(G77), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n209), .B1(new_n272), .B2(new_n273), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n536), .B1(new_n537), .B2(KEYINPUT71), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT6), .ZN(new_n539));
  INV_X1    g0339(.A(G97), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n540), .A2(new_n209), .ZN(new_n541));
  NOR2_X1   g0341(.A1(G97), .A2(G107), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n539), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n209), .A2(KEYINPUT6), .A3(G97), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(G20), .ZN(new_n546));
  INV_X1    g0346(.A(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT71), .ZN(new_n548));
  AOI211_X1 g0348(.A(new_n548), .B(new_n209), .C1(new_n272), .C2(new_n273), .ZN(new_n549));
  NOR3_X1   g0349(.A1(new_n538), .A2(new_n547), .A3(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(new_n262), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n440), .A2(G97), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n286), .A2(new_n540), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n532), .B(new_n535), .C1(new_n552), .C2(new_n555), .ZN(new_n556));
  AND2_X1   g0356(.A1(new_n483), .A2(new_n484), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(new_n459), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(G200), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n557), .A2(G190), .A3(new_n459), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n516), .A2(new_n559), .A3(new_n521), .A4(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n274), .A2(G107), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(new_n548), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n537), .A2(KEYINPUT71), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n563), .A2(new_n546), .A3(new_n564), .A4(new_n536), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n555), .B1(new_n565), .B2(new_n262), .ZN(new_n566));
  AOI21_X1  g0366(.A(G200), .B1(new_n530), .B2(new_n531), .ZN(new_n567));
  AND4_X1   g0367(.A1(new_n327), .A2(new_n533), .A3(new_n459), .A4(new_n531), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n566), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n207), .A2(new_n540), .A3(new_n209), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n349), .A2(new_n223), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n570), .A2(new_n571), .A3(KEYINPUT19), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n223), .B(G68), .C1(new_n301), .C2(new_n302), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT19), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n574), .B1(new_n362), .B2(new_n540), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n572), .A2(new_n573), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(new_n262), .ZN(new_n577));
  INV_X1    g0377(.A(new_n386), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n440), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n386), .A2(new_n286), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n577), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(KEYINPUT76), .ZN(new_n582));
  AOI22_X1  g0382(.A1(new_n576), .A2(new_n262), .B1(new_n386), .B2(new_n286), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT76), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n583), .A2(new_n584), .A3(new_n579), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n218), .A2(new_n346), .ZN(new_n586));
  OAI221_X1 g0386(.A(new_n586), .B1(G244), .B2(new_n346), .C1(new_n301), .C2(new_n302), .ZN(new_n587));
  NAND2_X1  g0387(.A1(G33), .A2(G116), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(new_n305), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT75), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n450), .A2(new_n591), .A3(G250), .ZN(new_n592));
  AOI21_X1  g0392(.A(G274), .B1(KEYINPUT75), .B2(G250), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n592), .B1(new_n450), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n296), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n590), .A2(new_n595), .ZN(new_n596));
  AOI22_X1  g0396(.A1(new_n582), .A2(new_n585), .B1(new_n357), .B2(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n590), .A2(new_n308), .A3(new_n595), .ZN(new_n598));
  AND3_X1   g0398(.A1(new_n440), .A2(KEYINPUT77), .A3(G87), .ZN(new_n599));
  AOI21_X1  g0399(.A(KEYINPUT77), .B1(new_n440), .B2(G87), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n583), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(new_n601), .ZN(new_n602));
  AND2_X1   g0402(.A1(new_n594), .A2(new_n296), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n344), .B1(new_n588), .B2(new_n587), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n396), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n590), .A2(G190), .A3(new_n595), .ZN(new_n606));
  AND2_X1   g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  AOI22_X1  g0407(.A1(new_n597), .A2(new_n598), .B1(new_n602), .B2(new_n607), .ZN(new_n608));
  AND4_X1   g0408(.A1(new_n556), .A2(new_n561), .A3(new_n569), .A4(new_n608), .ZN(new_n609));
  AND4_X1   g0409(.A1(new_n428), .A2(new_n467), .A3(new_n523), .A4(new_n609), .ZN(G372));
  NAND2_X1  g0410(.A1(new_n332), .A2(new_n335), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n337), .B1(new_n611), .B2(KEYINPUT17), .ZN(new_n612));
  INV_X1    g0412(.A(new_n394), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n378), .A2(new_n613), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n612), .B1(new_n375), .B2(new_n614), .ZN(new_n615));
  AND2_X1   g0415(.A1(new_n312), .A2(new_n313), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n422), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  AND2_X1   g0417(.A1(new_n617), .A2(new_n424), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n532), .A2(new_n535), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n619), .A2(new_n566), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n620), .A2(KEYINPUT26), .A3(new_n608), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT26), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n582), .A2(new_n585), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n596), .A2(new_n357), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n623), .A2(new_n624), .A3(new_n598), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n607), .A2(new_n602), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n622), .B1(new_n556), .B2(new_n627), .ZN(new_n628));
  AOI22_X1  g0428(.A1(new_n621), .A2(new_n628), .B1(new_n597), .B2(new_n598), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n556), .A2(new_n561), .A3(new_n569), .A4(new_n608), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n629), .B1(new_n523), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n428), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n618), .A2(new_n632), .ZN(G369));
  INV_X1    g0433(.A(G13), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n634), .A2(G20), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(new_n222), .ZN(new_n636));
  OR2_X1    g0436(.A1(new_n636), .A2(KEYINPUT27), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(KEYINPUT27), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n637), .A2(G213), .A3(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(G343), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n471), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g0443(.A(new_n478), .B(new_n643), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n644), .A2(new_n467), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(G330), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n516), .A2(new_n521), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(new_n641), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(new_n561), .ZN(new_n649));
  INV_X1    g0449(.A(new_n494), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n522), .A2(new_n642), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n646), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g0455(.A(new_n655), .B(KEYINPUT82), .Z(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n478), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n658), .A2(new_n641), .ZN(new_n659));
  AOI22_X1  g0459(.A1(new_n652), .A2(new_n659), .B1(new_n522), .B2(new_n642), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n657), .A2(new_n660), .ZN(G399));
  NAND2_X1  g0461(.A1(new_n228), .A2(new_n448), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(G1), .ZN(new_n663));
  OR2_X1    g0463(.A1(new_n570), .A2(G116), .ZN(new_n664));
  OAI22_X1  g0464(.A1(new_n663), .A2(new_n664), .B1(new_n240), .B2(new_n662), .ZN(new_n665));
  XNOR2_X1  g0465(.A(new_n665), .B(KEYINPUT28), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT29), .ZN(new_n667));
  AOI21_X1  g0467(.A(KEYINPUT85), .B1(new_n658), .B2(new_n651), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT85), .ZN(new_n669));
  NOR3_X1   g0469(.A1(new_n478), .A2(new_n522), .A3(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n609), .B1(new_n668), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(KEYINPUT86), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT86), .ZN(new_n673));
  OAI211_X1 g0473(.A(new_n673), .B(new_n609), .C1(new_n668), .C2(new_n670), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n672), .A2(new_n629), .A3(new_n674), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n667), .B1(new_n675), .B2(new_n642), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n631), .A2(new_n642), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n677), .A2(KEYINPUT29), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n534), .A2(new_n485), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n472), .A2(new_n596), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT30), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n534), .A2(new_n465), .A3(new_n596), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n558), .A2(new_n308), .ZN(new_n686));
  OR2_X1    g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(KEYINPUT83), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n680), .A2(KEYINPUT30), .A3(new_n681), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT83), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n684), .A2(new_n687), .A3(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n689), .A2(new_n690), .A3(new_n692), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n693), .A2(KEYINPUT31), .A3(new_n641), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  OAI21_X1  g0495(.A(KEYINPUT84), .B1(new_n685), .B2(new_n686), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(new_n690), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n685), .A2(new_n686), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT84), .ZN(new_n700));
  AOI22_X1  g0500(.A1(new_n699), .A2(new_n700), .B1(new_n682), .B2(new_n683), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n642), .B1(new_n698), .B2(new_n701), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n609), .A2(new_n467), .A3(new_n523), .A4(new_n642), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n702), .B1(new_n703), .B2(KEYINPUT31), .ZN(new_n704));
  OAI21_X1  g0504(.A(G330), .B1(new_n695), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n679), .A2(new_n705), .ZN(new_n706));
  XOR2_X1   g0506(.A(new_n706), .B(KEYINPUT87), .Z(new_n707));
  OAI21_X1  g0507(.A(new_n666), .B1(new_n707), .B2(G1), .ZN(G364));
  AOI21_X1  g0508(.A(new_n663), .B1(G45), .B2(new_n635), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n223), .A2(new_n327), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n396), .A2(new_n308), .A3(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(G303), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n223), .A2(new_n308), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n715), .A2(new_n327), .A3(G200), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(G317), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(KEYINPUT33), .ZN(new_n719));
  OR2_X1    g0519(.A1(new_n718), .A2(KEYINPUT33), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n717), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n308), .A2(G200), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n711), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n345), .B1(new_n724), .B2(G322), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n223), .A2(G190), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(new_n722), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(G311), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n721), .A2(new_n725), .A3(new_n729), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n715), .A2(G190), .A3(G200), .ZN(new_n731));
  OR2_X1    g0531(.A1(new_n731), .A2(KEYINPUT88), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(KEYINPUT88), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g0534(.A(new_n734), .B(KEYINPUT89), .ZN(new_n735));
  AOI211_X1 g0535(.A(new_n714), .B(new_n730), .C1(new_n735), .C2(G326), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n396), .A2(new_n308), .A3(new_n726), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(G179), .A2(G200), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n726), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  AOI22_X1  g0541(.A1(new_n738), .A2(G283), .B1(G329), .B2(new_n741), .ZN(new_n742));
  XOR2_X1   g0542(.A(new_n742), .B(KEYINPUT90), .Z(new_n743));
  AOI21_X1  g0543(.A(new_n223), .B1(new_n739), .B2(G190), .ZN(new_n744));
  OAI211_X1 g0544(.A(new_n736), .B(new_n743), .C1(new_n481), .C2(new_n744), .ZN(new_n745));
  XOR2_X1   g0545(.A(new_n745), .B(KEYINPUT91), .Z(new_n746));
  OAI22_X1  g0546(.A1(new_n716), .A2(new_n217), .B1(new_n744), .B2(new_n540), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n747), .B1(new_n734), .B2(G50), .ZN(new_n748));
  INV_X1    g0548(.A(G58), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n345), .B1(new_n723), .B2(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n750), .B1(G77), .B2(new_n728), .ZN(new_n751));
  INV_X1    g0551(.A(new_n712), .ZN(new_n752));
  AOI22_X1  g0552(.A1(G87), .A2(new_n752), .B1(new_n738), .B2(G107), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n748), .A2(new_n751), .A3(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n741), .A2(G159), .ZN(new_n755));
  XNOR2_X1  g0555(.A(new_n755), .B(KEYINPUT32), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n746), .B1(new_n754), .B2(new_n756), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n237), .B1(G20), .B2(new_n357), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n710), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n229), .A2(new_n345), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n241), .A2(new_n452), .ZN(new_n761));
  OAI211_X1 g0561(.A(new_n760), .B(new_n761), .C1(new_n256), .C2(new_n452), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n228), .A2(G355), .A3(new_n345), .ZN(new_n763));
  OAI211_X1 g0563(.A(new_n762), .B(new_n763), .C1(G116), .C2(new_n228), .ZN(new_n764));
  NOR2_X1   g0564(.A1(G13), .A2(G33), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(G20), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n758), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n764), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n767), .ZN(new_n770));
  OAI211_X1 g0570(.A(new_n759), .B(new_n769), .C1(new_n645), .C2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n645), .A2(G330), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n646), .A2(new_n710), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n771), .B1(new_n772), .B2(new_n773), .ZN(G396));
  NOR2_X1   g0574(.A1(new_n737), .A2(new_n207), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n775), .B1(G311), .B2(new_n741), .ZN(new_n776));
  XNOR2_X1  g0576(.A(new_n776), .B(KEYINPUT92), .ZN(new_n777));
  INV_X1    g0577(.A(new_n744), .ZN(new_n778));
  AOI22_X1  g0578(.A1(new_n717), .A2(G283), .B1(new_n778), .B2(G97), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n345), .B1(new_n724), .B2(G294), .ZN(new_n780));
  OAI211_X1 g0580(.A(new_n779), .B(new_n780), .C1(new_n209), .C2(new_n712), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n781), .B1(G303), .B2(new_n734), .ZN(new_n782));
  OAI211_X1 g0582(.A(new_n777), .B(new_n782), .C1(new_n431), .C2(new_n727), .ZN(new_n783));
  AOI22_X1  g0583(.A1(new_n717), .A2(G150), .B1(new_n724), .B2(G143), .ZN(new_n784));
  INV_X1    g0584(.A(new_n734), .ZN(new_n785));
  INV_X1    g0585(.A(G137), .ZN(new_n786));
  OAI221_X1 g0586(.A(new_n784), .B1(new_n277), .B2(new_n727), .C1(new_n785), .C2(new_n786), .ZN(new_n787));
  XNOR2_X1  g0587(.A(new_n787), .B(KEYINPUT34), .ZN(new_n788));
  AOI22_X1  g0588(.A1(new_n738), .A2(G68), .B1(G58), .B2(new_n778), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n316), .B1(new_n741), .B2(G132), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n791), .B1(new_n202), .B2(new_n712), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n783), .B1(new_n790), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n758), .A2(new_n765), .ZN(new_n794));
  AOI22_X1  g0594(.A1(new_n793), .A2(new_n758), .B1(new_n363), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n392), .A2(new_n641), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n403), .A2(new_n394), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n797), .A2(KEYINPUT93), .ZN(new_n798));
  INV_X1    g0598(.A(KEYINPUT93), .ZN(new_n799));
  NAND4_X1  g0599(.A1(new_n403), .A2(new_n799), .A3(new_n394), .A4(new_n796), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n613), .A2(new_n641), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  OAI211_X1 g0603(.A(new_n795), .B(new_n709), .C1(new_n803), .C2(new_n766), .ZN(new_n804));
  AND2_X1   g0604(.A1(new_n798), .A2(new_n800), .ZN(new_n805));
  AOI21_X1  g0605(.A(KEYINPUT26), .B1(new_n620), .B2(new_n608), .ZN(new_n806));
  NOR3_X1   g0606(.A1(new_n556), .A2(new_n627), .A3(new_n622), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n625), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n630), .A2(new_n523), .ZN(new_n809));
  OAI211_X1 g0609(.A(new_n642), .B(new_n805), .C1(new_n808), .C2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n677), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n810), .B1(new_n811), .B2(new_n803), .ZN(new_n812));
  XNOR2_X1  g0612(.A(new_n812), .B(new_n705), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n804), .B1(new_n813), .B2(new_n709), .ZN(G384));
  OAI21_X1  g0614(.A(new_n428), .B1(new_n676), .B2(new_n678), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n815), .A2(new_n618), .ZN(new_n816));
  XNOR2_X1  g0616(.A(new_n816), .B(KEYINPUT94), .ZN(new_n817));
  INV_X1    g0617(.A(KEYINPUT39), .ZN(new_n818));
  INV_X1    g0618(.A(new_n639), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n291), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n821), .B1(new_n612), .B2(new_n616), .ZN(new_n822));
  XNOR2_X1  g0622(.A(new_n333), .B(KEYINPUT70), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n310), .A2(new_n820), .ZN(new_n824));
  OAI21_X1  g0624(.A(KEYINPUT37), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  AND2_X1   g0625(.A1(new_n310), .A2(new_n820), .ZN(new_n826));
  INV_X1    g0626(.A(KEYINPUT37), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n826), .A2(new_n827), .A3(new_n611), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n825), .A2(new_n828), .ZN(new_n829));
  AND3_X1   g0629(.A1(new_n822), .A2(KEYINPUT38), .A3(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n333), .ZN(new_n831));
  OAI21_X1  g0631(.A(KEYINPUT37), .B1(new_n824), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n828), .A2(new_n832), .ZN(new_n833));
  AOI21_X1  g0633(.A(KEYINPUT38), .B1(new_n822), .B2(new_n833), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n818), .B1(new_n830), .B2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT38), .ZN(new_n836));
  INV_X1    g0636(.A(new_n337), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n837), .B1(new_n823), .B2(new_n315), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n820), .B1(new_n838), .B2(new_n314), .ZN(new_n839));
  NOR3_X1   g0639(.A1(new_n823), .A2(KEYINPUT37), .A3(new_n824), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n827), .B1(new_n826), .B2(new_n611), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n836), .B1(new_n839), .B2(new_n842), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n822), .A2(KEYINPUT38), .A3(new_n829), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n843), .A2(KEYINPUT39), .A3(new_n844), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n375), .A2(new_n641), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n835), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n616), .A2(new_n639), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n374), .A2(new_n641), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n375), .A2(new_n378), .A3(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n378), .ZN(new_n851));
  OAI211_X1 g0651(.A(new_n374), .B(new_n641), .C1(new_n851), .C2(new_n361), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n613), .A2(new_n642), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n810), .A2(new_n854), .ZN(new_n855));
  AOI21_X1  g0655(.A(KEYINPUT38), .B1(new_n822), .B2(new_n829), .ZN(new_n856));
  OAI211_X1 g0656(.A(new_n853), .B(new_n855), .C1(new_n830), .C2(new_n856), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n847), .A2(new_n848), .A3(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  XNOR2_X1  g0659(.A(new_n817), .B(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n853), .A2(new_n803), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n703), .A2(KEYINPUT31), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n684), .B1(new_n687), .B2(KEYINPUT84), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n641), .B1(new_n863), .B2(new_n697), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT31), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n861), .B1(new_n865), .B2(new_n868), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n869), .B1(new_n856), .B2(new_n830), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT40), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  AOI22_X1  g0672(.A1(new_n338), .A2(new_n821), .B1(new_n828), .B2(new_n832), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n844), .B1(KEYINPUT38), .B2(new_n873), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n874), .A2(new_n869), .A3(KEYINPUT40), .ZN(new_n875));
  AND2_X1   g0675(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n867), .B1(new_n862), .B2(new_n864), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n877), .A2(new_n427), .ZN(new_n878));
  XOR2_X1   g0678(.A(new_n876), .B(new_n878), .Z(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(G330), .ZN(new_n880));
  XNOR2_X1  g0680(.A(new_n860), .B(new_n880), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n881), .B1(new_n222), .B2(new_n635), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n431), .B1(new_n545), .B2(KEYINPUT35), .ZN(new_n883));
  OAI211_X1 g0683(.A(new_n883), .B(new_n238), .C1(KEYINPUT35), .C2(new_n545), .ZN(new_n884));
  XNOR2_X1  g0684(.A(new_n884), .B(KEYINPUT36), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n264), .A2(G77), .ZN(new_n886));
  OAI22_X1  g0686(.A1(new_n240), .A2(new_n886), .B1(G50), .B2(new_n217), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n887), .A2(G1), .A3(new_n634), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n882), .A2(new_n885), .A3(new_n888), .ZN(G367));
  AOI22_X1  g0689(.A1(new_n735), .A2(G311), .B1(G303), .B2(new_n724), .ZN(new_n890));
  XNOR2_X1  g0690(.A(new_n890), .B(KEYINPUT100), .ZN(new_n891));
  OAI221_X1 g0691(.A(new_n316), .B1(new_n718), .B2(new_n740), .C1(new_n737), .C2(new_n540), .ZN(new_n892));
  XOR2_X1   g0692(.A(new_n892), .B(KEYINPUT102), .Z(new_n893));
  INV_X1    g0693(.A(KEYINPUT101), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT46), .ZN(new_n895));
  NOR4_X1   g0695(.A1(new_n712), .A2(new_n894), .A3(new_n895), .A4(new_n431), .ZN(new_n896));
  AOI22_X1  g0696(.A1(new_n717), .A2(G294), .B1(new_n778), .B2(G107), .ZN(new_n897));
  OAI22_X1  g0697(.A1(new_n712), .A2(new_n431), .B1(new_n894), .B2(new_n895), .ZN(new_n898));
  OAI211_X1 g0698(.A(new_n897), .B(new_n898), .C1(KEYINPUT101), .C2(KEYINPUT46), .ZN(new_n899));
  NOR3_X1   g0699(.A1(new_n893), .A2(new_n896), .A3(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(G283), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n891), .B(new_n900), .C1(new_n901), .C2(new_n727), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n723), .A2(new_n406), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n735), .A2(G143), .ZN(new_n904));
  AOI22_X1  g0704(.A1(G58), .A2(new_n752), .B1(new_n738), .B2(G77), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n744), .A2(new_n217), .ZN(new_n906));
  OAI221_X1 g0706(.A(new_n345), .B1(new_n740), .B2(new_n786), .C1(new_n202), .C2(new_n727), .ZN(new_n907));
  AOI211_X1 g0707(.A(new_n906), .B(new_n907), .C1(G159), .C2(new_n717), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n904), .A2(new_n905), .A3(new_n908), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n902), .B1(new_n903), .B2(new_n909), .ZN(new_n910));
  XNOR2_X1  g0710(.A(new_n910), .B(KEYINPUT47), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n710), .B1(new_n911), .B2(new_n758), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n760), .A2(new_n252), .ZN(new_n913));
  OAI211_X1 g0713(.A(new_n913), .B(new_n768), .C1(new_n228), .C2(new_n386), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n914), .B(KEYINPUT99), .ZN(new_n915));
  NOR3_X1   g0715(.A1(new_n625), .A2(new_n602), .A3(new_n642), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT95), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n602), .A2(new_n642), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n917), .B1(new_n627), .B2(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n918), .B1(new_n921), .B2(new_n916), .ZN(new_n922));
  OAI211_X1 g0722(.A(new_n912), .B(new_n915), .C1(new_n770), .C2(new_n922), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n556), .B(new_n569), .C1(new_n566), .C2(new_n642), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n924), .B1(new_n556), .B2(new_n642), .ZN(new_n925));
  NAND4_X1  g0725(.A1(new_n925), .A2(new_n653), .A3(new_n652), .A4(new_n659), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n926), .B(KEYINPUT42), .ZN(new_n927));
  OR2_X1    g0727(.A1(new_n924), .A2(new_n651), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n641), .B1(new_n928), .B2(new_n556), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT96), .ZN(new_n931));
  OR3_X1    g0731(.A1(new_n930), .A2(new_n931), .A3(KEYINPUT43), .ZN(new_n932));
  OAI21_X1  g0732(.A(KEYINPUT43), .B1(new_n930), .B2(new_n931), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n934), .B1(new_n929), .B2(new_n927), .ZN(new_n935));
  MUX2_X1   g0735(.A(new_n934), .B(new_n935), .S(new_n922), .Z(new_n936));
  NAND2_X1  g0736(.A1(new_n656), .A2(new_n925), .ZN(new_n937));
  XOR2_X1   g0737(.A(new_n936), .B(new_n937), .Z(new_n938));
  NAND2_X1  g0738(.A1(new_n635), .A2(G45), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(G1), .ZN(new_n940));
  XOR2_X1   g0740(.A(new_n940), .B(KEYINPUT98), .Z(new_n941));
  NAND2_X1  g0741(.A1(new_n660), .A2(new_n925), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT97), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n942), .B(new_n943), .ZN(new_n944));
  OR2_X1    g0744(.A1(new_n944), .A2(KEYINPUT45), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n660), .A2(new_n925), .ZN(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  AOI22_X1  g0747(.A1(new_n944), .A2(KEYINPUT45), .B1(KEYINPUT44), .B2(new_n947), .ZN(new_n948));
  OR2_X1    g0748(.A1(new_n947), .A2(KEYINPUT44), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n945), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  OR2_X1    g0750(.A1(new_n950), .A2(new_n656), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(new_n656), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  XOR2_X1   g0753(.A(new_n654), .B(new_n659), .Z(new_n954));
  XNOR2_X1  g0754(.A(new_n954), .B(new_n646), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n707), .B1(new_n953), .B2(new_n955), .ZN(new_n956));
  XOR2_X1   g0756(.A(new_n662), .B(KEYINPUT41), .Z(new_n957));
  AOI21_X1  g0757(.A(new_n941), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n923), .B1(new_n938), .B2(new_n958), .ZN(G387));
  INV_X1    g0759(.A(new_n955), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n707), .A2(new_n960), .ZN(new_n961));
  XOR2_X1   g0761(.A(new_n662), .B(KEYINPUT105), .Z(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n964), .B(KEYINPUT106), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(new_n707), .B2(new_n960), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n960), .A2(new_n941), .ZN(new_n967));
  AOI22_X1  g0767(.A1(new_n717), .A2(G311), .B1(new_n724), .B2(G317), .ZN(new_n968));
  INV_X1    g0768(.A(new_n735), .ZN(new_n969));
  XOR2_X1   g0769(.A(KEYINPUT104), .B(G322), .Z(new_n970));
  OAI221_X1 g0770(.A(new_n968), .B1(new_n713), .B2(new_n727), .C1(new_n969), .C2(new_n970), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n971), .B(KEYINPUT48), .ZN(new_n972));
  OAI221_X1 g0772(.A(new_n972), .B1(new_n901), .B2(new_n744), .C1(new_n481), .C2(new_n712), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT49), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n973), .A2(new_n974), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n345), .B1(new_n738), .B2(G116), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  AOI211_X1 g0778(.A(new_n975), .B(new_n978), .C1(G326), .C2(new_n741), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n778), .A2(new_n578), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n980), .B1(new_n284), .B2(new_n716), .ZN(new_n981));
  OAI221_X1 g0781(.A(new_n345), .B1(new_n740), .B2(new_n406), .C1(new_n217), .C2(new_n727), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n737), .A2(new_n540), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n712), .A2(new_n363), .ZN(new_n984));
  NOR4_X1   g0784(.A1(new_n981), .A2(new_n982), .A3(new_n983), .A4(new_n984), .ZN(new_n985));
  OAI221_X1 g0785(.A(new_n985), .B1(new_n202), .B2(new_n723), .C1(new_n277), .C2(new_n785), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n986), .B(KEYINPUT103), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n758), .B1(new_n979), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n289), .A2(new_n202), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n664), .B1(new_n989), .B2(KEYINPUT50), .ZN(new_n990));
  OAI211_X1 g0790(.A(new_n990), .B(new_n452), .C1(KEYINPUT50), .C2(new_n989), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n991), .B1(G68), .B2(G77), .ZN(new_n992));
  INV_X1    g0792(.A(new_n248), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n760), .B1(new_n993), .B2(new_n452), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n228), .A2(new_n664), .A3(new_n345), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n992), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n228), .A2(G107), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n768), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n654), .A2(new_n767), .ZN(new_n999));
  NAND4_X1  g0799(.A1(new_n988), .A2(new_n709), .A3(new_n998), .A4(new_n999), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n966), .A2(new_n967), .A3(new_n1000), .ZN(G393));
  INV_X1    g0801(.A(new_n961), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n953), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n962), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1004), .B1(new_n1003), .B2(new_n1002), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1003), .A2(new_n941), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n316), .B1(new_n970), .B2(new_n740), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(new_n734), .A2(G317), .B1(G311), .B2(new_n724), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT52), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n716), .A2(new_n713), .B1(new_n744), .B2(new_n431), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1010), .B1(G294), .B2(new_n728), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n1011), .ZN(new_n1012));
  AOI211_X1 g0812(.A(new_n1007), .B(new_n1009), .C1(KEYINPUT107), .C2(new_n1012), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(G107), .A2(new_n738), .B1(new_n752), .B2(G283), .ZN(new_n1014));
  OAI211_X1 g0814(.A(new_n1013), .B(new_n1014), .C1(KEYINPUT107), .C2(new_n1012), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n734), .A2(G150), .B1(G159), .B2(new_n724), .ZN(new_n1016));
  XOR2_X1   g0816(.A(new_n1016), .B(KEYINPUT51), .Z(new_n1017));
  AOI21_X1  g0817(.A(new_n316), .B1(new_n741), .B2(G143), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n1018), .B1(new_n202), .B2(new_n716), .C1(new_n363), .C2(new_n744), .ZN(new_n1019));
  AOI211_X1 g0819(.A(new_n775), .B(new_n1019), .C1(G68), .C2(new_n752), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n1017), .B(new_n1020), .C1(new_n284), .C2(new_n727), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1015), .A2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n710), .B1(new_n1022), .B2(new_n758), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n760), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n768), .B1(new_n540), .B2(new_n228), .C1(new_n1024), .C2(new_n259), .ZN(new_n1025));
  OAI211_X1 g0825(.A(new_n1023), .B(new_n1025), .C1(new_n770), .C2(new_n925), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1005), .A2(new_n1006), .A3(new_n1026), .ZN(G390));
  INV_X1    g0827(.A(new_n853), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n803), .A2(G330), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1028), .B1(new_n877), .B2(new_n1029), .ZN(new_n1030));
  AND2_X1   g0830(.A1(new_n803), .A2(G330), .ZN(new_n1031));
  OAI211_X1 g0831(.A(new_n1031), .B(new_n853), .C1(new_n695), .C2(new_n704), .ZN(new_n1032));
  AND2_X1   g0832(.A1(new_n1030), .A2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n675), .A2(new_n642), .A3(new_n805), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1034), .A2(new_n854), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n1035), .ZN(new_n1036));
  OAI211_X1 g0836(.A(new_n1031), .B(new_n853), .C1(new_n704), .C2(new_n867), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1029), .B1(new_n865), .B2(new_n694), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1037), .B1(new_n1038), .B2(new_n853), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n1033), .A2(new_n1036), .B1(new_n1039), .B2(new_n855), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n878), .A2(G330), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n815), .A2(new_n618), .A3(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(KEYINPUT108), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n855), .A2(new_n853), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n846), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NOR3_X1   g0846(.A1(new_n830), .A2(new_n856), .A3(new_n818), .ZN(new_n1047));
  AND2_X1   g0847(.A1(new_n828), .A2(new_n832), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n836), .B1(new_n839), .B2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g0849(.A(KEYINPUT39), .B1(new_n1049), .B2(new_n844), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1046), .B1(new_n1047), .B2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1028), .B1(new_n1034), .B2(new_n854), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1045), .B1(new_n830), .B2(new_n834), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n1051), .B(new_n1032), .C1(new_n1052), .C2(new_n1053), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n1037), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1053), .B1(new_n1035), .B2(new_n853), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n846), .B1(new_n855), .B2(new_n853), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1057), .B1(new_n835), .B2(new_n845), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1055), .B1(new_n1056), .B2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1043), .A2(new_n1054), .A3(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1054), .A2(new_n1059), .ZN(new_n1061));
  INV_X1    g0861(.A(KEYINPUT108), .ZN(new_n1062));
  AND3_X1   g0862(.A1(new_n815), .A2(new_n618), .A3(new_n1041), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1039), .A2(new_n855), .ZN(new_n1064));
  NAND4_X1  g0864(.A1(new_n1030), .A2(new_n1034), .A3(new_n1032), .A4(new_n854), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1062), .B1(new_n1063), .B2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1061), .A2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1060), .A2(new_n1068), .A3(new_n963), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1054), .A2(new_n1059), .A3(new_n941), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n765), .B1(new_n1047), .B2(new_n1050), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n217), .A2(new_n737), .B1(new_n712), .B2(new_n207), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n316), .B1(new_n740), .B2(new_n481), .C1(new_n540), .C2(new_n727), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n716), .A2(new_n209), .B1(new_n744), .B2(new_n363), .ZN(new_n1074));
  NOR3_X1   g0874(.A1(new_n1072), .A2(new_n1073), .A3(new_n1074), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n1075), .B1(new_n431), .B2(new_n723), .C1(new_n901), .C2(new_n785), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n734), .A2(G128), .B1(G132), .B2(new_n724), .ZN(new_n1077));
  XOR2_X1   g0877(.A(new_n1077), .B(KEYINPUT109), .Z(new_n1078));
  NOR2_X1   g0878(.A1(new_n712), .A2(new_n406), .ZN(new_n1079));
  XNOR2_X1  g0879(.A(new_n1079), .B(KEYINPUT53), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n716), .A2(new_n786), .B1(new_n744), .B2(new_n277), .ZN(new_n1081));
  XOR2_X1   g0881(.A(KEYINPUT54), .B(G143), .Z(new_n1082));
  INV_X1    g0882(.A(new_n1082), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n345), .B1(new_n1083), .B2(new_n727), .ZN(new_n1084));
  AOI211_X1 g0884(.A(new_n1081), .B(new_n1084), .C1(G50), .C2(new_n738), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1078), .A2(new_n1080), .A3(new_n1085), .ZN(new_n1086));
  INV_X1    g0886(.A(G125), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n740), .A2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1076), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1089));
  XOR2_X1   g0889(.A(new_n1089), .B(KEYINPUT110), .Z(new_n1090));
  AOI21_X1  g0890(.A(new_n710), .B1(new_n1090), .B2(new_n758), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n794), .ZN(new_n1092));
  OAI211_X1 g0892(.A(new_n1071), .B(new_n1091), .C1(new_n289), .C2(new_n1092), .ZN(new_n1093));
  AND3_X1   g0893(.A1(new_n1069), .A2(new_n1070), .A3(new_n1093), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1094), .ZN(G378));
  NAND3_X1  g0895(.A1(new_n1054), .A2(new_n1059), .A3(new_n1066), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(new_n1063), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n850), .A2(new_n852), .B1(new_n801), .B2(new_n802), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1098), .B1(new_n704), .B2(new_n867), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1099), .B1(new_n843), .B2(new_n844), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n875), .B(G330), .C1(new_n1100), .C2(KEYINPUT40), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n425), .A2(KEYINPUT55), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n425), .A2(KEYINPUT55), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n410), .A2(new_n819), .ZN(new_n1105));
  XOR2_X1   g0905(.A(new_n1105), .B(KEYINPUT56), .Z(new_n1106));
  NAND3_X1  g0906(.A1(new_n1103), .A2(new_n1104), .A3(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1106), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1101), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(KEYINPUT116), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1112), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1106), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1104), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1114), .B1(new_n1115), .B2(new_n1102), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1116), .A2(new_n1107), .A3(KEYINPUT116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1113), .A2(new_n1117), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n872), .A2(new_n1118), .A3(G330), .A4(new_n875), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1111), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1120), .A2(new_n859), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1111), .A2(new_n858), .A3(new_n1119), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n1097), .A2(KEYINPUT57), .A3(new_n1121), .A4(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(KEYINPUT117), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(KEYINPUT57), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1097), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1126), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  AND3_X1   g0929(.A1(new_n1111), .A2(new_n858), .A3(new_n1119), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n858), .B1(new_n1111), .B2(new_n1119), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n1132), .A2(KEYINPUT117), .A3(KEYINPUT57), .A4(new_n1097), .ZN(new_n1133));
  NAND4_X1  g0933(.A1(new_n1125), .A2(new_n1129), .A3(new_n963), .A4(new_n1133), .ZN(new_n1134));
  OAI221_X1 g0934(.A(new_n316), .B1(new_n901), .B2(new_n740), .C1(new_n737), .C2(new_n749), .ZN(new_n1135));
  NOR3_X1   g0935(.A1(new_n1135), .A2(G41), .A3(new_n984), .ZN(new_n1136));
  XOR2_X1   g0936(.A(new_n1136), .B(KEYINPUT112), .Z(new_n1137));
  AOI21_X1  g0937(.A(new_n906), .B1(G107), .B2(new_n724), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1138), .B1(new_n540), .B2(new_n716), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1139), .B1(G116), .B2(new_n734), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n1137), .B(new_n1140), .C1(new_n386), .C2(new_n727), .ZN(new_n1141));
  INV_X1    g0941(.A(KEYINPUT58), .ZN(new_n1142));
  INV_X1    g0942(.A(KEYINPUT111), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n202), .B1(new_n301), .B2(G41), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n1141), .A2(new_n1142), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1145), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1146));
  XOR2_X1   g0946(.A(new_n1146), .B(KEYINPUT113), .Z(new_n1147));
  AOI22_X1  g0947(.A1(new_n717), .A2(G132), .B1(new_n724), .B2(G128), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1148), .B1(new_n406), .B2(new_n744), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1149), .B1(new_n752), .B2(new_n1082), .ZN(new_n1150));
  OAI221_X1 g0950(.A(new_n1150), .B1(new_n1087), .B2(new_n785), .C1(new_n786), .C2(new_n727), .ZN(new_n1151));
  XOR2_X1   g0951(.A(new_n1151), .B(KEYINPUT114), .Z(new_n1152));
  INV_X1    g0952(.A(KEYINPUT59), .ZN(new_n1153));
  OR2_X1    g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1155));
  AOI21_X1  g0955(.A(G33), .B1(new_n741), .B2(G124), .ZN(new_n1156));
  AOI21_X1  g0956(.A(G41), .B1(new_n738), .B2(G159), .ZN(new_n1157));
  NAND4_X1  g0957(.A1(new_n1154), .A2(new_n1155), .A3(new_n1156), .A4(new_n1157), .ZN(new_n1158));
  OAI211_X1 g0958(.A(new_n1147), .B(new_n1158), .C1(new_n1142), .C2(new_n1141), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT115), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(new_n1159), .B(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n710), .B1(new_n1161), .B2(new_n758), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n794), .A2(new_n202), .ZN(new_n1163));
  OAI211_X1 g0963(.A(new_n1162), .B(new_n1163), .C1(new_n766), .C2(new_n1118), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1121), .A2(new_n941), .A3(new_n1122), .ZN(new_n1165));
  AND2_X1   g0965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1134), .A2(new_n1166), .ZN(G375));
  NAND2_X1  g0967(.A1(new_n1063), .A2(new_n1066), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1168), .A2(new_n1169), .A3(new_n957), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1028), .A2(new_n765), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n734), .A2(G132), .ZN(new_n1172));
  XOR2_X1   g0972(.A(new_n1172), .B(KEYINPUT119), .Z(new_n1173));
  OAI21_X1  g0973(.A(new_n345), .B1(new_n723), .B2(new_n786), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n1083), .A2(new_n716), .B1(new_n202), .B2(new_n744), .ZN(new_n1175));
  AOI211_X1 g0975(.A(new_n1174), .B(new_n1175), .C1(G128), .C2(new_n741), .ZN(new_n1176));
  OAI221_X1 g0976(.A(new_n1176), .B1(new_n749), .B2(new_n737), .C1(new_n277), .C2(new_n712), .ZN(new_n1177));
  AOI211_X1 g0977(.A(new_n1173), .B(new_n1177), .C1(G150), .C2(new_n728), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n785), .A2(new_n481), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n345), .B1(new_n741), .B2(G303), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n717), .A2(G116), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n728), .A2(G107), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n1180), .A2(new_n1181), .A3(new_n980), .A4(new_n1182), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n723), .A2(new_n901), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n363), .A2(new_n737), .B1(new_n712), .B2(new_n540), .ZN(new_n1185));
  NOR4_X1   g0985(.A1(new_n1179), .A2(new_n1183), .A3(new_n1184), .A4(new_n1185), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n758), .B1(new_n1178), .B2(new_n1186), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n709), .B1(new_n1092), .B2(G68), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(new_n1188), .B(KEYINPUT118), .ZN(new_n1189));
  AND3_X1   g0989(.A1(new_n1171), .A2(new_n1187), .A3(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1190), .B1(new_n1066), .B2(new_n941), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1170), .A2(new_n1191), .ZN(G381));
  NOR2_X1   g0992(.A1(G375), .A2(G378), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  NOR3_X1   g0994(.A1(new_n1194), .A2(G387), .A3(G390), .ZN(new_n1195));
  NOR4_X1   g0995(.A1(G393), .A2(G396), .A3(G384), .A4(G381), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1195), .A2(new_n1196), .ZN(G407));
  OAI211_X1 g0997(.A(G407), .B(G213), .C1(G343), .C2(new_n1194), .ZN(G409));
  INV_X1    g0998(.A(KEYINPUT126), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n640), .A2(G213), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n1097), .A2(new_n957), .A3(new_n1121), .A4(new_n1122), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1201), .A2(new_n1165), .A3(new_n1164), .ZN(new_n1202));
  AND3_X1   g1002(.A1(new_n1094), .A2(KEYINPUT120), .A3(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(KEYINPUT120), .B1(new_n1094), .B2(new_n1202), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  AND3_X1   g1005(.A1(new_n1134), .A2(G378), .A3(new_n1166), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1200), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT123), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT60), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1169), .A2(new_n1210), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1040), .A2(KEYINPUT60), .A3(new_n1042), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n1211), .A2(new_n963), .A3(new_n1168), .A4(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1213), .A2(new_n1191), .ZN(new_n1214));
  XNOR2_X1  g1014(.A(new_n1214), .B(G384), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n640), .A2(G213), .A3(G2897), .ZN(new_n1216));
  XOR2_X1   g1016(.A(new_n1215), .B(new_n1216), .Z(new_n1217));
  NAND3_X1  g1017(.A1(new_n1134), .A2(G378), .A3(new_n1166), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1218), .B1(new_n1204), .B2(new_n1203), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1219), .A2(KEYINPUT123), .A3(new_n1200), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1209), .A2(new_n1217), .A3(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT125), .ZN(new_n1222));
  XNOR2_X1  g1022(.A(KEYINPUT124), .B(KEYINPUT61), .ZN(new_n1223));
  AND3_X1   g1023(.A1(new_n1221), .A2(new_n1222), .A3(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1222), .B1(new_n1221), .B2(new_n1223), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  XNOR2_X1  g1026(.A(new_n1219), .B(KEYINPUT121), .ZN(new_n1227));
  INV_X1    g1027(.A(KEYINPUT62), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1227), .A2(new_n1228), .A3(new_n1215), .A4(new_n1200), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1215), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1230), .B1(new_n1209), .B2(new_n1220), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1229), .B1(new_n1228), .B2(new_n1231), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1199), .B1(new_n1226), .B2(new_n1232), .ZN(new_n1233));
  XNOR2_X1  g1033(.A(G393), .B(G396), .ZN(new_n1234));
  NAND4_X1  g1034(.A1(G387), .A2(new_n1006), .A3(new_n1026), .A4(new_n1005), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1235), .A2(KEYINPUT122), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1234), .A2(new_n1236), .ZN(new_n1237));
  XNOR2_X1  g1037(.A(G387), .B(G390), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1238), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1237), .A2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1237), .A2(new_n1239), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(new_n1244));
  AND2_X1   g1044(.A1(new_n1219), .A2(KEYINPUT121), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n1219), .A2(KEYINPUT121), .ZN(new_n1246));
  OAI211_X1 g1046(.A(new_n1215), .B(new_n1200), .C1(new_n1245), .C2(new_n1246), .ZN(new_n1247));
  MUX2_X1   g1047(.A(new_n1247), .B(new_n1231), .S(KEYINPUT62), .Z(new_n1248));
  OAI211_X1 g1048(.A(new_n1248), .B(KEYINPUT126), .C1(new_n1225), .C2(new_n1224), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1233), .A2(new_n1244), .A3(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1227), .A2(new_n1200), .ZN(new_n1251));
  AND2_X1   g1051(.A1(new_n1251), .A2(new_n1217), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT63), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1247), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT61), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1231), .A2(KEYINPUT63), .ZN(new_n1256));
  NAND4_X1  g1056(.A1(new_n1254), .A2(new_n1243), .A3(new_n1255), .A4(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1250), .A2(new_n1257), .ZN(G405));
  NAND2_X1  g1058(.A1(G375), .A2(new_n1094), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1259), .A2(new_n1218), .ZN(new_n1260));
  XNOR2_X1  g1060(.A(new_n1260), .B(new_n1230), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1243), .A2(KEYINPUT127), .A3(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1243), .A2(KEYINPUT127), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT127), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1241), .A2(new_n1264), .A3(new_n1242), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1263), .A2(new_n1265), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1262), .B1(new_n1266), .B2(new_n1261), .ZN(G402));
endmodule


