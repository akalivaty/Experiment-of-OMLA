//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 1 0 1 0 1 0 0 1 0 1 0 1 0 0 1 0 1 0 1 0 1 0 1 0 1 0 1 0 1 0 1 1 0 1 1 1 0 1 0 0 0 1 1 0 0 1 0 0 1 1 1 0 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:01 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1282, new_n1283, new_n1284, new_n1285,
    new_n1286, new_n1287, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1353,
    new_n1354, new_n1355, new_n1356, new_n1357;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G68), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT64), .ZN(new_n213));
  OAI21_X1  g0013(.A(G50), .B1(G58), .B2(G68), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n215));
  INV_X1    g0015(.A(G77), .ZN(new_n216));
  INV_X1    g0016(.A(G244), .ZN(new_n217));
  INV_X1    g0017(.A(G107), .ZN(new_n218));
  INV_X1    g0018(.A(G264), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n221));
  INV_X1    g0021(.A(G232), .ZN(new_n222));
  INV_X1    g0022(.A(G97), .ZN(new_n223));
  INV_X1    g0023(.A(G257), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n221), .B1(new_n202), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n206), .B1(new_n220), .B2(new_n225), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n209), .B1(new_n213), .B2(new_n214), .C1(KEYINPUT1), .C2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XOR2_X1   g0028(.A(G250), .B(G257), .Z(new_n229));
  XNOR2_X1  g0029(.A(G264), .B(G270), .ZN(new_n230));
  XOR2_X1   g0030(.A(new_n229), .B(new_n230), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT65), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(new_n222), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n232), .B(new_n236), .ZN(G358));
  XOR2_X1   g0037(.A(G68), .B(G77), .Z(new_n238));
  XOR2_X1   g0038(.A(G50), .B(G58), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n240), .B(KEYINPUT66), .Z(new_n241));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G351));
  NAND2_X1  g0045(.A1(G33), .A2(G41), .ZN(new_n246));
  NAND3_X1  g0046(.A1(new_n246), .A2(G1), .A3(G13), .ZN(new_n247));
  OR2_X1    g0047(.A1(G223), .A2(G1698), .ZN(new_n248));
  INV_X1    g0048(.A(G1698), .ZN(new_n249));
  AND2_X1   g0049(.A1(KEYINPUT3), .A2(G33), .ZN(new_n250));
  NOR2_X1   g0050(.A1(KEYINPUT3), .A2(G33), .ZN(new_n251));
  OAI221_X1 g0051(.A(new_n248), .B1(G226), .B2(new_n249), .C1(new_n250), .C2(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(G33), .A2(G87), .ZN(new_n253));
  AOI21_X1  g0053(.A(new_n247), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G41), .ZN(new_n255));
  INV_X1    g0055(.A(G45), .ZN(new_n256));
  AOI21_X1  g0056(.A(G1), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n257), .A2(new_n247), .A3(G274), .ZN(new_n258));
  INV_X1    g0058(.A(G1), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n259), .B1(G41), .B2(G45), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n247), .A2(new_n260), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n258), .B1(new_n261), .B2(new_n222), .ZN(new_n262));
  INV_X1    g0062(.A(G179), .ZN(new_n263));
  NOR3_X1   g0063(.A1(new_n254), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  OR2_X1    g0064(.A1(new_n254), .A2(new_n262), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n264), .B1(G169), .B2(new_n265), .ZN(new_n266));
  NAND3_X1  g0066(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(new_n210), .ZN(new_n268));
  AND2_X1   g0068(.A1(G58), .A2(G68), .ZN(new_n269));
  NOR2_X1   g0069(.A1(G58), .A2(G68), .ZN(new_n270));
  OAI21_X1  g0070(.A(G20), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NOR2_X1   g0071(.A1(G20), .A2(G33), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G159), .ZN(new_n273));
  AND3_X1   g0073(.A1(new_n271), .A2(KEYINPUT77), .A3(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(KEYINPUT77), .B1(new_n271), .B2(new_n273), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT7), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n277), .A2(G20), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT3), .ZN(new_n279));
  INV_X1    g0079(.A(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(KEYINPUT3), .A2(G33), .ZN(new_n282));
  AND3_X1   g0082(.A1(new_n278), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  OAI21_X1  g0083(.A(KEYINPUT76), .B1(new_n250), .B2(new_n251), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT76), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n281), .A2(new_n285), .A3(new_n282), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n284), .A2(new_n286), .A3(new_n211), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n283), .B1(new_n287), .B2(new_n277), .ZN(new_n288));
  INV_X1    g0088(.A(G68), .ZN(new_n289));
  OAI211_X1 g0089(.A(new_n276), .B(KEYINPUT16), .C1(new_n288), .C2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n271), .A2(new_n273), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT77), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n271), .A2(KEYINPUT77), .A3(new_n273), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  OAI21_X1  g0095(.A(KEYINPUT67), .B1(new_n250), .B2(new_n251), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT67), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n281), .A2(new_n297), .A3(new_n282), .ZN(new_n298));
  AOI21_X1  g0098(.A(G20), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT78), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n250), .A2(new_n251), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n300), .B1(new_n301), .B2(new_n278), .ZN(new_n302));
  AND4_X1   g0102(.A1(new_n300), .A2(new_n278), .A3(new_n281), .A4(new_n282), .ZN(new_n303));
  OAI22_X1  g0103(.A1(new_n299), .A2(KEYINPUT7), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n295), .B1(new_n304), .B2(G68), .ZN(new_n305));
  OAI211_X1 g0105(.A(new_n268), .B(new_n290), .C1(new_n305), .C2(KEYINPUT16), .ZN(new_n306));
  NAND2_X1  g0106(.A1(KEYINPUT69), .A2(G58), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT8), .ZN(new_n308));
  XNOR2_X1  g0108(.A(new_n307), .B(new_n308), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n309), .B1(new_n259), .B2(G20), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n259), .A2(G13), .A3(G20), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n311), .A2(new_n210), .A3(new_n267), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(new_n311), .ZN(new_n314));
  AOI22_X1  g0114(.A1(new_n310), .A2(new_n313), .B1(new_n314), .B2(new_n309), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n266), .B1(new_n306), .B2(new_n315), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n316), .A2(KEYINPUT18), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT18), .ZN(new_n318));
  AOI211_X1 g0118(.A(new_n318), .B(new_n266), .C1(new_n306), .C2(new_n315), .ZN(new_n319));
  NOR3_X1   g0119(.A1(new_n317), .A2(new_n319), .A3(KEYINPUT79), .ZN(new_n320));
  INV_X1    g0120(.A(new_n315), .ZN(new_n321));
  AND2_X1   g0121(.A1(new_n290), .A2(new_n268), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT16), .ZN(new_n323));
  NOR3_X1   g0123(.A1(new_n250), .A2(new_n251), .A3(KEYINPUT67), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n297), .B1(new_n281), .B2(new_n282), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n211), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(new_n277), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n301), .A2(new_n278), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(KEYINPUT78), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n283), .A2(new_n300), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n289), .B1(new_n327), .B2(new_n331), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n323), .B1(new_n332), .B2(new_n295), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n321), .B1(new_n322), .B2(new_n333), .ZN(new_n334));
  OAI211_X1 g0134(.A(KEYINPUT79), .B(new_n318), .C1(new_n334), .C2(new_n266), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n254), .A2(new_n262), .ZN(new_n336));
  INV_X1    g0136(.A(G190), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n338), .B1(G200), .B2(new_n336), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n306), .A2(new_n315), .A3(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT17), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n306), .A2(KEYINPUT17), .A3(new_n315), .A4(new_n339), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n335), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n320), .A2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(new_n258), .ZN(new_n346));
  INV_X1    g0146(.A(new_n261), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n346), .B1(G226), .B2(new_n347), .ZN(new_n348));
  NAND4_X1  g0148(.A1(new_n296), .A2(new_n298), .A3(G223), .A4(G1698), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n324), .A2(new_n325), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n349), .B1(new_n350), .B2(new_n216), .ZN(new_n351));
  NAND4_X1  g0151(.A1(new_n296), .A2(new_n298), .A3(G222), .A4(new_n249), .ZN(new_n352));
  OR2_X1    g0152(.A1(new_n352), .A2(KEYINPUT68), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(KEYINPUT68), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n351), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n348), .B1(new_n355), .B2(new_n247), .ZN(new_n356));
  INV_X1    g0156(.A(G169), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  OAI21_X1  g0158(.A(G20), .B1(new_n203), .B2(G68), .ZN(new_n359));
  INV_X1    g0159(.A(G150), .ZN(new_n360));
  INV_X1    g0160(.A(new_n272), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n211), .A2(G33), .ZN(new_n362));
  OAI221_X1 g0162(.A(new_n359), .B1(new_n360), .B2(new_n361), .C1(new_n309), .C2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(new_n268), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n201), .B1(new_n259), .B2(G20), .ZN(new_n365));
  AOI22_X1  g0165(.A1(new_n313), .A2(new_n365), .B1(new_n201), .B2(new_n314), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  OAI211_X1 g0167(.A(new_n263), .B(new_n348), .C1(new_n355), .C2(new_n247), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n358), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT71), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n216), .B1(new_n259), .B2(G20), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n313), .A2(new_n372), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n373), .B1(G77), .B2(new_n311), .ZN(new_n374));
  NAND2_X1  g0174(.A1(G20), .A2(G77), .ZN(new_n375));
  XNOR2_X1  g0175(.A(KEYINPUT8), .B(G58), .ZN(new_n376));
  XNOR2_X1  g0176(.A(KEYINPUT15), .B(G87), .ZN(new_n377));
  OAI221_X1 g0177(.A(new_n375), .B1(new_n376), .B2(new_n361), .C1(new_n362), .C2(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n374), .B1(new_n378), .B2(new_n268), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n296), .A2(new_n298), .ZN(new_n380));
  XNOR2_X1  g0180(.A(KEYINPUT70), .B(G107), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n247), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NOR2_X1   g0182(.A1(G232), .A2(G1698), .ZN(new_n383));
  INV_X1    g0183(.A(G238), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n383), .B1(new_n384), .B2(G1698), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n382), .B1(new_n380), .B2(new_n385), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n346), .B1(G244), .B2(new_n347), .ZN(new_n387));
  AND2_X1   g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(G200), .ZN(new_n389));
  OAI211_X1 g0189(.A(new_n371), .B(new_n379), .C1(new_n388), .C2(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n389), .B1(new_n386), .B2(new_n387), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n378), .A2(new_n268), .ZN(new_n392));
  OAI211_X1 g0192(.A(new_n392), .B(new_n373), .C1(G77), .C2(new_n311), .ZN(new_n393));
  OAI21_X1  g0193(.A(KEYINPUT71), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n388), .A2(G190), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n390), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n386), .A2(new_n387), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n379), .B1(new_n397), .B2(new_n357), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n398), .B1(G179), .B2(new_n397), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n396), .A2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT9), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n367), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n364), .A2(KEYINPUT9), .A3(new_n366), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n404), .B1(G200), .B2(new_n356), .ZN(new_n405));
  OAI211_X1 g0205(.A(G190), .B(new_n348), .C1(new_n355), .C2(new_n247), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT10), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT72), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n408), .B1(new_n356), .B2(G200), .ZN(new_n409));
  OAI211_X1 g0209(.A(new_n405), .B(new_n406), .C1(new_n407), .C2(new_n409), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n409), .A2(new_n407), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n356), .A2(G200), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n412), .A2(new_n406), .A3(new_n403), .A4(new_n402), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  AOI211_X1 g0214(.A(new_n370), .B(new_n400), .C1(new_n410), .C2(new_n414), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n361), .A2(new_n201), .ZN(new_n416));
  OAI22_X1  g0216(.A1(new_n362), .A2(new_n216), .B1(new_n211), .B2(G68), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n268), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  XNOR2_X1  g0218(.A(new_n418), .B(KEYINPUT11), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT73), .ZN(new_n420));
  OR2_X1    g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n419), .A2(new_n420), .ZN(new_n422));
  OAI21_X1  g0222(.A(KEYINPUT12), .B1(new_n311), .B2(G68), .ZN(new_n423));
  OR3_X1    g0223(.A1(new_n311), .A2(KEYINPUT12), .A3(G68), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n289), .B1(new_n259), .B2(G20), .ZN(new_n425));
  AOI22_X1  g0225(.A1(new_n423), .A2(new_n424), .B1(new_n313), .B2(new_n425), .ZN(new_n426));
  AND3_X1   g0226(.A1(new_n421), .A2(new_n422), .A3(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT14), .ZN(new_n429));
  NOR2_X1   g0229(.A1(G226), .A2(G1698), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n430), .B1(new_n222), .B2(G1698), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n296), .A2(new_n431), .A3(new_n298), .ZN(new_n432));
  NAND2_X1  g0232(.A1(G33), .A2(G97), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n210), .B1(G33), .B2(G41), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT13), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n258), .B1(new_n261), .B2(new_n384), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n436), .A2(new_n437), .A3(new_n439), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n247), .B1(new_n432), .B2(new_n433), .ZN(new_n441));
  OAI21_X1  g0241(.A(KEYINPUT13), .B1(new_n441), .B2(new_n438), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n429), .B1(new_n443), .B2(G169), .ZN(new_n444));
  AOI211_X1 g0244(.A(KEYINPUT14), .B(new_n357), .C1(new_n440), .C2(new_n442), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n440), .A2(G179), .A3(new_n442), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT74), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n440), .A2(new_n442), .A3(KEYINPUT74), .A4(G179), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  AND3_X1   g0251(.A1(new_n446), .A2(KEYINPUT75), .A3(new_n451), .ZN(new_n452));
  AOI21_X1  g0252(.A(KEYINPUT75), .B1(new_n446), .B2(new_n451), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n428), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n443), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(G190), .ZN(new_n456));
  OAI211_X1 g0256(.A(new_n427), .B(new_n456), .C1(new_n455), .C2(new_n389), .ZN(new_n457));
  AND4_X1   g0257(.A1(new_n345), .A2(new_n415), .A3(new_n454), .A4(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n211), .A2(G87), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT22), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(KEYINPUT87), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT87), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(KEYINPUT22), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n459), .B1(new_n461), .B2(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n464), .A2(new_n296), .A3(new_n298), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n211), .B1(new_n250), .B2(new_n251), .ZN(new_n466));
  INV_X1    g0266(.A(G87), .ZN(new_n467));
  OAI21_X1  g0267(.A(KEYINPUT22), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT23), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n470), .A2(new_n218), .A3(G20), .ZN(new_n471));
  INV_X1    g0271(.A(G116), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n471), .B1(new_n472), .B2(new_n362), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n381), .A2(G20), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n473), .B1(new_n474), .B2(KEYINPUT23), .ZN(new_n475));
  XNOR2_X1  g0275(.A(KEYINPUT88), .B(KEYINPUT24), .ZN(new_n476));
  AND3_X1   g0276(.A1(new_n469), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n476), .B1(new_n469), .B2(new_n475), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n268), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(KEYINPUT89), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT89), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n481), .B(new_n268), .C1(new_n477), .C2(new_n478), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  OAI21_X1  g0283(.A(KEYINPUT81), .B1(new_n280), .B2(G1), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT81), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n485), .A2(new_n259), .A3(G33), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n313), .A2(new_n488), .A3(KEYINPUT82), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT82), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n490), .B1(new_n487), .B2(new_n312), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n489), .A2(G107), .A3(new_n491), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n311), .A2(G107), .ZN(new_n493));
  XNOR2_X1  g0293(.A(new_n493), .B(KEYINPUT25), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n483), .A2(new_n496), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n256), .A2(G1), .ZN(new_n498));
  XNOR2_X1  g0298(.A(KEYINPUT5), .B(G41), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n435), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(G274), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n435), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n259), .A2(G45), .ZN(new_n503));
  NOR2_X1   g0303(.A1(KEYINPUT5), .A2(G41), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(KEYINPUT5), .A2(G41), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n503), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  AOI22_X1  g0307(.A1(new_n500), .A2(G264), .B1(new_n502), .B2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(G250), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(new_n249), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n224), .A2(G1698), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n510), .B(new_n511), .C1(new_n250), .C2(new_n251), .ZN(new_n512));
  NAND2_X1  g0312(.A1(G33), .A2(G294), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(new_n435), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n508), .A2(new_n515), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n516), .A2(new_n263), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n515), .A2(KEYINPUT90), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n247), .B1(new_n512), .B2(new_n513), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT90), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n518), .A2(new_n508), .A3(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n517), .B1(G169), .B2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n497), .A2(new_n524), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n518), .A2(new_n508), .A3(new_n337), .A4(new_n521), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n507), .A2(G274), .A3(new_n247), .ZN(new_n527));
  INV_X1    g0327(.A(new_n506), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n498), .B1(new_n528), .B2(new_n504), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(new_n247), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n527), .B1(new_n219), .B2(new_n530), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n389), .B1(new_n531), .B2(new_n519), .ZN(new_n532));
  AND2_X1   g0332(.A1(new_n526), .A2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n483), .A2(new_n496), .A3(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n529), .A2(G270), .A3(new_n247), .ZN(new_n536));
  AND2_X1   g0336(.A1(new_n527), .A2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(G303), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n538), .B1(new_n296), .B2(new_n298), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n219), .A2(G1698), .ZN(new_n540));
  OAI221_X1 g0340(.A(new_n540), .B1(G257), .B2(G1698), .C1(new_n250), .C2(new_n251), .ZN(new_n541));
  INV_X1    g0341(.A(new_n541), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n435), .B1(new_n539), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n537), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n488), .A2(new_n313), .A3(G116), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n314), .A2(new_n472), .ZN(new_n546));
  AOI22_X1  g0346(.A1(new_n267), .A2(new_n210), .B1(G20), .B2(new_n472), .ZN(new_n547));
  NAND2_X1  g0347(.A1(G33), .A2(G283), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n548), .B(new_n211), .C1(G33), .C2(new_n223), .ZN(new_n549));
  AND3_X1   g0349(.A1(new_n547), .A2(KEYINPUT20), .A3(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(KEYINPUT20), .B1(new_n547), .B2(new_n549), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n545), .B(new_n546), .C1(new_n550), .C2(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n544), .A2(G169), .A3(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT21), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n537), .A2(new_n543), .A3(G179), .ZN(new_n556));
  INV_X1    g0356(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(new_n552), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n537), .A2(new_n543), .A3(G190), .ZN(new_n559));
  INV_X1    g0359(.A(new_n552), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n527), .A2(new_n536), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n541), .B1(new_n350), .B2(new_n538), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n561), .B1(new_n562), .B2(new_n435), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n559), .B(new_n560), .C1(new_n563), .C2(new_n389), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n544), .A2(KEYINPUT21), .A3(G169), .A4(new_n552), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n555), .A2(new_n558), .A3(new_n564), .A4(new_n565), .ZN(new_n566));
  NOR2_X1   g0366(.A1(G87), .A2(G97), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n381), .A2(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT19), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(KEYINPUT86), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT86), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(KEYINPUT19), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n433), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n568), .B1(new_n573), .B2(G20), .ZN(new_n574));
  AOI21_X1  g0374(.A(G20), .B1(new_n281), .B2(new_n282), .ZN(new_n575));
  XNOR2_X1  g0375(.A(KEYINPUT86), .B(KEYINPUT19), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n211), .A2(G33), .A3(G97), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n575), .A2(G68), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n574), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n268), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n489), .A2(new_n491), .A3(G87), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n377), .A2(new_n314), .ZN(new_n582));
  AND3_X1   g0382(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n384), .A2(new_n249), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n217), .A2(G1698), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n584), .B(new_n585), .C1(new_n250), .C2(new_n251), .ZN(new_n586));
  NAND2_X1  g0386(.A1(G33), .A2(G116), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT85), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n586), .A2(KEYINPUT85), .A3(new_n587), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n590), .A2(new_n435), .A3(new_n591), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n435), .B1(new_n509), .B2(new_n503), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n498), .A2(new_n501), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(G200), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n247), .B1(new_n588), .B2(new_n589), .ZN(new_n598));
  AOI22_X1  g0398(.A1(new_n598), .A2(new_n591), .B1(new_n594), .B2(new_n593), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(G190), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n583), .A2(new_n597), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n596), .A2(new_n357), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n599), .A2(new_n263), .ZN(new_n603));
  INV_X1    g0403(.A(new_n377), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n489), .A2(new_n491), .A3(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n580), .A2(new_n605), .A3(new_n582), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n602), .A2(new_n603), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n601), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n566), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n525), .A2(new_n535), .A3(new_n609), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n314), .A2(G97), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n489), .A2(new_n491), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n611), .B1(new_n612), .B2(G97), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT6), .ZN(new_n614));
  NOR3_X1   g0414(.A1(new_n614), .A2(new_n223), .A3(G107), .ZN(new_n615));
  XNOR2_X1  g0415(.A(G97), .B(G107), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n615), .B1(new_n614), .B2(new_n616), .ZN(new_n617));
  OAI22_X1  g0417(.A1(new_n617), .A2(new_n211), .B1(new_n216), .B2(new_n361), .ZN(new_n618));
  INV_X1    g0418(.A(new_n381), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n618), .B1(new_n304), .B2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(new_n268), .ZN(new_n621));
  OAI21_X1  g0421(.A(KEYINPUT80), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT80), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n381), .B1(new_n327), .B2(new_n331), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n623), .B(new_n268), .C1(new_n624), .C2(new_n618), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n613), .B1(new_n622), .B2(new_n625), .ZN(new_n626));
  NOR3_X1   g0426(.A1(new_n380), .A2(new_n509), .A3(new_n249), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT4), .ZN(new_n628));
  NOR3_X1   g0428(.A1(new_n628), .A2(new_n217), .A3(G1698), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n296), .A2(new_n298), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n249), .A2(G244), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n628), .B1(new_n301), .B2(new_n631), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n630), .A2(new_n632), .A3(new_n548), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n435), .B1(new_n627), .B2(new_n633), .ZN(new_n634));
  OAI21_X1  g0434(.A(KEYINPUT83), .B1(new_n530), .B2(new_n224), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT83), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n529), .A2(new_n636), .A3(G257), .A4(new_n247), .ZN(new_n637));
  AOI22_X1  g0437(.A1(new_n635), .A2(new_n637), .B1(new_n502), .B2(new_n507), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n634), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(G190), .ZN(new_n640));
  OAI211_X1 g0440(.A(new_n626), .B(new_n640), .C1(new_n389), .C2(new_n639), .ZN(new_n641));
  INV_X1    g0441(.A(new_n613), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n304), .A2(new_n619), .ZN(new_n643));
  INV_X1    g0443(.A(new_n618), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n623), .B1(new_n645), .B2(new_n268), .ZN(new_n646));
  NOR3_X1   g0446(.A1(new_n620), .A2(KEYINPUT80), .A3(new_n621), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n642), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  AND3_X1   g0448(.A1(new_n634), .A2(new_n638), .A3(G179), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n357), .B1(new_n634), .B2(new_n638), .ZN(new_n650));
  OR2_X1    g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT84), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n648), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n649), .A2(new_n650), .ZN(new_n654));
  OAI21_X1  g0454(.A(KEYINPUT84), .B1(new_n626), .B2(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n641), .A2(new_n653), .A3(new_n655), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n610), .A2(new_n656), .ZN(new_n657));
  AND2_X1   g0457(.A1(new_n458), .A2(new_n657), .ZN(G372));
  NOR2_X1   g0458(.A1(new_n317), .A2(new_n319), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  OAI211_X1 g0460(.A(new_n457), .B(new_n398), .C1(G179), .C2(new_n397), .ZN(new_n661));
  AND2_X1   g0461(.A1(new_n454), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n342), .A2(new_n343), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n660), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n410), .A2(new_n414), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n370), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  AND3_X1   g0466(.A1(new_n602), .A2(new_n603), .A3(new_n606), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n555), .A2(new_n558), .A3(new_n565), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n668), .B1(new_n497), .B2(new_n524), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n596), .A2(new_n337), .ZN(new_n670));
  AOI22_X1  g0470(.A1(new_n579), .A2(new_n268), .B1(new_n314), .B2(new_n377), .ZN(new_n671));
  OAI211_X1 g0471(.A(new_n671), .B(new_n581), .C1(new_n599), .C2(new_n389), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n670), .B1(new_n672), .B2(KEYINPUT91), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT91), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n583), .A2(new_n597), .A3(new_n674), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n667), .B1(new_n673), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(new_n535), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n669), .A2(new_n677), .ZN(new_n678));
  AND3_X1   g0478(.A1(new_n641), .A2(new_n653), .A3(new_n655), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n667), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n626), .A2(new_n654), .ZN(new_n681));
  AOI21_X1  g0481(.A(KEYINPUT26), .B1(new_n676), .B2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n653), .A2(new_n655), .ZN(new_n684));
  INV_X1    g0484(.A(new_n608), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT26), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n683), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n680), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n458), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n666), .A2(new_n690), .ZN(new_n691));
  XOR2_X1   g0491(.A(new_n691), .B(KEYINPUT92), .Z(G369));
  NAND3_X1  g0492(.A1(new_n259), .A2(new_n211), .A3(G13), .ZN(new_n693));
  XNOR2_X1  g0493(.A(new_n693), .B(KEYINPUT93), .ZN(new_n694));
  AND2_X1   g0494(.A1(new_n694), .A2(KEYINPUT27), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n694), .A2(KEYINPUT27), .ZN(new_n696));
  INV_X1    g0496(.A(G213), .ZN(new_n697));
  NOR3_X1   g0497(.A1(new_n695), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(G343), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n699), .A2(new_n560), .ZN(new_n700));
  OR2_X1    g0500(.A1(new_n566), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n668), .A2(new_n700), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  XOR2_X1   g0503(.A(new_n703), .B(KEYINPUT94), .Z(new_n704));
  AND2_X1   g0504(.A1(new_n704), .A2(G330), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n525), .A2(new_n535), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n699), .B1(new_n483), .B2(new_n496), .ZN(new_n707));
  OAI22_X1  g0507(.A1(new_n706), .A2(new_n707), .B1(new_n525), .B2(new_n699), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n705), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n668), .A2(new_n699), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n525), .A2(new_n711), .A3(new_n535), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n523), .B1(new_n483), .B2(new_n496), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(new_n699), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n709), .A2(new_n716), .ZN(G399));
  INV_X1    g0517(.A(new_n207), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n718), .A2(G41), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n568), .A2(G116), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n720), .A2(new_n721), .A3(G1), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n722), .B1(new_n214), .B2(new_n720), .ZN(new_n723));
  XNOR2_X1  g0523(.A(new_n723), .B(KEYINPUT28), .ZN(new_n724));
  AND3_X1   g0524(.A1(new_n676), .A2(new_n681), .A3(KEYINPUT26), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n725), .B1(new_n686), .B2(new_n687), .ZN(new_n726));
  OAI211_X1 g0526(.A(new_n535), .B(new_n676), .C1(new_n713), .C2(new_n668), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n607), .B1(new_n727), .B2(new_n656), .ZN(new_n728));
  OAI211_X1 g0528(.A(KEYINPUT29), .B(new_n699), .C1(new_n726), .C2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n699), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n730), .B1(new_n680), .B2(new_n688), .ZN(new_n731));
  XNOR2_X1  g0531(.A(KEYINPUT96), .B(KEYINPUT29), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n729), .B1(new_n731), .B2(new_n733), .ZN(new_n734));
  OR2_X1    g0534(.A1(new_n566), .A2(new_n608), .ZN(new_n735));
  AOI211_X1 g0535(.A(new_n495), .B(new_n533), .C1(new_n480), .C2(new_n482), .ZN(new_n736));
  NOR3_X1   g0536(.A1(new_n735), .A2(new_n713), .A3(new_n736), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n737), .A2(new_n679), .A3(new_n699), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n519), .B1(G264), .B2(new_n500), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n592), .A2(new_n739), .A3(new_n595), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(KEYINPUT95), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT95), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n599), .A2(new_n742), .A3(new_n739), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n741), .A2(new_n639), .A3(new_n557), .A4(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT30), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n634), .A2(new_n638), .ZN(new_n747));
  AOI21_X1  g0547(.A(G179), .B1(new_n508), .B2(new_n515), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n747), .A2(new_n596), .A3(new_n544), .A4(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n747), .A2(new_n556), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n750), .A2(KEYINPUT30), .A3(new_n743), .A4(new_n741), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n746), .A2(new_n749), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(new_n730), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT31), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n752), .A2(KEYINPUT31), .A3(new_n730), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n738), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(G330), .ZN(new_n758));
  AND2_X1   g0558(.A1(new_n734), .A2(new_n758), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n724), .B1(new_n759), .B2(G1), .ZN(G364));
  INV_X1    g0560(.A(G13), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(G20), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n259), .B1(new_n762), .B2(G45), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n719), .A2(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n705), .A2(new_n765), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n766), .B1(G330), .B2(new_n704), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n350), .A2(new_n207), .ZN(new_n768));
  INV_X1    g0568(.A(G355), .ZN(new_n769));
  OAI22_X1  g0569(.A1(new_n768), .A2(new_n769), .B1(G116), .B2(new_n207), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n284), .A2(new_n286), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(new_n718), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n772), .B1(G45), .B2(new_n214), .ZN(new_n773));
  OR2_X1    g0573(.A1(new_n773), .A2(KEYINPUT97), .ZN(new_n774));
  AOI22_X1  g0574(.A1(new_n773), .A2(KEYINPUT97), .B1(G45), .B2(new_n240), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n770), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  OAI211_X1 g0576(.A(G1), .B(G13), .C1(new_n211), .C2(G169), .ZN(new_n777));
  OR2_X1    g0577(.A1(new_n777), .A2(KEYINPUT98), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n777), .A2(KEYINPUT98), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(G13), .A2(G33), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(G20), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n780), .A2(new_n783), .ZN(new_n784));
  XOR2_X1   g0584(.A(new_n784), .B(KEYINPUT99), .Z(new_n785));
  OAI21_X1  g0585(.A(new_n765), .B1(new_n776), .B2(new_n785), .ZN(new_n786));
  NOR4_X1   g0586(.A1(new_n211), .A2(new_n389), .A3(G179), .A4(G190), .ZN(new_n787));
  XOR2_X1   g0587(.A(new_n787), .B(KEYINPUT101), .Z(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(new_n218), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(G20), .A2(G179), .ZN(new_n792));
  XOR2_X1   g0592(.A(new_n792), .B(KEYINPUT100), .Z(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(G190), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(G200), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n794), .A2(new_n389), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  OAI221_X1 g0598(.A(new_n791), .B1(new_n796), .B2(new_n202), .C1(new_n201), .C2(new_n798), .ZN(new_n799));
  AND3_X1   g0599(.A1(new_n793), .A2(new_n337), .A3(G200), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(KEYINPUT102), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n800), .A2(KEYINPUT102), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n804), .A2(new_n289), .ZN(new_n805));
  NOR2_X1   g0605(.A1(G179), .A2(G200), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n211), .B1(new_n806), .B2(G190), .ZN(new_n807));
  NOR4_X1   g0607(.A1(new_n211), .A2(new_n337), .A3(new_n389), .A4(G179), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  OAI221_X1 g0609(.A(new_n350), .B1(new_n223), .B2(new_n807), .C1(new_n809), .C2(new_n467), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n806), .A2(G20), .A3(new_n337), .ZN(new_n811));
  INV_X1    g0611(.A(G159), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n813), .B(KEYINPUT32), .ZN(new_n814));
  NOR2_X1   g0614(.A1(G190), .A2(G200), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n793), .A2(new_n815), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n814), .B1(new_n216), .B2(new_n816), .ZN(new_n817));
  OR3_X1    g0617(.A1(new_n805), .A2(new_n810), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n795), .A2(G322), .ZN(new_n819));
  INV_X1    g0619(.A(G326), .ZN(new_n820));
  INV_X1    g0620(.A(G283), .ZN(new_n821));
  OAI221_X1 g0621(.A(new_n819), .B1(new_n798), .B2(new_n820), .C1(new_n821), .C2(new_n789), .ZN(new_n822));
  INV_X1    g0622(.A(G329), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n380), .B1(new_n823), .B2(new_n811), .ZN(new_n824));
  INV_X1    g0624(.A(G294), .ZN(new_n825));
  OAI22_X1  g0625(.A1(new_n809), .A2(new_n538), .B1(new_n825), .B2(new_n807), .ZN(new_n826));
  INV_X1    g0626(.A(new_n816), .ZN(new_n827));
  AOI211_X1 g0627(.A(new_n824), .B(new_n826), .C1(G311), .C2(new_n827), .ZN(new_n828));
  XOR2_X1   g0628(.A(KEYINPUT33), .B(G317), .Z(new_n829));
  OAI21_X1  g0629(.A(new_n828), .B1(new_n804), .B2(new_n829), .ZN(new_n830));
  OAI22_X1  g0630(.A1(new_n799), .A2(new_n818), .B1(new_n822), .B2(new_n830), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n786), .B1(new_n831), .B2(new_n780), .ZN(new_n832));
  INV_X1    g0632(.A(new_n783), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n832), .B1(new_n703), .B2(new_n833), .ZN(new_n834));
  AND2_X1   g0634(.A1(new_n767), .A2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(G396));
  OR3_X1    g0636(.A1(new_n399), .A2(KEYINPUT104), .A3(new_n699), .ZN(new_n837));
  OAI21_X1  g0637(.A(KEYINPUT104), .B1(new_n399), .B2(new_n699), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  OAI211_X1 g0639(.A(new_n396), .B(new_n399), .C1(new_n379), .C2(new_n699), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  XNOR2_X1  g0641(.A(new_n731), .B(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n765), .B1(new_n842), .B2(new_n758), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n843), .B1(new_n758), .B2(new_n842), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n780), .A2(new_n781), .ZN(new_n845));
  XOR2_X1   g0645(.A(new_n845), .B(KEYINPUT103), .Z(new_n846));
  OAI21_X1  g0646(.A(new_n765), .B1(new_n846), .B2(G77), .ZN(new_n847));
  INV_X1    g0647(.A(G143), .ZN(new_n848));
  OAI22_X1  g0648(.A1(new_n796), .A2(new_n848), .B1(new_n816), .B2(new_n812), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n849), .B1(G137), .B2(new_n797), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n850), .B1(new_n360), .B2(new_n804), .ZN(new_n851));
  XOR2_X1   g0651(.A(new_n851), .B(KEYINPUT34), .Z(new_n852));
  NOR2_X1   g0652(.A1(new_n789), .A2(new_n289), .ZN(new_n853));
  INV_X1    g0653(.A(G132), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n771), .B1(new_n854), .B2(new_n811), .ZN(new_n855));
  OAI22_X1  g0655(.A1(new_n809), .A2(new_n201), .B1(new_n202), .B2(new_n807), .ZN(new_n856));
  OR3_X1    g0656(.A1(new_n853), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n789), .A2(new_n467), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  OAI221_X1 g0659(.A(new_n859), .B1(new_n796), .B2(new_n825), .C1(new_n538), .C2(new_n798), .ZN(new_n860));
  INV_X1    g0660(.A(G311), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n380), .B1(new_n861), .B2(new_n811), .ZN(new_n862));
  OAI22_X1  g0662(.A1(new_n809), .A2(new_n218), .B1(new_n223), .B2(new_n807), .ZN(new_n863));
  AOI211_X1 g0663(.A(new_n862), .B(new_n863), .C1(G116), .C2(new_n827), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n864), .B1(new_n804), .B2(new_n821), .ZN(new_n865));
  OAI22_X1  g0665(.A1(new_n852), .A2(new_n857), .B1(new_n860), .B2(new_n865), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n847), .B1(new_n866), .B2(new_n780), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n867), .B1(new_n782), .B2(new_n841), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n844), .A2(new_n868), .ZN(G384));
  INV_X1    g0669(.A(new_n617), .ZN(new_n870));
  AND2_X1   g0670(.A1(new_n870), .A2(KEYINPUT35), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n870), .A2(KEYINPUT35), .ZN(new_n872));
  NOR4_X1   g0672(.A1(new_n871), .A2(new_n872), .A3(new_n472), .A4(new_n213), .ZN(new_n873));
  XOR2_X1   g0673(.A(new_n873), .B(KEYINPUT36), .Z(new_n874));
  OAI21_X1  g0674(.A(G77), .B1(new_n202), .B2(new_n289), .ZN(new_n875));
  OAI22_X1  g0675(.A1(new_n875), .A2(new_n214), .B1(G50), .B2(new_n289), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n876), .A2(G1), .A3(new_n761), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g0678(.A(new_n878), .B(KEYINPUT105), .ZN(new_n879));
  AND2_X1   g0679(.A1(new_n287), .A2(new_n277), .ZN(new_n880));
  OAI21_X1  g0680(.A(G68), .B1(new_n880), .B2(new_n283), .ZN(new_n881));
  AOI21_X1  g0681(.A(KEYINPUT16), .B1(new_n881), .B2(new_n276), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n290), .A2(new_n268), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n315), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(new_n698), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n886), .B1(new_n320), .B2(new_n344), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT37), .ZN(new_n888));
  INV_X1    g0688(.A(new_n266), .ZN(new_n889));
  AOI22_X1  g0689(.A1(new_n334), .A2(new_n339), .B1(new_n884), .B2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT106), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n886), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(new_n340), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n276), .B1(new_n288), .B2(new_n289), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n323), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n895), .A2(new_n268), .A3(new_n290), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n266), .B1(new_n896), .B2(new_n315), .ZN(new_n897));
  OAI21_X1  g0697(.A(KEYINPUT106), .B1(new_n893), .B2(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n888), .B1(new_n892), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n306), .A2(new_n315), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(new_n889), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n698), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n901), .A2(new_n902), .A3(new_n340), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n903), .A2(KEYINPUT37), .ZN(new_n904));
  OAI211_X1 g0704(.A(new_n887), .B(KEYINPUT38), .C1(new_n899), .C2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(KEYINPUT107), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n659), .A2(new_n663), .ZN(new_n907));
  AND2_X1   g0707(.A1(new_n903), .A2(KEYINPUT37), .ZN(new_n908));
  OAI22_X1  g0708(.A1(new_n907), .A2(new_n902), .B1(new_n908), .B2(new_n904), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT38), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n321), .B1(new_n322), .B2(new_n895), .ZN(new_n912));
  OAI211_X1 g0712(.A(new_n891), .B(new_n340), .C1(new_n912), .C2(new_n266), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n885), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n884), .A2(new_n889), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n891), .B1(new_n915), .B2(new_n340), .ZN(new_n916));
  OAI21_X1  g0716(.A(KEYINPUT37), .B1(new_n914), .B2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(new_n904), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT107), .ZN(new_n920));
  NAND4_X1  g0720(.A1(new_n919), .A2(new_n920), .A3(KEYINPUT38), .A4(new_n887), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n906), .A2(new_n911), .A3(new_n921), .ZN(new_n922));
  AND2_X1   g0722(.A1(new_n839), .A2(new_n840), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n428), .A2(new_n730), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n454), .A2(new_n457), .A3(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT75), .ZN(new_n926));
  INV_X1    g0726(.A(new_n451), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n437), .B1(new_n436), .B2(new_n439), .ZN(new_n928));
  NOR3_X1   g0728(.A1(new_n441), .A2(KEYINPUT13), .A3(new_n438), .ZN(new_n929));
  OAI21_X1  g0729(.A(G169), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(KEYINPUT14), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n443), .A2(new_n429), .A3(G169), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n926), .B1(new_n927), .B2(new_n933), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n446), .A2(KEYINPUT75), .A3(new_n451), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(new_n457), .ZN(new_n937));
  OAI211_X1 g0737(.A(new_n428), .B(new_n730), .C1(new_n936), .C2(new_n937), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n923), .B1(new_n925), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n753), .A2(KEYINPUT108), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT108), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n752), .A2(new_n941), .A3(new_n730), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n940), .A2(new_n754), .A3(new_n942), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n943), .A2(new_n738), .A3(new_n756), .ZN(new_n944));
  AND3_X1   g0744(.A1(new_n939), .A2(KEYINPUT40), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n922), .A2(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT40), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n898), .A2(new_n913), .A3(new_n885), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n904), .B1(new_n948), .B2(KEYINPUT37), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT79), .ZN(new_n950));
  NOR3_X1   g0750(.A1(new_n316), .A2(new_n950), .A3(KEYINPUT18), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n663), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n901), .A2(new_n318), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n316), .A2(KEYINPUT18), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n953), .A2(new_n950), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n885), .B1(new_n952), .B2(new_n955), .ZN(new_n956));
  NOR3_X1   g0756(.A1(new_n949), .A2(new_n956), .A3(new_n910), .ZN(new_n957));
  AOI21_X1  g0757(.A(KEYINPUT38), .B1(new_n919), .B2(new_n887), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n939), .A2(new_n944), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n947), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  AND2_X1   g0761(.A1(new_n946), .A2(new_n961), .ZN(new_n962));
  AND2_X1   g0762(.A1(new_n458), .A2(new_n944), .ZN(new_n963));
  AND2_X1   g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n962), .A2(new_n963), .ZN(new_n965));
  INV_X1    g0765(.A(G330), .ZN(new_n966));
  NOR3_X1   g0766(.A1(new_n964), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  XOR2_X1   g0767(.A(new_n967), .B(KEYINPUT109), .Z(new_n968));
  AOI21_X1  g0768(.A(new_n608), .B1(new_n653), .B2(new_n655), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n682), .B1(new_n969), .B2(KEYINPUT26), .ZN(new_n970));
  OAI211_X1 g0770(.A(new_n699), .B(new_n841), .C1(new_n728), .C2(new_n970), .ZN(new_n971));
  OR2_X1    g0771(.A1(new_n399), .A2(new_n730), .ZN(new_n972));
  AOI22_X1  g0772(.A1(new_n971), .A2(new_n972), .B1(new_n925), .B2(new_n938), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n910), .B1(new_n949), .B2(new_n956), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n974), .A2(new_n905), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  OR2_X1    g0776(.A1(new_n660), .A2(new_n698), .ZN(new_n977));
  AOI21_X1  g0777(.A(KEYINPUT39), .B1(new_n909), .B2(new_n910), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n906), .A2(new_n921), .A3(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n975), .A2(KEYINPUT39), .ZN(new_n980));
  AND2_X1   g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n454), .A2(new_n730), .ZN(new_n982));
  INV_X1    g0782(.A(new_n982), .ZN(new_n983));
  OAI211_X1 g0783(.A(new_n976), .B(new_n977), .C1(new_n981), .C2(new_n983), .ZN(new_n984));
  OAI211_X1 g0784(.A(new_n458), .B(new_n729), .C1(new_n731), .C2(new_n733), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n985), .A2(new_n666), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n984), .B(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(new_n987), .ZN(new_n988));
  OAI22_X1  g0788(.A1(new_n968), .A2(new_n988), .B1(new_n259), .B2(new_n762), .ZN(new_n989));
  INV_X1    g0789(.A(new_n968), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n990), .A2(new_n987), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n879), .B1(new_n989), .B2(new_n991), .ZN(G367));
  AOI211_X1 g0792(.A(new_n783), .B(new_n780), .C1(new_n718), .C2(new_n604), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n231), .A2(new_n772), .ZN(new_n994));
  AOI211_X1 g0794(.A(new_n719), .B(new_n764), .C1(new_n993), .C2(new_n994), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n676), .B1(new_n583), .B2(new_n699), .ZN(new_n996));
  OR3_X1    g0796(.A1(new_n607), .A2(new_n583), .A3(new_n699), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT46), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n999), .B1(new_n809), .B2(new_n472), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n808), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1001));
  OAI211_X1 g0801(.A(new_n1000), .B(new_n1001), .C1(new_n821), .C2(new_n816), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n787), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n1003), .A2(new_n223), .B1(new_n381), .B2(new_n807), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n811), .ZN(new_n1005));
  AOI211_X1 g0805(.A(new_n771), .B(new_n1004), .C1(G317), .C2(new_n1005), .ZN(new_n1006));
  OAI221_X1 g0806(.A(new_n1006), .B1(new_n538), .B2(new_n796), .C1(new_n861), .C2(new_n798), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n804), .ZN(new_n1008));
  AOI211_X1 g0808(.A(new_n1002), .B(new_n1007), .C1(G294), .C2(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(KEYINPUT112), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n807), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(G68), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n1012), .B1(new_n796), .B2(new_n360), .C1(new_n848), .C2(new_n798), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT113), .ZN(new_n1014));
  OR2_X1    g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1008), .A2(G159), .ZN(new_n1017));
  OAI22_X1  g0817(.A1(new_n809), .A2(new_n202), .B1(new_n1003), .B2(new_n216), .ZN(new_n1018));
  INV_X1    g0818(.A(G137), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n350), .B1(new_n1019), .B2(new_n811), .ZN(new_n1020));
  AOI211_X1 g0820(.A(new_n1018), .B(new_n1020), .C1(G50), .C2(new_n827), .ZN(new_n1021));
  NAND4_X1  g0821(.A1(new_n1015), .A2(new_n1016), .A3(new_n1017), .A4(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1010), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n1023), .ZN(new_n1024));
  AND2_X1   g0824(.A1(new_n1024), .A2(KEYINPUT47), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n780), .B1(new_n1024), .B2(KEYINPUT47), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n995), .B1(new_n833), .B2(new_n998), .C1(new_n1025), .C2(new_n1026), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n679), .B1(new_n626), .B2(new_n699), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n681), .A2(new_n730), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT110), .ZN(new_n1030));
  AND2_X1   g0830(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n1031), .A2(new_n712), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1032), .B(KEYINPUT42), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n1031), .A2(new_n525), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n699), .B1(new_n1034), .B2(new_n684), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1033), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n998), .ZN(new_n1037));
  INV_X1    g0837(.A(KEYINPUT43), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n998), .A2(KEYINPUT43), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1036), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  NAND4_X1  g0841(.A1(new_n1033), .A2(new_n1035), .A3(new_n1038), .A4(new_n1037), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n709), .A2(new_n1031), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1043), .A2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1041), .A2(new_n1044), .A3(new_n1042), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g0848(.A(KEYINPUT111), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1050), .A2(KEYINPUT45), .A3(new_n716), .ZN(new_n1051));
  INV_X1    g0851(.A(KEYINPUT45), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1052), .B1(new_n1031), .B2(new_n715), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1031), .A2(KEYINPUT44), .A3(new_n715), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT44), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1055), .B1(new_n1050), .B2(new_n716), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n1051), .A2(new_n1053), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1049), .B1(new_n1057), .B2(new_n709), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1053), .A2(new_n1051), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1054), .A2(new_n1056), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n709), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1061), .A2(KEYINPUT111), .A3(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1058), .A2(new_n1063), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n712), .B1(new_n708), .B2(new_n711), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n705), .B(new_n1065), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n1066), .B(new_n759), .C1(new_n1061), .C2(new_n1062), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n759), .B1(new_n1064), .B2(new_n1067), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n719), .B(KEYINPUT41), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n764), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1027), .B1(new_n1048), .B2(new_n1070), .ZN(G387));
  OAI22_X1  g0871(.A1(new_n768), .A2(new_n721), .B1(G107), .B2(new_n207), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n772), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n721), .ZN(new_n1074));
  AOI211_X1 g0874(.A(G45), .B(new_n1074), .C1(G68), .C2(G77), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n376), .A2(G50), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT50), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1073), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n236), .A2(G45), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1072), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n765), .B1(new_n1080), .B2(new_n785), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n201), .A2(new_n796), .B1(new_n798), .B2(new_n812), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1082), .B1(G97), .B2(new_n788), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n771), .B1(new_n360), .B2(new_n811), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n808), .A2(G77), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1085), .B1(new_n377), .B2(new_n807), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n1084), .B(new_n1086), .C1(G68), .C2(new_n827), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n1083), .B(new_n1087), .C1(new_n309), .C2(new_n804), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n809), .A2(new_n825), .B1(new_n821), .B2(new_n807), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n795), .A2(G317), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1090), .B1(new_n538), .B2(new_n816), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1091), .B1(G322), .B2(new_n797), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1092), .B1(new_n861), .B2(new_n804), .ZN(new_n1093));
  INV_X1    g0893(.A(KEYINPUT48), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1089), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1095), .B1(new_n1094), .B2(new_n1093), .ZN(new_n1096));
  XOR2_X1   g0896(.A(new_n1096), .B(KEYINPUT49), .Z(new_n1097));
  INV_X1    g0897(.A(new_n771), .ZN(new_n1098));
  OAI221_X1 g0898(.A(new_n1098), .B1(new_n820), .B2(new_n811), .C1(new_n472), .C2(new_n1003), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1088), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1081), .B1(new_n1100), .B2(new_n780), .ZN(new_n1101));
  OR2_X1    g0901(.A1(new_n708), .A2(new_n833), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n1066), .A2(new_n764), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1066), .A2(new_n759), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(new_n719), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n1066), .A2(new_n759), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1103), .B1(new_n1105), .B2(new_n1106), .ZN(G393));
  OAI21_X1  g0907(.A(new_n784), .B1(new_n223), .B2(new_n207), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n1073), .A2(new_n244), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n765), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(G311), .A2(new_n795), .B1(new_n797), .B2(G317), .ZN(new_n1111));
  XNOR2_X1  g0911(.A(new_n1111), .B(KEYINPUT52), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1008), .A2(G303), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n827), .A2(G294), .ZN(new_n1114));
  OAI22_X1  g0914(.A1(new_n809), .A2(new_n821), .B1(new_n472), .B2(new_n807), .ZN(new_n1115));
  AOI211_X1 g0915(.A(new_n350), .B(new_n1115), .C1(G322), .C2(new_n1005), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n1113), .A2(new_n791), .A3(new_n1114), .A4(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1008), .A2(G50), .ZN(new_n1118));
  OR2_X1    g0918(.A1(new_n816), .A2(new_n376), .ZN(new_n1119));
  OAI22_X1  g0919(.A1(new_n809), .A2(new_n289), .B1(new_n216), .B2(new_n807), .ZN(new_n1120));
  AOI211_X1 g0920(.A(new_n1098), .B(new_n1120), .C1(G143), .C2(new_n1005), .ZN(new_n1121));
  NAND4_X1  g0921(.A1(new_n1118), .A2(new_n859), .A3(new_n1119), .A4(new_n1121), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(G150), .A2(new_n797), .B1(new_n795), .B2(G159), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(new_n1123), .B(KEYINPUT51), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n1112), .A2(new_n1117), .B1(new_n1122), .B2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1110), .B1(new_n1125), .B2(new_n780), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1126), .B1(new_n1050), .B2(new_n833), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(new_n1057), .B(new_n709), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1127), .B1(new_n1128), .B2(new_n763), .ZN(new_n1129));
  OR2_X1    g0929(.A1(new_n1064), .A2(new_n1067), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n720), .B1(new_n1128), .B2(new_n1104), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1129), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1132), .ZN(G390));
  OAI211_X1 g0933(.A(new_n979), .B(new_n980), .C1(new_n982), .C2(new_n973), .ZN(new_n1134));
  OAI211_X1 g0934(.A(new_n699), .B(new_n841), .C1(new_n726), .C2(new_n728), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1135), .A2(new_n972), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n925), .A2(new_n938), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1138), .A2(new_n922), .A3(new_n983), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1134), .A2(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n756), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1141), .B1(new_n657), .B2(new_n699), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n966), .B1(new_n1142), .B2(new_n943), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(new_n939), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1140), .A2(new_n1145), .ZN(new_n1146));
  NAND4_X1  g0946(.A1(new_n757), .A2(new_n1137), .A3(G330), .A4(new_n841), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1134), .A2(new_n1139), .A3(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1137), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n757), .A2(G330), .A3(new_n841), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(new_n1150), .A2(new_n1151), .B1(new_n1143), .B2(new_n939), .ZN(new_n1152));
  AND2_X1   g0952(.A1(new_n971), .A2(new_n972), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1147), .A2(new_n972), .A3(new_n1135), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1137), .B1(new_n1143), .B2(new_n841), .ZN(new_n1155));
  OAI22_X1  g0955(.A1(new_n1152), .A2(new_n1153), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT114), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n458), .A2(G330), .A3(new_n944), .ZN(new_n1158));
  NAND4_X1  g0958(.A1(new_n985), .A2(new_n666), .A3(new_n1157), .A4(new_n1158), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n985), .A2(new_n666), .A3(new_n1158), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1160), .A2(KEYINPUT114), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1156), .A2(new_n1159), .A3(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n720), .B1(new_n1149), .B2(new_n1162), .ZN(new_n1163));
  AND3_X1   g0963(.A1(new_n1134), .A2(new_n1139), .A3(new_n1147), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1144), .B1(new_n1134), .B2(new_n1139), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1162), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1163), .A2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1146), .A2(new_n764), .A3(new_n1148), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n981), .A2(new_n781), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n309), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n765), .B1(new_n846), .B2(new_n1172), .ZN(new_n1173));
  OR3_X1    g0973(.A1(new_n809), .A2(KEYINPUT53), .A3(new_n360), .ZN(new_n1174));
  OAI21_X1  g0974(.A(KEYINPUT53), .B1(new_n809), .B2(new_n360), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(KEYINPUT54), .B(G143), .ZN(new_n1176));
  OAI211_X1 g0976(.A(new_n1174), .B(new_n1175), .C1(new_n816), .C2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1177), .B1(new_n1008), .B2(G137), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n1003), .A2(new_n201), .B1(new_n812), .B2(new_n807), .ZN(new_n1179));
  INV_X1    g0979(.A(G125), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n350), .B1(new_n1180), .B2(new_n811), .ZN(new_n1181));
  AOI211_X1 g0981(.A(new_n1179), .B(new_n1181), .C1(new_n795), .C2(G132), .ZN(new_n1182));
  INV_X1    g0982(.A(G128), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1178), .B(new_n1182), .C1(new_n1183), .C2(new_n798), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n853), .B1(G116), .B2(new_n795), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1185), .B1(new_n821), .B2(new_n798), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n380), .B1(new_n825), .B2(new_n811), .ZN(new_n1187));
  OAI22_X1  g0987(.A1(new_n809), .A2(new_n467), .B1(new_n216), .B2(new_n807), .ZN(new_n1188));
  AOI211_X1 g0988(.A(new_n1187), .B(new_n1188), .C1(G97), .C2(new_n827), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1189), .B1(new_n804), .B2(new_n381), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1184), .B1(new_n1186), .B2(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1173), .B1(new_n1191), .B2(new_n780), .ZN(new_n1192));
  XOR2_X1   g0992(.A(new_n1192), .B(KEYINPUT115), .Z(new_n1193));
  NAND2_X1  g0993(.A1(new_n1171), .A2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1170), .A2(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1169), .A2(new_n1196), .ZN(G378));
  NAND2_X1  g0997(.A1(new_n665), .A2(new_n369), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n367), .A2(new_n698), .ZN(new_n1199));
  XOR2_X1   g0999(.A(new_n1199), .B(KEYINPUT55), .Z(new_n1200));
  XNOR2_X1  g1000(.A(new_n1198), .B(new_n1200), .ZN(new_n1201));
  XOR2_X1   g1001(.A(KEYINPUT117), .B(KEYINPUT56), .Z(new_n1202));
  INV_X1    g1002(.A(new_n1202), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(new_n1201), .B(new_n1203), .ZN(new_n1204));
  AND4_X1   g1004(.A1(G330), .A2(new_n946), .A3(new_n961), .A4(new_n1204), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n939), .B(new_n944), .C1(new_n957), .C2(new_n958), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n966), .B1(new_n1206), .B2(new_n947), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1204), .B1(new_n1207), .B2(new_n946), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n984), .B1(new_n1205), .B2(new_n1208), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n946), .A2(new_n961), .A3(G330), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1204), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n976), .A2(new_n977), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n983), .B1(new_n979), .B2(new_n980), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1207), .A2(new_n946), .A3(new_n1204), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1212), .A2(new_n1215), .A3(new_n1216), .ZN(new_n1217));
  AND2_X1   g1017(.A1(new_n1209), .A2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1204), .A2(new_n781), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n765), .B1(new_n846), .B2(G50), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1098), .A2(new_n255), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n787), .A2(G58), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1005), .A2(G283), .ZN(new_n1223));
  NAND4_X1  g1023(.A1(new_n1085), .A2(new_n1012), .A3(new_n1222), .A4(new_n1223), .ZN(new_n1224));
  AOI211_X1 g1024(.A(new_n1221), .B(new_n1224), .C1(new_n604), .C2(new_n827), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(G107), .A2(new_n795), .B1(new_n797), .B2(G116), .ZN(new_n1226));
  OAI211_X1 g1026(.A(new_n1225), .B(new_n1226), .C1(new_n804), .C2(new_n223), .ZN(new_n1227));
  INV_X1    g1027(.A(KEYINPUT58), .ZN(new_n1228));
  AOI21_X1  g1028(.A(G50), .B1(new_n280), .B2(new_n255), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n1227), .A2(new_n1228), .B1(new_n1221), .B2(new_n1229), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(new_n827), .A2(G137), .B1(G150), .B2(new_n1011), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1231), .B1(new_n1180), .B2(new_n798), .ZN(new_n1232));
  OAI22_X1  g1032(.A1(new_n796), .A2(new_n1183), .B1(new_n809), .B2(new_n1176), .ZN(new_n1233));
  XOR2_X1   g1033(.A(new_n1233), .B(KEYINPUT116), .Z(new_n1234));
  AOI211_X1 g1034(.A(new_n1232), .B(new_n1234), .C1(G132), .C2(new_n1008), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(KEYINPUT59), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n787), .A2(G159), .ZN(new_n1238));
  AOI211_X1 g1038(.A(G33), .B(G41), .C1(new_n1005), .C2(G124), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1237), .A2(new_n1238), .A3(new_n1239), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1236), .A2(KEYINPUT59), .ZN(new_n1241));
  OAI221_X1 g1041(.A(new_n1230), .B1(new_n1228), .B2(new_n1227), .C1(new_n1240), .C2(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1220), .B1(new_n1242), .B2(new_n780), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(new_n1218), .A2(new_n764), .B1(new_n1219), .B2(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1156), .ZN(new_n1245));
  OAI211_X1 g1045(.A(new_n1159), .B(new_n1161), .C1(new_n1149), .C2(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(KEYINPUT57), .B1(new_n1246), .B2(new_n1218), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1161), .A2(new_n1159), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1248), .B1(new_n1166), .B2(new_n1156), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1209), .A2(new_n1217), .A3(KEYINPUT57), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n719), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1244), .B1(new_n1247), .B2(new_n1251), .ZN(G375));
  NAND2_X1  g1052(.A1(new_n1248), .A2(new_n1245), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1253), .A2(new_n1069), .A3(new_n1162), .ZN(new_n1254));
  XNOR2_X1  g1054(.A(new_n1254), .B(KEYINPUT118), .ZN(new_n1255));
  XNOR2_X1  g1055(.A(new_n763), .B(KEYINPUT119), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1156), .A2(new_n1257), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n765), .B1(new_n846), .B2(G68), .ZN(new_n1259));
  OAI22_X1  g1059(.A1(new_n821), .A2(new_n796), .B1(new_n798), .B2(new_n825), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1260), .B1(G77), .B2(new_n788), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n380), .B1(new_n538), .B2(new_n811), .ZN(new_n1262));
  OAI22_X1  g1062(.A1(new_n809), .A2(new_n223), .B1(new_n377), .B2(new_n807), .ZN(new_n1263));
  AOI211_X1 g1063(.A(new_n1262), .B(new_n1263), .C1(new_n619), .C2(new_n827), .ZN(new_n1264));
  OAI211_X1 g1064(.A(new_n1261), .B(new_n1264), .C1(new_n472), .C2(new_n804), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n771), .B1(new_n1183), .B2(new_n811), .ZN(new_n1266));
  OAI221_X1 g1066(.A(new_n1222), .B1(new_n201), .B2(new_n807), .C1(new_n809), .C2(new_n812), .ZN(new_n1267));
  AOI211_X1 g1067(.A(new_n1266), .B(new_n1267), .C1(G150), .C2(new_n827), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(G132), .A2(new_n797), .B1(new_n795), .B2(G137), .ZN(new_n1269));
  OAI211_X1 g1069(.A(new_n1268), .B(new_n1269), .C1(new_n804), .C2(new_n1176), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1265), .A2(new_n1270), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1259), .B1(new_n1271), .B2(new_n780), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1272), .B1(new_n1137), .B2(new_n782), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1258), .A2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1255), .A2(new_n1275), .ZN(G381));
  NOR3_X1   g1076(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1277));
  XNOR2_X1  g1077(.A(new_n1277), .B(KEYINPUT120), .ZN(new_n1278));
  OAI211_X1 g1078(.A(new_n1027), .B(new_n1132), .C1(new_n1048), .C2(new_n1070), .ZN(new_n1279));
  NOR4_X1   g1079(.A1(new_n1278), .A2(G381), .A3(G378), .A4(new_n1279), .ZN(new_n1280));
  OAI211_X1 g1080(.A(new_n1280), .B(new_n1244), .C1(new_n1247), .C2(new_n1251), .ZN(G407));
  AOI21_X1  g1081(.A(new_n1195), .B1(new_n1163), .B2(new_n1168), .ZN(new_n1282));
  OR3_X1    g1082(.A1(new_n697), .A2(KEYINPUT121), .A3(G343), .ZN(new_n1283));
  OAI21_X1  g1083(.A(KEYINPUT121), .B1(new_n697), .B2(G343), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1282), .A2(new_n1286), .ZN(new_n1287));
  OAI211_X1 g1087(.A(G407), .B(G213), .C1(G375), .C2(new_n1287), .ZN(G409));
  NAND3_X1  g1088(.A1(new_n1209), .A2(new_n1217), .A3(new_n1069), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1249), .A2(new_n1289), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1209), .A2(new_n1217), .A3(new_n1257), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1243), .A2(new_n1219), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1282), .B1(new_n1290), .B2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1294), .A2(KEYINPUT122), .ZN(new_n1295));
  OAI211_X1 g1095(.A(G378), .B(new_n1244), .C1(new_n1247), .C2(new_n1251), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT122), .ZN(new_n1297));
  OAI211_X1 g1097(.A(new_n1282), .B(new_n1297), .C1(new_n1290), .C2(new_n1293), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1295), .A2(new_n1296), .A3(new_n1298), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1156), .B1(new_n1159), .B2(new_n1161), .ZN(new_n1300));
  OAI211_X1 g1100(.A(new_n719), .B(new_n1162), .C1(new_n1300), .C2(KEYINPUT60), .ZN(new_n1301));
  AND3_X1   g1101(.A1(new_n1248), .A2(new_n1245), .A3(KEYINPUT60), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1275), .B1(new_n1301), .B2(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(G384), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  OAI211_X1 g1105(.A(new_n1275), .B(G384), .C1(new_n1301), .C2(new_n1302), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1307), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1299), .A2(new_n1285), .A3(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1309), .A2(KEYINPUT62), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1286), .A2(KEYINPUT124), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1305), .A2(new_n1306), .A3(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1286), .A2(G2897), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1312), .A2(new_n1314), .ZN(new_n1315));
  NAND4_X1  g1115(.A1(new_n1305), .A2(new_n1306), .A3(new_n1313), .A4(new_n1311), .ZN(new_n1316));
  AND2_X1   g1116(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1299), .A2(new_n1285), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1317), .A2(new_n1318), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT61), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT62), .ZN(new_n1321));
  NAND4_X1  g1121(.A1(new_n1299), .A2(new_n1308), .A3(new_n1321), .A4(new_n1285), .ZN(new_n1322));
  NAND4_X1  g1122(.A1(new_n1310), .A2(new_n1319), .A3(new_n1320), .A4(new_n1322), .ZN(new_n1323));
  XNOR2_X1  g1123(.A(G393), .B(new_n835), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT127), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(G387), .A2(new_n1325), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1324), .B1(new_n1326), .B2(G390), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(G387), .A2(new_n1325), .A3(new_n1132), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1327), .A2(new_n1328), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(G387), .A2(G390), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1330), .A2(new_n1279), .A3(new_n1324), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1331), .A2(KEYINPUT126), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT126), .ZN(new_n1333));
  NAND4_X1  g1133(.A1(new_n1330), .A2(new_n1279), .A3(new_n1333), .A4(new_n1324), .ZN(new_n1334));
  AND3_X1   g1134(.A1(new_n1329), .A2(new_n1332), .A3(new_n1334), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1323), .A2(new_n1335), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1318), .A2(KEYINPUT123), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT123), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1299), .A2(new_n1338), .A3(new_n1285), .ZN(new_n1339));
  NAND3_X1  g1139(.A1(new_n1315), .A2(KEYINPUT125), .A3(new_n1316), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1341));
  INV_X1    g1141(.A(KEYINPUT125), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1341), .A2(new_n1342), .ZN(new_n1343));
  NAND4_X1  g1143(.A1(new_n1337), .A2(new_n1339), .A3(new_n1340), .A4(new_n1343), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1309), .A2(KEYINPUT63), .ZN(new_n1345));
  INV_X1    g1145(.A(KEYINPUT63), .ZN(new_n1346));
  NAND4_X1  g1146(.A1(new_n1299), .A2(new_n1308), .A3(new_n1346), .A4(new_n1285), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1345), .A2(new_n1347), .ZN(new_n1348));
  AOI22_X1  g1148(.A1(new_n1328), .A2(new_n1327), .B1(new_n1331), .B2(KEYINPUT126), .ZN(new_n1349));
  AOI21_X1  g1149(.A(KEYINPUT61), .B1(new_n1349), .B2(new_n1334), .ZN(new_n1350));
  NAND3_X1  g1150(.A1(new_n1344), .A2(new_n1348), .A3(new_n1350), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1336), .A2(new_n1351), .ZN(G405));
  NAND2_X1  g1152(.A1(G375), .A2(new_n1282), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1353), .A2(new_n1296), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1354), .A2(new_n1308), .ZN(new_n1355));
  NAND3_X1  g1155(.A1(new_n1353), .A2(new_n1307), .A3(new_n1296), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1355), .A2(new_n1356), .ZN(new_n1357));
  XNOR2_X1  g1157(.A(new_n1335), .B(new_n1357), .ZN(G402));
endmodule


