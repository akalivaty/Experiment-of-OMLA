//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1 0 0 0 0 0 0 0 0 0 0 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 0 0 1 0 0 1 1 1 1 1 1 0 0 1 0 0 0 0 1 0 1 0 1 0 0 1 1 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:35 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1212, new_n1213,
    new_n1214, new_n1215, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1292, new_n1293,
    new_n1294, new_n1295;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  OR3_X1    g0006(.A1(new_n206), .A2(KEYINPUT64), .A3(G13), .ZN(new_n207));
  OAI21_X1  g0007(.A(KEYINPUT64), .B1(new_n206), .B2(G13), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  AND2_X1   g0011(.A1(new_n211), .A2(KEYINPUT0), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(KEYINPUT0), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n214));
  INV_X1    g0014(.A(G58), .ZN(new_n215));
  INV_X1    g0015(.A(G232), .ZN(new_n216));
  INV_X1    g0016(.A(G97), .ZN(new_n217));
  INV_X1    g0017(.A(G257), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n214), .B1(new_n215), .B2(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n206), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  AND2_X1   g0023(.A1(new_n223), .A2(KEYINPUT1), .ZN(new_n224));
  INV_X1    g0024(.A(new_n201), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n225), .A2(G50), .ZN(new_n226));
  INV_X1    g0026(.A(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  INV_X1    g0028(.A(G20), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n227), .A2(new_n230), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n231), .B1(new_n223), .B2(KEYINPUT1), .ZN(new_n232));
  NOR4_X1   g0032(.A1(new_n212), .A2(new_n213), .A3(new_n224), .A4(new_n232), .ZN(G361));
  XOR2_X1   g0033(.A(G238), .B(G244), .Z(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT65), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XOR2_X1   g0042(.A(G107), .B(G116), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(KEYINPUT66), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G87), .B(G97), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G50), .B(G68), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G58), .B(G77), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(new_n246), .B(new_n249), .Z(G351));
  OR2_X1    g0050(.A1(KEYINPUT3), .A2(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(KEYINPUT3), .A2(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n253), .A2(G232), .A3(G1698), .ZN(new_n254));
  INV_X1    g0054(.A(G33), .ZN(new_n255));
  INV_X1    g0055(.A(G1698), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n253), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G226), .ZN(new_n258));
  OAI221_X1 g0058(.A(new_n254), .B1(new_n255), .B2(new_n217), .C1(new_n257), .C2(new_n258), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n228), .B1(G33), .B2(G41), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G1), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n262), .B1(G41), .B2(G45), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(KEYINPUT67), .ZN(new_n264));
  NAND2_X1  g0064(.A1(G33), .A2(G41), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n265), .A2(G1), .A3(G13), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT67), .ZN(new_n267));
  OAI211_X1 g0067(.A(new_n267), .B(new_n262), .C1(G41), .C2(G45), .ZN(new_n268));
  NAND4_X1  g0068(.A1(new_n264), .A2(G274), .A3(new_n266), .A4(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n266), .A2(new_n263), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n270), .B1(G238), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n261), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(KEYINPUT13), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT72), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT13), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n261), .A2(new_n273), .A3(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n275), .A2(new_n276), .A3(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(new_n274), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n280), .A2(KEYINPUT72), .A3(new_n277), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n279), .A2(G169), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(KEYINPUT14), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT73), .ZN(new_n284));
  AND3_X1   g0084(.A1(new_n275), .A2(new_n284), .A3(new_n278), .ZN(new_n285));
  NOR3_X1   g0085(.A1(new_n280), .A2(new_n284), .A3(new_n277), .ZN(new_n286));
  OAI21_X1  g0086(.A(G179), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT14), .ZN(new_n288));
  NAND4_X1  g0088(.A1(new_n279), .A2(new_n281), .A3(new_n288), .A4(G169), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n283), .A2(new_n287), .A3(new_n289), .ZN(new_n290));
  NAND3_X1  g0090(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(new_n228), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n293), .B1(G1), .B2(new_n229), .ZN(new_n294));
  INV_X1    g0094(.A(G68), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  XNOR2_X1  g0096(.A(new_n296), .B(KEYINPUT74), .ZN(new_n297));
  INV_X1    g0097(.A(G13), .ZN(new_n298));
  NOR3_X1   g0098(.A1(new_n298), .A2(new_n229), .A3(G1), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(new_n295), .ZN(new_n300));
  XNOR2_X1  g0100(.A(new_n300), .B(KEYINPUT12), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n297), .A2(new_n301), .ZN(new_n302));
  XNOR2_X1  g0102(.A(new_n302), .B(KEYINPUT75), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n255), .A2(G20), .ZN(new_n304));
  AOI22_X1  g0104(.A1(new_n304), .A2(G77), .B1(G20), .B2(new_n295), .ZN(new_n305));
  NOR2_X1   g0105(.A1(G20), .A2(G33), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n305), .B1(new_n202), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(new_n292), .ZN(new_n309));
  XNOR2_X1  g0109(.A(new_n309), .B(KEYINPUT11), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n303), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n290), .A2(new_n311), .ZN(new_n312));
  OAI21_X1  g0112(.A(G190), .B1(new_n285), .B2(new_n286), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n279), .A2(G200), .A3(new_n281), .ZN(new_n314));
  NAND4_X1  g0114(.A1(new_n313), .A2(new_n303), .A3(new_n310), .A4(new_n314), .ZN(new_n315));
  AND2_X1   g0115(.A1(new_n312), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT68), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT8), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n317), .B1(new_n318), .B2(G58), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n215), .A2(KEYINPUT68), .A3(KEYINPUT8), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n318), .A2(G58), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n319), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n294), .A2(new_n322), .ZN(new_n323));
  OR2_X1    g0123(.A1(new_n322), .A2(new_n299), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT77), .ZN(new_n325));
  AND3_X1   g0125(.A1(new_n323), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n325), .B1(new_n323), .B2(new_n324), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  OR2_X1    g0128(.A1(G223), .A2(G1698), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n258), .A2(G1698), .ZN(new_n330));
  AND2_X1   g0130(.A1(KEYINPUT3), .A2(G33), .ZN(new_n331));
  NOR2_X1   g0131(.A1(KEYINPUT3), .A2(G33), .ZN(new_n332));
  OAI211_X1 g0132(.A(new_n329), .B(new_n330), .C1(new_n331), .C2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(G33), .A2(G87), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(new_n260), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n272), .A2(G232), .ZN(new_n337));
  NAND4_X1  g0137(.A1(new_n336), .A2(new_n269), .A3(G190), .A4(new_n337), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n268), .A2(new_n266), .A3(G274), .ZN(new_n339));
  AND2_X1   g0139(.A1(new_n263), .A2(KEYINPUT67), .ZN(new_n340));
  OAI22_X1  g0140(.A1(new_n339), .A2(new_n340), .B1(new_n271), .B2(new_n216), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n266), .B1(new_n333), .B2(new_n334), .ZN(new_n342));
  OAI21_X1  g0142(.A(G200), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  AND2_X1   g0143(.A1(new_n338), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n251), .A2(new_n229), .A3(new_n252), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT7), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND4_X1  g0147(.A1(new_n251), .A2(KEYINPUT7), .A3(new_n229), .A4(new_n252), .ZN(new_n348));
  AOI21_X1  g0148(.A(KEYINPUT76), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT76), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n350), .B1(new_n345), .B2(new_n346), .ZN(new_n351));
  OAI21_X1  g0151(.A(G68), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n215), .A2(new_n295), .ZN(new_n353));
  OAI21_X1  g0153(.A(G20), .B1(new_n353), .B2(new_n201), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n306), .A2(G159), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  AOI21_X1  g0157(.A(KEYINPUT16), .B1(new_n352), .B2(new_n357), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n331), .A2(new_n332), .ZN(new_n359));
  AOI21_X1  g0159(.A(KEYINPUT7), .B1(new_n359), .B2(new_n229), .ZN(new_n360));
  NOR4_X1   g0160(.A1(new_n331), .A2(new_n332), .A3(new_n346), .A4(G20), .ZN(new_n361));
  OAI21_X1  g0161(.A(G68), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n362), .A2(KEYINPUT16), .A3(new_n357), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(new_n292), .ZN(new_n364));
  OAI211_X1 g0164(.A(new_n328), .B(new_n344), .C1(new_n358), .C2(new_n364), .ZN(new_n365));
  XNOR2_X1  g0165(.A(new_n365), .B(KEYINPUT17), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n328), .B1(new_n358), .B2(new_n364), .ZN(new_n367));
  INV_X1    g0167(.A(G179), .ZN(new_n368));
  NAND4_X1  g0168(.A1(new_n336), .A2(new_n269), .A3(new_n368), .A4(new_n337), .ZN(new_n369));
  INV_X1    g0169(.A(G169), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n370), .B1(new_n341), .B2(new_n342), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(KEYINPUT78), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT78), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n369), .A2(new_n371), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n367), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(KEYINPUT18), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT18), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n367), .A2(new_n376), .A3(new_n379), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n366), .A2(new_n378), .A3(new_n380), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n269), .B1(new_n258), .B2(new_n271), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n253), .A2(G223), .A3(G1698), .ZN(new_n383));
  INV_X1    g0183(.A(G77), .ZN(new_n384));
  INV_X1    g0184(.A(G222), .ZN(new_n385));
  OAI221_X1 g0185(.A(new_n383), .B1(new_n384), .B2(new_n253), .C1(new_n257), .C2(new_n385), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n382), .B1(new_n386), .B2(new_n260), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT70), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n388), .A2(new_n389), .A3(G200), .ZN(new_n390));
  INV_X1    g0190(.A(G200), .ZN(new_n391));
  OAI21_X1  g0191(.A(KEYINPUT70), .B1(new_n387), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(new_n393), .ZN(new_n394));
  OAI21_X1  g0194(.A(G50), .B1(new_n229), .B2(G1), .ZN(new_n395));
  XNOR2_X1  g0195(.A(new_n395), .B(KEYINPUT69), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n299), .A2(new_n292), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(new_n299), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n398), .B1(G50), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n322), .A2(new_n304), .ZN(new_n401));
  AOI22_X1  g0201(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n306), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n293), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n400), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(KEYINPUT9), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT9), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n406), .B1(new_n400), .B2(new_n403), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n387), .A2(G190), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n405), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT71), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n394), .A2(new_n410), .A3(new_n411), .A4(KEYINPUT10), .ZN(new_n412));
  OR2_X1    g0212(.A1(new_n411), .A2(KEYINPUT10), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n411), .A2(KEYINPUT10), .ZN(new_n414));
  OAI211_X1 g0214(.A(new_n413), .B(new_n414), .C1(new_n393), .C2(new_n409), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n412), .A2(new_n415), .ZN(new_n416));
  AND2_X1   g0216(.A1(new_n272), .A2(G244), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n253), .A2(G232), .A3(new_n256), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n253), .A2(G238), .A3(G1698), .ZN(new_n419));
  INV_X1    g0219(.A(G107), .ZN(new_n420));
  OAI211_X1 g0220(.A(new_n418), .B(new_n419), .C1(new_n420), .C2(new_n253), .ZN(new_n421));
  AOI211_X1 g0221(.A(new_n270), .B(new_n417), .C1(new_n260), .C2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(new_n368), .ZN(new_n423));
  XNOR2_X1  g0223(.A(KEYINPUT8), .B(G58), .ZN(new_n424));
  OAI22_X1  g0224(.A1(new_n424), .A2(new_n307), .B1(new_n229), .B2(new_n384), .ZN(new_n425));
  XNOR2_X1  g0225(.A(KEYINPUT15), .B(G87), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n425), .B1(new_n427), .B2(new_n304), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n428), .A2(new_n293), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n299), .A2(new_n384), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n430), .B1(new_n294), .B2(new_n384), .ZN(new_n431));
  OAI221_X1 g0231(.A(new_n423), .B1(G169), .B2(new_n422), .C1(new_n429), .C2(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n404), .B1(new_n388), .B2(new_n370), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n433), .B1(G179), .B2(new_n388), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n422), .A2(G190), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n429), .A2(new_n431), .ZN(new_n436));
  OAI211_X1 g0236(.A(new_n435), .B(new_n436), .C1(new_n391), .C2(new_n422), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n432), .A2(new_n434), .A3(new_n437), .ZN(new_n438));
  NOR3_X1   g0238(.A1(new_n381), .A2(new_n416), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n316), .A2(new_n439), .ZN(new_n440));
  AOI211_X1 g0240(.A(new_n292), .B(new_n299), .C1(new_n262), .C2(G33), .ZN(new_n441));
  OR2_X1    g0241(.A1(KEYINPUT85), .A2(G116), .ZN(new_n442));
  NAND2_X1  g0242(.A1(KEYINPUT85), .A2(G116), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  AOI22_X1  g0245(.A1(new_n441), .A2(G116), .B1(new_n299), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(G33), .A2(G283), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n447), .B(new_n229), .C1(G33), .C2(new_n217), .ZN(new_n448));
  XNOR2_X1  g0248(.A(new_n448), .B(KEYINPUT89), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n293), .B1(new_n445), .B2(G20), .ZN(new_n450));
  AND3_X1   g0250(.A1(new_n449), .A2(KEYINPUT20), .A3(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(KEYINPUT20), .B1(new_n449), .B2(new_n450), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n446), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(G303), .ZN(new_n454));
  OAI22_X1  g0254(.A1(new_n257), .A2(new_n218), .B1(new_n454), .B2(new_n253), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n253), .A2(G264), .A3(G1698), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n260), .B1(new_n455), .B2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT81), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT5), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n459), .B1(new_n460), .B2(G41), .ZN(new_n461));
  INV_X1    g0261(.A(G41), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n462), .A2(KEYINPUT81), .A3(KEYINPUT5), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n462), .A2(KEYINPUT5), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n262), .A2(G45), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n464), .A2(new_n467), .A3(G274), .A4(new_n266), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n260), .B1(new_n464), .B2(new_n467), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(G270), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n458), .A2(new_n468), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n453), .B1(G200), .B2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(G190), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n472), .B1(new_n473), .B2(new_n471), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n453), .A2(KEYINPUT21), .A3(G169), .A4(new_n471), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n453), .A2(G169), .A3(new_n471), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT21), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n471), .A2(new_n368), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(new_n453), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n474), .A2(new_n475), .A3(new_n478), .A4(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT91), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT25), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n483), .B1(new_n399), .B2(G107), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n299), .A2(KEYINPUT25), .A3(new_n420), .ZN(new_n485));
  AOI22_X1  g0285(.A1(new_n441), .A2(G107), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  OAI21_X1  g0287(.A(KEYINPUT23), .B1(new_n229), .B2(G107), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT23), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n489), .A2(new_n420), .A3(G20), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n255), .B1(new_n442), .B2(new_n443), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n491), .B1(new_n492), .B2(new_n229), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n229), .B(G87), .C1(new_n331), .C2(new_n332), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT90), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(KEYINPUT22), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  AND2_X1   g0297(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n494), .A2(new_n497), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n493), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(KEYINPUT24), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n494), .A2(new_n497), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n253), .A2(new_n229), .A3(G87), .A4(new_n496), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT24), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n504), .A2(new_n505), .A3(new_n493), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n501), .A2(new_n506), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n487), .B1(new_n507), .B2(new_n292), .ZN(new_n508));
  OAI211_X1 g0308(.A(G250), .B(new_n256), .C1(new_n331), .C2(new_n332), .ZN(new_n509));
  OAI211_X1 g0309(.A(G257), .B(G1698), .C1(new_n331), .C2(new_n332), .ZN(new_n510));
  INV_X1    g0310(.A(G294), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n509), .B(new_n510), .C1(new_n255), .C2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(new_n260), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n469), .A2(G264), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n513), .A2(new_n468), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(new_n370), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n516), .B1(G179), .B2(new_n515), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n482), .B1(new_n508), .B2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(new_n506), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n505), .B1(new_n504), .B2(new_n493), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n292), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(new_n486), .ZN(new_n522));
  AOI22_X1  g0322(.A1(new_n512), .A2(new_n260), .B1(new_n469), .B2(G264), .ZN(new_n523));
  AOI21_X1  g0323(.A(G169), .B1(new_n523), .B2(new_n468), .ZN(new_n524));
  AND4_X1   g0324(.A1(new_n368), .A2(new_n513), .A3(new_n468), .A4(new_n514), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n522), .A2(new_n526), .A3(KEYINPUT91), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n523), .A2(G190), .A3(new_n468), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n515), .A2(G200), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n508), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n518), .A2(new_n527), .A3(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT92), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n518), .A2(new_n527), .A3(new_n530), .A4(KEYINPUT92), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n481), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n350), .B1(new_n360), .B2(new_n361), .ZN(new_n536));
  INV_X1    g0336(.A(new_n351), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n420), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT6), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n217), .A2(new_n420), .ZN(new_n540));
  NOR2_X1   g0340(.A1(G97), .A2(G107), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n420), .A2(KEYINPUT6), .A3(G97), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AOI22_X1  g0344(.A1(new_n544), .A2(G20), .B1(G77), .B2(new_n306), .ZN(new_n545));
  INV_X1    g0345(.A(new_n545), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n292), .B1(new_n538), .B2(new_n546), .ZN(new_n547));
  OAI21_X1  g0347(.A(KEYINPUT79), .B1(new_n399), .B2(G97), .ZN(new_n548));
  OR3_X1    g0348(.A1(new_n399), .A2(KEYINPUT79), .A3(G97), .ZN(new_n549));
  AOI22_X1  g0349(.A1(new_n548), .A2(new_n549), .B1(new_n441), .B2(G97), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n547), .A2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(G45), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n552), .A2(G1), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n460), .A2(G41), .ZN(new_n554));
  AND3_X1   g0354(.A1(new_n462), .A2(KEYINPUT81), .A3(KEYINPUT5), .ZN(new_n555));
  AOI21_X1  g0355(.A(KEYINPUT81), .B1(new_n462), .B2(KEYINPUT5), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n553), .B(new_n554), .C1(new_n555), .C2(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT82), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n557), .A2(new_n558), .A3(G257), .A4(new_n266), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(new_n468), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n558), .B1(new_n469), .B2(G257), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  OAI211_X1 g0362(.A(G244), .B(new_n256), .C1(new_n331), .C2(new_n332), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT4), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n253), .A2(KEYINPUT4), .A3(G244), .A4(new_n256), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n253), .A2(G250), .A3(G1698), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n565), .A2(new_n566), .A3(new_n447), .A4(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT80), .ZN(new_n569));
  AND3_X1   g0369(.A1(new_n568), .A2(new_n569), .A3(new_n260), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n569), .B1(new_n568), .B2(new_n260), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n562), .B(new_n368), .C1(new_n570), .C2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n469), .A2(G257), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(KEYINPUT82), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n574), .A2(new_n559), .A3(new_n468), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n568), .A2(new_n260), .ZN(new_n576));
  INV_X1    g0376(.A(new_n576), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n370), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n551), .A2(new_n572), .A3(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT83), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n551), .A2(new_n572), .A3(new_n578), .A4(KEYINPUT83), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n562), .B1(new_n570), .B2(new_n571), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(G200), .ZN(new_n584));
  OAI21_X1  g0384(.A(G107), .B1(new_n349), .B2(new_n351), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n293), .B1(new_n585), .B2(new_n545), .ZN(new_n586));
  INV_X1    g0386(.A(new_n550), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n562), .A2(G190), .A3(new_n576), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n584), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(G250), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n553), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n266), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT84), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n592), .A2(KEYINPUT84), .A3(new_n266), .ZN(new_n596));
  AOI22_X1  g0396(.A1(new_n595), .A2(new_n596), .B1(G274), .B2(new_n553), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n253), .A2(G244), .A3(G1698), .ZN(new_n598));
  OAI211_X1 g0398(.A(G238), .B(new_n256), .C1(new_n331), .C2(new_n332), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n444), .A2(G33), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n598), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n260), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n597), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(new_n370), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n253), .A2(new_n229), .A3(G68), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(KEYINPUT86), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT19), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n304), .A2(new_n607), .A3(G97), .ZN(new_n608));
  AOI21_X1  g0408(.A(G20), .B1(G33), .B2(G97), .ZN(new_n609));
  INV_X1    g0409(.A(G87), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n609), .B1(new_n610), .B2(new_n541), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n608), .B1(new_n611), .B2(new_n607), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT86), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n253), .A2(new_n613), .A3(new_n229), .A4(G68), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n606), .A2(new_n612), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n292), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n426), .A2(new_n299), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n441), .A2(new_n427), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n616), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n597), .A2(new_n368), .A3(new_n602), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n604), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  AND2_X1   g0421(.A1(new_n601), .A2(new_n260), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n553), .A2(G274), .ZN(new_n623));
  INV_X1    g0423(.A(new_n596), .ZN(new_n624));
  AOI21_X1  g0424(.A(KEYINPUT84), .B1(new_n592), .B2(new_n266), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n623), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  OAI21_X1  g0426(.A(G200), .B1(new_n622), .B2(new_n626), .ZN(new_n627));
  AOI22_X1  g0427(.A1(new_n615), .A2(new_n292), .B1(new_n299), .B2(new_n426), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n441), .A2(KEYINPUT87), .A3(G87), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT87), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n397), .B1(G1), .B2(new_n255), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n630), .B1(new_n631), .B2(new_n610), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n629), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n597), .A2(G190), .A3(new_n602), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n627), .A2(new_n628), .A3(new_n633), .A4(new_n634), .ZN(new_n635));
  AND2_X1   g0435(.A1(new_n621), .A2(new_n635), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n581), .A2(new_n582), .A3(new_n590), .A4(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT88), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n637), .A2(new_n638), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n535), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n440), .A2(new_n641), .ZN(G372));
  INV_X1    g0442(.A(new_n434), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n312), .A2(new_n432), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n644), .A2(new_n315), .A3(new_n366), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n378), .A2(new_n380), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT93), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n416), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n412), .A2(new_n415), .A3(KEYINPUT93), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n643), .B1(new_n647), .B2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n621), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n621), .A2(new_n635), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n654), .A2(new_n579), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT26), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n653), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n654), .B1(new_n581), .B2(new_n582), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n657), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n522), .A2(new_n526), .ZN(new_n660));
  AND4_X1   g0460(.A1(new_n660), .A2(new_n478), .A3(new_n475), .A4(new_n480), .ZN(new_n661));
  INV_X1    g0461(.A(new_n530), .ZN(new_n662));
  NOR3_X1   g0462(.A1(new_n637), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n659), .A2(new_n663), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n652), .B1(new_n440), .B2(new_n664), .ZN(G369));
  NAND3_X1  g0465(.A1(new_n478), .A2(new_n475), .A3(new_n480), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n262), .A2(new_n229), .A3(G13), .ZN(new_n668));
  OR2_X1    g0468(.A1(new_n668), .A2(KEYINPUT27), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(KEYINPUT27), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n669), .A2(new_n670), .A3(G213), .ZN(new_n671));
  INV_X1    g0471(.A(G343), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n453), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n667), .A2(new_n474), .A3(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n675), .B1(new_n667), .B2(new_n674), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(G330), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n673), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n660), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n533), .A2(new_n534), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n522), .A2(new_n673), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n682), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n680), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n667), .A2(new_n673), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n683), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n660), .A2(new_n673), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n687), .A2(new_n692), .ZN(G399));
  INV_X1    g0493(.A(new_n209), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n694), .A2(G41), .ZN(new_n695));
  INV_X1    g0495(.A(G116), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n541), .A2(new_n610), .A3(new_n696), .ZN(new_n697));
  NOR3_X1   g0497(.A1(new_n695), .A2(new_n262), .A3(new_n697), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n698), .B1(new_n227), .B2(new_n695), .ZN(new_n699));
  XNOR2_X1  g0499(.A(KEYINPUT94), .B(KEYINPUT28), .ZN(new_n700));
  XNOR2_X1  g0500(.A(new_n699), .B(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n681), .B1(new_n659), .B2(new_n663), .ZN(new_n702));
  AND2_X1   g0502(.A1(new_n581), .A2(new_n582), .ZN(new_n703));
  OAI211_X1 g0503(.A(KEYINPUT96), .B(new_n656), .C1(new_n703), .C2(new_n654), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT96), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n705), .B1(new_n658), .B2(KEYINPUT26), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n655), .A2(KEYINPUT26), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n704), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n637), .A2(new_n662), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n518), .A2(new_n527), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(new_n667), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n653), .B1(new_n709), .B2(new_n712), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n673), .B1(new_n708), .B2(new_n713), .ZN(new_n714));
  MUX2_X1   g0514(.A(new_n702), .B(new_n714), .S(KEYINPUT29), .Z(new_n715));
  OAI211_X1 g0515(.A(new_n535), .B(new_n681), .C1(new_n639), .C2(new_n640), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n575), .A2(new_n577), .ZN(new_n717));
  INV_X1    g0517(.A(new_n523), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n603), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n479), .A2(new_n717), .A3(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT30), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n479), .A2(new_n717), .A3(KEYINPUT30), .A4(new_n719), .ZN(new_n723));
  AOI21_X1  g0523(.A(G179), .B1(new_n597), .B2(new_n602), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n583), .A2(new_n515), .A3(new_n471), .A4(new_n724), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n722), .A2(new_n723), .A3(new_n725), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n726), .A2(KEYINPUT31), .A3(new_n673), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT95), .ZN(new_n728));
  XNOR2_X1  g0528(.A(new_n727), .B(new_n728), .ZN(new_n729));
  AND2_X1   g0529(.A1(new_n726), .A2(new_n673), .ZN(new_n730));
  OR2_X1    g0530(.A1(new_n730), .A2(KEYINPUT31), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n716), .A2(new_n729), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(G330), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n715), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n701), .B1(new_n735), .B2(G1), .ZN(G364));
  XNOR2_X1  g0536(.A(new_n679), .B(KEYINPUT97), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n298), .A2(G20), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n262), .B1(new_n738), .B2(G45), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n695), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  OAI211_X1 g0542(.A(new_n737), .B(new_n742), .C1(G330), .C2(new_n676), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n209), .A2(G355), .A3(new_n253), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n744), .B1(G116), .B2(new_n209), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n209), .A2(new_n359), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n746), .B1(new_n552), .B2(new_n227), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n249), .A2(G45), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n745), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(G13), .A2(G33), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(G20), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n228), .B1(G20), .B2(new_n370), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g0554(.A(new_n754), .B(KEYINPUT98), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n741), .B1(new_n749), .B2(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n229), .A2(new_n368), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(G200), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(G190), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  XOR2_X1   g0560(.A(KEYINPUT33), .B(G317), .Z(new_n761));
  NOR2_X1   g0561(.A1(new_n229), .A2(G179), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n762), .A2(new_n473), .A3(G200), .ZN(new_n763));
  INV_X1    g0563(.A(G283), .ZN(new_n764));
  OAI22_X1  g0564(.A1(new_n760), .A2(new_n761), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n758), .A2(new_n473), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(G326), .ZN(new_n767));
  NOR2_X1   g0567(.A1(G179), .A2(G200), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n229), .B1(new_n768), .B2(G190), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n767), .B1(new_n511), .B2(new_n769), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n768), .A2(G20), .A3(new_n473), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n253), .B1(new_n772), .B2(G329), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n762), .A2(G190), .A3(G200), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n773), .B1(new_n454), .B2(new_n774), .ZN(new_n775));
  NOR3_X1   g0575(.A1(new_n765), .A2(new_n770), .A3(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(G311), .ZN(new_n777));
  INV_X1    g0577(.A(new_n757), .ZN(new_n778));
  AOI21_X1  g0578(.A(G200), .B1(new_n778), .B2(KEYINPUT99), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n779), .B1(KEYINPUT99), .B2(new_n778), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(G190), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(G322), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n780), .A2(new_n473), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  OAI221_X1 g0585(.A(new_n776), .B1(new_n777), .B2(new_n782), .C1(new_n783), .C2(new_n785), .ZN(new_n786));
  OAI22_X1  g0586(.A1(new_n610), .A2(new_n774), .B1(new_n763), .B2(new_n420), .ZN(new_n787));
  INV_X1    g0587(.A(new_n769), .ZN(new_n788));
  AOI211_X1 g0588(.A(new_n359), .B(new_n787), .C1(G97), .C2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(G159), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n771), .A2(new_n790), .ZN(new_n791));
  XNOR2_X1  g0591(.A(new_n791), .B(KEYINPUT32), .ZN(new_n792));
  AOI22_X1  g0592(.A1(new_n759), .A2(G68), .B1(new_n766), .B2(G50), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n789), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  OAI22_X1  g0594(.A1(new_n215), .A2(new_n785), .B1(new_n782), .B2(new_n384), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n786), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n756), .B1(new_n796), .B2(new_n753), .ZN(new_n797));
  INV_X1    g0597(.A(new_n752), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n797), .B1(new_n676), .B2(new_n798), .ZN(new_n799));
  AND2_X1   g0599(.A1(new_n743), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(G396));
  NOR2_X1   g0601(.A1(new_n432), .A2(new_n673), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n437), .B1(new_n436), .B2(new_n681), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n802), .B1(new_n432), .B2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n702), .A2(new_n805), .ZN(new_n806));
  OAI211_X1 g0606(.A(new_n681), .B(new_n804), .C1(new_n659), .C2(new_n663), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n741), .B1(new_n733), .B2(new_n808), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n809), .B1(new_n733), .B2(new_n808), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n753), .A2(new_n750), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n742), .B1(new_n384), .B2(new_n811), .ZN(new_n812));
  OAI22_X1  g0612(.A1(new_n511), .A2(new_n785), .B1(new_n782), .B2(new_n445), .ZN(new_n813));
  OAI221_X1 g0613(.A(new_n359), .B1(new_n771), .B2(new_n777), .C1(new_n217), .C2(new_n769), .ZN(new_n814));
  OAI22_X1  g0614(.A1(new_n760), .A2(new_n764), .B1(new_n763), .B2(new_n610), .ZN(new_n815));
  INV_X1    g0615(.A(new_n766), .ZN(new_n816));
  OAI22_X1  g0616(.A1(new_n816), .A2(new_n454), .B1(new_n420), .B2(new_n774), .ZN(new_n817));
  NOR4_X1   g0617(.A1(new_n813), .A2(new_n814), .A3(new_n815), .A4(new_n817), .ZN(new_n818));
  AOI22_X1  g0618(.A1(new_n759), .A2(G150), .B1(new_n766), .B2(G137), .ZN(new_n819));
  XNOR2_X1  g0619(.A(new_n819), .B(KEYINPUT100), .ZN(new_n820));
  INV_X1    g0620(.A(G143), .ZN(new_n821));
  OAI221_X1 g0621(.A(new_n820), .B1(new_n821), .B2(new_n785), .C1(new_n790), .C2(new_n782), .ZN(new_n822));
  XNOR2_X1  g0622(.A(new_n822), .B(KEYINPUT34), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n763), .A2(new_n295), .ZN(new_n824));
  INV_X1    g0624(.A(G132), .ZN(new_n825));
  OAI221_X1 g0625(.A(new_n253), .B1(new_n771), .B2(new_n825), .C1(new_n215), .C2(new_n769), .ZN(new_n826));
  INV_X1    g0626(.A(new_n774), .ZN(new_n827));
  AOI211_X1 g0627(.A(new_n824), .B(new_n826), .C1(G50), .C2(new_n827), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n818), .B1(new_n823), .B2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n753), .ZN(new_n830));
  OAI221_X1 g0630(.A(new_n812), .B1(new_n804), .B2(new_n751), .C1(new_n829), .C2(new_n830), .ZN(new_n831));
  AND2_X1   g0631(.A1(new_n810), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(G384));
  OR2_X1    g0633(.A1(new_n544), .A2(KEYINPUT35), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n544), .A2(KEYINPUT35), .ZN(new_n835));
  NAND4_X1  g0635(.A1(new_n834), .A2(G116), .A3(new_n230), .A4(new_n835), .ZN(new_n836));
  XOR2_X1   g0636(.A(new_n836), .B(KEYINPUT36), .Z(new_n837));
  OR3_X1    g0637(.A1(new_n226), .A2(new_n384), .A3(new_n353), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n202), .A2(G68), .ZN(new_n839));
  AOI211_X1 g0639(.A(new_n262), .B(G13), .C1(new_n838), .C2(new_n839), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n837), .A2(new_n840), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n652), .B1(new_n715), .B2(new_n440), .ZN(new_n842));
  XNOR2_X1  g0642(.A(new_n842), .B(KEYINPUT106), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT38), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n323), .A2(new_n324), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n845), .A2(KEYINPUT77), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n323), .A2(new_n324), .A3(new_n325), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT16), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n295), .B1(new_n536), .B2(new_n537), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n849), .B1(new_n850), .B2(new_n356), .ZN(new_n851));
  AND2_X1   g0651(.A1(new_n363), .A2(new_n292), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n848), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  AND3_X1   g0653(.A1(new_n369), .A2(new_n371), .A3(new_n374), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n374), .B1(new_n369), .B2(new_n371), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n365), .B1(new_n853), .B2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT103), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT37), .ZN(new_n860));
  INV_X1    g0660(.A(new_n671), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n367), .A2(new_n861), .ZN(new_n862));
  NAND4_X1  g0662(.A1(new_n858), .A2(new_n859), .A3(new_n860), .A4(new_n862), .ZN(new_n863));
  NAND4_X1  g0663(.A1(new_n377), .A2(new_n862), .A3(new_n860), .A4(new_n365), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(KEYINPUT103), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n377), .A2(new_n862), .A3(new_n365), .ZN(new_n866));
  AOI22_X1  g0666(.A1(new_n863), .A2(new_n865), .B1(KEYINPUT37), .B2(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n862), .B1(new_n646), .B2(new_n366), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n844), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n295), .B1(new_n347), .B2(new_n348), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n849), .B1(new_n870), .B2(new_n356), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n871), .A2(new_n363), .A3(new_n292), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n328), .A2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT102), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n328), .A2(new_n872), .A3(KEYINPUT102), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n875), .A2(new_n861), .A3(new_n876), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n875), .A2(new_n376), .A3(new_n876), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n877), .A2(new_n878), .A3(new_n365), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(KEYINPUT37), .ZN(new_n880));
  AND2_X1   g0680(.A1(new_n864), .A2(KEYINPUT103), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n864), .A2(KEYINPUT103), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n880), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  AND2_X1   g0683(.A1(new_n875), .A2(new_n876), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n381), .A2(new_n861), .A3(new_n884), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n883), .A2(KEYINPUT38), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n869), .A2(new_n886), .ZN(new_n887));
  OAI21_X1  g0687(.A(KEYINPUT105), .B1(new_n887), .B2(KEYINPUT39), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT105), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT39), .ZN(new_n890));
  NAND4_X1  g0690(.A1(new_n869), .A2(new_n886), .A3(new_n889), .A4(new_n890), .ZN(new_n891));
  AOI22_X1  g0691(.A1(new_n863), .A2(new_n865), .B1(KEYINPUT37), .B2(new_n879), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n877), .B1(new_n646), .B2(new_n366), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n844), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n886), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(KEYINPUT39), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n888), .A2(new_n891), .A3(new_n896), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n290), .A2(new_n311), .A3(new_n681), .ZN(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  XOR2_X1   g0700(.A(new_n802), .B(KEYINPUT101), .Z(new_n901));
  NAND2_X1  g0701(.A1(new_n807), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n311), .A2(new_n673), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n312), .A2(new_n315), .A3(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n290), .A2(new_n311), .A3(new_n673), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n895), .A2(new_n902), .A3(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT104), .ZN(new_n908));
  OR2_X1    g0708(.A1(new_n646), .A2(new_n861), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n907), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n907), .A2(new_n909), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(KEYINPUT104), .ZN(new_n912));
  AND3_X1   g0712(.A1(new_n900), .A2(new_n910), .A3(new_n912), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n843), .B(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n716), .A2(new_n731), .A3(new_n727), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n805), .B1(new_n904), .B2(new_n905), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n887), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(KEYINPUT40), .ZN(new_n918));
  AOI21_X1  g0718(.A(KEYINPUT40), .B1(new_n894), .B2(new_n886), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n919), .A2(new_n915), .A3(new_n916), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(new_n440), .ZN(new_n922));
  AND2_X1   g0722(.A1(new_n922), .A2(new_n915), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n678), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n924), .B1(new_n923), .B2(new_n921), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n914), .A2(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n926), .B1(new_n262), .B2(new_n738), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n914), .A2(new_n925), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n841), .B1(new_n927), .B2(new_n928), .ZN(G367));
  INV_X1    g0729(.A(new_n755), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n930), .B1(new_n209), .B2(new_n426), .ZN(new_n931));
  AND3_X1   g0731(.A1(new_n241), .A2(new_n209), .A3(new_n359), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n741), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(G317), .ZN(new_n934));
  OAI221_X1 g0734(.A(new_n359), .B1(new_n771), .B2(new_n934), .C1(new_n816), .C2(new_n777), .ZN(new_n935));
  AOI22_X1  g0735(.A1(new_n759), .A2(G294), .B1(G107), .B2(new_n788), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n827), .A2(KEYINPUT46), .A3(G116), .ZN(new_n937));
  INV_X1    g0737(.A(new_n763), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(G97), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n936), .A2(new_n937), .A3(new_n939), .ZN(new_n940));
  AOI21_X1  g0740(.A(KEYINPUT46), .B1(new_n827), .B2(new_n444), .ZN(new_n941));
  NOR3_X1   g0741(.A1(new_n935), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  AOI22_X1  g0742(.A1(G283), .A2(new_n781), .B1(new_n784), .B2(G303), .ZN(new_n943));
  INV_X1    g0743(.A(G137), .ZN(new_n944));
  OAI221_X1 g0744(.A(new_n253), .B1(new_n771), .B2(new_n944), .C1(new_n760), .C2(new_n790), .ZN(new_n945));
  OAI22_X1  g0745(.A1(new_n215), .A2(new_n774), .B1(new_n763), .B2(new_n384), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n788), .A2(G68), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(new_n816), .B2(new_n821), .ZN(new_n948));
  NOR3_X1   g0748(.A1(new_n945), .A2(new_n946), .A3(new_n948), .ZN(new_n949));
  AOI22_X1  g0749(.A1(G50), .A2(new_n781), .B1(new_n784), .B2(G150), .ZN(new_n950));
  AOI22_X1  g0750(.A1(new_n942), .A2(new_n943), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  XOR2_X1   g0751(.A(new_n951), .B(KEYINPUT47), .Z(new_n952));
  AOI21_X1  g0752(.A(new_n933), .B1(new_n952), .B2(new_n753), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n628), .A2(new_n633), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(new_n673), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n636), .A2(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n956), .B1(new_n621), .B2(new_n955), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n953), .B1(new_n957), .B2(new_n798), .ZN(new_n958));
  OAI211_X1 g0758(.A(new_n703), .B(new_n590), .C1(new_n588), .C2(new_n681), .ZN(new_n959));
  OR2_X1    g0759(.A1(new_n579), .A2(new_n681), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n703), .B1(new_n962), .B2(new_n711), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(new_n681), .ZN(new_n964));
  OAI21_X1  g0764(.A(KEYINPUT42), .B1(new_n962), .B2(new_n689), .ZN(new_n965));
  OR3_X1    g0765(.A1(new_n962), .A2(KEYINPUT42), .A3(new_n689), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n964), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  OR3_X1    g0767(.A1(new_n967), .A2(KEYINPUT43), .A3(new_n957), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n968), .B(KEYINPUT107), .ZN(new_n969));
  XOR2_X1   g0769(.A(new_n957), .B(KEYINPUT43), .Z(new_n970));
  NAND2_X1  g0770(.A1(new_n967), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n972), .B1(new_n687), .B2(new_n962), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n969), .A2(new_n686), .A3(new_n961), .A4(new_n971), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  XOR2_X1   g0775(.A(new_n695), .B(KEYINPUT41), .Z(new_n976));
  NAND2_X1  g0776(.A1(new_n692), .A2(new_n961), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT45), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n977), .B(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n962), .B1(new_n690), .B2(new_n691), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT44), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n980), .B(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n979), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(new_n686), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n979), .A2(new_n687), .A3(new_n982), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(new_n688), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n690), .B1(new_n685), .B2(new_n988), .ZN(new_n989));
  MUX2_X1   g0789(.A(new_n737), .B(new_n679), .S(new_n989), .Z(new_n990));
  NOR2_X1   g0790(.A1(new_n990), .A2(new_n734), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n987), .A2(new_n991), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n976), .B1(new_n992), .B2(new_n735), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n993), .A2(new_n740), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n958), .B1(new_n975), .B2(new_n994), .ZN(G387));
  INV_X1    g0795(.A(new_n991), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n990), .A2(new_n734), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n996), .A2(new_n997), .A3(new_n695), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n788), .A2(new_n427), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n999), .B1(new_n785), .B2(new_n202), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(KEYINPUT109), .ZN(new_n1001));
  OAI211_X1 g0801(.A(new_n253), .B(new_n939), .C1(new_n816), .C2(new_n790), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n1002), .B1(new_n322), .B2(new_n759), .ZN(new_n1003));
  INV_X1    g0803(.A(G150), .ZN(new_n1004));
  OAI22_X1  g0804(.A1(new_n774), .A2(new_n384), .B1(new_n1004), .B2(new_n771), .ZN(new_n1005));
  XOR2_X1   g0805(.A(new_n1005), .B(KEYINPUT108), .Z(new_n1006));
  AOI21_X1  g0806(.A(new_n1006), .B1(G68), .B2(new_n781), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n1001), .A2(new_n1003), .A3(new_n1007), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n253), .B1(new_n772), .B2(G326), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(new_n759), .A2(G311), .B1(new_n766), .B2(G322), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n1010), .B1(new_n782), .B2(new_n454), .C1(new_n934), .C2(new_n785), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT48), .ZN(new_n1012));
  OR2_X1    g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(new_n827), .A2(G294), .B1(new_n788), .B2(G283), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1013), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT49), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n1009), .B1(new_n445), .B2(new_n763), .C1(new_n1016), .C2(new_n1017), .ZN(new_n1018));
  AND2_X1   g0818(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1008), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1020), .A2(new_n753), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n238), .A2(G45), .A3(new_n359), .ZN(new_n1022));
  OAI21_X1  g0822(.A(KEYINPUT50), .B1(new_n424), .B2(G50), .ZN(new_n1023));
  OAI211_X1 g0823(.A(new_n1023), .B(new_n552), .C1(new_n295), .C2(new_n384), .ZN(new_n1024));
  NOR3_X1   g0824(.A1(new_n424), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n359), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n697), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n694), .B1(new_n1022), .B2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n930), .B1(new_n420), .B2(new_n209), .ZN(new_n1030));
  OAI211_X1 g0830(.A(new_n1021), .B(new_n741), .C1(new_n1029), .C2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1031), .B1(new_n685), .B2(new_n752), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1032), .B(KEYINPUT110), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n998), .B(new_n1033), .C1(new_n739), .C2(new_n990), .ZN(G393));
  NAND2_X1  g0834(.A1(new_n987), .A2(new_n740), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n246), .A2(new_n746), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n930), .B1(new_n217), .B2(new_n209), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n741), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n359), .B1(new_n771), .B2(new_n783), .C1(new_n763), .C2(new_n420), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n760), .A2(new_n454), .B1(new_n445), .B2(new_n769), .ZN(new_n1040));
  AOI211_X1 g0840(.A(new_n1039), .B(new_n1040), .C1(G283), .C2(new_n827), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1041), .B1(new_n511), .B2(new_n782), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n784), .A2(G311), .B1(G317), .B2(new_n766), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT52), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n784), .A2(G159), .B1(G150), .B2(new_n766), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT51), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n253), .B1(new_n771), .B2(new_n821), .C1(new_n763), .C2(new_n610), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n760), .A2(new_n202), .B1(new_n295), .B2(new_n774), .ZN(new_n1048));
  AOI211_X1 g0848(.A(new_n1047), .B(new_n1048), .C1(G77), .C2(new_n788), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1049), .B1(new_n424), .B2(new_n782), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n1042), .A2(new_n1044), .B1(new_n1046), .B2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1038), .B1(new_n1051), .B2(new_n753), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1052), .B1(new_n961), .B2(new_n798), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1035), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1054), .A2(KEYINPUT111), .ZN(new_n1055));
  INV_X1    g0855(.A(KEYINPUT111), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1035), .A2(new_n1056), .A3(new_n1053), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1055), .A2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n996), .A2(new_n986), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n992), .A2(new_n695), .A3(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1058), .A2(new_n1060), .ZN(G390));
  INV_X1    g0861(.A(new_n811), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n741), .B1(new_n322), .B2(new_n1062), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1063), .B(KEYINPUT112), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n759), .A2(G137), .B1(new_n766), .B2(G128), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1065), .B1(new_n202), .B2(new_n763), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(KEYINPUT54), .B(G143), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1066), .B1(new_n781), .B2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n827), .A2(G150), .ZN(new_n1070));
  OR2_X1    g0870(.A1(new_n1070), .A2(KEYINPUT53), .ZN(new_n1071));
  INV_X1    g0871(.A(G125), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n253), .B1(new_n771), .B2(new_n1072), .C1(new_n790), .C2(new_n769), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1073), .B1(KEYINPUT53), .B2(new_n1070), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n784), .A2(G132), .ZN(new_n1075));
  NAND4_X1  g0875(.A1(new_n1069), .A2(new_n1071), .A3(new_n1074), .A4(new_n1075), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n782), .A2(new_n217), .B1(new_n420), .B2(new_n760), .ZN(new_n1077));
  INV_X1    g0877(.A(KEYINPUT113), .ZN(new_n1078));
  OR2_X1    g0878(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n359), .B1(new_n771), .B2(new_n511), .C1(new_n774), .C2(new_n610), .ZN(new_n1081));
  AOI211_X1 g0881(.A(new_n824), .B(new_n1081), .C1(G283), .C2(new_n766), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1079), .A2(new_n1080), .A3(new_n1082), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n784), .A2(G116), .B1(G77), .B2(new_n788), .ZN(new_n1084));
  XOR2_X1   g0884(.A(new_n1084), .B(KEYINPUT114), .Z(new_n1085));
  OAI21_X1  g0885(.A(new_n1076), .B1(new_n1083), .B2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1064), .B1(new_n1086), .B2(new_n753), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1087), .B1(new_n897), .B2(new_n751), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n803), .A2(new_n432), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n802), .B1(new_n714), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n906), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n898), .B(new_n887), .C1(new_n1090), .C2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n899), .B1(new_n902), .B2(new_n906), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1092), .B1(new_n897), .B2(new_n1093), .ZN(new_n1094));
  AND2_X1   g0894(.A1(new_n915), .A2(G330), .ZN(new_n1095));
  AND2_X1   g0895(.A1(new_n1095), .A2(new_n916), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n732), .A2(G330), .A3(new_n916), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n1092), .B(new_n1098), .C1(new_n897), .C2(new_n1093), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1088), .B1(new_n1100), .B2(new_n739), .ZN(new_n1101));
  AND2_X1   g0901(.A1(new_n1095), .A2(new_n922), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n842), .A2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n915), .A2(G330), .A3(new_n804), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(new_n1091), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1105), .A2(new_n1090), .A3(new_n1098), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n732), .A2(G330), .A3(new_n804), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n916), .A2(new_n1095), .B1(new_n1107), .B2(new_n1091), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n902), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1106), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  NAND4_X1  g0910(.A1(new_n1097), .A2(new_n1103), .A3(new_n1099), .A4(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n695), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1103), .A2(new_n1110), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1112), .B1(new_n1100), .B2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1101), .B1(new_n1111), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1115), .ZN(G378));
  AOI21_X1  g0916(.A(new_n678), .B1(new_n918), .B2(new_n920), .ZN(new_n1117));
  AND3_X1   g0917(.A1(new_n412), .A2(KEYINPUT93), .A3(new_n415), .ZN(new_n1118));
  AOI21_X1  g0918(.A(KEYINPUT93), .B1(new_n412), .B2(new_n415), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n434), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n404), .A2(new_n671), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1121), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n434), .B(new_n1123), .C1(new_n1118), .C2(new_n1119), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1125));
  AND3_X1   g0925(.A1(new_n1122), .A2(new_n1124), .A3(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1125), .B1(new_n1122), .B2(new_n1124), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  OAI21_X1  g0929(.A(KEYINPUT117), .B1(new_n1117), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(KEYINPUT117), .ZN(new_n1131));
  AND2_X1   g0931(.A1(new_n915), .A2(new_n916), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n1132), .A2(new_n919), .B1(new_n917), .B2(KEYINPUT40), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n1131), .B(new_n1128), .C1(new_n1133), .C2(new_n678), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1125), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1123), .B1(new_n651), .B2(new_n434), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1124), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1135), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1122), .A2(new_n1124), .A3(new_n1125), .ZN(new_n1139));
  AND3_X1   g0939(.A1(new_n1138), .A2(KEYINPUT116), .A3(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(KEYINPUT116), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1142), .A2(new_n1117), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1130), .A2(new_n1134), .A3(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n913), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  NAND4_X1  g0946(.A1(new_n913), .A2(new_n1130), .A3(new_n1134), .A4(new_n1143), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1148), .A2(new_n740), .ZN(new_n1149));
  AOI211_X1 g0949(.A(G41), .B(new_n253), .C1(new_n772), .C2(G283), .ZN(new_n1150));
  OAI221_X1 g0950(.A(new_n1150), .B1(new_n215), .B2(new_n763), .C1(new_n384), .C2(new_n774), .ZN(new_n1151));
  XOR2_X1   g0951(.A(new_n1151), .B(KEYINPUT115), .Z(new_n1152));
  NOR2_X1   g0952(.A1(new_n785), .A2(new_n420), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n782), .A2(new_n426), .ZN(new_n1154));
  OAI221_X1 g0954(.A(new_n947), .B1(new_n816), .B2(new_n696), .C1(new_n217), .C2(new_n760), .ZN(new_n1155));
  NOR4_X1   g0955(.A1(new_n1152), .A2(new_n1153), .A3(new_n1154), .A4(new_n1155), .ZN(new_n1156));
  OR2_X1    g0956(.A1(new_n1156), .A2(KEYINPUT58), .ZN(new_n1157));
  OAI22_X1  g0957(.A1(new_n774), .A2(new_n1067), .B1(new_n769), .B2(new_n1004), .ZN(new_n1158));
  OAI22_X1  g0958(.A1(new_n760), .A2(new_n825), .B1(new_n816), .B2(new_n1072), .ZN(new_n1159));
  AOI211_X1 g0959(.A(new_n1158), .B(new_n1159), .C1(G137), .C2(new_n781), .ZN(new_n1160));
  INV_X1    g0960(.A(G128), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1160), .B1(new_n1161), .B2(new_n785), .ZN(new_n1162));
  OR2_X1    g0962(.A1(new_n1162), .A2(KEYINPUT59), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1162), .A2(KEYINPUT59), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n938), .A2(G159), .ZN(new_n1165));
  AOI211_X1 g0965(.A(G33), .B(G41), .C1(new_n772), .C2(G124), .ZN(new_n1166));
  NAND4_X1  g0966(.A1(new_n1163), .A2(new_n1164), .A3(new_n1165), .A4(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1156), .A2(KEYINPUT58), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n202), .B1(new_n331), .B2(G41), .ZN(new_n1169));
  NAND4_X1  g0969(.A1(new_n1157), .A2(new_n1167), .A3(new_n1168), .A4(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1170), .A2(new_n753), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n742), .B1(new_n202), .B2(new_n811), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n1171), .B(new_n1172), .C1(new_n1142), .C2(new_n751), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1149), .A2(new_n1173), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n1146), .A2(new_n1147), .B1(new_n1103), .B2(new_n1111), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1112), .B1(new_n1175), .B2(KEYINPUT57), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1111), .A2(new_n1103), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1148), .A2(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT57), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1174), .B1(new_n1176), .B2(new_n1180), .ZN(new_n1181));
  XNOR2_X1  g0981(.A(new_n1181), .B(KEYINPUT118), .ZN(G375));
  OAI221_X1 g0982(.A(new_n1106), .B1(new_n1108), .B2(new_n1109), .C1(new_n842), .C2(new_n1102), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n976), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1183), .A2(new_n1113), .A3(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n742), .B1(new_n295), .B2(new_n811), .ZN(new_n1186));
  OAI22_X1  g0986(.A1(new_n420), .A2(new_n782), .B1(new_n785), .B2(new_n764), .ZN(new_n1187));
  OAI221_X1 g0987(.A(new_n359), .B1(new_n771), .B2(new_n454), .C1(new_n763), .C2(new_n384), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(new_n766), .A2(G294), .B1(new_n827), .B2(G97), .ZN(new_n1189));
  OAI211_X1 g0989(.A(new_n1189), .B(new_n999), .C1(new_n445), .C2(new_n760), .ZN(new_n1190));
  NOR3_X1   g0990(.A1(new_n1187), .A2(new_n1188), .A3(new_n1190), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n253), .B1(new_n771), .B2(new_n1161), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1192), .B1(G58), .B2(new_n938), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n827), .A2(G159), .B1(new_n788), .B2(G50), .ZN(new_n1194));
  OAI211_X1 g0994(.A(new_n1193), .B(new_n1194), .C1(new_n782), .C2(new_n1004), .ZN(new_n1195));
  XOR2_X1   g0995(.A(new_n1195), .B(KEYINPUT120), .Z(new_n1196));
  AOI22_X1  g0996(.A1(G132), .A2(new_n766), .B1(new_n759), .B2(new_n1068), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1197), .B1(new_n785), .B2(new_n944), .ZN(new_n1198));
  XOR2_X1   g0998(.A(new_n1198), .B(KEYINPUT119), .Z(new_n1199));
  AOI21_X1  g0999(.A(new_n1191), .B1(new_n1196), .B2(new_n1199), .ZN(new_n1200));
  OAI221_X1 g1000(.A(new_n1186), .B1(new_n830), .B2(new_n1200), .C1(new_n906), .C2(new_n751), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(new_n1110), .B2(new_n740), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1185), .A2(new_n1203), .ZN(new_n1204));
  XNOR2_X1  g1004(.A(new_n1204), .B(KEYINPUT121), .ZN(G381));
  NOR2_X1   g1005(.A1(G375), .A2(G378), .ZN(new_n1206));
  INV_X1    g1006(.A(G390), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1207), .A2(new_n832), .ZN(new_n1208));
  OR2_X1    g1008(.A1(G393), .A2(G396), .ZN(new_n1209));
  NOR4_X1   g1009(.A1(new_n1208), .A2(G387), .A3(G381), .A4(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1206), .A2(new_n1210), .ZN(G407));
  INV_X1    g1011(.A(G213), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n1212), .A2(G343), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1206), .A2(new_n1213), .ZN(new_n1214));
  XOR2_X1   g1014(.A(new_n1214), .B(KEYINPUT122), .Z(new_n1215));
  NAND3_X1  g1015(.A1(new_n1215), .A2(G213), .A3(G407), .ZN(G409));
  XNOR2_X1  g1016(.A(G393), .B(new_n800), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1207), .A2(G387), .ZN(new_n1218));
  OAI211_X1 g1018(.A(G390), .B(new_n958), .C1(new_n994), .C2(new_n975), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1217), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1220), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1218), .A2(new_n1219), .A3(new_n1217), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(KEYINPUT61), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT125), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1113), .A2(new_n695), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT124), .ZN(new_n1227));
  AOI21_X1  g1027(.A(KEYINPUT60), .B1(new_n1183), .B2(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1183), .A2(new_n1227), .A3(KEYINPUT60), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1226), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1203), .ZN(new_n1232));
  NOR3_X1   g1032(.A1(new_n1231), .A2(new_n832), .A3(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1230), .ZN(new_n1234));
  OAI211_X1 g1034(.A(new_n695), .B(new_n1113), .C1(new_n1234), .C2(new_n1228), .ZN(new_n1235));
  AOI21_X1  g1035(.A(G384), .B1(new_n1235), .B2(new_n1203), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1225), .B1(new_n1233), .B2(new_n1236), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n832), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1235), .A2(G384), .A3(new_n1203), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1238), .A2(new_n1239), .A3(KEYINPUT125), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1213), .A2(G2897), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1237), .A2(new_n1240), .A3(new_n1241), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n1233), .A2(new_n1236), .ZN(new_n1243));
  OR2_X1    g1043(.A1(new_n1243), .A2(new_n1241), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1175), .A2(new_n1184), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1173), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1246), .B1(new_n1148), .B2(new_n740), .ZN(new_n1247));
  AOI21_X1  g1047(.A(G378), .B1(new_n1245), .B2(new_n1247), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1129), .B1(new_n921), .B2(G330), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(new_n1249), .A2(new_n1131), .B1(new_n1117), .B2(new_n1142), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n913), .B1(new_n1250), .B2(new_n1130), .ZN(new_n1251));
  AND4_X1   g1051(.A1(new_n913), .A2(new_n1130), .A3(new_n1134), .A4(new_n1143), .ZN(new_n1252));
  OAI211_X1 g1052(.A(KEYINPUT57), .B(new_n1177), .C1(new_n1251), .C2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1253), .A2(new_n695), .ZN(new_n1254));
  AOI21_X1  g1054(.A(KEYINPUT57), .B1(new_n1148), .B2(new_n1177), .ZN(new_n1255));
  OAI211_X1 g1055(.A(G378), .B(new_n1247), .C1(new_n1254), .C2(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT123), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1176), .A2(new_n1180), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1259), .A2(KEYINPUT123), .A3(G378), .A4(new_n1247), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1248), .B1(new_n1258), .B2(new_n1260), .ZN(new_n1261));
  OAI211_X1 g1061(.A(new_n1242), .B(new_n1244), .C1(new_n1261), .C2(new_n1213), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1258), .A2(new_n1260), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1248), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1213), .B1(new_n1263), .B2(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1237), .A2(new_n1240), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT62), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(KEYINPUT127), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1265), .A2(new_n1267), .A3(new_n1269), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1268), .A2(KEYINPUT127), .ZN(new_n1271));
  OAI211_X1 g1071(.A(new_n1224), .B(new_n1262), .C1(new_n1270), .C2(new_n1271), .ZN(new_n1272));
  NOR3_X1   g1072(.A1(new_n1261), .A2(new_n1213), .A3(new_n1266), .ZN(new_n1273));
  NOR3_X1   g1073(.A1(new_n1273), .A2(KEYINPUT127), .A3(new_n1268), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1223), .B1(new_n1272), .B2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT126), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1244), .A2(new_n1242), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1224), .B1(new_n1265), .B2(new_n1277), .ZN(new_n1278));
  AOI21_X1  g1078(.A(KEYINPUT63), .B1(new_n1265), .B2(new_n1267), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1213), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1281), .A2(KEYINPUT63), .A3(new_n1282), .A4(new_n1267), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1222), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1284), .A2(new_n1220), .ZN(new_n1285));
  AND2_X1   g1085(.A1(new_n1283), .A2(new_n1285), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1276), .B1(new_n1280), .B2(new_n1286), .ZN(new_n1287));
  OAI211_X1 g1087(.A(new_n1262), .B(new_n1224), .C1(new_n1273), .C2(KEYINPUT63), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1283), .A2(new_n1285), .ZN(new_n1289));
  NOR3_X1   g1089(.A1(new_n1288), .A2(new_n1289), .A3(KEYINPUT126), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1275), .B1(new_n1287), .B2(new_n1290), .ZN(G405));
  NAND2_X1  g1091(.A1(G375), .A2(new_n1115), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1292), .A2(new_n1263), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1293), .A2(new_n1267), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1294), .B1(new_n1243), .B2(new_n1293), .ZN(new_n1295));
  XNOR2_X1  g1095(.A(new_n1295), .B(new_n1223), .ZN(G402));
endmodule


