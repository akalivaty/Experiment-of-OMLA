//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 1 0 1 0 1 1 1 0 1 0 1 0 0 1 0 0 0 0 1 0 0 1 0 1 1 0 1 0 0 1 1 1 0 0 0 1 1 0 0 1 1 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:41 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n715,
    new_n716, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n736, new_n737, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n776, new_n777,
    new_n778, new_n779, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n788, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n818, new_n819, new_n820, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n900, new_n901, new_n903, new_n904, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n964, new_n965, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n981, new_n982, new_n983,
    new_n984, new_n986, new_n987, new_n988, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1010, new_n1011, new_n1012;
  INV_X1    g000(.A(KEYINPUT74), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT22), .ZN(new_n203));
  AOI22_X1  g002(.A1(new_n202), .A2(new_n203), .B1(G211gat), .B2(G218gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n204), .B1(new_n202), .B2(new_n203), .ZN(new_n205));
  XNOR2_X1  g004(.A(G197gat), .B(G204gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G211gat), .B(G218gat), .ZN(new_n208));
  XNOR2_X1  g007(.A(new_n207), .B(new_n208), .ZN(new_n209));
  XNOR2_X1  g008(.A(new_n209), .B(KEYINPUT75), .ZN(new_n210));
  XNOR2_X1  g009(.A(KEYINPUT76), .B(KEYINPUT29), .ZN(new_n211));
  XOR2_X1   g010(.A(G141gat), .B(G148gat), .Z(new_n212));
  INV_X1    g011(.A(G155gat), .ZN(new_n213));
  INV_X1    g012(.A(G162gat), .ZN(new_n214));
  OAI21_X1  g013(.A(KEYINPUT2), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n212), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g015(.A(G155gat), .B(G162gat), .ZN(new_n217));
  INV_X1    g016(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n212), .A2(new_n217), .A3(new_n215), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n211), .B1(new_n221), .B2(KEYINPUT3), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n210), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(G228gat), .A2(G233gat), .ZN(new_n224));
  INV_X1    g023(.A(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT3), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n226), .B1(new_n209), .B2(KEYINPUT29), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(new_n221), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n223), .A2(new_n225), .A3(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(new_n211), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n226), .B1(new_n209), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n222), .A2(new_n209), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT86), .ZN(new_n234));
  AOI22_X1  g033(.A1(new_n221), .A2(new_n232), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n222), .A2(KEYINPUT86), .A3(new_n209), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n225), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  OAI21_X1  g036(.A(G22gat), .B1(new_n230), .B2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(G22gat), .ZN(new_n239));
  AND2_X1   g038(.A1(new_n235), .A2(new_n236), .ZN(new_n240));
  OAI211_X1 g039(.A(new_n239), .B(new_n229), .C1(new_n240), .C2(new_n225), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n238), .A2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT87), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n229), .B1(new_n240), .B2(new_n225), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n243), .B1(new_n244), .B2(G22gat), .ZN(new_n245));
  XNOR2_X1  g044(.A(G78gat), .B(G106gat), .ZN(new_n246));
  XNOR2_X1  g045(.A(KEYINPUT31), .B(G50gat), .ZN(new_n247));
  XOR2_X1   g046(.A(new_n246), .B(new_n247), .Z(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n242), .B1(new_n245), .B2(new_n249), .ZN(new_n250));
  NAND4_X1  g049(.A1(new_n238), .A2(new_n241), .A3(new_n243), .A4(new_n248), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  AND2_X1   g051(.A1(new_n219), .A2(new_n220), .ZN(new_n253));
  XNOR2_X1  g052(.A(KEYINPUT69), .B(G134gat), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(G127gat), .ZN(new_n255));
  XNOR2_X1  g054(.A(KEYINPUT70), .B(G127gat), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(G134gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(G113gat), .A2(G120gat), .ZN(new_n258));
  INV_X1    g057(.A(G113gat), .ZN(new_n259));
  INV_X1    g058(.A(G120gat), .ZN(new_n260));
  AOI21_X1  g059(.A(KEYINPUT1), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  AOI22_X1  g060(.A1(new_n255), .A2(new_n257), .B1(new_n258), .B2(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(KEYINPUT71), .B(G113gat), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n263), .A2(new_n260), .ZN(new_n264));
  INV_X1    g063(.A(G127gat), .ZN(new_n265));
  OR2_X1    g064(.A1(new_n265), .A2(G134gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(G134gat), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n266), .A2(new_n261), .A3(new_n267), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n264), .A2(new_n268), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n262), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n253), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(KEYINPUT81), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT81), .ZN(new_n274));
  NAND4_X1  g073(.A1(new_n253), .A2(new_n270), .A3(new_n274), .A4(new_n271), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n253), .A2(new_n270), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(KEYINPUT4), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n273), .A2(new_n275), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(G225gat), .A2(G233gat), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n262), .ZN(new_n281));
  INV_X1    g080(.A(new_n269), .ZN(new_n282));
  AOI22_X1  g081(.A1(new_n281), .A2(new_n282), .B1(new_n221), .B2(KEYINPUT3), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n253), .A2(new_n226), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n280), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n278), .A2(KEYINPUT82), .A3(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(KEYINPUT84), .B(KEYINPUT5), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n281), .A2(new_n282), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(new_n221), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT83), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n289), .A2(new_n290), .A3(new_n276), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n288), .A2(KEYINPUT83), .A3(new_n221), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n291), .A2(new_n280), .A3(new_n292), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n286), .A2(new_n287), .A3(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(KEYINPUT82), .B1(new_n278), .B2(new_n285), .ZN(new_n295));
  OAI21_X1  g094(.A(KEYINPUT85), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n295), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT85), .ZN(new_n298));
  AND2_X1   g097(.A1(new_n293), .A2(new_n287), .ZN(new_n299));
  NAND4_X1  g098(.A1(new_n297), .A2(new_n298), .A3(new_n299), .A4(new_n286), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n296), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n285), .ZN(new_n302));
  INV_X1    g101(.A(new_n272), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n271), .B1(new_n253), .B2(new_n270), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NOR3_X1   g104(.A1(new_n302), .A2(new_n305), .A3(new_n287), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n301), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT89), .ZN(new_n309));
  XNOR2_X1  g108(.A(G1gat), .B(G29gat), .ZN(new_n310));
  XNOR2_X1  g109(.A(new_n310), .B(KEYINPUT0), .ZN(new_n311));
  XNOR2_X1  g110(.A(G57gat), .B(G85gat), .ZN(new_n312));
  XOR2_X1   g111(.A(new_n311), .B(new_n312), .Z(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n308), .A2(new_n309), .A3(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT88), .ZN(new_n316));
  AOI22_X1  g115(.A1(new_n277), .A2(new_n272), .B1(new_n284), .B2(new_n283), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n316), .B1(new_n317), .B2(new_n279), .ZN(new_n318));
  AND2_X1   g117(.A1(new_n283), .A2(new_n284), .ZN(new_n319));
  OAI211_X1 g118(.A(KEYINPUT88), .B(new_n280), .C1(new_n305), .C2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT39), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n314), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n291), .A2(new_n292), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n322), .B1(new_n324), .B2(new_n279), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n325), .A2(new_n318), .A3(new_n320), .ZN(new_n326));
  AND3_X1   g125(.A1(new_n323), .A2(KEYINPUT40), .A3(new_n326), .ZN(new_n327));
  AOI21_X1  g126(.A(KEYINPUT40), .B1(new_n323), .B2(new_n326), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n306), .B1(new_n296), .B2(new_n300), .ZN(new_n330));
  OAI21_X1  g129(.A(KEYINPUT89), .B1(new_n330), .B2(new_n313), .ZN(new_n331));
  AND3_X1   g130(.A1(new_n315), .A2(new_n329), .A3(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT80), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT77), .ZN(new_n334));
  NAND2_X1  g133(.A1(G226gat), .A2(G233gat), .ZN(new_n335));
  INV_X1    g134(.A(G169gat), .ZN(new_n336));
  INV_X1    g135(.A(G176gat), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  NOR2_X1   g138(.A1(G169gat), .A2(G176gat), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT66), .ZN(new_n341));
  XNOR2_X1  g140(.A(new_n340), .B(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT23), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n339), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT67), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  XNOR2_X1  g145(.A(new_n340), .B(KEYINPUT66), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(KEYINPUT23), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n348), .A2(KEYINPUT67), .A3(new_n339), .ZN(new_n349));
  OAI21_X1  g148(.A(KEYINPUT25), .B1(new_n340), .B2(KEYINPUT23), .ZN(new_n350));
  XOR2_X1   g149(.A(KEYINPUT68), .B(G183gat), .Z(new_n351));
  INV_X1    g150(.A(G190gat), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(G183gat), .ZN(new_n354));
  OAI21_X1  g153(.A(KEYINPUT24), .B1(new_n354), .B2(new_n352), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT24), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n356), .A2(G183gat), .A3(G190gat), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n350), .B1(new_n353), .B2(new_n358), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n346), .A2(new_n349), .A3(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT25), .ZN(new_n361));
  INV_X1    g160(.A(new_n340), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n338), .B1(new_n362), .B2(new_n343), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n363), .B1(new_n343), .B2(new_n362), .ZN(new_n364));
  AOI22_X1  g163(.A1(new_n355), .A2(new_n357), .B1(new_n354), .B2(new_n352), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n361), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  OR2_X1    g165(.A1(new_n342), .A2(KEYINPUT26), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n338), .B1(KEYINPUT26), .B2(new_n362), .ZN(new_n368));
  AOI22_X1  g167(.A1(new_n367), .A2(new_n368), .B1(G183gat), .B2(G190gat), .ZN(new_n369));
  XNOR2_X1  g168(.A(KEYINPUT27), .B(G183gat), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n370), .A2(KEYINPUT28), .A3(new_n352), .ZN(new_n371));
  NOR2_X1   g170(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n372));
  XNOR2_X1  g171(.A(KEYINPUT68), .B(G183gat), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n372), .B1(new_n373), .B2(KEYINPUT27), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n374), .A2(G190gat), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n371), .B1(new_n375), .B2(KEYINPUT28), .ZN(new_n376));
  AOI22_X1  g175(.A1(new_n360), .A2(new_n366), .B1(new_n369), .B2(new_n376), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n335), .B1(new_n377), .B2(new_n231), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n359), .B1(new_n344), .B2(new_n345), .ZN(new_n379));
  AOI21_X1  g178(.A(KEYINPUT67), .B1(new_n348), .B2(new_n339), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n366), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n369), .A2(new_n376), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(new_n335), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n334), .B1(new_n378), .B2(new_n385), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n384), .B1(new_n383), .B2(new_n211), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n387), .A2(KEYINPUT77), .ZN(new_n388));
  OAI211_X1 g187(.A(KEYINPUT78), .B(new_n210), .C1(new_n386), .C2(new_n388), .ZN(new_n389));
  OR3_X1    g188(.A1(new_n377), .A2(KEYINPUT79), .A3(new_n335), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n385), .A2(KEYINPUT79), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT29), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n384), .B1(new_n383), .B2(new_n392), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n390), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(new_n209), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n389), .A2(new_n396), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n377), .A2(new_n335), .ZN(new_n398));
  OAI21_X1  g197(.A(KEYINPUT77), .B1(new_n387), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n378), .A2(new_n334), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(KEYINPUT78), .B1(new_n401), .B2(new_n210), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n333), .B1(new_n397), .B2(new_n402), .ZN(new_n403));
  XNOR2_X1  g202(.A(G8gat), .B(G36gat), .ZN(new_n404));
  XNOR2_X1  g203(.A(G64gat), .B(G92gat), .ZN(new_n405));
  XOR2_X1   g204(.A(new_n404), .B(new_n405), .Z(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n210), .B1(new_n386), .B2(new_n388), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT78), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND4_X1  g209(.A1(new_n410), .A2(KEYINPUT80), .A3(new_n396), .A4(new_n389), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n403), .A2(new_n407), .A3(new_n411), .ZN(new_n412));
  NAND4_X1  g211(.A1(new_n410), .A2(new_n406), .A3(new_n396), .A4(new_n389), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT30), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n397), .A2(new_n402), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n416), .A2(KEYINPUT30), .A3(new_n406), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n412), .A2(new_n415), .A3(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n252), .B1(new_n332), .B2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT37), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n410), .A2(new_n420), .A3(new_n396), .A4(new_n389), .ZN(new_n421));
  INV_X1    g220(.A(new_n210), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n399), .A2(new_n400), .A3(new_n422), .ZN(new_n423));
  OAI211_X1 g222(.A(new_n209), .B(new_n390), .C1(new_n391), .C2(new_n393), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(KEYINPUT38), .B1(new_n425), .B2(KEYINPUT37), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n421), .A2(new_n426), .A3(new_n407), .ZN(new_n427));
  AND2_X1   g226(.A1(new_n427), .A2(new_n413), .ZN(new_n428));
  AOI21_X1  g227(.A(KEYINPUT6), .B1(new_n330), .B2(new_n313), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n315), .A2(new_n429), .A3(new_n331), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n308), .A2(KEYINPUT6), .A3(new_n314), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT90), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n330), .A2(new_n313), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n434), .A2(KEYINPUT90), .A3(KEYINPUT6), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n428), .A2(new_n430), .A3(new_n433), .A4(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT38), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n403), .A2(KEYINPUT37), .A3(new_n411), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n406), .B1(new_n416), .B2(new_n420), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n437), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n419), .B1(new_n436), .B2(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n301), .A2(new_n313), .A3(new_n307), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT6), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n431), .B1(new_n444), .B2(new_n434), .ZN(new_n445));
  XNOR2_X1  g244(.A(new_n413), .B(KEYINPUT30), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n445), .A2(new_n446), .A3(new_n412), .ZN(new_n447));
  XNOR2_X1  g246(.A(KEYINPUT72), .B(G71gat), .ZN(new_n448));
  INV_X1    g247(.A(G99gat), .ZN(new_n449));
  XNOR2_X1  g248(.A(new_n448), .B(new_n449), .ZN(new_n450));
  XOR2_X1   g249(.A(G15gat), .B(G43gat), .Z(new_n451));
  XNOR2_X1  g250(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n383), .A2(new_n270), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n377), .A2(new_n288), .ZN(new_n454));
  NAND2_X1  g253(.A1(G227gat), .A2(G233gat), .ZN(new_n455));
  XOR2_X1   g254(.A(new_n455), .B(KEYINPUT64), .Z(new_n456));
  XOR2_X1   g255(.A(new_n456), .B(KEYINPUT65), .Z(new_n457));
  NAND3_X1  g256(.A1(new_n453), .A2(new_n454), .A3(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT33), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n452), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n458), .A2(KEYINPUT32), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  OAI211_X1 g261(.A(new_n458), .B(KEYINPUT32), .C1(new_n459), .C2(new_n452), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n453), .A2(new_n454), .ZN(new_n465));
  INV_X1    g264(.A(new_n456), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n457), .A2(KEYINPUT34), .ZN(new_n468));
  AOI22_X1  g267(.A1(new_n467), .A2(KEYINPUT34), .B1(new_n465), .B2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n464), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n462), .A2(new_n469), .A3(new_n463), .ZN(new_n472));
  NOR2_X1   g271(.A1(KEYINPUT73), .A2(KEYINPUT36), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT73), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT36), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  OAI211_X1 g275(.A(new_n471), .B(new_n472), .C1(new_n473), .C2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(new_n472), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n469), .B1(new_n462), .B2(new_n463), .ZN(new_n479));
  OAI22_X1  g278(.A1(new_n478), .A2(new_n479), .B1(new_n474), .B2(new_n475), .ZN(new_n480));
  AOI22_X1  g279(.A1(new_n447), .A2(new_n252), .B1(new_n477), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n441), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n471), .A2(new_n472), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n252), .A2(new_n483), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n445), .A2(new_n446), .A3(new_n484), .A4(new_n412), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(KEYINPUT35), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n430), .A2(new_n433), .A3(new_n435), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT35), .ZN(new_n488));
  AND3_X1   g287(.A1(new_n412), .A2(new_n415), .A3(new_n417), .ZN(new_n489));
  NAND4_X1  g288(.A1(new_n487), .A2(new_n488), .A3(new_n489), .A4(new_n484), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n486), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n482), .A2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(G57gat), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(G64gat), .ZN(new_n494));
  INV_X1    g293(.A(G64gat), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(G57gat), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(G71gat), .A2(G78gat), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT9), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n497), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n498), .A2(KEYINPUT97), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT96), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n503), .B1(G71gat), .B2(G78gat), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT97), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n505), .A2(G71gat), .A3(G78gat), .ZN(new_n506));
  AND3_X1   g305(.A1(new_n502), .A2(new_n504), .A3(new_n506), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n504), .B1(new_n502), .B2(new_n506), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n501), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  AND2_X1   g308(.A1(G71gat), .A2(G78gat), .ZN(new_n510));
  NOR2_X1   g309(.A1(G71gat), .A2(G78gat), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AND3_X1   g311(.A1(new_n497), .A2(new_n512), .A3(new_n500), .ZN(new_n513));
  INV_X1    g312(.A(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n509), .A2(new_n514), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n515), .A2(KEYINPUT21), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n516), .B(KEYINPUT98), .ZN(new_n517));
  XOR2_X1   g316(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n518));
  XNOR2_X1  g317(.A(new_n517), .B(new_n518), .ZN(new_n519));
  XOR2_X1   g318(.A(G183gat), .B(G211gat), .Z(new_n520));
  XOR2_X1   g319(.A(new_n519), .B(new_n520), .Z(new_n521));
  NAND2_X1  g320(.A1(new_n239), .A2(G15gat), .ZN(new_n522));
  INV_X1    g321(.A(G15gat), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(G22gat), .ZN(new_n524));
  INV_X1    g323(.A(G1gat), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(KEYINPUT16), .ZN(new_n526));
  AND3_X1   g325(.A1(new_n522), .A2(new_n524), .A3(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(G8gat), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n522), .A2(new_n524), .ZN(new_n530));
  AOI22_X1  g329(.A1(new_n530), .A2(new_n525), .B1(KEYINPUT93), .B2(G8gat), .ZN(new_n531));
  AND2_X1   g330(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT92), .ZN(new_n533));
  AOI21_X1  g332(.A(G1gat), .B1(new_n522), .B2(new_n524), .ZN(new_n534));
  AOI22_X1  g333(.A1(new_n527), .A2(new_n533), .B1(new_n534), .B2(KEYINPUT93), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n522), .A2(new_n524), .A3(new_n526), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(KEYINPUT92), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n528), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  AOI211_X1 g337(.A(new_n532), .B(new_n538), .C1(KEYINPUT21), .C2(new_n515), .ZN(new_n539));
  XNOR2_X1  g338(.A(G127gat), .B(G155gat), .ZN(new_n540));
  NAND2_X1  g339(.A1(G231gat), .A2(G233gat), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n540), .B(new_n541), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n539), .B(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n521), .A2(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n519), .B(new_n520), .ZN(new_n545));
  INV_X1    g344(.A(new_n543), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(G36gat), .ZN(new_n549));
  AND2_X1   g348(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n550));
  NOR2_X1   g349(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n549), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(G29gat), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n553), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(G50gat), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(G43gat), .ZN(new_n557));
  INV_X1    g356(.A(G43gat), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n558), .A2(G50gat), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n557), .A2(new_n559), .A3(KEYINPUT15), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n555), .A2(new_n561), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n556), .A2(G43gat), .ZN(new_n563));
  AOI21_X1  g362(.A(KEYINPUT15), .B1(new_n563), .B2(KEYINPUT91), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT91), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n557), .A2(new_n559), .A3(new_n565), .ZN(new_n566));
  AOI22_X1  g365(.A1(new_n564), .A2(new_n566), .B1(new_n552), .B2(new_n554), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n562), .B1(new_n567), .B2(new_n561), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n568), .A2(KEYINPUT17), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT17), .ZN(new_n570));
  OAI211_X1 g369(.A(new_n570), .B(new_n562), .C1(new_n567), .C2(new_n561), .ZN(new_n571));
  NAND2_X1  g370(.A1(G99gat), .A2(G106gat), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(KEYINPUT8), .ZN(new_n573));
  NAND2_X1  g372(.A1(G85gat), .A2(G92gat), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT7), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(G85gat), .ZN(new_n577));
  INV_X1    g376(.A(G92gat), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g378(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n580));
  NAND4_X1  g379(.A1(new_n573), .A2(new_n576), .A3(new_n579), .A4(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n572), .ZN(new_n582));
  NOR2_X1   g381(.A1(G99gat), .A2(G106gat), .ZN(new_n583));
  OR2_X1    g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  AND3_X1   g384(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n586));
  AOI21_X1  g385(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n582), .A2(new_n583), .ZN(new_n589));
  AOI22_X1  g388(.A1(KEYINPUT8), .A2(new_n572), .B1(new_n577), .B2(new_n578), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  NAND4_X1  g390(.A1(new_n569), .A2(new_n571), .A3(new_n585), .A4(new_n591), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n560), .B1(new_n552), .B2(new_n554), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n564), .A2(new_n566), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n594), .A2(new_n555), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n593), .B1(new_n595), .B2(new_n560), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n585), .A2(new_n591), .ZN(new_n597));
  AND2_X1   g396(.A1(G232gat), .A2(G233gat), .ZN(new_n598));
  AOI22_X1  g397(.A1(new_n596), .A2(new_n597), .B1(KEYINPUT41), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n592), .A2(new_n599), .ZN(new_n600));
  XOR2_X1   g399(.A(G190gat), .B(G218gat), .Z(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n600), .B(new_n602), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n598), .A2(KEYINPUT41), .ZN(new_n604));
  XNOR2_X1  g403(.A(G134gat), .B(G162gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n604), .B(new_n605), .ZN(new_n606));
  OR2_X1    g405(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n603), .A2(new_n606), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n548), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n502), .A2(new_n506), .ZN(new_n611));
  INV_X1    g410(.A(new_n504), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n502), .A2(new_n504), .A3(new_n506), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n513), .B1(new_n615), .B2(new_n501), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n581), .A2(new_n584), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n589), .B1(new_n588), .B2(new_n590), .ZN(new_n618));
  OAI21_X1  g417(.A(KEYINPUT10), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n616), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n597), .A2(new_n509), .A3(new_n514), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT99), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n581), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(new_n589), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n581), .A2(new_n584), .A3(new_n622), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n621), .B1(new_n626), .B2(new_n616), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT10), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n620), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(G230gat), .A2(G233gat), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  OAI21_X1  g430(.A(KEYINPUT100), .B1(new_n629), .B2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT100), .ZN(new_n633));
  AOI22_X1  g432(.A1(new_n494), .A2(new_n496), .B1(new_n499), .B2(new_n498), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n634), .B1(new_n613), .B2(new_n614), .ZN(new_n635));
  OAI211_X1 g434(.A(new_n624), .B(new_n625), .C1(new_n635), .C2(new_n513), .ZN(new_n636));
  AOI21_X1  g435(.A(KEYINPUT10), .B1(new_n636), .B2(new_n621), .ZN(new_n637));
  OAI211_X1 g436(.A(new_n633), .B(new_n630), .C1(new_n637), .C2(new_n620), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n636), .A2(new_n631), .A3(new_n621), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(G120gat), .B(G148gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(KEYINPUT101), .ZN(new_n642));
  XNOR2_X1  g441(.A(G176gat), .B(G204gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n642), .B(new_n643), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n640), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n632), .A2(new_n638), .A3(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT102), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND4_X1  g447(.A1(new_n632), .A2(KEYINPUT102), .A3(new_n638), .A4(new_n645), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n629), .A2(new_n631), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n644), .B1(new_n651), .B2(new_n640), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n610), .A2(new_n653), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n596), .B1(new_n538), .B2(new_n532), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT94), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n530), .A2(KEYINPUT93), .A3(new_n525), .ZN(new_n657));
  NAND4_X1  g456(.A1(new_n522), .A2(new_n524), .A3(new_n526), .A4(new_n533), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n537), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  AOI22_X1  g458(.A1(new_n659), .A2(G8gat), .B1(new_n529), .B2(new_n531), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n660), .A2(new_n568), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n655), .A2(new_n656), .A3(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(G229gat), .A2(G233gat), .ZN(new_n663));
  XOR2_X1   g462(.A(new_n663), .B(KEYINPUT13), .Z(new_n664));
  NAND3_X1  g463(.A1(new_n660), .A2(KEYINPUT94), .A3(new_n568), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n662), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT95), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND4_X1  g467(.A1(new_n662), .A2(KEYINPUT95), .A3(new_n664), .A4(new_n665), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n569), .A2(new_n660), .A3(new_n571), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n671), .A2(new_n663), .A3(new_n655), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(KEYINPUT18), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g473(.A(G113gat), .B(G141gat), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n675), .B(G197gat), .ZN(new_n676));
  XOR2_X1   g475(.A(KEYINPUT11), .B(G169gat), .Z(new_n677));
  XNOR2_X1  g476(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n678), .B(KEYINPUT12), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n674), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n670), .A2(new_n673), .A3(new_n679), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n654), .A2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  AOI21_X1  g484(.A(KEYINPUT103), .B1(new_n492), .B2(new_n685), .ZN(new_n686));
  AOI22_X1  g485(.A1(new_n441), .A2(new_n481), .B1(new_n486), .B2(new_n490), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT103), .ZN(new_n688));
  NOR3_X1   g487(.A1(new_n687), .A2(new_n688), .A3(new_n684), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n690), .A2(new_n445), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(new_n525), .ZN(G1324gat));
  OAI21_X1  g491(.A(new_n418), .B1(new_n686), .B2(new_n689), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT104), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  OAI211_X1 g494(.A(KEYINPUT104), .B(new_n418), .C1(new_n686), .C2(new_n689), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n695), .A2(G8gat), .A3(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n690), .ZN(new_n698));
  XOR2_X1   g497(.A(KEYINPUT16), .B(G8gat), .Z(new_n699));
  NAND4_X1  g498(.A1(new_n698), .A2(KEYINPUT42), .A3(new_n418), .A4(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n699), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n701), .B1(new_n695), .B2(new_n696), .ZN(new_n702));
  OAI211_X1 g501(.A(new_n697), .B(new_n700), .C1(new_n702), .C2(KEYINPUT42), .ZN(G1325gat));
  NAND2_X1  g502(.A1(new_n477), .A2(new_n480), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(KEYINPUT106), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT106), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n477), .A2(new_n480), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  NOR3_X1   g507(.A1(new_n690), .A2(new_n523), .A3(new_n708), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n523), .B1(new_n690), .B2(new_n483), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT105), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  OAI211_X1 g511(.A(KEYINPUT105), .B(new_n523), .C1(new_n690), .C2(new_n483), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n709), .B1(new_n712), .B2(new_n713), .ZN(G1326gat));
  NAND2_X1  g513(.A1(new_n698), .A2(new_n252), .ZN(new_n715));
  XNOR2_X1  g514(.A(KEYINPUT43), .B(G22gat), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n715), .B(new_n716), .ZN(G1327gat));
  NOR2_X1   g516(.A1(new_n687), .A2(new_n609), .ZN(new_n718));
  INV_X1    g517(.A(new_n683), .ZN(new_n719));
  NOR3_X1   g518(.A1(new_n548), .A2(new_n719), .A3(new_n653), .ZN(new_n720));
  AND2_X1   g519(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(new_n445), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n721), .A2(new_n553), .A3(new_n722), .ZN(new_n723));
  XOR2_X1   g522(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n724));
  XNOR2_X1  g523(.A(new_n723), .B(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(new_n609), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n492), .A2(KEYINPUT44), .A3(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT44), .ZN(new_n728));
  AOI22_X1  g527(.A1(new_n447), .A2(new_n252), .B1(new_n705), .B2(new_n707), .ZN(new_n729));
  AOI22_X1  g528(.A1(new_n441), .A2(new_n729), .B1(new_n486), .B2(new_n490), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n728), .B1(new_n730), .B2(new_n609), .ZN(new_n731));
  AND2_X1   g530(.A1(new_n727), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(new_n720), .ZN(new_n733));
  OAI21_X1  g532(.A(G29gat), .B1(new_n733), .B2(new_n445), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n725), .A2(new_n734), .ZN(G1328gat));
  NAND3_X1  g534(.A1(new_n721), .A2(new_n549), .A3(new_n418), .ZN(new_n736));
  OR2_X1    g535(.A1(new_n736), .A2(KEYINPUT46), .ZN(new_n737));
  OAI21_X1  g536(.A(G36gat), .B1(new_n733), .B2(new_n489), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n736), .A2(KEYINPUT46), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n737), .A2(new_n738), .A3(new_n739), .ZN(G1329gat));
  NOR2_X1   g539(.A1(new_n483), .A2(G43gat), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n492), .A2(new_n726), .A3(new_n720), .A4(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(KEYINPUT109), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT109), .ZN(new_n744));
  NAND4_X1  g543(.A1(new_n718), .A2(new_n744), .A3(new_n720), .A4(new_n741), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  AOI21_X1  g545(.A(KEYINPUT47), .B1(new_n746), .B2(KEYINPUT108), .ZN(new_n747));
  INV_X1    g546(.A(new_n708), .ZN(new_n748));
  NAND4_X1  g547(.A1(new_n727), .A2(new_n731), .A3(new_n748), .A4(new_n720), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(G43gat), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(new_n746), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n747), .A2(new_n751), .ZN(new_n752));
  OAI211_X1 g551(.A(new_n750), .B(new_n746), .C1(KEYINPUT108), .C2(KEYINPUT47), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(G1330gat));
  NAND4_X1  g553(.A1(new_n727), .A2(new_n731), .A3(new_n252), .A4(new_n720), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(G50gat), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT110), .ZN(new_n757));
  AOI21_X1  g556(.A(KEYINPUT48), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n721), .A2(new_n556), .A3(new_n252), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n756), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  OAI211_X1 g560(.A(new_n756), .B(new_n759), .C1(new_n757), .C2(KEYINPUT48), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(G1331gat));
  NAND2_X1  g562(.A1(new_n441), .A2(new_n729), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(new_n491), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT111), .ZN(new_n766));
  INV_X1    g565(.A(new_n652), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n767), .B1(new_n648), .B2(new_n649), .ZN(new_n768));
  NOR3_X1   g567(.A1(new_n610), .A2(new_n683), .A3(new_n768), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n765), .A2(new_n766), .A3(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(new_n769), .ZN(new_n771));
  OAI21_X1  g570(.A(KEYINPUT111), .B1(new_n730), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n773), .A2(new_n445), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n774), .B(new_n493), .ZN(G1332gat));
  INV_X1    g574(.A(new_n773), .ZN(new_n776));
  XNOR2_X1  g575(.A(KEYINPUT49), .B(G64gat), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n776), .A2(new_n418), .A3(new_n777), .ZN(new_n778));
  OAI22_X1  g577(.A1(new_n773), .A2(new_n489), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n778), .A2(new_n779), .ZN(G1333gat));
  OAI21_X1  g579(.A(G71gat), .B1(new_n773), .B2(new_n708), .ZN(new_n781));
  OR2_X1    g580(.A1(new_n483), .A2(G71gat), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n781), .B1(new_n773), .B2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT50), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  OAI211_X1 g584(.A(new_n781), .B(KEYINPUT50), .C1(new_n773), .C2(new_n782), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(G1334gat));
  NAND2_X1  g586(.A1(new_n776), .A2(new_n252), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n788), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g588(.A1(new_n548), .A2(new_n683), .ZN(new_n790));
  INV_X1    g589(.A(new_n790), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n791), .A2(new_n768), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n732), .A2(new_n792), .ZN(new_n793));
  OAI21_X1  g592(.A(G85gat), .B1(new_n793), .B2(new_n445), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT51), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n791), .B1(KEYINPUT112), .B2(new_n795), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n765), .A2(new_n726), .A3(new_n796), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n795), .A2(KEYINPUT112), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(new_n798), .ZN(new_n800));
  NAND4_X1  g599(.A1(new_n765), .A2(new_n726), .A3(new_n796), .A4(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n799), .A2(new_n653), .A3(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n722), .A2(new_n577), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n794), .B1(new_n802), .B2(new_n803), .ZN(G1336gat));
  NOR2_X1   g603(.A1(new_n489), .A2(G92gat), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n799), .A2(new_n653), .A3(new_n801), .A4(new_n805), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n727), .A2(new_n731), .A3(new_n418), .A4(new_n792), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(G92gat), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT113), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT52), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n809), .A2(new_n810), .ZN(new_n813));
  AND4_X1   g612(.A1(new_n806), .A2(new_n808), .A3(new_n812), .A4(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n811), .B1(new_n807), .B2(G92gat), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n813), .B1(new_n815), .B2(new_n806), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n814), .A2(new_n816), .ZN(G1337gat));
  OAI21_X1  g616(.A(G99gat), .B1(new_n793), .B2(new_n708), .ZN(new_n818));
  NOR3_X1   g617(.A1(new_n483), .A2(G99gat), .A3(new_n768), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n799), .A2(new_n801), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n818), .A2(new_n820), .ZN(G1338gat));
  NAND4_X1  g620(.A1(new_n727), .A2(new_n731), .A3(new_n252), .A4(new_n792), .ZN(new_n822));
  XOR2_X1   g621(.A(KEYINPUT114), .B(G106gat), .Z(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(new_n252), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n825), .A2(G106gat), .ZN(new_n826));
  NAND4_X1  g625(.A1(new_n799), .A2(new_n653), .A3(new_n801), .A4(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n824), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(KEYINPUT53), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT53), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n824), .A2(new_n827), .A3(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n829), .A2(new_n831), .ZN(G1339gat));
  INV_X1    g631(.A(KEYINPUT121), .ZN(new_n833));
  INV_X1    g632(.A(new_n548), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT118), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n664), .B1(new_n662), .B2(new_n665), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n663), .B1(new_n671), .B2(new_n655), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n678), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(KEYINPUT117), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT117), .ZN(new_n840));
  OAI211_X1 g639(.A(new_n840), .B(new_n678), .C1(new_n836), .C2(new_n837), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n653), .A2(new_n835), .A3(new_n682), .A4(new_n842), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n682), .A2(new_n841), .A3(new_n839), .ZN(new_n844));
  OAI21_X1  g643(.A(KEYINPUT118), .B1(new_n844), .B2(new_n768), .ZN(new_n845));
  AND2_X1   g644(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT54), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n847), .B1(new_n629), .B2(new_n631), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n632), .A2(new_n848), .A3(new_n638), .ZN(new_n849));
  OAI211_X1 g648(.A(new_n847), .B(new_n630), .C1(new_n637), .C2(new_n620), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n850), .A2(KEYINPUT115), .A3(new_n644), .ZN(new_n851));
  INV_X1    g650(.A(new_n851), .ZN(new_n852));
  AOI21_X1  g651(.A(KEYINPUT115), .B1(new_n850), .B2(new_n644), .ZN(new_n853));
  OAI211_X1 g652(.A(new_n849), .B(KEYINPUT55), .C1(new_n852), .C2(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n650), .A2(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(new_n853), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(new_n851), .ZN(new_n857));
  AOI21_X1  g656(.A(KEYINPUT55), .B1(new_n857), .B2(new_n849), .ZN(new_n858));
  OAI21_X1  g657(.A(KEYINPUT116), .B1(new_n855), .B2(new_n858), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n849), .B1(new_n852), .B2(new_n853), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT55), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT116), .ZN(new_n863));
  NAND4_X1  g662(.A1(new_n862), .A2(new_n863), .A3(new_n650), .A4(new_n854), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n859), .A2(new_n683), .A3(new_n864), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n726), .B1(new_n846), .B2(new_n865), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n609), .A2(new_n844), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n859), .A2(new_n867), .A3(new_n864), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n834), .B1(new_n866), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n654), .A2(new_n719), .ZN(new_n871));
  AND3_X1   g670(.A1(new_n870), .A2(KEYINPUT119), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(KEYINPUT119), .B1(new_n870), .B2(new_n871), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n722), .A2(new_n489), .ZN(new_n875));
  INV_X1    g674(.A(new_n875), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n874), .A2(new_n825), .A3(new_n876), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n877), .A2(new_n483), .A3(new_n719), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT119), .ZN(new_n879));
  AND3_X1   g678(.A1(new_n859), .A2(new_n683), .A3(new_n864), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n843), .A2(new_n845), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n609), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n548), .B1(new_n882), .B2(new_n868), .ZN(new_n883));
  NOR3_X1   g682(.A1(new_n610), .A2(new_n683), .A3(new_n653), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n879), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n870), .A2(KEYINPUT119), .A3(new_n871), .ZN(new_n886));
  NAND4_X1  g685(.A1(new_n885), .A2(new_n722), .A3(new_n484), .A4(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT120), .ZN(new_n888));
  AND2_X1   g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n887), .A2(new_n888), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n489), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n683), .A2(new_n263), .ZN(new_n892));
  OAI221_X1 g691(.A(new_n833), .B1(new_n878), .B2(new_n259), .C1(new_n891), .C2(new_n892), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n878), .A2(new_n259), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n874), .A2(KEYINPUT120), .A3(new_n722), .A4(new_n484), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n887), .A2(new_n888), .ZN(new_n896));
  AOI211_X1 g695(.A(new_n418), .B(new_n892), .C1(new_n895), .C2(new_n896), .ZN(new_n897));
  OAI21_X1  g696(.A(KEYINPUT121), .B1(new_n894), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n893), .A2(new_n898), .ZN(G1340gat));
  NOR4_X1   g698(.A1(new_n877), .A2(new_n260), .A3(new_n483), .A4(new_n768), .ZN(new_n900));
  OR2_X1    g699(.A1(new_n891), .A2(new_n768), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n900), .B1(new_n901), .B2(new_n260), .ZN(G1341gat));
  NAND2_X1  g701(.A1(new_n548), .A2(new_n256), .ZN(new_n903));
  NOR3_X1   g702(.A1(new_n877), .A2(new_n483), .A3(new_n834), .ZN(new_n904));
  OAI22_X1  g703(.A1(new_n891), .A2(new_n903), .B1(new_n904), .B2(new_n256), .ZN(G1342gat));
  INV_X1    g704(.A(KEYINPUT122), .ZN(new_n906));
  NOR3_X1   g705(.A1(new_n872), .A2(new_n873), .A3(new_n252), .ZN(new_n907));
  INV_X1    g706(.A(new_n483), .ZN(new_n908));
  NAND4_X1  g707(.A1(new_n907), .A2(new_n908), .A3(new_n726), .A4(new_n876), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(G134gat), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n489), .A2(new_n254), .A3(new_n726), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n911), .B1(new_n895), .B2(new_n896), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT56), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n910), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  AOI211_X1 g713(.A(KEYINPUT56), .B(new_n911), .C1(new_n895), .C2(new_n896), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n906), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  INV_X1    g715(.A(new_n911), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n917), .B1(new_n889), .B2(new_n890), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(KEYINPUT56), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n912), .A2(new_n913), .ZN(new_n920));
  NAND4_X1  g719(.A1(new_n919), .A2(KEYINPUT122), .A3(new_n920), .A4(new_n910), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n916), .A2(new_n921), .ZN(G1343gat));
  INV_X1    g721(.A(KEYINPUT57), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n874), .A2(new_n923), .A3(new_n252), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n876), .A2(new_n708), .ZN(new_n925));
  INV_X1    g724(.A(new_n860), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n861), .B1(new_n926), .B2(KEYINPUT123), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n927), .B1(KEYINPUT123), .B2(new_n926), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n683), .A2(new_n650), .A3(new_n854), .ZN(new_n929));
  OAI22_X1  g728(.A1(new_n928), .A2(new_n929), .B1(new_n768), .B2(new_n844), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n930), .A2(new_n609), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n548), .B1(new_n931), .B2(new_n868), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n252), .B1(new_n932), .B2(new_n884), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n925), .B1(new_n933), .B2(KEYINPUT57), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n924), .A2(new_n934), .ZN(new_n935));
  OAI21_X1  g734(.A(G141gat), .B1(new_n935), .B2(new_n719), .ZN(new_n936));
  NOR3_X1   g735(.A1(new_n748), .A2(new_n825), .A3(new_n418), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n874), .A2(new_n722), .A3(new_n937), .ZN(new_n938));
  OR3_X1    g737(.A1(new_n938), .A2(G141gat), .A3(new_n719), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n936), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(KEYINPUT58), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT58), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n936), .A2(new_n942), .A3(new_n939), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n941), .A2(new_n943), .ZN(G1344gat));
  XOR2_X1   g743(.A(KEYINPUT124), .B(KEYINPUT59), .Z(new_n945));
  NAND2_X1  g744(.A1(new_n874), .A2(new_n252), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n946), .A2(KEYINPUT57), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n884), .B(KEYINPUT125), .ZN(new_n948));
  NAND4_X1  g747(.A1(new_n867), .A2(new_n650), .A3(new_n854), .A4(new_n862), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n548), .B1(new_n931), .B2(new_n949), .ZN(new_n950));
  OAI211_X1 g749(.A(new_n923), .B(new_n252), .C1(new_n948), .C2(new_n950), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n925), .A2(new_n768), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n947), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n945), .B1(new_n953), .B2(G148gat), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n935), .A2(new_n768), .ZN(new_n955));
  INV_X1    g754(.A(G148gat), .ZN(new_n956));
  OR2_X1    g755(.A1(new_n956), .A2(KEYINPUT59), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n653), .A2(new_n956), .ZN(new_n959));
  OAI22_X1  g758(.A1(new_n954), .A2(new_n958), .B1(new_n938), .B2(new_n959), .ZN(G1345gat));
  OAI21_X1  g759(.A(G155gat), .B1(new_n935), .B2(new_n834), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n548), .A2(new_n213), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n961), .B1(new_n938), .B2(new_n962), .ZN(G1346gat));
  NOR3_X1   g762(.A1(new_n935), .A2(new_n214), .A3(new_n609), .ZN(new_n964));
  OR2_X1    g763(.A1(new_n938), .A2(new_n609), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n964), .B1(new_n214), .B2(new_n965), .ZN(G1347gat));
  NAND2_X1  g765(.A1(new_n418), .A2(new_n445), .ZN(new_n967));
  NOR2_X1   g766(.A1(new_n967), .A2(new_n483), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n907), .A2(new_n968), .ZN(new_n969));
  NOR3_X1   g768(.A1(new_n969), .A2(new_n336), .A3(new_n719), .ZN(new_n970));
  NOR3_X1   g769(.A1(new_n872), .A2(new_n873), .A3(new_n722), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n971), .A2(new_n418), .A3(new_n484), .ZN(new_n972));
  OR2_X1    g771(.A1(new_n972), .A2(new_n719), .ZN(new_n973));
  AOI21_X1  g772(.A(new_n970), .B1(new_n973), .B2(new_n336), .ZN(G1348gat));
  NAND4_X1  g773(.A1(new_n907), .A2(G176gat), .A3(new_n653), .A4(new_n968), .ZN(new_n975));
  INV_X1    g774(.A(KEYINPUT126), .ZN(new_n976));
  OR2_X1    g775(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  OAI21_X1  g776(.A(new_n337), .B1(new_n972), .B2(new_n768), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n975), .A2(new_n976), .ZN(new_n979));
  AND3_X1   g778(.A1(new_n977), .A2(new_n978), .A3(new_n979), .ZN(G1349gat));
  OAI21_X1  g779(.A(new_n373), .B1(new_n969), .B2(new_n834), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n548), .A2(new_n370), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n981), .B1(new_n972), .B2(new_n982), .ZN(new_n983));
  AND2_X1   g782(.A1(KEYINPUT127), .A2(KEYINPUT60), .ZN(new_n984));
  XNOR2_X1  g783(.A(new_n983), .B(new_n984), .ZN(G1350gat));
  OAI21_X1  g784(.A(G190gat), .B1(new_n969), .B2(new_n609), .ZN(new_n986));
  XNOR2_X1  g785(.A(new_n986), .B(KEYINPUT61), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n726), .A2(new_n352), .ZN(new_n988));
  OAI21_X1  g787(.A(new_n987), .B1(new_n972), .B2(new_n988), .ZN(G1351gat));
  NAND3_X1  g788(.A1(new_n708), .A2(new_n252), .A3(new_n418), .ZN(new_n990));
  INV_X1    g789(.A(new_n990), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n971), .A2(new_n991), .ZN(new_n992));
  INV_X1    g791(.A(new_n992), .ZN(new_n993));
  AOI21_X1  g792(.A(G197gat), .B1(new_n993), .B2(new_n683), .ZN(new_n994));
  AND2_X1   g793(.A1(new_n947), .A2(new_n951), .ZN(new_n995));
  NOR2_X1   g794(.A1(new_n748), .A2(new_n967), .ZN(new_n996));
  AND2_X1   g795(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  AND2_X1   g796(.A1(new_n683), .A2(G197gat), .ZN(new_n998));
  AOI21_X1  g797(.A(new_n994), .B1(new_n997), .B2(new_n998), .ZN(G1352gat));
  NAND3_X1  g798(.A1(new_n995), .A2(new_n653), .A3(new_n996), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n1000), .A2(G204gat), .ZN(new_n1001));
  NOR3_X1   g800(.A1(new_n992), .A2(G204gat), .A3(new_n768), .ZN(new_n1002));
  XNOR2_X1  g801(.A(new_n1002), .B(KEYINPUT62), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n1001), .A2(new_n1003), .ZN(G1353gat));
  OR3_X1    g803(.A1(new_n992), .A2(G211gat), .A3(new_n834), .ZN(new_n1005));
  NAND4_X1  g804(.A1(new_n947), .A2(new_n548), .A3(new_n951), .A4(new_n996), .ZN(new_n1006));
  AND3_X1   g805(.A1(new_n1006), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1007));
  AOI21_X1  g806(.A(KEYINPUT63), .B1(new_n1006), .B2(G211gat), .ZN(new_n1008));
  OAI21_X1  g807(.A(new_n1005), .B1(new_n1007), .B2(new_n1008), .ZN(G1354gat));
  NAND3_X1  g808(.A1(new_n995), .A2(new_n726), .A3(new_n996), .ZN(new_n1010));
  NAND2_X1  g809(.A1(new_n1010), .A2(G218gat), .ZN(new_n1011));
  OR3_X1    g810(.A1(new_n992), .A2(G218gat), .A3(new_n609), .ZN(new_n1012));
  NAND2_X1  g811(.A1(new_n1011), .A2(new_n1012), .ZN(G1355gat));
endmodule


