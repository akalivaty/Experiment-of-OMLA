

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737;

  BUF_X1 U371 ( .A(n691), .Z(n703) );
  OR2_X1 U372 ( .A1(n564), .A2(n446), .ZN(n449) );
  XNOR2_X1 U373 ( .A(n459), .B(n723), .ZN(n488) );
  XNOR2_X1 U374 ( .A(n429), .B(n428), .ZN(n366) );
  XNOR2_X1 U375 ( .A(n489), .B(n488), .ZN(n686) );
  XOR2_X1 U376 ( .A(n533), .B(KEYINPUT80), .Z(n349) );
  NOR2_X1 U377 ( .A1(n353), .A2(n354), .ZN(n372) );
  XNOR2_X1 U378 ( .A(n538), .B(KEYINPUT40), .ZN(n736) );
  XNOR2_X1 U379 ( .A(n449), .B(n448), .ZN(n562) );
  XNOR2_X1 U380 ( .A(n551), .B(KEYINPUT19), .ZN(n516) );
  XNOR2_X1 U381 ( .A(n399), .B(n356), .ZN(n510) );
  XNOR2_X1 U382 ( .A(n458), .B(n457), .ZN(n723) );
  XNOR2_X1 U383 ( .A(n385), .B(n384), .ZN(n452) );
  XNOR2_X1 U384 ( .A(n357), .B(G122), .ZN(n433) );
  XNOR2_X1 U385 ( .A(n381), .B(G101), .ZN(n383) );
  INV_X1 U386 ( .A(KEYINPUT88), .ZN(n381) );
  NOR2_X1 U387 ( .A1(G953), .A2(G237), .ZN(n450) );
  NAND2_X1 U388 ( .A1(n523), .A2(n522), .ZN(n351) );
  NAND2_X1 U389 ( .A1(n350), .A2(KEYINPUT71), .ZN(n352) );
  NAND2_X1 U390 ( .A1(n351), .A2(n352), .ZN(n527) );
  INV_X1 U391 ( .A(n523), .ZN(n350) );
  XNOR2_X1 U392 ( .A(n545), .B(KEYINPUT46), .ZN(n353) );
  NAND2_X1 U393 ( .A1(n549), .A2(n349), .ZN(n354) );
  BUF_X1 U394 ( .A(n584), .Z(n355) );
  XNOR2_X1 U395 ( .A(n580), .B(KEYINPUT35), .ZN(n584) );
  XNOR2_X1 U396 ( .A(n575), .B(KEYINPUT33), .ZN(n640) );
  NOR2_X1 U397 ( .A1(n574), .A2(n573), .ZN(n575) );
  NOR2_X1 U398 ( .A1(n640), .A2(n564), .ZN(n576) );
  NOR2_X4 U399 ( .A1(n602), .A2(n601), .ZN(n691) );
  OR2_X1 U400 ( .A1(n562), .A2(n568), .ZN(n586) );
  INV_X1 U401 ( .A(KEYINPUT48), .ZN(n367) );
  NAND2_X1 U402 ( .A1(n372), .A2(n369), .ZN(n368) );
  XNOR2_X1 U403 ( .A(n430), .B(G134), .ZN(n458) );
  NAND2_X1 U404 ( .A1(n595), .A2(n594), .ZN(n362) );
  XNOR2_X1 U405 ( .A(n365), .B(n364), .ZN(n363) );
  INV_X1 U406 ( .A(KEYINPUT84), .ZN(n364) );
  NAND2_X1 U407 ( .A1(n510), .A2(n641), .ZN(n551) );
  INV_X1 U408 ( .A(G107), .ZN(n357) );
  INV_X1 U409 ( .A(G146), .ZN(n459) );
  XNOR2_X1 U410 ( .A(n425), .B(n424), .ZN(n427) );
  XNOR2_X1 U411 ( .A(n442), .B(n441), .ZN(n530) );
  XNOR2_X1 U412 ( .A(n582), .B(n581), .ZN(n583) );
  INV_X1 U413 ( .A(KEYINPUT85), .ZN(n581) );
  XNOR2_X1 U414 ( .A(G125), .B(G146), .ZN(n411) );
  XNOR2_X1 U415 ( .A(n417), .B(n416), .ZN(n419) );
  INV_X1 U416 ( .A(G122), .ZN(n416) );
  INV_X1 U417 ( .A(KEYINPUT45), .ZN(n358) );
  NAND2_X1 U418 ( .A1(n362), .A2(n361), .ZN(n360) );
  OR2_X1 U419 ( .A1(n611), .A2(n596), .ZN(n399) );
  XNOR2_X1 U420 ( .A(G119), .B(G128), .ZN(n463) );
  XNOR2_X1 U421 ( .A(n477), .B(n476), .ZN(n478) );
  INV_X1 U422 ( .A(KEYINPUT64), .ZN(n391) );
  XNOR2_X1 U423 ( .A(n440), .B(n439), .ZN(n699) );
  XNOR2_X1 U424 ( .A(n693), .B(n692), .ZN(n694) );
  OR2_X1 U425 ( .A1(n725), .A2(G952), .ZN(n685) );
  XNOR2_X1 U426 ( .A(n371), .B(n370), .ZN(n734) );
  INV_X1 U427 ( .A(KEYINPUT114), .ZN(n370) );
  NOR2_X2 U428 ( .A1(n505), .A2(n530), .ZN(n629) );
  XNOR2_X1 U429 ( .A(n374), .B(n373), .ZN(n732) );
  INV_X1 U430 ( .A(KEYINPUT111), .ZN(n373) );
  INV_X1 U431 ( .A(n577), .ZN(n531) );
  XNOR2_X1 U432 ( .A(n689), .B(n688), .ZN(n690) );
  XOR2_X1 U433 ( .A(n398), .B(KEYINPUT78), .Z(n356) );
  XNOR2_X2 U434 ( .A(n359), .B(n358), .ZN(n670) );
  NAND2_X1 U435 ( .A1(n363), .A2(n360), .ZN(n359) );
  NAND2_X1 U436 ( .A1(n593), .A2(n592), .ZN(n361) );
  NAND2_X1 U437 ( .A1(n583), .A2(n378), .ZN(n365) );
  NAND2_X1 U438 ( .A1(n366), .A2(G221), .ZN(n470) );
  NAND2_X1 U439 ( .A1(n366), .A2(G217), .ZN(n432) );
  XNOR2_X2 U440 ( .A(n368), .B(n367), .ZN(n599) );
  INV_X1 U441 ( .A(n734), .ZN(n369) );
  NAND2_X1 U442 ( .A1(n555), .A2(n568), .ZN(n371) );
  NAND2_X1 U443 ( .A1(n532), .A2(n732), .ZN(n533) );
  NAND2_X1 U444 ( .A1(n375), .A2(n531), .ZN(n374) );
  XNOR2_X1 U445 ( .A(n528), .B(KEYINPUT110), .ZN(n375) );
  INV_X1 U446 ( .A(n411), .ZN(n410) );
  XNOR2_X2 U447 ( .A(n427), .B(n426), .ZN(n529) );
  AND2_X1 U448 ( .A1(n572), .A2(n571), .ZN(n376) );
  XOR2_X1 U449 ( .A(n509), .B(KEYINPUT43), .Z(n377) );
  NOR2_X1 U450 ( .A1(n617), .A2(n376), .ZN(n378) );
  INV_X1 U451 ( .A(KEYINPUT8), .ZN(n428) );
  INV_X1 U452 ( .A(KEYINPUT82), .ZN(n560) );
  XNOR2_X1 U453 ( .A(n419), .B(n418), .ZN(n421) );
  XNOR2_X1 U454 ( .A(n561), .B(n560), .ZN(n668) );
  XNOR2_X1 U455 ( .A(n432), .B(n431), .ZN(n440) );
  INV_X1 U456 ( .A(KEYINPUT125), .ZN(n704) );
  XNOR2_X1 U457 ( .A(n524), .B(KEYINPUT6), .ZN(n573) );
  XNOR2_X1 U458 ( .A(n686), .B(n687), .ZN(n688) );
  XNOR2_X1 U459 ( .A(n537), .B(KEYINPUT39), .ZN(n556) );
  XNOR2_X1 U460 ( .A(n433), .B(KEYINPUT16), .ZN(n380) );
  XNOR2_X1 U461 ( .A(KEYINPUT87), .B(G110), .ZN(n379) );
  XNOR2_X1 U462 ( .A(n379), .B(G104), .ZN(n482) );
  XNOR2_X1 U463 ( .A(n380), .B(n482), .ZN(n386) );
  XNOR2_X1 U464 ( .A(G116), .B(G113), .ZN(n382) );
  XNOR2_X1 U465 ( .A(n383), .B(n382), .ZN(n385) );
  XNOR2_X1 U466 ( .A(KEYINPUT3), .B(G119), .ZN(n384) );
  XNOR2_X1 U467 ( .A(n386), .B(n452), .ZN(n717) );
  XNOR2_X1 U468 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n387) );
  XNOR2_X1 U469 ( .A(n410), .B(n387), .ZN(n390) );
  XNOR2_X1 U470 ( .A(KEYINPUT90), .B(KEYINPUT4), .ZN(n388) );
  XNOR2_X1 U471 ( .A(n388), .B(KEYINPUT89), .ZN(n389) );
  XNOR2_X1 U472 ( .A(n390), .B(n389), .ZN(n395) );
  XNOR2_X2 U473 ( .A(n391), .B(G953), .ZN(n725) );
  NAND2_X1 U474 ( .A1(n725), .A2(G224), .ZN(n393) );
  INV_X1 U475 ( .A(G143), .ZN(n392) );
  XNOR2_X1 U476 ( .A(n392), .B(G128), .ZN(n430) );
  XNOR2_X1 U477 ( .A(n393), .B(n430), .ZN(n394) );
  XNOR2_X1 U478 ( .A(n395), .B(n394), .ZN(n396) );
  XNOR2_X1 U479 ( .A(n717), .B(n396), .ZN(n611) );
  XNOR2_X1 U480 ( .A(KEYINPUT15), .B(G902), .ZN(n443) );
  INV_X1 U481 ( .A(n443), .ZN(n596) );
  INV_X1 U482 ( .A(G902), .ZN(n461) );
  INV_X1 U483 ( .A(G237), .ZN(n397) );
  NAND2_X1 U484 ( .A1(n461), .A2(n397), .ZN(n400) );
  NAND2_X1 U485 ( .A1(n400), .A2(G210), .ZN(n398) );
  NAND2_X1 U486 ( .A1(n400), .A2(G214), .ZN(n641) );
  NAND2_X1 U487 ( .A1(G234), .A2(G237), .ZN(n401) );
  XNOR2_X1 U488 ( .A(n401), .B(KEYINPUT14), .ZN(n403) );
  NAND2_X1 U489 ( .A1(G952), .A2(n403), .ZN(n402) );
  XOR2_X1 U490 ( .A(KEYINPUT91), .B(n402), .Z(n667) );
  NOR2_X1 U491 ( .A1(G953), .A2(n667), .ZN(n503) );
  INV_X1 U492 ( .A(G953), .ZN(n710) );
  NOR2_X1 U493 ( .A1(G898), .A2(n710), .ZN(n719) );
  AND2_X1 U494 ( .A1(G902), .A2(n403), .ZN(n499) );
  AND2_X1 U495 ( .A1(n719), .A2(n499), .ZN(n404) );
  OR2_X1 U496 ( .A1(n503), .A2(n404), .ZN(n405) );
  XNOR2_X1 U497 ( .A(n405), .B(KEYINPUT92), .ZN(n406) );
  NAND2_X1 U498 ( .A1(n516), .A2(n406), .ZN(n409) );
  INV_X1 U499 ( .A(KEYINPUT65), .ZN(n407) );
  XNOR2_X1 U500 ( .A(n407), .B(KEYINPUT0), .ZN(n408) );
  XNOR2_X1 U501 ( .A(n409), .B(n408), .ZN(n564) );
  XNOR2_X1 U502 ( .A(KEYINPUT13), .B(KEYINPUT101), .ZN(n425) );
  XOR2_X1 U503 ( .A(KEYINPUT10), .B(n411), .Z(n471) );
  INV_X1 U504 ( .A(n471), .ZN(n415) );
  XOR2_X1 U505 ( .A(KEYINPUT100), .B(G104), .Z(n413) );
  XNOR2_X1 U506 ( .A(G113), .B(G131), .ZN(n412) );
  XNOR2_X1 U507 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U508 ( .A(n415), .B(n414), .ZN(n423) );
  NAND2_X1 U509 ( .A1(G214), .A2(n450), .ZN(n417) );
  XOR2_X1 U510 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n418) );
  XNOR2_X1 U511 ( .A(G143), .B(G140), .ZN(n420) );
  XNOR2_X1 U512 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U513 ( .A(n423), .B(n422), .ZN(n693) );
  NOR2_X1 U514 ( .A1(G902), .A2(n693), .ZN(n424) );
  INV_X1 U515 ( .A(G475), .ZN(n426) );
  NAND2_X1 U516 ( .A1(n725), .A2(G234), .ZN(n429) );
  INV_X1 U517 ( .A(n458), .ZN(n431) );
  XNOR2_X1 U518 ( .A(KEYINPUT104), .B(KEYINPUT9), .ZN(n434) );
  XNOR2_X1 U519 ( .A(n434), .B(n433), .ZN(n438) );
  XOR2_X1 U520 ( .A(KEYINPUT103), .B(KEYINPUT102), .Z(n436) );
  XNOR2_X1 U521 ( .A(G116), .B(KEYINPUT7), .ZN(n435) );
  XNOR2_X1 U522 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U523 ( .A(n438), .B(n437), .Z(n439) );
  NOR2_X1 U524 ( .A1(n699), .A2(G902), .ZN(n442) );
  INV_X1 U525 ( .A(G478), .ZN(n441) );
  NOR2_X1 U526 ( .A1(n529), .A2(n530), .ZN(n539) );
  NAND2_X1 U527 ( .A1(G234), .A2(n443), .ZN(n444) );
  XNOR2_X1 U528 ( .A(KEYINPUT20), .B(n444), .ZN(n473) );
  AND2_X1 U529 ( .A1(n473), .A2(G221), .ZN(n445) );
  XNOR2_X1 U530 ( .A(n445), .B(KEYINPUT21), .ZN(n652) );
  NAND2_X1 U531 ( .A1(n539), .A2(n652), .ZN(n446) );
  INV_X1 U532 ( .A(KEYINPUT69), .ZN(n447) );
  XNOR2_X1 U533 ( .A(n447), .B(KEYINPUT22), .ZN(n448) );
  INV_X1 U534 ( .A(n562), .ZN(n495) );
  NAND2_X1 U535 ( .A1(n450), .A2(G210), .ZN(n451) );
  XNOR2_X1 U536 ( .A(n452), .B(n451), .ZN(n456) );
  XOR2_X1 U537 ( .A(KEYINPUT5), .B(KEYINPUT98), .Z(n454) );
  XNOR2_X1 U538 ( .A(G137), .B(KEYINPUT97), .ZN(n453) );
  XNOR2_X1 U539 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U540 ( .A(n456), .B(n455), .ZN(n460) );
  XNOR2_X1 U541 ( .A(G131), .B(KEYINPUT4), .ZN(n457) );
  XNOR2_X1 U542 ( .A(n460), .B(n488), .ZN(n603) );
  NAND2_X1 U543 ( .A1(n603), .A2(n461), .ZN(n462) );
  XNOR2_X2 U544 ( .A(n462), .B(G472), .ZN(n524) );
  XNOR2_X1 U545 ( .A(n573), .B(KEYINPUT77), .ZN(n493) );
  XOR2_X1 U546 ( .A(KEYINPUT68), .B(G110), .Z(n464) );
  XNOR2_X1 U547 ( .A(n464), .B(n463), .ZN(n468) );
  XOR2_X1 U548 ( .A(KEYINPUT23), .B(KEYINPUT94), .Z(n466) );
  XNOR2_X1 U549 ( .A(KEYINPUT24), .B(KEYINPUT95), .ZN(n465) );
  XNOR2_X1 U550 ( .A(n466), .B(n465), .ZN(n467) );
  XOR2_X1 U551 ( .A(n468), .B(n467), .Z(n469) );
  XNOR2_X1 U552 ( .A(n470), .B(n469), .ZN(n472) );
  XOR2_X1 U553 ( .A(G137), .B(G140), .Z(n483) );
  XNOR2_X1 U554 ( .A(n483), .B(n471), .ZN(n722) );
  XNOR2_X1 U555 ( .A(n472), .B(n722), .ZN(n705) );
  NOR2_X1 U556 ( .A1(n705), .A2(G902), .ZN(n479) );
  AND2_X1 U557 ( .A1(G217), .A2(n473), .ZN(n477) );
  XOR2_X1 U558 ( .A(KEYINPUT72), .B(KEYINPUT96), .Z(n475) );
  XNOR2_X1 U559 ( .A(KEYINPUT73), .B(KEYINPUT25), .ZN(n474) );
  XNOR2_X1 U560 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X2 U561 ( .A(n479), .B(n478), .ZN(n588) );
  XNOR2_X1 U562 ( .A(n588), .B(KEYINPUT107), .ZN(n651) );
  XOR2_X1 U563 ( .A(KEYINPUT74), .B(KEYINPUT93), .Z(n481) );
  NAND2_X1 U564 ( .A1(G227), .A2(n725), .ZN(n480) );
  XNOR2_X1 U565 ( .A(n481), .B(n480), .ZN(n487) );
  XNOR2_X1 U566 ( .A(G101), .B(n482), .ZN(n485) );
  XOR2_X1 U567 ( .A(n483), .B(G107), .Z(n484) );
  XNOR2_X1 U568 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U569 ( .A(n487), .B(n486), .ZN(n489) );
  NOR2_X2 U570 ( .A1(G902), .A2(n686), .ZN(n491) );
  XNOR2_X1 U571 ( .A(KEYINPUT67), .B(G469), .ZN(n490) );
  XNOR2_X2 U572 ( .A(n491), .B(n490), .ZN(n520) );
  XNOR2_X2 U573 ( .A(n520), .B(KEYINPUT1), .ZN(n568) );
  INV_X1 U574 ( .A(n568), .ZN(n554) );
  OR2_X1 U575 ( .A1(n651), .A2(n554), .ZN(n492) );
  NOR2_X1 U576 ( .A1(n493), .A2(n492), .ZN(n494) );
  NAND2_X1 U577 ( .A1(n495), .A2(n494), .ZN(n498) );
  INV_X1 U578 ( .A(KEYINPUT76), .ZN(n496) );
  XNOR2_X1 U579 ( .A(n496), .B(KEYINPUT32), .ZN(n497) );
  XNOR2_X1 U580 ( .A(n498), .B(n497), .ZN(n591) );
  XOR2_X1 U581 ( .A(G119), .B(n591), .Z(G21) );
  INV_X1 U582 ( .A(n725), .ZN(n500) );
  NAND2_X1 U583 ( .A1(n500), .A2(n499), .ZN(n501) );
  NOR2_X1 U584 ( .A1(G900), .A2(n501), .ZN(n502) );
  NOR2_X1 U585 ( .A1(n503), .A2(n502), .ZN(n521) );
  NAND2_X1 U586 ( .A1(n588), .A2(n652), .ZN(n504) );
  NOR2_X1 U587 ( .A1(n521), .A2(n504), .ZN(n513) );
  INV_X1 U588 ( .A(n529), .ZN(n505) );
  INV_X1 U589 ( .A(n629), .ZN(n633) );
  NOR2_X1 U590 ( .A1(n573), .A2(n633), .ZN(n506) );
  NAND2_X1 U591 ( .A1(n513), .A2(n506), .ZN(n507) );
  XNOR2_X1 U592 ( .A(KEYINPUT109), .B(n507), .ZN(n550) );
  NAND2_X1 U593 ( .A1(n550), .A2(n641), .ZN(n508) );
  NOR2_X1 U594 ( .A1(n568), .A2(n508), .ZN(n509) );
  INV_X1 U595 ( .A(n510), .ZN(n534) );
  NAND2_X1 U596 ( .A1(n377), .A2(n534), .ZN(n558) );
  XNOR2_X1 U597 ( .A(n558), .B(G140), .ZN(G42) );
  INV_X1 U598 ( .A(n530), .ZN(n511) );
  NOR2_X1 U599 ( .A1(n511), .A2(n529), .ZN(n619) );
  XOR2_X1 U600 ( .A(KEYINPUT105), .B(n619), .Z(n557) );
  OR2_X1 U601 ( .A1(n629), .A2(n557), .ZN(n512) );
  XNOR2_X1 U602 ( .A(KEYINPUT106), .B(n512), .ZN(n571) );
  AND2_X1 U603 ( .A1(n524), .A2(n513), .ZN(n514) );
  XNOR2_X1 U604 ( .A(KEYINPUT28), .B(n514), .ZN(n515) );
  NAND2_X1 U605 ( .A1(n515), .A2(n520), .ZN(n542) );
  INV_X1 U606 ( .A(n516), .ZN(n517) );
  NOR2_X1 U607 ( .A1(n542), .A2(n517), .ZN(n630) );
  NAND2_X1 U608 ( .A1(n571), .A2(n630), .ZN(n518) );
  NAND2_X1 U609 ( .A1(n518), .A2(KEYINPUT47), .ZN(n532) );
  INV_X1 U610 ( .A(n652), .ZN(n519) );
  NOR2_X2 U611 ( .A1(n519), .A2(n588), .ZN(n654) );
  NAND2_X1 U612 ( .A1(n520), .A2(n654), .ZN(n565) );
  NOR2_X2 U613 ( .A1(n565), .A2(n521), .ZN(n523) );
  INV_X1 U614 ( .A(KEYINPUT71), .ZN(n522) );
  NAND2_X1 U615 ( .A1(n524), .A2(n641), .ZN(n525) );
  XOR2_X1 U616 ( .A(KEYINPUT30), .B(n525), .Z(n526) );
  NAND2_X1 U617 ( .A1(n527), .A2(n526), .ZN(n535) );
  NOR2_X1 U618 ( .A1(n535), .A2(n534), .ZN(n528) );
  NAND2_X1 U619 ( .A1(n530), .A2(n529), .ZN(n577) );
  XNOR2_X1 U620 ( .A(n534), .B(KEYINPUT38), .ZN(n642) );
  INV_X1 U621 ( .A(n535), .ZN(n536) );
  NAND2_X1 U622 ( .A1(n642), .A2(n536), .ZN(n537) );
  NAND2_X1 U623 ( .A1(n629), .A2(n556), .ZN(n538) );
  INV_X1 U624 ( .A(n539), .ZN(n644) );
  NAND2_X1 U625 ( .A1(n642), .A2(n641), .ZN(n646) );
  NOR2_X1 U626 ( .A1(n644), .A2(n646), .ZN(n541) );
  XNOR2_X1 U627 ( .A(KEYINPUT41), .B(KEYINPUT112), .ZN(n540) );
  XNOR2_X1 U628 ( .A(n541), .B(n540), .ZN(n679) );
  NOR2_X1 U629 ( .A1(n679), .A2(n542), .ZN(n544) );
  XNOR2_X1 U630 ( .A(KEYINPUT113), .B(KEYINPUT42), .ZN(n543) );
  XNOR2_X1 U631 ( .A(n544), .B(n543), .ZN(n737) );
  NAND2_X1 U632 ( .A1(n736), .A2(n737), .ZN(n545) );
  INV_X1 U633 ( .A(n571), .ZN(n645) );
  XNOR2_X1 U634 ( .A(KEYINPUT47), .B(KEYINPUT66), .ZN(n546) );
  NOR2_X1 U635 ( .A1(n645), .A2(n546), .ZN(n547) );
  XNOR2_X1 U636 ( .A(KEYINPUT70), .B(n547), .ZN(n548) );
  NAND2_X1 U637 ( .A1(n548), .A2(n630), .ZN(n549) );
  INV_X1 U638 ( .A(n550), .ZN(n552) );
  NOR2_X1 U639 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U640 ( .A(n553), .B(KEYINPUT36), .ZN(n555) );
  NAND2_X1 U641 ( .A1(n557), .A2(n556), .ZN(n639) );
  AND2_X1 U642 ( .A1(n558), .A2(n639), .ZN(n598) );
  AND2_X1 U643 ( .A1(KEYINPUT2), .A2(n598), .ZN(n559) );
  NAND2_X1 U644 ( .A1(n599), .A2(n559), .ZN(n561) );
  NAND2_X1 U645 ( .A1(n651), .A2(n573), .ZN(n563) );
  NOR2_X1 U646 ( .A1(n586), .A2(n563), .ZN(n617) );
  INV_X1 U647 ( .A(n564), .ZN(n567) );
  NOR2_X1 U648 ( .A1(n524), .A2(n565), .ZN(n566) );
  NAND2_X1 U649 ( .A1(n567), .A2(n566), .ZN(n620) );
  NAND2_X1 U650 ( .A1(n654), .A2(n568), .ZN(n574) );
  INV_X1 U651 ( .A(n524), .ZN(n587) );
  NOR2_X1 U652 ( .A1(n574), .A2(n587), .ZN(n569) );
  XNOR2_X1 U653 ( .A(n569), .B(KEYINPUT99), .ZN(n659) );
  NOR2_X1 U654 ( .A1(n659), .A2(n564), .ZN(n570) );
  XNOR2_X1 U655 ( .A(n570), .B(KEYINPUT31), .ZN(n636) );
  NAND2_X1 U656 ( .A1(n620), .A2(n636), .ZN(n572) );
  XNOR2_X1 U657 ( .A(n576), .B(KEYINPUT34), .ZN(n579) );
  XNOR2_X1 U658 ( .A(n577), .B(KEYINPUT75), .ZN(n578) );
  NAND2_X1 U659 ( .A1(n579), .A2(n578), .ZN(n580) );
  NAND2_X1 U660 ( .A1(n584), .A2(KEYINPUT44), .ZN(n582) );
  OR2_X1 U661 ( .A1(n355), .A2(KEYINPUT44), .ZN(n592) );
  INV_X1 U662 ( .A(KEYINPUT108), .ZN(n585) );
  XNOR2_X1 U663 ( .A(n586), .B(n585), .ZN(n590) );
  AND2_X1 U664 ( .A1(n588), .A2(n587), .ZN(n589) );
  AND2_X1 U665 ( .A1(n590), .A2(n589), .ZN(n625) );
  NOR2_X2 U666 ( .A1(n625), .A2(n591), .ZN(n593) );
  INV_X1 U667 ( .A(n593), .ZN(n595) );
  INV_X1 U668 ( .A(KEYINPUT44), .ZN(n594) );
  INV_X1 U669 ( .A(n670), .ZN(n711) );
  NAND2_X1 U670 ( .A1(n668), .A2(n711), .ZN(n597) );
  NAND2_X1 U671 ( .A1(n597), .A2(n596), .ZN(n602) );
  NAND2_X1 U672 ( .A1(n599), .A2(n598), .ZN(n671) );
  NOR2_X1 U673 ( .A1(n670), .A2(n671), .ZN(n600) );
  NOR2_X1 U674 ( .A1(n600), .A2(KEYINPUT2), .ZN(n601) );
  NAND2_X1 U675 ( .A1(n691), .A2(G472), .ZN(n606) );
  XNOR2_X1 U676 ( .A(KEYINPUT86), .B(KEYINPUT62), .ZN(n604) );
  XNOR2_X1 U677 ( .A(n603), .B(n604), .ZN(n605) );
  XNOR2_X1 U678 ( .A(n606), .B(n605), .ZN(n607) );
  NAND2_X1 U679 ( .A1(n607), .A2(n685), .ZN(n608) );
  XNOR2_X1 U680 ( .A(n608), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U681 ( .A1(n691), .A2(G210), .ZN(n613) );
  XOR2_X1 U682 ( .A(KEYINPUT79), .B(KEYINPUT54), .Z(n609) );
  XNOR2_X1 U683 ( .A(n609), .B(KEYINPUT55), .ZN(n610) );
  XNOR2_X1 U684 ( .A(n611), .B(n610), .ZN(n612) );
  XNOR2_X1 U685 ( .A(n613), .B(n612), .ZN(n614) );
  NAND2_X1 U686 ( .A1(n614), .A2(n685), .ZN(n616) );
  XNOR2_X1 U687 ( .A(KEYINPUT83), .B(KEYINPUT56), .ZN(n615) );
  XNOR2_X1 U688 ( .A(n616), .B(n615), .ZN(G51) );
  XOR2_X1 U689 ( .A(G101), .B(n617), .Z(G3) );
  NOR2_X1 U690 ( .A1(n633), .A2(n620), .ZN(n618) );
  XOR2_X1 U691 ( .A(G104), .B(n618), .Z(G6) );
  INV_X1 U692 ( .A(n619), .ZN(n637) );
  NOR2_X1 U693 ( .A1(n620), .A2(n637), .ZN(n624) );
  XOR2_X1 U694 ( .A(KEYINPUT26), .B(KEYINPUT115), .Z(n622) );
  XNOR2_X1 U695 ( .A(G107), .B(KEYINPUT27), .ZN(n621) );
  XNOR2_X1 U696 ( .A(n622), .B(n621), .ZN(n623) );
  XNOR2_X1 U697 ( .A(n624), .B(n623), .ZN(G9) );
  XOR2_X1 U698 ( .A(G110), .B(n625), .Z(n626) );
  XNOR2_X1 U699 ( .A(KEYINPUT116), .B(n626), .ZN(G12) );
  XOR2_X1 U700 ( .A(G128), .B(KEYINPUT29), .Z(n628) );
  NAND2_X1 U701 ( .A1(n630), .A2(n619), .ZN(n627) );
  XNOR2_X1 U702 ( .A(n628), .B(n627), .ZN(G30) );
  XOR2_X1 U703 ( .A(G146), .B(KEYINPUT117), .Z(n632) );
  NAND2_X1 U704 ( .A1(n630), .A2(n629), .ZN(n631) );
  XNOR2_X1 U705 ( .A(n632), .B(n631), .ZN(G48) );
  NOR2_X1 U706 ( .A1(n633), .A2(n636), .ZN(n634) );
  XOR2_X1 U707 ( .A(KEYINPUT118), .B(n634), .Z(n635) );
  XNOR2_X1 U708 ( .A(G113), .B(n635), .ZN(G15) );
  NOR2_X1 U709 ( .A1(n637), .A2(n636), .ZN(n638) );
  XOR2_X1 U710 ( .A(G116), .B(n638), .Z(G18) );
  XNOR2_X1 U711 ( .A(G134), .B(n639), .ZN(G36) );
  NOR2_X1 U712 ( .A1(n642), .A2(n641), .ZN(n643) );
  NOR2_X1 U713 ( .A1(n644), .A2(n643), .ZN(n648) );
  NOR2_X1 U714 ( .A1(n646), .A2(n645), .ZN(n647) );
  NOR2_X1 U715 ( .A1(n648), .A2(n647), .ZN(n649) );
  XNOR2_X1 U716 ( .A(n649), .B(KEYINPUT120), .ZN(n650) );
  NOR2_X1 U717 ( .A1(n640), .A2(n650), .ZN(n664) );
  NOR2_X1 U718 ( .A1(n652), .A2(n651), .ZN(n653) );
  XNOR2_X1 U719 ( .A(n653), .B(KEYINPUT49), .ZN(n658) );
  OR2_X1 U720 ( .A1(n568), .A2(n654), .ZN(n655) );
  XOR2_X1 U721 ( .A(KEYINPUT50), .B(n655), .Z(n656) );
  NOR2_X1 U722 ( .A1(n524), .A2(n656), .ZN(n657) );
  NAND2_X1 U723 ( .A1(n658), .A2(n657), .ZN(n660) );
  NAND2_X1 U724 ( .A1(n660), .A2(n659), .ZN(n661) );
  XNOR2_X1 U725 ( .A(KEYINPUT51), .B(n661), .ZN(n662) );
  NOR2_X1 U726 ( .A1(n679), .A2(n662), .ZN(n663) );
  NOR2_X1 U727 ( .A1(n664), .A2(n663), .ZN(n665) );
  XNOR2_X1 U728 ( .A(n665), .B(KEYINPUT52), .ZN(n666) );
  NOR2_X1 U729 ( .A1(n667), .A2(n666), .ZN(n678) );
  AND2_X1 U730 ( .A1(n668), .A2(n711), .ZN(n676) );
  INV_X1 U731 ( .A(KEYINPUT2), .ZN(n669) );
  NAND2_X1 U732 ( .A1(n670), .A2(n669), .ZN(n674) );
  INV_X1 U733 ( .A(n671), .ZN(n724) );
  NOR2_X1 U734 ( .A1(n724), .A2(KEYINPUT2), .ZN(n672) );
  XNOR2_X1 U735 ( .A(n672), .B(KEYINPUT81), .ZN(n673) );
  NAND2_X1 U736 ( .A1(n674), .A2(n673), .ZN(n675) );
  NOR2_X1 U737 ( .A1(n676), .A2(n675), .ZN(n677) );
  NOR2_X1 U738 ( .A1(n678), .A2(n677), .ZN(n682) );
  NOR2_X1 U739 ( .A1(n679), .A2(n640), .ZN(n680) );
  XNOR2_X1 U740 ( .A(n680), .B(KEYINPUT121), .ZN(n681) );
  NAND2_X1 U741 ( .A1(n682), .A2(n681), .ZN(n683) );
  NOR2_X1 U742 ( .A1(n683), .A2(G953), .ZN(n684) );
  XNOR2_X1 U743 ( .A(n684), .B(KEYINPUT53), .ZN(G75) );
  INV_X1 U744 ( .A(n685), .ZN(n709) );
  NAND2_X1 U745 ( .A1(n703), .A2(G469), .ZN(n689) );
  XOR2_X1 U746 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n687) );
  NOR2_X1 U747 ( .A1(n709), .A2(n690), .ZN(G54) );
  NAND2_X1 U748 ( .A1(n691), .A2(G475), .ZN(n695) );
  XOR2_X1 U749 ( .A(KEYINPUT122), .B(KEYINPUT59), .Z(n692) );
  XNOR2_X1 U750 ( .A(n695), .B(n694), .ZN(n696) );
  NOR2_X2 U751 ( .A1(n696), .A2(n709), .ZN(n698) );
  XOR2_X1 U752 ( .A(KEYINPUT123), .B(KEYINPUT60), .Z(n697) );
  XNOR2_X1 U753 ( .A(n698), .B(n697), .ZN(G60) );
  NAND2_X1 U754 ( .A1(n703), .A2(G478), .ZN(n701) );
  XNOR2_X1 U755 ( .A(n699), .B(KEYINPUT124), .ZN(n700) );
  XNOR2_X1 U756 ( .A(n701), .B(n700), .ZN(n702) );
  NOR2_X1 U757 ( .A1(n709), .A2(n702), .ZN(G63) );
  NAND2_X1 U758 ( .A1(n703), .A2(G217), .ZN(n707) );
  XNOR2_X1 U759 ( .A(n705), .B(n704), .ZN(n706) );
  XNOR2_X1 U760 ( .A(n707), .B(n706), .ZN(n708) );
  NOR2_X1 U761 ( .A1(n709), .A2(n708), .ZN(G66) );
  NAND2_X1 U762 ( .A1(n711), .A2(n710), .ZN(n715) );
  NAND2_X1 U763 ( .A1(G953), .A2(G224), .ZN(n712) );
  XNOR2_X1 U764 ( .A(KEYINPUT61), .B(n712), .ZN(n713) );
  NAND2_X1 U765 ( .A1(n713), .A2(G898), .ZN(n714) );
  NAND2_X1 U766 ( .A1(n715), .A2(n714), .ZN(n721) );
  XNOR2_X1 U767 ( .A(KEYINPUT126), .B(KEYINPUT127), .ZN(n716) );
  XNOR2_X1 U768 ( .A(n717), .B(n716), .ZN(n718) );
  NOR2_X1 U769 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U770 ( .A(n721), .B(n720), .ZN(G69) );
  XNOR2_X1 U771 ( .A(n723), .B(n722), .ZN(n727) );
  XOR2_X1 U772 ( .A(n727), .B(n724), .Z(n726) );
  NAND2_X1 U773 ( .A1(n726), .A2(n725), .ZN(n731) );
  XNOR2_X1 U774 ( .A(G227), .B(n727), .ZN(n728) );
  NAND2_X1 U775 ( .A1(n728), .A2(G900), .ZN(n729) );
  NAND2_X1 U776 ( .A1(n729), .A2(G953), .ZN(n730) );
  NAND2_X1 U777 ( .A1(n731), .A2(n730), .ZN(G72) );
  XOR2_X1 U778 ( .A(n355), .B(G122), .Z(G24) );
  XNOR2_X1 U779 ( .A(G143), .B(n732), .ZN(G45) );
  XOR2_X1 U780 ( .A(KEYINPUT37), .B(KEYINPUT119), .Z(n733) );
  XNOR2_X1 U781 ( .A(n734), .B(n733), .ZN(n735) );
  XNOR2_X1 U782 ( .A(G125), .B(n735), .ZN(G27) );
  XNOR2_X1 U783 ( .A(G131), .B(n736), .ZN(G33) );
  XNOR2_X1 U784 ( .A(G137), .B(n737), .ZN(G39) );
endmodule

