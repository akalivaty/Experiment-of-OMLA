//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 0 1 1 1 1 0 1 0 0 1 0 0 0 1 0 0 0 0 1 1 1 1 1 1 1 1 1 0 1 0 0 1 0 1 1 0 1 0 0 1 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:28 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n698, new_n699,
    new_n700, new_n701, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984;
  NAND2_X1  g000(.A1(G234), .A2(G237), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n187), .A2(G952), .A3(new_n188), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n189), .B(KEYINPUT91), .ZN(new_n190));
  XOR2_X1   g004(.A(KEYINPUT21), .B(G898), .Z(new_n191));
  AND3_X1   g005(.A1(new_n187), .A2(G902), .A3(G953), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n190), .B1(new_n191), .B2(new_n193), .ZN(new_n194));
  OAI21_X1  g008(.A(G214), .B1(G237), .B2(G902), .ZN(new_n195));
  INV_X1    g009(.A(G902), .ZN(new_n196));
  INV_X1    g010(.A(G119), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G116), .ZN(new_n198));
  INV_X1    g012(.A(G116), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G119), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n198), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G113), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(KEYINPUT2), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT2), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G113), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n201), .A2(new_n203), .A3(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n203), .A2(new_n205), .ZN(new_n207));
  XNOR2_X1  g021(.A(G116), .B(G119), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  AND3_X1   g023(.A1(new_n206), .A2(new_n209), .A3(KEYINPUT66), .ZN(new_n210));
  AOI21_X1  g024(.A(KEYINPUT66), .B1(new_n206), .B2(new_n209), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G104), .ZN(new_n213));
  OAI21_X1  g027(.A(KEYINPUT3), .B1(new_n213), .B2(G107), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(KEYINPUT80), .ZN(new_n215));
  OR3_X1    g029(.A1(new_n213), .A2(KEYINPUT3), .A3(G107), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT80), .ZN(new_n217));
  OAI211_X1 g031(.A(new_n217), .B(KEYINPUT3), .C1(new_n213), .C2(G107), .ZN(new_n218));
  INV_X1    g032(.A(G107), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n219), .A2(G104), .ZN(new_n220));
  INV_X1    g034(.A(new_n220), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n215), .A2(new_n216), .A3(new_n218), .A4(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G101), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n220), .B1(new_n214), .B2(KEYINPUT80), .ZN(new_n224));
  INV_X1    g038(.A(G101), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n224), .A2(new_n225), .A3(new_n216), .A4(new_n218), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n223), .A2(KEYINPUT4), .A3(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT4), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n222), .A2(new_n228), .A3(G101), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n212), .A2(new_n227), .A3(new_n229), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n213), .A2(G107), .ZN(new_n231));
  OAI21_X1  g045(.A(G101), .B1(new_n231), .B2(new_n220), .ZN(new_n232));
  AND2_X1   g046(.A1(new_n226), .A2(new_n232), .ZN(new_n233));
  XNOR2_X1  g047(.A(KEYINPUT83), .B(KEYINPUT5), .ZN(new_n234));
  OR2_X1    g048(.A1(new_n201), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(new_n198), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n202), .B1(new_n234), .B2(new_n236), .ZN(new_n237));
  AOI22_X1  g051(.A1(new_n235), .A2(new_n237), .B1(new_n208), .B2(new_n207), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n233), .A2(new_n238), .ZN(new_n239));
  AND2_X1   g053(.A1(new_n230), .A2(new_n239), .ZN(new_n240));
  XNOR2_X1  g054(.A(G110), .B(G122), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  AND2_X1   g056(.A1(KEYINPUT64), .A2(G146), .ZN(new_n243));
  NOR2_X1   g057(.A1(KEYINPUT64), .A2(G146), .ZN(new_n244));
  OAI21_X1  g058(.A(G143), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(G146), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n246), .A2(G143), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(G128), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n249), .A2(KEYINPUT1), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n245), .A2(new_n248), .A3(new_n250), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n249), .B1(new_n245), .B2(KEYINPUT1), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n246), .A2(G143), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n243), .A2(new_n244), .ZN(new_n255));
  INV_X1    g069(.A(G143), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n254), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n251), .B1(new_n252), .B2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(G125), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  XNOR2_X1  g074(.A(KEYINPUT64), .B(G146), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n253), .B1(new_n261), .B2(G143), .ZN(new_n262));
  NAND2_X1  g076(.A1(KEYINPUT0), .A2(G128), .ZN(new_n263));
  OR2_X1    g077(.A1(KEYINPUT0), .A2(G128), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n262), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  NAND4_X1  g079(.A1(new_n245), .A2(KEYINPUT0), .A3(G128), .A4(new_n248), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n265), .A2(G125), .A3(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n188), .A2(G224), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(KEYINPUT7), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n260), .A2(new_n267), .A3(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(new_n233), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(new_n238), .ZN(new_n272));
  XNOR2_X1  g086(.A(new_n241), .B(KEYINPUT8), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n208), .A2(KEYINPUT5), .ZN(new_n274));
  AOI22_X1  g088(.A1(new_n237), .A2(new_n274), .B1(new_n208), .B2(new_n207), .ZN(new_n275));
  OAI211_X1 g089(.A(new_n272), .B(new_n273), .C1(new_n275), .C2(new_n271), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n260), .A2(new_n267), .ZN(new_n277));
  XOR2_X1   g091(.A(new_n268), .B(KEYINPUT86), .Z(new_n278));
  NAND3_X1  g092(.A1(new_n277), .A2(KEYINPUT7), .A3(new_n278), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n242), .A2(new_n270), .A3(new_n276), .A4(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n230), .A2(new_n239), .ZN(new_n281));
  XOR2_X1   g095(.A(new_n241), .B(KEYINPUT84), .Z(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT85), .ZN(new_n284));
  AOI22_X1  g098(.A1(new_n281), .A2(new_n283), .B1(new_n284), .B2(KEYINPUT6), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(KEYINPUT6), .ZN(new_n286));
  AOI211_X1 g100(.A(new_n286), .B(new_n282), .C1(new_n230), .C2(new_n239), .ZN(new_n287));
  AND4_X1   g101(.A1(KEYINPUT6), .A2(new_n230), .A3(new_n241), .A4(new_n239), .ZN(new_n288));
  NOR3_X1   g102(.A1(new_n285), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  XOR2_X1   g103(.A(new_n277), .B(new_n268), .Z(new_n290));
  OAI211_X1 g104(.A(new_n196), .B(new_n280), .C1(new_n289), .C2(new_n290), .ZN(new_n291));
  OAI21_X1  g105(.A(G210), .B1(G237), .B2(G902), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n281), .A2(new_n283), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(new_n286), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n240), .A2(KEYINPUT6), .A3(new_n241), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n281), .A2(new_n284), .A3(KEYINPUT6), .A4(new_n283), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n296), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(new_n290), .ZN(new_n300));
  AOI21_X1  g114(.A(G902), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n292), .B1(new_n301), .B2(new_n280), .ZN(new_n302));
  OAI211_X1 g116(.A(new_n194), .B(new_n195), .C1(new_n294), .C2(new_n302), .ZN(new_n303));
  XOR2_X1   g117(.A(KEYINPUT9), .B(G234), .Z(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(new_n196), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(G221), .ZN(new_n306));
  XOR2_X1   g120(.A(new_n306), .B(KEYINPUT79), .Z(new_n307));
  INV_X1    g121(.A(G469), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT82), .ZN(new_n309));
  XNOR2_X1  g123(.A(G110), .B(G140), .ZN(new_n310));
  INV_X1    g124(.A(G227), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n311), .A2(G953), .ZN(new_n312));
  XOR2_X1   g126(.A(new_n310), .B(new_n312), .Z(new_n313));
  AOI21_X1  g127(.A(new_n249), .B1(new_n253), .B2(KEYINPUT1), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n314), .B1(new_n245), .B2(new_n248), .ZN(new_n315));
  AND3_X1   g129(.A1(new_n245), .A2(new_n248), .A3(new_n250), .ZN(new_n316));
  OAI211_X1 g130(.A(new_n226), .B(new_n232), .C1(new_n315), .C2(new_n316), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n317), .B1(new_n233), .B2(new_n258), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT11), .ZN(new_n319));
  INV_X1    g133(.A(G134), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n319), .B1(new_n320), .B2(G137), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(G137), .ZN(new_n322));
  INV_X1    g136(.A(G137), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n323), .A2(KEYINPUT11), .A3(G134), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n321), .A2(new_n322), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(G131), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT65), .ZN(new_n327));
  INV_X1    g141(.A(G131), .ZN(new_n328));
  NAND4_X1  g142(.A1(new_n321), .A2(new_n324), .A3(new_n328), .A4(new_n322), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n326), .A2(new_n327), .A3(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n325), .A2(KEYINPUT65), .A3(G131), .ZN(new_n331));
  AND2_X1   g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n318), .A2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT12), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n318), .A2(KEYINPUT12), .A3(new_n332), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT81), .ZN(new_n338));
  AND3_X1   g152(.A1(new_n330), .A2(new_n338), .A3(new_n331), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n338), .B1(new_n330), .B2(new_n331), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT10), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n317), .A2(new_n342), .ZN(new_n343));
  NAND4_X1  g157(.A1(new_n227), .A2(new_n266), .A3(new_n265), .A4(new_n229), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n233), .A2(KEYINPUT10), .A3(new_n258), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n341), .A2(new_n343), .A3(new_n344), .A4(new_n345), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n313), .B1(new_n337), .B2(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n344), .A2(new_n343), .A3(new_n345), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(new_n332), .ZN(new_n349));
  AND3_X1   g163(.A1(new_n349), .A2(new_n346), .A3(new_n313), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n309), .B1(new_n347), .B2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(new_n313), .ZN(new_n352));
  AND3_X1   g166(.A1(new_n318), .A2(KEYINPUT12), .A3(new_n332), .ZN(new_n353));
  AOI21_X1  g167(.A(KEYINPUT12), .B1(new_n318), .B2(new_n332), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(new_n346), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n352), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n349), .A2(new_n346), .A3(new_n313), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n357), .A2(KEYINPUT82), .A3(new_n358), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n308), .B1(new_n351), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n346), .A2(new_n313), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n355), .A2(new_n361), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n313), .B1(new_n349), .B2(new_n346), .ZN(new_n363));
  OAI211_X1 g177(.A(new_n308), .B(new_n196), .C1(new_n362), .C2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(G469), .A2(G902), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n307), .B1(new_n360), .B2(new_n366), .ZN(new_n367));
  XNOR2_X1  g181(.A(G113), .B(G122), .ZN(new_n368));
  XNOR2_X1  g182(.A(KEYINPUT87), .B(G104), .ZN(new_n369));
  XOR2_X1   g183(.A(new_n368), .B(new_n369), .Z(new_n370));
  NOR3_X1   g184(.A1(new_n259), .A2(KEYINPUT16), .A3(G140), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  XOR2_X1   g186(.A(G125), .B(G140), .Z(new_n373));
  INV_X1    g187(.A(KEYINPUT16), .ZN(new_n374));
  OAI211_X1 g188(.A(G146), .B(new_n372), .C1(new_n373), .C2(new_n374), .ZN(new_n375));
  NOR2_X1   g189(.A1(G237), .A2(G953), .ZN(new_n376));
  AND3_X1   g190(.A1(new_n376), .A2(G143), .A3(G214), .ZN(new_n377));
  AOI21_X1  g191(.A(G143), .B1(new_n376), .B2(G214), .ZN(new_n378));
  OAI211_X1 g192(.A(KEYINPUT17), .B(G131), .C1(new_n377), .C2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(G140), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n259), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(G125), .A2(G140), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n374), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n246), .B1(new_n383), .B2(new_n371), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n375), .A2(new_n379), .A3(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(KEYINPUT88), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n377), .A2(new_n378), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(new_n328), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT17), .ZN(new_n389));
  OAI21_X1  g203(.A(G131), .B1(new_n377), .B2(new_n378), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n388), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT88), .ZN(new_n392));
  NAND4_X1  g206(.A1(new_n375), .A2(new_n379), .A3(new_n384), .A4(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n386), .A2(new_n391), .A3(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(new_n373), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(new_n261), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n396), .B1(new_n246), .B2(new_n395), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT18), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n387), .B1(new_n398), .B2(new_n328), .ZN(new_n399));
  OAI211_X1 g213(.A(new_n397), .B(new_n399), .C1(new_n398), .C2(new_n390), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n370), .B1(new_n394), .B2(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n394), .A2(new_n400), .A3(new_n370), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(KEYINPUT89), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT89), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n394), .A2(new_n404), .A3(new_n400), .A4(new_n370), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n401), .B1(new_n403), .B2(new_n405), .ZN(new_n406));
  OAI21_X1  g220(.A(G475), .B1(new_n406), .B2(G902), .ZN(new_n407));
  INV_X1    g221(.A(G122), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(G116), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n199), .A2(G122), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(G107), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n409), .A2(new_n410), .A3(new_n219), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n256), .A2(G128), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n249), .A2(G143), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n415), .A2(new_n416), .A3(KEYINPUT13), .ZN(new_n417));
  OAI211_X1 g231(.A(new_n417), .B(G134), .C1(KEYINPUT13), .C2(new_n415), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n415), .A2(new_n416), .A3(new_n320), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n414), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n415), .A2(new_n416), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(G134), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(new_n419), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n199), .A2(KEYINPUT14), .A3(G122), .ZN(new_n424));
  OAI211_X1 g238(.A(G107), .B(new_n424), .C1(new_n411), .C2(KEYINPUT14), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n423), .A2(new_n425), .A3(new_n413), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n420), .A2(new_n426), .ZN(new_n427));
  XOR2_X1   g241(.A(KEYINPUT69), .B(G217), .Z(new_n428));
  NAND3_X1  g242(.A1(new_n428), .A2(new_n304), .A3(new_n188), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n429), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n420), .A2(new_n426), .A3(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n430), .A2(KEYINPUT90), .A3(new_n432), .ZN(new_n433));
  OR3_X1    g247(.A1(new_n427), .A2(KEYINPUT90), .A3(new_n429), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n433), .A2(new_n434), .A3(new_n196), .ZN(new_n435));
  INV_X1    g249(.A(G478), .ZN(new_n436));
  OR2_X1    g250(.A1(new_n436), .A2(KEYINPUT15), .ZN(new_n437));
  XNOR2_X1  g251(.A(new_n435), .B(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT20), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n403), .A2(new_n405), .ZN(new_n440));
  XOR2_X1   g254(.A(new_n373), .B(KEYINPUT19), .Z(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(new_n261), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(new_n375), .ZN(new_n443));
  AND2_X1   g257(.A1(new_n388), .A2(new_n390), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n400), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n370), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  AOI21_X1  g261(.A(G475), .B1(new_n440), .B2(new_n447), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n439), .B1(new_n448), .B2(new_n196), .ZN(new_n449));
  AOI22_X1  g263(.A1(new_n403), .A2(new_n405), .B1(new_n446), .B2(new_n445), .ZN(new_n450));
  NOR4_X1   g264(.A1(new_n450), .A2(KEYINPUT20), .A3(G475), .A4(G902), .ZN(new_n451));
  OAI211_X1 g265(.A(new_n407), .B(new_n438), .C1(new_n449), .C2(new_n451), .ZN(new_n452));
  NOR3_X1   g266(.A1(new_n303), .A2(new_n367), .A3(new_n452), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n330), .A2(new_n265), .A3(new_n266), .A4(new_n331), .ZN(new_n454));
  INV_X1    g268(.A(new_n322), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n320), .A2(G137), .ZN(new_n456));
  OAI21_X1  g270(.A(G131), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  AND2_X1   g271(.A1(new_n457), .A2(new_n329), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n258), .A2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT30), .ZN(new_n460));
  AND3_X1   g274(.A1(new_n454), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n460), .B1(new_n454), .B2(new_n459), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n212), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n206), .A2(new_n209), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT66), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n206), .A2(new_n209), .A3(KEYINPUT66), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n454), .A2(new_n459), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n376), .A2(G210), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n470), .B(G101), .ZN(new_n471));
  XNOR2_X1  g285(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n471), .B(new_n472), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n463), .A2(KEYINPUT31), .A3(new_n469), .A4(new_n473), .ZN(new_n474));
  AND2_X1   g288(.A1(new_n474), .A2(new_n196), .ZN(new_n475));
  INV_X1    g289(.A(new_n473), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT28), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n454), .A2(new_n459), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(new_n212), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n477), .B1(new_n479), .B2(new_n469), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n469), .A2(new_n477), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n476), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT31), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n463), .A2(new_n469), .A3(new_n473), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(G472), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n475), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT32), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n475), .A2(new_n486), .A3(KEYINPUT32), .A4(new_n487), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n490), .A2(KEYINPUT67), .A3(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT67), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n488), .A2(new_n493), .A3(new_n489), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  AND3_X1   g309(.A1(new_n454), .A2(new_n459), .A3(new_n468), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n468), .B1(new_n454), .B2(new_n459), .ZN(new_n497));
  OAI21_X1  g311(.A(KEYINPUT28), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n498), .A2(KEYINPUT29), .A3(new_n481), .A4(new_n473), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n498), .A2(new_n481), .A3(new_n473), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT29), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n473), .B1(new_n463), .B2(new_n469), .ZN(new_n503));
  OAI211_X1 g317(.A(new_n196), .B(new_n499), .C1(new_n502), .C2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(G472), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT68), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n504), .A2(KEYINPUT68), .A3(G472), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n495), .A2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT25), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(KEYINPUT77), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n249), .A2(KEYINPUT23), .A3(G119), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n513), .B(KEYINPUT70), .ZN(new_n514));
  OAI21_X1  g328(.A(KEYINPUT23), .B1(new_n249), .B2(G119), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT71), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n249), .A2(G119), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n197), .A2(G128), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n519), .A2(KEYINPUT71), .A3(KEYINPUT23), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n517), .A2(new_n518), .A3(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(G110), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n514), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(KEYINPUT73), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT73), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n514), .A2(new_n521), .A3(new_n525), .A4(new_n522), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n518), .A2(new_n519), .ZN(new_n528));
  XNOR2_X1  g342(.A(KEYINPUT24), .B(G110), .ZN(new_n529));
  AND3_X1   g343(.A1(new_n528), .A2(new_n529), .A3(KEYINPUT74), .ZN(new_n530));
  AOI21_X1  g344(.A(KEYINPUT74), .B1(new_n528), .B2(new_n529), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(KEYINPUT75), .B1(new_n527), .B2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT75), .ZN(new_n535));
  AOI211_X1 g349(.A(new_n535), .B(new_n532), .C1(new_n524), .C2(new_n526), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n396), .A2(new_n375), .ZN(new_n537));
  NOR3_X1   g351(.A1(new_n534), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n514), .A2(new_n521), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(G110), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n375), .A2(new_n384), .ZN(new_n541));
  OAI211_X1 g355(.A(new_n540), .B(new_n541), .C1(new_n528), .C2(new_n529), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT72), .ZN(new_n543));
  XNOR2_X1  g357(.A(new_n542), .B(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n545), .B(G137), .ZN(new_n546));
  XNOR2_X1  g360(.A(KEYINPUT76), .B(KEYINPUT22), .ZN(new_n547));
  XNOR2_X1  g361(.A(new_n546), .B(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  NOR3_X1   g363(.A1(new_n538), .A2(new_n544), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n527), .A2(new_n533), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(new_n535), .ZN(new_n552));
  INV_X1    g366(.A(new_n537), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n527), .A2(KEYINPUT75), .A3(new_n533), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n542), .B(KEYINPUT72), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n548), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  OAI211_X1 g371(.A(new_n196), .B(new_n512), .C1(new_n550), .C2(new_n557), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n511), .A2(KEYINPUT77), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(new_n428), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n561), .B1(G234), .B2(new_n196), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n549), .B1(new_n538), .B2(new_n544), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n555), .A2(new_n556), .A3(new_n548), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n559), .ZN(new_n566));
  NAND4_X1  g380(.A1(new_n565), .A2(new_n196), .A3(new_n566), .A4(new_n512), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n560), .A2(new_n562), .A3(new_n567), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n562), .A2(G902), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n565), .A2(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(KEYINPUT78), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n568), .A2(KEYINPUT78), .A3(new_n570), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  OAI211_X1 g387(.A(new_n453), .B(new_n510), .C1(new_n571), .C2(new_n573), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n574), .B(G101), .ZN(G3));
  OAI21_X1  g389(.A(new_n407), .B1(new_n449), .B2(new_n451), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT33), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n433), .A2(new_n434), .A3(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n430), .A2(KEYINPUT33), .A3(new_n432), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n578), .A2(new_n196), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(G478), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT92), .ZN(new_n582));
  OR2_X1    g396(.A1(new_n435), .A2(G478), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n582), .B1(new_n581), .B2(new_n583), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n576), .A2(new_n587), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n303), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n475), .A2(new_n486), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(G472), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(new_n488), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n367), .A2(new_n592), .ZN(new_n593));
  OAI211_X1 g407(.A(new_n589), .B(new_n593), .C1(new_n573), .C2(new_n571), .ZN(new_n594));
  XOR2_X1   g408(.A(KEYINPUT34), .B(G104), .Z(new_n595));
  XNOR2_X1  g409(.A(new_n594), .B(new_n595), .ZN(G6));
  INV_X1    g410(.A(new_n367), .ZN(new_n597));
  INV_X1    g411(.A(new_n592), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n568), .A2(new_n570), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT78), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n599), .B1(new_n602), .B2(new_n572), .ZN(new_n603));
  INV_X1    g417(.A(new_n438), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n407), .B(KEYINPUT94), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n440), .A2(new_n447), .ZN(new_n606));
  INV_X1    g420(.A(G475), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n606), .A2(new_n607), .A3(new_n196), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(KEYINPUT20), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n448), .A2(new_n439), .A3(new_n196), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  AND2_X1   g425(.A1(new_n611), .A2(KEYINPUT93), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n611), .A2(KEYINPUT93), .ZN(new_n613));
  OAI211_X1 g427(.A(new_n604), .B(new_n605), .C1(new_n612), .C2(new_n613), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n614), .A2(new_n303), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n603), .A2(new_n615), .ZN(new_n616));
  XOR2_X1   g430(.A(KEYINPUT35), .B(G107), .Z(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(G9));
  NAND2_X1  g432(.A1(new_n555), .A2(new_n556), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n548), .A2(KEYINPUT36), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n619), .B(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(new_n569), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n568), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(new_n598), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT95), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n623), .A2(KEYINPUT95), .A3(new_n598), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(new_n453), .ZN(new_n629));
  XOR2_X1   g443(.A(KEYINPUT37), .B(G110), .Z(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(G12));
  AOI22_X1  g445(.A1(new_n492), .A2(new_n494), .B1(new_n507), .B2(new_n508), .ZN(new_n632));
  AND2_X1   g446(.A1(new_n568), .A2(new_n622), .ZN(new_n633));
  INV_X1    g447(.A(new_n195), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n291), .A2(new_n293), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n301), .A2(new_n292), .A3(new_n280), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n634), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  NOR4_X1   g452(.A1(new_n632), .A2(new_n633), .A3(new_n367), .A4(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n190), .ZN(new_n640));
  INV_X1    g454(.A(G900), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n640), .B1(new_n641), .B2(new_n192), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n614), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n639), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(G128), .ZN(G30));
  XOR2_X1   g459(.A(new_n642), .B(KEYINPUT39), .Z(new_n646));
  NAND2_X1  g460(.A1(new_n597), .A2(new_n646), .ZN(new_n647));
  XOR2_X1   g461(.A(new_n647), .B(KEYINPUT40), .Z(new_n648));
  NAND2_X1  g462(.A1(new_n635), .A2(new_n636), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT38), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n576), .A2(new_n604), .A3(new_n195), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n463), .A2(new_n469), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n655), .A2(new_n476), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n496), .A2(new_n497), .ZN(new_n657));
  AOI21_X1  g471(.A(G902), .B1(new_n657), .B2(new_n476), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  OAI21_X1  g473(.A(G472), .B1(new_n656), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n495), .A2(new_n660), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n648), .A2(new_n633), .A3(new_n653), .A4(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(G143), .ZN(G45));
  INV_X1    g477(.A(new_n588), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT96), .ZN(new_n665));
  INV_X1    g479(.A(new_n642), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n664), .A2(new_n665), .A3(new_n637), .A4(new_n666), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n576), .A2(new_n587), .A3(new_n666), .ZN(new_n668));
  OAI21_X1  g482(.A(KEYINPUT96), .B1(new_n638), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  NOR3_X1   g484(.A1(new_n632), .A2(new_n633), .A3(new_n367), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(KEYINPUT97), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT97), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n670), .A2(new_n671), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G146), .ZN(G48));
  AOI21_X1  g491(.A(new_n632), .B1(new_n602), .B2(new_n572), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n196), .B1(new_n362), .B2(new_n363), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(KEYINPUT98), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT98), .ZN(new_n681));
  OAI211_X1 g495(.A(new_n681), .B(new_n196), .C1(new_n362), .C2(new_n363), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n680), .A2(G469), .A3(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n364), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n683), .B1(KEYINPUT99), .B2(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT99), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n680), .A2(new_n686), .A3(G469), .A4(new_n682), .ZN(new_n687));
  AND3_X1   g501(.A1(new_n685), .A2(new_n306), .A3(new_n687), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n678), .A2(new_n589), .A3(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(KEYINPUT41), .B(G113), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n689), .B(new_n690), .ZN(G15));
  NAND3_X1  g505(.A1(new_n615), .A2(new_n678), .A3(new_n688), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(KEYINPUT100), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT100), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n615), .A2(new_n678), .A3(new_n694), .A4(new_n688), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G116), .ZN(G18));
  NOR3_X1   g511(.A1(new_n632), .A2(new_n633), .A3(new_n638), .ZN(new_n698));
  INV_X1    g512(.A(new_n194), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n452), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n698), .A2(new_n688), .A3(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G119), .ZN(G21));
  OAI21_X1  g516(.A(KEYINPUT101), .B1(new_n600), .B2(new_n592), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT101), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n598), .A2(new_n568), .A3(new_n704), .A4(new_n570), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(new_n649), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n652), .A2(new_n707), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n706), .A2(new_n194), .A3(new_n688), .A4(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G122), .ZN(G24));
  INV_X1    g524(.A(KEYINPUT102), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n668), .A2(new_n711), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n576), .A2(new_n587), .A3(KEYINPUT102), .A4(new_n666), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n624), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  AND4_X1   g528(.A1(new_n306), .A2(new_n685), .A3(new_n637), .A4(new_n687), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G125), .ZN(G27));
  INV_X1    g531(.A(KEYINPUT42), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n602), .A2(new_n572), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n707), .A2(new_n195), .ZN(new_n720));
  NOR3_X1   g534(.A1(new_n347), .A2(new_n350), .A3(new_n308), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n306), .B1(new_n366), .B2(new_n721), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n719), .A2(new_n510), .A3(new_n723), .ZN(new_n724));
  AND2_X1   g538(.A1(new_n712), .A2(new_n713), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n718), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  AOI211_X1 g540(.A(new_n722), .B(new_n720), .C1(new_n712), .C2(new_n713), .ZN(new_n727));
  AND2_X1   g541(.A1(new_n490), .A2(new_n491), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n600), .B1(new_n728), .B2(new_n509), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n727), .A2(KEYINPUT42), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n726), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G131), .ZN(G33));
  NAND3_X1  g546(.A1(new_n643), .A2(new_n678), .A3(new_n723), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G134), .ZN(G36));
  INV_X1    g548(.A(KEYINPUT45), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n351), .A2(new_n359), .A3(new_n735), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n357), .A2(KEYINPUT45), .A3(new_n358), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n736), .A2(new_n737), .A3(G469), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n738), .A2(KEYINPUT46), .A3(new_n365), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(new_n364), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(KEYINPUT103), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n738), .A2(new_n365), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT46), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT103), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n739), .A2(new_n745), .A3(new_n364), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n741), .A2(new_n744), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(new_n306), .ZN(new_n748));
  INV_X1    g562(.A(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT104), .ZN(new_n750));
  INV_X1    g564(.A(new_n586), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(new_n584), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n750), .B1(new_n576), .B2(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT43), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  OAI211_X1 g569(.A(new_n750), .B(KEYINPUT43), .C1(new_n576), .C2(new_n752), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n755), .A2(new_n592), .A3(new_n623), .A4(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT44), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n749), .A2(new_n759), .A3(new_n646), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n649), .A2(new_n634), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n761), .B1(new_n757), .B2(new_n758), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(new_n323), .ZN(G39));
  INV_X1    g578(.A(KEYINPUT47), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n748), .A2(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n747), .A2(KEYINPUT47), .A3(new_n306), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n719), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NOR3_X1   g582(.A1(new_n510), .A2(new_n668), .A3(new_n720), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G140), .ZN(G42));
  INV_X1    g585(.A(KEYINPUT114), .ZN(new_n772));
  NOR2_X1   g586(.A1(G952), .A2(G953), .ZN(new_n773));
  XOR2_X1   g587(.A(KEYINPUT110), .B(KEYINPUT54), .Z(new_n774));
  INV_X1    g588(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n604), .A2(new_n642), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n510), .A2(new_n597), .A3(new_n623), .A4(new_n776), .ZN(new_n777));
  OAI211_X1 g591(.A(new_n761), .B(new_n605), .C1(new_n612), .C2(new_n613), .ZN(new_n778));
  OR3_X1    g592(.A1(new_n777), .A2(KEYINPUT108), .A3(new_n778), .ZN(new_n779));
  OAI21_X1  g593(.A(KEYINPUT108), .B1(new_n777), .B2(new_n778), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(new_n624), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n727), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n781), .A2(new_n733), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n574), .A2(new_n594), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT106), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(new_n576), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n788), .A2(new_n604), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n789), .A2(new_n303), .ZN(new_n790));
  AOI22_X1  g604(.A1(new_n453), .A2(new_n628), .B1(new_n603), .B2(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n574), .A2(KEYINPUT106), .A3(new_n594), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n787), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(KEYINPUT107), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT107), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n787), .A2(new_n791), .A3(new_n795), .A4(new_n792), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n784), .B1(new_n794), .B2(new_n796), .ZN(new_n797));
  AOI22_X1  g611(.A1(new_n639), .A2(new_n643), .B1(new_n714), .B2(new_n715), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n652), .A2(new_n707), .A3(new_n722), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n799), .A2(new_n661), .A3(new_n633), .A4(new_n666), .ZN(new_n800));
  INV_X1    g614(.A(new_n675), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n674), .B1(new_n670), .B2(new_n671), .ZN(new_n802));
  OAI211_X1 g616(.A(new_n798), .B(new_n800), .C1(new_n801), .C2(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT52), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n676), .A2(KEYINPUT52), .A3(new_n798), .A4(new_n800), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  AND2_X1   g621(.A1(new_n797), .A2(new_n807), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n709), .A2(new_n689), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n696), .A2(new_n731), .A3(new_n701), .A4(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n810), .A2(KEYINPUT109), .ZN(new_n811));
  INV_X1    g625(.A(new_n701), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n812), .B1(new_n693), .B2(new_n695), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT109), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n813), .A2(new_n814), .A3(new_n731), .A4(new_n809), .ZN(new_n815));
  AND3_X1   g629(.A1(new_n811), .A2(KEYINPUT53), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n794), .A2(new_n796), .ZN(new_n817));
  AND4_X1   g631(.A1(new_n696), .A2(new_n701), .A3(new_n731), .A4(new_n809), .ZN(new_n818));
  INV_X1    g632(.A(new_n784), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n807), .A2(new_n817), .A3(new_n818), .A4(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT53), .ZN(new_n821));
  AOI22_X1  g635(.A1(new_n808), .A2(new_n816), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n820), .A2(new_n821), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n797), .A2(KEYINPUT53), .A3(new_n807), .A4(new_n818), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  AOI22_X1  g639(.A1(new_n775), .A2(new_n822), .B1(new_n825), .B2(KEYINPUT54), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n688), .A2(new_n761), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n755), .A2(new_n640), .A3(new_n756), .ZN(new_n828));
  AND2_X1   g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n829), .A2(new_n729), .ZN(new_n830));
  XNOR2_X1  g644(.A(new_n830), .B(KEYINPUT48), .ZN(new_n831));
  AND2_X1   g645(.A1(new_n828), .A2(new_n706), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n832), .A2(new_n715), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n188), .A2(G952), .ZN(new_n834));
  INV_X1    g648(.A(new_n661), .ZN(new_n835));
  AND4_X1   g649(.A1(new_n719), .A2(new_n827), .A3(new_n640), .A4(new_n835), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n834), .B1(new_n836), .B2(new_n664), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n831), .A2(new_n833), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n836), .A2(new_n788), .A3(new_n752), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n829), .A2(new_n782), .ZN(new_n841));
  OR2_X1    g655(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n840), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(new_n307), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n685), .A2(new_n844), .A3(new_n687), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n766), .A2(new_n845), .A3(new_n767), .ZN(new_n846));
  AND2_X1   g660(.A1(new_n846), .A2(new_n832), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n843), .B1(new_n847), .B2(new_n761), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n651), .A2(new_n634), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n828), .A2(new_n849), .A3(new_n688), .A4(new_n706), .ZN(new_n850));
  OR2_X1    g664(.A1(new_n850), .A2(KEYINPUT111), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT50), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n850), .A2(KEYINPUT111), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT112), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  OR2_X1    g670(.A1(new_n850), .A2(new_n852), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n851), .A2(KEYINPUT112), .A3(new_n853), .A4(new_n852), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n856), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n839), .B1(new_n848), .B2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n848), .A2(new_n859), .A3(new_n839), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n838), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n773), .B1(new_n826), .B2(new_n863), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n600), .A2(new_n844), .A3(new_n634), .ZN(new_n865));
  XOR2_X1   g679(.A(new_n865), .B(KEYINPUT105), .Z(new_n866));
  NAND2_X1  g680(.A1(new_n685), .A2(new_n687), .ZN(new_n867));
  AOI211_X1 g681(.A(new_n576), .B(new_n752), .C1(new_n867), .C2(KEYINPUT49), .ZN(new_n868));
  OR2_X1    g682(.A1(new_n867), .A2(KEYINPUT49), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n868), .A2(new_n651), .A3(new_n835), .A4(new_n869), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n866), .A2(new_n870), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n772), .B1(new_n864), .B2(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(new_n871), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n821), .B1(new_n810), .B2(KEYINPUT109), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n874), .A2(new_n797), .A3(new_n807), .A4(new_n815), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n823), .A2(new_n875), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n876), .A2(new_n774), .ZN(new_n877));
  INV_X1    g691(.A(new_n838), .ZN(new_n878));
  AND3_X1   g692(.A1(new_n848), .A2(new_n859), .A3(new_n839), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n878), .B1(new_n879), .B2(new_n860), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT54), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n881), .B1(new_n823), .B2(new_n824), .ZN(new_n882));
  NOR3_X1   g696(.A1(new_n877), .A2(new_n880), .A3(new_n882), .ZN(new_n883));
  OAI211_X1 g697(.A(KEYINPUT114), .B(new_n873), .C1(new_n883), .C2(new_n773), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n872), .A2(new_n884), .ZN(G75));
  INV_X1    g699(.A(KEYINPUT116), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n188), .A2(G952), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n876), .A2(G210), .A3(G902), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n299), .B(new_n290), .ZN(new_n889));
  XOR2_X1   g703(.A(new_n889), .B(KEYINPUT55), .Z(new_n890));
  XNOR2_X1  g704(.A(KEYINPUT115), .B(KEYINPUT56), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n887), .B1(new_n888), .B2(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(new_n890), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT56), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n895), .B1(new_n888), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n886), .B1(new_n894), .B2(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(new_n897), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n899), .A2(KEYINPUT116), .A3(new_n893), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n898), .A2(new_n900), .ZN(G51));
  NOR2_X1   g715(.A1(new_n822), .A2(new_n775), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n902), .A2(new_n877), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n365), .B(KEYINPUT57), .ZN(new_n904));
  OAI22_X1  g718(.A1(new_n903), .A2(new_n904), .B1(new_n363), .B2(new_n362), .ZN(new_n905));
  OR3_X1    g719(.A1(new_n822), .A2(new_n196), .A3(new_n738), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n887), .B1(new_n905), .B2(new_n906), .ZN(G54));
  INV_X1    g721(.A(KEYINPUT58), .ZN(new_n908));
  OAI21_X1  g722(.A(KEYINPUT117), .B1(new_n908), .B2(new_n607), .ZN(new_n909));
  OR3_X1    g723(.A1(new_n908), .A2(new_n607), .A3(KEYINPUT117), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n876), .A2(G902), .A3(new_n909), .A4(new_n910), .ZN(new_n911));
  AND2_X1   g725(.A1(new_n911), .A2(new_n450), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n911), .A2(new_n450), .ZN(new_n913));
  NOR3_X1   g727(.A1(new_n912), .A2(new_n913), .A3(new_n887), .ZN(G60));
  AND2_X1   g728(.A1(new_n578), .A2(new_n579), .ZN(new_n915));
  XNOR2_X1  g729(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n436), .A2(new_n196), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n916), .B(new_n917), .Z(new_n918));
  OAI211_X1 g732(.A(new_n915), .B(new_n918), .C1(new_n902), .C2(new_n877), .ZN(new_n919));
  INV_X1    g733(.A(new_n887), .ZN(new_n920));
  INV_X1    g734(.A(new_n918), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n826), .A2(new_n921), .ZN(new_n922));
  OAI211_X1 g736(.A(new_n919), .B(new_n920), .C1(new_n922), .C2(new_n915), .ZN(new_n923));
  INV_X1    g737(.A(new_n923), .ZN(G63));
  NAND2_X1  g738(.A1(G217), .A2(G902), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n925), .B(KEYINPUT60), .Z(new_n926));
  NAND3_X1  g740(.A1(new_n876), .A2(new_n621), .A3(new_n926), .ZN(new_n927));
  AND2_X1   g741(.A1(new_n927), .A2(new_n920), .ZN(new_n928));
  NAND2_X1  g742(.A1(KEYINPUT119), .A2(KEYINPUT61), .ZN(new_n929));
  OR2_X1    g743(.A1(KEYINPUT119), .A2(KEYINPUT61), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n565), .B1(new_n876), .B2(new_n926), .ZN(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n928), .A2(new_n929), .A3(new_n930), .A4(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n927), .A2(new_n920), .ZN(new_n934));
  OAI211_X1 g748(.A(KEYINPUT119), .B(KEYINPUT61), .C1(new_n934), .C2(new_n931), .ZN(new_n935));
  AND2_X1   g749(.A1(new_n933), .A2(new_n935), .ZN(G66));
  AOI21_X1  g750(.A(new_n188), .B1(new_n191), .B2(G224), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n817), .A2(new_n809), .A3(new_n813), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n937), .B1(new_n938), .B2(new_n188), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n289), .B1(G898), .B2(new_n188), .ZN(new_n940));
  XOR2_X1   g754(.A(new_n940), .B(KEYINPUT120), .Z(new_n941));
  XNOR2_X1  g755(.A(new_n939), .B(new_n941), .ZN(G69));
  NOR2_X1   g756(.A1(new_n461), .A2(new_n462), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(KEYINPUT121), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n944), .B(new_n441), .Z(new_n945));
  NAND2_X1  g759(.A1(G900), .A2(G953), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n731), .A2(new_n733), .ZN(new_n947));
  XOR2_X1   g761(.A(new_n947), .B(KEYINPUT123), .Z(new_n948));
  AOI21_X1  g762(.A(new_n763), .B1(new_n768), .B2(new_n769), .ZN(new_n949));
  AND2_X1   g763(.A1(new_n676), .A2(new_n798), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n749), .A2(new_n646), .A3(new_n708), .A4(new_n729), .ZN(new_n951));
  NAND4_X1  g765(.A1(new_n948), .A2(new_n949), .A3(new_n950), .A4(new_n951), .ZN(new_n952));
  OAI211_X1 g766(.A(new_n945), .B(new_n946), .C1(new_n952), .C2(G953), .ZN(new_n953));
  OAI21_X1  g767(.A(G953), .B1(new_n311), .B2(new_n641), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n950), .A2(new_n662), .ZN(new_n955));
  XOR2_X1   g769(.A(KEYINPUT122), .B(KEYINPUT62), .Z(new_n956));
  NAND2_X1  g770(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(new_n647), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n789), .A2(new_n588), .ZN(new_n959));
  NAND4_X1  g773(.A1(new_n678), .A2(new_n958), .A3(new_n761), .A4(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT62), .ZN(new_n961));
  OAI211_X1 g775(.A(new_n950), .B(new_n662), .C1(KEYINPUT122), .C2(new_n961), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n949), .A2(new_n957), .A3(new_n960), .A4(new_n962), .ZN(new_n963));
  AND2_X1   g777(.A1(new_n963), .A2(new_n188), .ZN(new_n964));
  OAI221_X1 g778(.A(new_n953), .B1(KEYINPUT124), .B2(new_n954), .C1(new_n964), .C2(new_n945), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n954), .A2(KEYINPUT124), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n965), .B(new_n966), .ZN(G72));
  NAND2_X1  g781(.A1(G472), .A2(G902), .ZN(new_n968));
  XOR2_X1   g782(.A(new_n968), .B(KEYINPUT63), .Z(new_n969));
  OAI21_X1  g783(.A(new_n969), .B1(new_n963), .B2(new_n938), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT125), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  OAI211_X1 g786(.A(KEYINPUT125), .B(new_n969), .C1(new_n963), .C2(new_n938), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n972), .A2(new_n656), .A3(new_n973), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n969), .B1(new_n952), .B2(new_n938), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n655), .A2(new_n476), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n976), .B(KEYINPUT126), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n887), .B1(new_n975), .B2(new_n977), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n656), .B1(new_n823), .B2(new_n824), .ZN(new_n979));
  INV_X1    g793(.A(KEYINPUT127), .ZN(new_n980));
  AND2_X1   g794(.A1(new_n976), .A2(new_n969), .ZN(new_n981));
  AND3_X1   g795(.A1(new_n979), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n980), .B1(new_n979), .B2(new_n981), .ZN(new_n983));
  OAI211_X1 g797(.A(new_n974), .B(new_n978), .C1(new_n982), .C2(new_n983), .ZN(new_n984));
  INV_X1    g798(.A(new_n984), .ZN(G57));
endmodule


