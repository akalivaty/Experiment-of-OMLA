//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 0 1 1 1 0 1 0 0 0 1 1 1 1 1 0 0 0 0 0 0 1 1 0 0 0 0 1 0 1 1 1 1 1 0 0 0 1 1 1 1 1 1 1 0 0 0 1 0 0 0 1 1 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:36 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n557, new_n558, new_n559,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n574, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n620, new_n623, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n849, new_n850,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  XNOR2_X1  g032(.A(KEYINPUT3), .B(G2104), .ZN(new_n458));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  NAND3_X1  g034(.A1(new_n458), .A2(G137), .A3(new_n459), .ZN(new_n460));
  AND2_X1   g035(.A1(new_n459), .A2(G2104), .ZN(new_n461));
  AND3_X1   g036(.A1(new_n461), .A2(KEYINPUT66), .A3(G101), .ZN(new_n462));
  AOI21_X1  g037(.A(KEYINPUT66), .B1(new_n461), .B2(G101), .ZN(new_n463));
  OAI21_X1  g038(.A(new_n460), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT65), .ZN(new_n466));
  OR2_X1    g041(.A1(new_n458), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n458), .A2(new_n466), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G125), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n465), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n464), .B1(new_n471), .B2(G2105), .ZN(G160));
  AND2_X1   g047(.A1(new_n458), .A2(KEYINPUT67), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n458), .A2(KEYINPUT67), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n459), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G136), .ZN(new_n477));
  OAI21_X1  g052(.A(G2105), .B1(new_n473), .B2(new_n474), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n459), .A2(G112), .ZN(new_n481));
  OAI21_X1  g056(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n477), .B(new_n480), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G162));
  INV_X1    g059(.A(G114), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(KEYINPUT68), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT68), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G114), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n459), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  XNOR2_X1  g064(.A(new_n489), .B(KEYINPUT69), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n490), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n491));
  AND3_X1   g066(.A1(new_n458), .A2(G126), .A3(G2105), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  AND2_X1   g068(.A1(new_n459), .A2(G138), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n467), .A2(new_n493), .A3(new_n468), .A4(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n458), .A2(new_n494), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n492), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n491), .A2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  NAND2_X1  g075(.A1(G75), .A2(G543), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT5), .ZN(new_n502));
  OAI21_X1  g077(.A(KEYINPUT70), .B1(new_n502), .B2(G543), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT70), .ZN(new_n504));
  INV_X1    g079(.A(G543), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n504), .A2(new_n505), .A3(KEYINPUT5), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n503), .A2(new_n506), .ZN(new_n507));
  OAI21_X1  g082(.A(KEYINPUT71), .B1(new_n505), .B2(KEYINPUT5), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT71), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n509), .A2(new_n502), .A3(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n507), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G62), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n501), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G651), .ZN(new_n515));
  XNOR2_X1  g090(.A(KEYINPUT6), .B(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G543), .ZN(new_n517));
  INV_X1    g092(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G50), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n515), .A2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT72), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n503), .A2(new_n506), .B1(new_n508), .B2(new_n510), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n521), .B1(new_n522), .B2(new_n516), .ZN(new_n523));
  AND4_X1   g098(.A1(new_n521), .A2(new_n507), .A3(new_n511), .A4(new_n516), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n520), .B1(G88), .B2(new_n525), .ZN(G166));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n527), .B(KEYINPUT7), .ZN(new_n528));
  INV_X1    g103(.A(G51), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n528), .B1(new_n517), .B2(new_n529), .ZN(new_n530));
  AND2_X1   g105(.A1(G63), .A2(G651), .ZN(new_n531));
  AOI21_X1  g106(.A(new_n530), .B1(new_n522), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n507), .A2(new_n511), .A3(new_n516), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(KEYINPUT72), .ZN(new_n534));
  NAND4_X1  g109(.A1(new_n507), .A2(new_n511), .A3(new_n521), .A4(new_n516), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n534), .A2(G89), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n532), .A2(new_n536), .ZN(G286));
  INV_X1    g112(.A(G286), .ZN(G168));
  NAND2_X1  g113(.A1(G77), .A2(G543), .ZN(new_n539));
  INV_X1    g114(.A(G64), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n539), .B1(new_n512), .B2(new_n540), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n541), .A2(G651), .B1(G52), .B2(new_n518), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n534), .A2(G90), .A3(new_n535), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n542), .A2(new_n543), .ZN(G301));
  INV_X1    g119(.A(G301), .ZN(G171));
  NAND3_X1  g120(.A1(new_n516), .A2(G43), .A3(G543), .ZN(new_n546));
  INV_X1    g121(.A(new_n546), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n507), .A2(new_n511), .A3(G56), .ZN(new_n548));
  NAND2_X1  g123(.A1(G68), .A2(G543), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  AOI21_X1  g125(.A(new_n547), .B1(new_n550), .B2(G651), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n534), .A2(G81), .A3(new_n535), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  NAND4_X1  g130(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g131(.A(KEYINPUT73), .B(KEYINPUT8), .Z(new_n557));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n557), .B(new_n558), .ZN(new_n559));
  NAND4_X1  g134(.A1(G319), .A2(G483), .A3(G661), .A4(new_n559), .ZN(G188));
  NAND2_X1  g135(.A1(G78), .A2(G543), .ZN(new_n561));
  INV_X1    g136(.A(G65), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n561), .B1(new_n512), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G651), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n516), .A2(G53), .A3(G543), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT9), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT74), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n568), .B1(new_n523), .B2(new_n524), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n534), .A2(KEYINPUT74), .A3(new_n535), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n567), .B1(new_n571), .B2(G91), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(G299));
  NAND2_X1  g148(.A1(new_n525), .A2(G88), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n574), .A2(new_n515), .A3(new_n519), .ZN(G303));
  NAND2_X1  g150(.A1(new_n571), .A2(G87), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n518), .A2(KEYINPUT75), .A3(G49), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT75), .ZN(new_n578));
  INV_X1    g153(.A(G49), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n578), .B1(new_n517), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  OAI21_X1  g156(.A(G651), .B1(new_n522), .B2(G74), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n576), .A2(new_n584), .ZN(G288));
  INV_X1    g160(.A(G86), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n586), .B1(new_n569), .B2(new_n570), .ZN(new_n587));
  NAND2_X1  g162(.A1(G73), .A2(G543), .ZN(new_n588));
  INV_X1    g163(.A(G61), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n512), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n590), .A2(G651), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n518), .A2(KEYINPUT76), .A3(G48), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT76), .ZN(new_n593));
  INV_X1    g168(.A(G48), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n517), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n591), .A2(new_n596), .ZN(new_n597));
  OR2_X1    g172(.A1(new_n587), .A2(new_n597), .ZN(G305));
  NAND2_X1  g173(.A1(G72), .A2(G543), .ZN(new_n599));
  INV_X1    g174(.A(G60), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n512), .B2(new_n600), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n601), .A2(G651), .B1(G47), .B2(new_n518), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n534), .A2(G85), .A3(new_n535), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(new_n603), .ZN(G290));
  NAND2_X1  g179(.A1(G301), .A2(G868), .ZN(new_n605));
  XOR2_X1   g180(.A(new_n605), .B(KEYINPUT77), .Z(new_n606));
  NAND2_X1  g181(.A1(G79), .A2(G543), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n607), .B(KEYINPUT78), .ZN(new_n608));
  INV_X1    g183(.A(G66), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n512), .B2(new_n609), .ZN(new_n610));
  AOI22_X1  g185(.A1(new_n610), .A2(G651), .B1(G54), .B2(new_n518), .ZN(new_n611));
  AOI21_X1  g186(.A(KEYINPUT10), .B1(new_n571), .B2(G92), .ZN(new_n612));
  INV_X1    g187(.A(KEYINPUT10), .ZN(new_n613));
  INV_X1    g188(.A(G92), .ZN(new_n614));
  AOI211_X1 g189(.A(new_n613), .B(new_n614), .C1(new_n569), .C2(new_n570), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n611), .B1(new_n612), .B2(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(new_n616), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n606), .B1(new_n617), .B2(G868), .ZN(G284));
  OAI21_X1  g193(.A(new_n606), .B1(new_n617), .B2(G868), .ZN(G321));
  NAND2_X1  g194(.A1(G286), .A2(G868), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n620), .B1(new_n572), .B2(G868), .ZN(G297));
  OAI21_X1  g196(.A(new_n620), .B1(new_n572), .B2(G868), .ZN(G280));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n617), .B1(new_n623), .B2(G860), .ZN(G148));
  INV_X1    g199(.A(KEYINPUT79), .ZN(new_n625));
  AOI21_X1  g200(.A(new_n625), .B1(new_n617), .B2(new_n623), .ZN(new_n626));
  NOR3_X1   g201(.A1(new_n523), .A2(new_n524), .A3(new_n568), .ZN(new_n627));
  AOI21_X1  g202(.A(KEYINPUT74), .B1(new_n534), .B2(new_n535), .ZN(new_n628));
  OAI21_X1  g203(.A(G92), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n629), .A2(new_n613), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n571), .A2(KEYINPUT10), .A3(G92), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n632), .A2(new_n623), .A3(new_n611), .ZN(new_n633));
  NOR2_X1   g208(.A1(new_n633), .A2(KEYINPUT79), .ZN(new_n634));
  INV_X1    g209(.A(G868), .ZN(new_n635));
  NOR3_X1   g210(.A1(new_n626), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  AOI21_X1  g211(.A(new_n636), .B1(new_n635), .B2(new_n554), .ZN(G323));
  XNOR2_X1  g212(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g213(.A1(new_n467), .A2(new_n468), .A3(new_n461), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(KEYINPUT12), .Z(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(KEYINPUT13), .Z(new_n641));
  INV_X1    g216(.A(G2100), .ZN(new_n642));
  OR2_X1    g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n641), .A2(new_n642), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n476), .A2(G135), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n479), .A2(G123), .ZN(new_n646));
  NOR2_X1   g221(.A1(new_n459), .A2(G111), .ZN(new_n647));
  OAI21_X1  g222(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n648));
  OAI211_X1 g223(.A(new_n645), .B(new_n646), .C1(new_n647), .C2(new_n648), .ZN(new_n649));
  INV_X1    g224(.A(G2096), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n643), .A2(new_n644), .A3(new_n651), .ZN(G156));
  XNOR2_X1  g227(.A(KEYINPUT15), .B(G2435), .ZN(new_n653));
  XNOR2_X1  g228(.A(KEYINPUT80), .B(G2438), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2427), .B(G2430), .ZN(new_n656));
  OR2_X1    g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n655), .A2(new_n656), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n657), .A2(KEYINPUT14), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2451), .B(G2454), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT16), .ZN(new_n661));
  XOR2_X1   g236(.A(G1341), .B(G1348), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n659), .B(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(G2443), .B(G2446), .Z(new_n665));
  OAI21_X1  g240(.A(G14), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n666), .B1(new_n665), .B2(new_n664), .ZN(G401));
  INV_X1    g242(.A(KEYINPUT18), .ZN(new_n668));
  XOR2_X1   g243(.A(G2084), .B(G2090), .Z(new_n669));
  XNOR2_X1  g244(.A(G2067), .B(G2678), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n671), .A2(KEYINPUT17), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n669), .A2(new_n670), .ZN(new_n673));
  OAI21_X1  g248(.A(new_n668), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(KEYINPUT81), .B(G2100), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(G2072), .B(G2078), .Z(new_n677));
  AOI21_X1  g252(.A(new_n677), .B1(new_n671), .B2(KEYINPUT18), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(new_n650), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n676), .B(new_n679), .ZN(G227));
  XOR2_X1   g255(.A(G1956), .B(G2474), .Z(new_n681));
  XOR2_X1   g256(.A(G1961), .B(G1966), .Z(new_n682));
  NAND2_X1  g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n683), .A2(KEYINPUT82), .ZN(new_n684));
  XOR2_X1   g259(.A(G1971), .B(G1976), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT19), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n683), .A2(KEYINPUT82), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n684), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  XOR2_X1   g263(.A(KEYINPUT83), .B(KEYINPUT20), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n681), .A2(new_n682), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n686), .A2(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(new_n691), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n693), .A2(new_n683), .ZN(new_n694));
  OAI211_X1 g269(.A(new_n690), .B(new_n692), .C1(new_n686), .C2(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XOR2_X1   g272(.A(G1991), .B(G1996), .Z(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  OR2_X1    g274(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1981), .B(G1986), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n697), .A2(new_n699), .ZN(new_n702));
  AND3_X1   g277(.A1(new_n700), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n701), .B1(new_n700), .B2(new_n702), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n703), .A2(new_n704), .ZN(G229));
  NOR2_X1   g280(.A1(G29), .A2(G33), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT94), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n459), .A2(G103), .A3(G2104), .ZN(new_n708));
  XOR2_X1   g283(.A(new_n708), .B(KEYINPUT25), .Z(new_n709));
  INV_X1    g284(.A(G139), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n709), .B1(new_n475), .B2(new_n710), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n467), .A2(G127), .A3(new_n468), .ZN(new_n712));
  NAND2_X1  g287(.A1(G115), .A2(G2104), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n459), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n711), .A2(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(G29), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n707), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT95), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(G2072), .Z(new_n720));
  NAND2_X1  g295(.A1(new_n717), .A2(G35), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(G162), .B2(new_n717), .ZN(new_n722));
  INV_X1    g297(.A(KEYINPUT29), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(new_n724), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n720), .B1(G2090), .B2(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(G16), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n727), .A2(G20), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT23), .Z(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(G299), .B2(G16), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(G1956), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n476), .A2(G141), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n479), .A2(G129), .ZN(new_n733));
  NAND3_X1  g308(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n734));
  INV_X1    g309(.A(KEYINPUT26), .ZN(new_n735));
  OR2_X1    g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n734), .A2(new_n735), .ZN(new_n737));
  AOI22_X1  g312(.A1(new_n736), .A2(new_n737), .B1(G105), .B2(new_n461), .ZN(new_n738));
  NAND3_X1  g313(.A1(new_n732), .A2(new_n733), .A3(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n740), .A2(new_n717), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(new_n717), .B2(G32), .ZN(new_n742));
  XNOR2_X1  g317(.A(KEYINPUT27), .B(G1996), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  XOR2_X1   g319(.A(new_n744), .B(KEYINPUT98), .Z(new_n745));
  NAND2_X1  g320(.A1(new_n727), .A2(G19), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(new_n554), .B2(new_n727), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(G1341), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n745), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g324(.A(KEYINPUT30), .B(G28), .ZN(new_n750));
  OR2_X1    g325(.A1(KEYINPUT31), .A2(G11), .ZN(new_n751));
  NAND2_X1  g326(.A1(KEYINPUT31), .A2(G11), .ZN(new_n752));
  AOI22_X1  g327(.A1(new_n750), .A2(new_n717), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(new_n649), .B2(new_n717), .ZN(new_n754));
  NAND2_X1  g329(.A1(G164), .A2(G29), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(G27), .B2(G29), .ZN(new_n756));
  INV_X1    g331(.A(G2078), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n754), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(G1966), .ZN(new_n759));
  NOR2_X1   g334(.A1(G168), .A2(new_n727), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(new_n727), .B2(G21), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n758), .B1(new_n759), .B2(new_n761), .ZN(new_n762));
  OAI22_X1  g337(.A1(new_n742), .A2(new_n743), .B1(new_n757), .B2(new_n756), .ZN(new_n763));
  XNOR2_X1  g338(.A(KEYINPUT96), .B(KEYINPUT24), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n764), .A2(G34), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n717), .B1(new_n764), .B2(G34), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n765), .B1(new_n766), .B2(KEYINPUT97), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(KEYINPUT97), .B2(new_n766), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(G160), .B2(G29), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(G2084), .ZN(new_n770));
  NOR3_X1   g345(.A1(new_n762), .A2(new_n763), .A3(new_n770), .ZN(new_n771));
  NAND4_X1  g346(.A1(new_n726), .A2(new_n731), .A3(new_n749), .A4(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(G2090), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n724), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT99), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n617), .A2(G16), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(G4), .B2(G16), .ZN(new_n777));
  INV_X1    g352(.A(G1348), .ZN(new_n778));
  OR2_X1    g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n777), .A2(new_n778), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n717), .A2(G26), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT28), .ZN(new_n782));
  OR2_X1    g357(.A1(G104), .A2(G2105), .ZN(new_n783));
  OAI211_X1 g358(.A(new_n783), .B(G2104), .C1(G116), .C2(new_n459), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n784), .B(KEYINPUT92), .Z(new_n785));
  INV_X1    g360(.A(G140), .ZN(new_n786));
  INV_X1    g361(.A(G128), .ZN(new_n787));
  OAI221_X1 g362(.A(new_n785), .B1(new_n475), .B2(new_n786), .C1(new_n787), .C2(new_n478), .ZN(new_n788));
  AND3_X1   g363(.A1(new_n788), .A2(KEYINPUT93), .A3(G29), .ZN(new_n789));
  AOI21_X1  g364(.A(KEYINPUT93), .B1(new_n788), .B2(G29), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n782), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  INV_X1    g366(.A(G2067), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  NOR2_X1   g368(.A1(G171), .A2(new_n727), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(G5), .B2(new_n727), .ZN(new_n795));
  INV_X1    g370(.A(G1961), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n761), .A2(new_n759), .ZN(new_n798));
  OR2_X1    g373(.A1(new_n795), .A2(new_n796), .ZN(new_n799));
  AND4_X1   g374(.A1(new_n793), .A2(new_n797), .A3(new_n798), .A4(new_n799), .ZN(new_n800));
  NAND4_X1  g375(.A1(new_n775), .A2(new_n779), .A3(new_n780), .A4(new_n800), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n772), .A2(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(new_n802), .ZN(new_n803));
  NOR2_X1   g378(.A1(G16), .A2(G23), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT88), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(G288), .B2(new_n727), .ZN(new_n806));
  XNOR2_X1  g381(.A(KEYINPUT33), .B(G1976), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(KEYINPUT89), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n587), .A2(new_n597), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n811), .A2(new_n727), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(G6), .B2(new_n727), .ZN(new_n813));
  XNOR2_X1  g388(.A(KEYINPUT32), .B(G1981), .ZN(new_n814));
  INV_X1    g389(.A(new_n814), .ZN(new_n815));
  OR2_X1    g390(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n813), .A2(new_n815), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n727), .A2(G22), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n818), .B1(G166), .B2(new_n727), .ZN(new_n819));
  INV_X1    g394(.A(G1971), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  NAND4_X1  g396(.A1(new_n810), .A2(new_n816), .A3(new_n817), .A4(new_n821), .ZN(new_n822));
  XOR2_X1   g397(.A(KEYINPUT90), .B(KEYINPUT34), .Z(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n717), .A2(G25), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n476), .A2(G131), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n479), .A2(G119), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n459), .A2(G107), .ZN(new_n828));
  OAI21_X1  g403(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n829));
  OAI211_X1 g404(.A(new_n826), .B(new_n827), .C1(new_n828), .C2(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT84), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n825), .B1(new_n831), .B2(new_n717), .ZN(new_n832));
  XOR2_X1   g407(.A(KEYINPUT35), .B(G1991), .Z(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT85), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n832), .B(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n727), .A2(G24), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT86), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n837), .B1(G290), .B2(G16), .ZN(new_n838));
  XNOR2_X1  g413(.A(KEYINPUT87), .B(G1986), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n838), .B(new_n839), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n835), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n824), .A2(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT36), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n843), .A2(KEYINPUT91), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(new_n844), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n824), .A2(new_n846), .A3(new_n841), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n803), .B1(new_n845), .B2(new_n847), .ZN(G311));
  AND3_X1   g423(.A1(new_n824), .A2(new_n846), .A3(new_n841), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n846), .B1(new_n824), .B2(new_n841), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n802), .B1(new_n849), .B2(new_n850), .ZN(G150));
  INV_X1    g426(.A(KEYINPUT100), .ZN(new_n852));
  AND3_X1   g427(.A1(new_n551), .A2(new_n852), .A3(new_n552), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n852), .B1(new_n551), .B2(new_n552), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n516), .A2(G55), .A3(G543), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(G80), .A2(G543), .ZN(new_n857));
  INV_X1    g432(.A(G67), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n857), .B1(new_n512), .B2(new_n858), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n856), .B1(new_n859), .B2(G651), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n534), .A2(G93), .A3(new_n535), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NOR3_X1   g437(.A1(new_n853), .A2(new_n854), .A3(new_n862), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n862), .A2(new_n553), .A3(KEYINPUT100), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(KEYINPUT38), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n616), .A2(new_n623), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n867), .B(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT39), .ZN(new_n870));
  AOI21_X1  g445(.A(G860), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n871), .B1(new_n870), .B2(new_n869), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n862), .A2(G860), .ZN(new_n873));
  XOR2_X1   g448(.A(new_n873), .B(KEYINPUT37), .Z(new_n874));
  NAND2_X1  g449(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(KEYINPUT101), .ZN(G145));
  XOR2_X1   g451(.A(new_n483), .B(new_n649), .Z(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(G160), .ZN(new_n878));
  OR2_X1    g453(.A1(G106), .A2(G2105), .ZN(new_n879));
  OAI211_X1 g454(.A(new_n879), .B(G2104), .C1(G118), .C2(new_n459), .ZN(new_n880));
  INV_X1    g455(.A(G142), .ZN(new_n881));
  INV_X1    g456(.A(G130), .ZN(new_n882));
  OAI221_X1 g457(.A(new_n880), .B1(new_n475), .B2(new_n881), .C1(new_n882), .C2(new_n478), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(KEYINPUT102), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(new_n640), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(new_n831), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n886), .A2(KEYINPUT103), .ZN(new_n887));
  INV_X1    g462(.A(new_n831), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n885), .B(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT103), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n788), .B(new_n499), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(new_n739), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n893), .B(new_n716), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  AND3_X1   g470(.A1(new_n887), .A2(new_n891), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n895), .B1(new_n887), .B2(new_n891), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n878), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n887), .A2(new_n891), .A3(new_n895), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n878), .B1(new_n894), .B2(new_n889), .ZN(new_n900));
  AOI21_X1  g475(.A(G37), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n898), .A2(new_n901), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n902), .B(KEYINPUT40), .ZN(G395));
  OAI22_X1  g478(.A1(new_n626), .A2(new_n634), .B1(new_n865), .B2(new_n863), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n617), .A2(new_n625), .A3(new_n623), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n633), .A2(KEYINPUT79), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n905), .A2(new_n906), .A3(new_n866), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n904), .A2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT104), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n572), .B1(new_n632), .B2(new_n611), .ZN(new_n910));
  OAI211_X1 g485(.A(new_n572), .B(new_n611), .C1(new_n612), .C2(new_n615), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n909), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n616), .A2(G299), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n914), .A2(KEYINPUT104), .A3(new_n911), .ZN(new_n915));
  AND2_X1   g490(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n908), .A2(new_n916), .ZN(new_n917));
  XOR2_X1   g492(.A(KEYINPUT106), .B(KEYINPUT41), .Z(new_n918));
  AOI21_X1  g493(.A(new_n918), .B1(new_n914), .B2(new_n911), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT41), .ZN(new_n920));
  AND3_X1   g495(.A1(new_n914), .A2(new_n920), .A3(new_n911), .ZN(new_n921));
  OAI211_X1 g496(.A(new_n904), .B(new_n907), .C1(new_n919), .C2(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n917), .A2(KEYINPUT105), .A3(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT105), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n908), .A2(new_n924), .A3(new_n916), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n602), .A2(KEYINPUT107), .A3(new_n603), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(KEYINPUT107), .B1(new_n602), .B2(new_n603), .ZN(new_n929));
  OAI211_X1 g504(.A(new_n576), .B(new_n584), .C1(new_n928), .C2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT107), .ZN(new_n931));
  NAND2_X1  g506(.A1(G290), .A2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(G87), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n933), .B1(new_n569), .B2(new_n570), .ZN(new_n934));
  OAI211_X1 g509(.A(new_n932), .B(new_n927), .C1(new_n934), .C2(new_n583), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n930), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n811), .A2(G303), .ZN(new_n937));
  OAI21_X1  g512(.A(G166), .B1(new_n597), .B2(new_n587), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n936), .A2(new_n939), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n930), .A2(new_n935), .A3(new_n937), .A4(new_n938), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n942), .B(KEYINPUT42), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n926), .A2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(new_n943), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n923), .A2(new_n925), .A3(new_n945), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n944), .A2(G868), .A3(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT108), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n948), .B1(new_n862), .B2(new_n635), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n944), .A2(new_n948), .A3(G868), .A4(new_n946), .ZN(new_n951));
  AND2_X1   g526(.A1(new_n950), .A2(new_n951), .ZN(G295));
  AND2_X1   g527(.A1(new_n950), .A2(new_n951), .ZN(G331));
  INV_X1    g528(.A(KEYINPUT44), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n553), .A2(KEYINPUT100), .ZN(new_n955));
  AND2_X1   g530(.A1(new_n860), .A2(new_n861), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n551), .A2(new_n852), .A3(new_n552), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n955), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(G301), .A2(G286), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n542), .A2(new_n536), .A3(new_n532), .A4(new_n543), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n958), .A2(new_n864), .A3(new_n959), .A4(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT110), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n959), .A2(new_n960), .ZN(new_n964));
  INV_X1    g539(.A(new_n964), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n965), .A2(KEYINPUT110), .A3(new_n864), .A4(new_n958), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n964), .B1(new_n863), .B2(new_n865), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n963), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  AND3_X1   g543(.A1(new_n914), .A2(new_n911), .A3(new_n918), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n920), .B1(new_n914), .B2(new_n911), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n968), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n967), .A2(KEYINPUT109), .A3(new_n961), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT109), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n866), .A2(new_n973), .A3(new_n965), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n975), .A2(new_n913), .A3(new_n915), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n971), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(new_n942), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT43), .ZN(new_n979));
  AND2_X1   g554(.A1(new_n963), .A2(new_n966), .ZN(new_n980));
  AND3_X1   g555(.A1(new_n914), .A2(new_n911), .A3(new_n967), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n942), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  OAI211_X1 g557(.A(new_n974), .B(new_n972), .C1(new_n921), .C2(new_n919), .ZN(new_n983));
  AOI21_X1  g558(.A(G37), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  AND3_X1   g559(.A1(new_n978), .A2(new_n979), .A3(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(new_n919), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n914), .A2(new_n920), .A3(new_n911), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n975), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  AND2_X1   g563(.A1(new_n980), .A2(new_n981), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n942), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n979), .B1(new_n990), .B2(new_n984), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n954), .B1(new_n985), .B2(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n990), .A2(new_n984), .A3(new_n979), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n979), .B1(new_n978), .B2(new_n984), .ZN(new_n994));
  OAI211_X1 g569(.A(KEYINPUT44), .B(new_n993), .C1(new_n994), .C2(KEYINPUT111), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT111), .ZN(new_n996));
  AOI211_X1 g571(.A(new_n996), .B(new_n979), .C1(new_n978), .C2(new_n984), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n992), .B1(new_n995), .B2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT112), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  OAI211_X1 g575(.A(new_n992), .B(KEYINPUT112), .C1(new_n995), .C2(new_n997), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(G397));
  INV_X1    g577(.A(G40), .ZN(new_n1003));
  AOI211_X1 g578(.A(new_n1003), .B(new_n464), .C1(new_n471), .C2(G2105), .ZN(new_n1004));
  AOI21_X1  g579(.A(G1384), .B1(new_n491), .B2(new_n498), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(G1976), .ZN(new_n1007));
  OAI211_X1 g582(.A(G8), .B(new_n1006), .C1(G288), .C2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(KEYINPUT52), .ZN(new_n1009));
  AOI21_X1  g584(.A(G1976), .B1(new_n576), .B2(new_n584), .ZN(new_n1010));
  OR2_X1    g585(.A1(new_n1010), .A2(KEYINPUT52), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1009), .B1(new_n1008), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1006), .A2(G8), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT117), .ZN(new_n1014));
  XOR2_X1   g589(.A(KEYINPUT116), .B(G1981), .Z(new_n1015));
  NOR2_X1   g590(.A1(G305), .A2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n597), .B1(G86), .B2(new_n525), .ZN(new_n1017));
  INV_X1    g592(.A(G1981), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1014), .B1(new_n1016), .B2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1013), .B1(new_n1020), .B2(KEYINPUT49), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT49), .ZN(new_n1022));
  OAI211_X1 g597(.A(new_n1014), .B(new_n1022), .C1(new_n1016), .C2(new_n1019), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1012), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(G303), .A2(G8), .ZN(new_n1025));
  XNOR2_X1  g600(.A(new_n1025), .B(KEYINPUT55), .ZN(new_n1026));
  NAND2_X1  g601(.A1(G160), .A2(G40), .ZN(new_n1027));
  INV_X1    g602(.A(G1384), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n499), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT45), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1027), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  XNOR2_X1  g606(.A(KEYINPUT113), .B(G1384), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n499), .A2(KEYINPUT45), .A3(new_n1032), .ZN(new_n1033));
  AOI21_X1  g608(.A(G1971), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT50), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1005), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1036), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1004), .B1(new_n1005), .B2(new_n1035), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1034), .B1(new_n773), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(G8), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1026), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1026), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1039), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n1044), .A2(G2090), .ZN(new_n1045));
  OAI211_X1 g620(.A(G8), .B(new_n1043), .C1(new_n1045), .C2(new_n1034), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1004), .B1(new_n1005), .B2(KEYINPUT45), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n759), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1029), .A2(KEYINPUT50), .ZN(new_n1050));
  INV_X1    g625(.A(G2084), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1050), .A2(new_n1051), .A3(new_n1004), .A4(new_n1036), .ZN(new_n1052));
  AOI211_X1 g627(.A(new_n1041), .B(G286), .C1(new_n1049), .C2(new_n1052), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1024), .A2(new_n1042), .A3(new_n1046), .A4(new_n1053), .ZN(new_n1054));
  AND2_X1   g629(.A1(new_n1054), .A2(KEYINPUT118), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT63), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1056), .B1(new_n1054), .B2(KEYINPUT118), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1024), .A2(new_n1042), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(KEYINPUT119), .ZN(new_n1059));
  AND3_X1   g634(.A1(new_n1046), .A2(KEYINPUT63), .A3(new_n1053), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1058), .A2(KEYINPUT119), .ZN(new_n1062));
  OAI22_X1  g637(.A1(new_n1055), .A2(new_n1057), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  XNOR2_X1  g638(.A(KEYINPUT120), .B(KEYINPUT56), .ZN(new_n1064));
  XNOR2_X1  g639(.A(new_n1064), .B(G2072), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1031), .A2(new_n1033), .A3(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(G1956), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1067), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1068));
  OR2_X1    g643(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1069));
  NAND2_X1  g644(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1066), .A2(new_n1068), .A3(new_n1069), .A4(new_n1070), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n778), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT121), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1004), .A2(new_n1005), .A3(new_n792), .ZN(new_n1074));
  AND3_X1   g649(.A1(new_n1072), .A2(new_n1073), .A3(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1073), .B1(new_n1072), .B2(new_n1074), .ZN(new_n1076));
  NOR3_X1   g651(.A1(new_n1075), .A2(new_n1076), .A3(new_n616), .ZN(new_n1077));
  AOI22_X1  g652(.A1(new_n1068), .A2(new_n1066), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1071), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(KEYINPUT122), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT122), .ZN(new_n1081));
  OAI211_X1 g656(.A(new_n1081), .B(new_n1071), .C1(new_n1077), .C2(new_n1078), .ZN(new_n1082));
  NOR3_X1   g657(.A1(new_n1075), .A2(new_n1076), .A3(KEYINPUT60), .ZN(new_n1083));
  OAI21_X1  g658(.A(KEYINPUT60), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(new_n617), .ZN(new_n1085));
  OAI211_X1 g660(.A(KEYINPUT60), .B(new_n616), .C1(new_n1075), .C2(new_n1076), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1083), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  XNOR2_X1  g662(.A(KEYINPUT123), .B(G1996), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1031), .A2(new_n1033), .A3(new_n1089), .ZN(new_n1090));
  XOR2_X1   g665(.A(KEYINPUT58), .B(G1341), .Z(new_n1091));
  NAND2_X1  g666(.A1(new_n1006), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(new_n554), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(KEYINPUT124), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT59), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n553), .B1(new_n1090), .B2(new_n1092), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT124), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1096), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1095), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT61), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1071), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1101), .B1(new_n1102), .B2(new_n1078), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1094), .A2(KEYINPUT124), .A3(new_n1096), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1066), .A2(new_n1068), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1107), .A2(KEYINPUT61), .A3(new_n1071), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1100), .A2(new_n1103), .A3(new_n1104), .A4(new_n1108), .ZN(new_n1109));
  OAI211_X1 g684(.A(new_n1080), .B(new_n1082), .C1(new_n1087), .C2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1049), .A2(new_n1052), .ZN(new_n1111));
  OAI21_X1  g686(.A(G8), .B1(new_n1111), .B2(G286), .ZN(new_n1112));
  AOI21_X1  g687(.A(G168), .B1(new_n1049), .B2(new_n1052), .ZN(new_n1113));
  OAI21_X1  g688(.A(KEYINPUT51), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT51), .ZN(new_n1115));
  OAI211_X1 g690(.A(new_n1115), .B(G8), .C1(new_n1111), .C2(G286), .ZN(new_n1116));
  AND2_X1   g691(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1044), .A2(new_n796), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT53), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1119), .B1(new_n1120), .B2(G2078), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1031), .B1(new_n1030), .B2(new_n1029), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n757), .A2(KEYINPUT53), .ZN(new_n1123));
  OAI211_X1 g698(.A(new_n1118), .B(new_n1121), .C1(new_n1122), .C2(new_n1123), .ZN(new_n1124));
  XOR2_X1   g699(.A(G301), .B(KEYINPUT54), .Z(new_n1125));
  INV_X1    g700(.A(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(KEYINPUT45), .B1(new_n499), .B2(new_n1032), .ZN(new_n1128));
  NOR3_X1   g703(.A1(new_n1128), .A2(new_n1027), .A3(new_n1123), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1126), .B1(new_n1033), .B2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1130), .A2(new_n1121), .A3(new_n1118), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1127), .A2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1024), .A2(new_n1046), .A3(new_n1042), .ZN(new_n1133));
  NOR3_X1   g708(.A1(new_n1117), .A2(new_n1132), .A3(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1110), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1136));
  NOR2_X1   g711(.A1(G288), .A2(G1976), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1016), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1024), .ZN(new_n1139));
  OAI22_X1  g714(.A1(new_n1138), .A2(new_n1013), .B1(new_n1139), .B2(new_n1046), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT62), .ZN(new_n1141));
  AND3_X1   g716(.A1(new_n1114), .A2(new_n1141), .A3(new_n1116), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1141), .B1(new_n1114), .B2(new_n1116), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1124), .A2(G171), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1133), .A2(new_n1145), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1140), .B1(new_n1144), .B2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1063), .A2(new_n1135), .A3(new_n1147), .ZN(new_n1148));
  AND2_X1   g723(.A1(new_n1128), .A2(new_n1004), .ZN(new_n1149));
  XNOR2_X1  g724(.A(new_n739), .B(G1996), .ZN(new_n1150));
  XNOR2_X1  g725(.A(new_n788), .B(G2067), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1149), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  XNOR2_X1  g727(.A(new_n1152), .B(KEYINPUT114), .ZN(new_n1153));
  XNOR2_X1  g728(.A(new_n831), .B(new_n833), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1153), .B1(new_n1149), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1149), .ZN(new_n1156));
  XOR2_X1   g731(.A(G290), .B(G1986), .Z(new_n1157));
  OAI21_X1  g732(.A(new_n1155), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  XOR2_X1   g733(.A(new_n1158), .B(KEYINPUT115), .Z(new_n1159));
  NAND2_X1  g734(.A1(new_n1148), .A2(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(G1996), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1149), .A2(new_n1161), .ZN(new_n1162));
  XNOR2_X1  g737(.A(new_n1162), .B(KEYINPUT46), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1149), .B1(new_n1151), .B2(new_n739), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  XOR2_X1   g740(.A(new_n1165), .B(KEYINPUT47), .Z(new_n1166));
  NOR3_X1   g741(.A1(new_n1156), .A2(G1986), .A3(G290), .ZN(new_n1167));
  XOR2_X1   g742(.A(new_n1167), .B(KEYINPUT48), .Z(new_n1168));
  AOI21_X1  g743(.A(new_n1166), .B1(new_n1155), .B2(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT126), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n831), .A2(new_n833), .ZN(new_n1171));
  NOR2_X1   g746(.A1(new_n1153), .A2(new_n1171), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n788), .A2(G2067), .ZN(new_n1173));
  NOR2_X1   g748(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n1174), .A2(KEYINPUT125), .ZN(new_n1175));
  OAI221_X1 g750(.A(KEYINPUT125), .B1(G2067), .B2(new_n788), .C1(new_n1153), .C2(new_n1171), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1176), .A2(new_n1149), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1170), .B1(new_n1175), .B2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1169), .A2(new_n1178), .ZN(new_n1179));
  NOR3_X1   g754(.A1(new_n1175), .A2(new_n1177), .A3(new_n1170), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1160), .A2(new_n1181), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g757(.A(G319), .ZN(new_n1184));
  NOR3_X1   g758(.A1(G401), .A2(new_n1184), .A3(G227), .ZN(new_n1185));
  OAI21_X1  g759(.A(new_n1185), .B1(new_n703), .B2(new_n704), .ZN(new_n1186));
  XNOR2_X1  g760(.A(new_n1186), .B(KEYINPUT127), .ZN(new_n1187));
  OR2_X1    g761(.A1(new_n985), .A2(new_n991), .ZN(new_n1188));
  NAND3_X1  g762(.A1(new_n902), .A2(new_n1187), .A3(new_n1188), .ZN(G225));
  INV_X1    g763(.A(G225), .ZN(G308));
endmodule


