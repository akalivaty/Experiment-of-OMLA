//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 0 1 0 0 1 0 0 1 0 0 1 0 0 0 1 1 1 0 1 1 0 0 1 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 1 1 1 0 0 0 0 1 1 1 1 0 1 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n698, new_n699, new_n700,
    new_n701, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n771, new_n772, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n782, new_n783, new_n784,
    new_n785, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n796, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n827, new_n828, new_n829, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n905, new_n906, new_n908, new_n909, new_n911, new_n912, new_n913,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n940, new_n941, new_n943, new_n944, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1017, new_n1018;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT16), .ZN(new_n203));
  OAI21_X1  g002(.A(new_n202), .B1(new_n203), .B2(G1gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n204), .B1(G1gat), .B2(new_n202), .ZN(new_n205));
  OR2_X1    g004(.A1(new_n205), .A2(G8gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(G8gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT21), .ZN(new_n208));
  XOR2_X1   g007(.A(G57gat), .B(G64gat), .Z(new_n209));
  INV_X1    g008(.A(KEYINPUT9), .ZN(new_n210));
  INV_X1    g009(.A(G71gat), .ZN(new_n211));
  INV_X1    g010(.A(G78gat), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n210), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n209), .A2(new_n213), .ZN(new_n214));
  XOR2_X1   g013(.A(G71gat), .B(G78gat), .Z(new_n215));
  XNOR2_X1  g014(.A(new_n214), .B(new_n215), .ZN(new_n216));
  OAI211_X1 g015(.A(new_n206), .B(new_n207), .C1(new_n208), .C2(new_n216), .ZN(new_n217));
  AND2_X1   g016(.A1(new_n217), .A2(KEYINPUT92), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n217), .A2(KEYINPUT92), .ZN(new_n219));
  XNOR2_X1  g018(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n220));
  OR3_X1    g019(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n220), .B1(new_n218), .B2(new_n219), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n216), .A2(new_n208), .ZN(new_n224));
  NAND2_X1  g023(.A1(G231gat), .A2(G233gat), .ZN(new_n225));
  INV_X1    g024(.A(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n224), .B(new_n226), .ZN(new_n227));
  XNOR2_X1  g026(.A(G127gat), .B(G155gat), .ZN(new_n228));
  XOR2_X1   g027(.A(new_n228), .B(KEYINPUT20), .Z(new_n229));
  NAND2_X1  g028(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(new_n224), .B(new_n225), .ZN(new_n231));
  INV_X1    g030(.A(new_n229), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  XOR2_X1   g032(.A(G183gat), .B(G211gat), .Z(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n230), .A2(new_n233), .A3(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n235), .B1(new_n230), .B2(new_n233), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n223), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n230), .A2(new_n233), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(new_n234), .ZN(new_n241));
  NAND4_X1  g040(.A1(new_n241), .A2(new_n221), .A3(new_n222), .A4(new_n236), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n239), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT96), .ZN(new_n244));
  XNOR2_X1  g043(.A(KEYINPUT94), .B(G92gat), .ZN(new_n245));
  INV_X1    g044(.A(G85gat), .ZN(new_n246));
  NAND2_X1  g045(.A1(G99gat), .A2(G106gat), .ZN(new_n247));
  AOI22_X1  g046(.A1(new_n245), .A2(new_n246), .B1(KEYINPUT8), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(G85gat), .A2(G92gat), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n249), .B(KEYINPUT7), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  XNOR2_X1  g050(.A(G99gat), .B(G106gat), .ZN(new_n252));
  XNOR2_X1  g051(.A(new_n252), .B(KEYINPUT95), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n251), .A2(new_n253), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n244), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  OR2_X1    g056(.A1(new_n251), .A2(new_n253), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n258), .A2(new_n254), .A3(KEYINPUT96), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  XNOR2_X1  g059(.A(KEYINPUT14), .B(G29gat), .ZN(new_n261));
  INV_X1    g060(.A(G36gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(G43gat), .B(G50gat), .ZN(new_n264));
  INV_X1    g063(.A(G29gat), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n265), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n266));
  NAND4_X1  g065(.A1(new_n263), .A2(KEYINPUT15), .A3(new_n264), .A4(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(new_n267), .B(KEYINPUT87), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT17), .ZN(new_n269));
  XOR2_X1   g068(.A(new_n264), .B(KEYINPUT15), .Z(new_n270));
  NAND2_X1  g069(.A1(new_n263), .A2(new_n266), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  AND3_X1   g071(.A1(new_n268), .A2(new_n269), .A3(new_n272), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n269), .B1(new_n268), .B2(new_n272), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n260), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n268), .A2(new_n272), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n276), .A2(new_n257), .A3(new_n259), .ZN(new_n277));
  NAND2_X1  g076(.A1(G232gat), .A2(G233gat), .ZN(new_n278));
  XOR2_X1   g077(.A(new_n278), .B(KEYINPUT93), .Z(new_n279));
  INV_X1    g078(.A(KEYINPUT41), .ZN(new_n280));
  OR2_X1    g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n275), .A2(new_n277), .A3(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(G190gat), .B(G218gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(KEYINPUT97), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n279), .A2(new_n280), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n286), .B(G134gat), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n287), .B(G162gat), .ZN(new_n288));
  INV_X1    g087(.A(new_n283), .ZN(new_n289));
  NAND4_X1  g088(.A1(new_n275), .A2(new_n289), .A3(new_n277), .A4(new_n281), .ZN(new_n290));
  AOI22_X1  g089(.A1(new_n285), .A2(new_n288), .B1(new_n284), .B2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT97), .ZN(new_n292));
  NAND4_X1  g091(.A1(new_n284), .A2(new_n292), .A3(new_n290), .A4(new_n288), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n243), .B1(new_n291), .B2(new_n294), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n216), .B1(new_n255), .B2(new_n256), .ZN(new_n296));
  INV_X1    g095(.A(new_n215), .ZN(new_n297));
  XNOR2_X1  g096(.A(new_n214), .B(new_n297), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n258), .A2(new_n254), .A3(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT10), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n296), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n216), .A2(new_n300), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n257), .A2(new_n259), .A3(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(G230gat), .A2(G233gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n296), .A2(new_n299), .ZN(new_n307));
  INV_X1    g106(.A(new_n305), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  XNOR2_X1  g108(.A(G120gat), .B(G148gat), .ZN(new_n310));
  XNOR2_X1  g109(.A(G176gat), .B(G204gat), .ZN(new_n311));
  XOR2_X1   g110(.A(new_n310), .B(new_n311), .Z(new_n312));
  NAND3_X1  g111(.A1(new_n306), .A2(new_n309), .A3(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT98), .ZN(new_n314));
  OR2_X1    g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n313), .A2(new_n314), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n306), .A2(new_n309), .ZN(new_n318));
  INV_X1    g117(.A(new_n312), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n317), .A2(new_n320), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n295), .A2(new_n321), .ZN(new_n322));
  XNOR2_X1  g121(.A(G113gat), .B(G141gat), .ZN(new_n323));
  XNOR2_X1  g122(.A(new_n323), .B(G197gat), .ZN(new_n324));
  XOR2_X1   g123(.A(KEYINPUT11), .B(G169gat), .Z(new_n325));
  XNOR2_X1  g124(.A(new_n324), .B(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n326), .B(KEYINPUT12), .ZN(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n206), .A2(new_n207), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n330), .B1(new_n273), .B2(new_n274), .ZN(new_n331));
  NAND2_X1  g130(.A1(G229gat), .A2(G233gat), .ZN(new_n332));
  XOR2_X1   g131(.A(new_n332), .B(KEYINPUT88), .Z(new_n333));
  AOI22_X1  g132(.A1(new_n268), .A2(new_n272), .B1(new_n206), .B2(new_n207), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n331), .A2(new_n333), .A3(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT18), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(KEYINPUT89), .ZN(new_n339));
  XOR2_X1   g138(.A(new_n333), .B(KEYINPUT13), .Z(new_n340));
  NOR2_X1   g139(.A1(new_n276), .A2(new_n329), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n340), .B1(new_n341), .B2(new_n334), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT89), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n336), .A2(new_n343), .A3(new_n337), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n339), .A2(new_n342), .A3(new_n344), .ZN(new_n345));
  NAND4_X1  g144(.A1(new_n331), .A2(KEYINPUT18), .A3(new_n333), .A4(new_n335), .ZN(new_n346));
  AND2_X1   g145(.A1(new_n346), .A2(KEYINPUT90), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n346), .A2(KEYINPUT90), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n328), .B1(new_n345), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n342), .A2(new_n327), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n351), .B1(new_n337), .B2(new_n336), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n352), .B1(new_n347), .B2(new_n348), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n350), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n322), .A2(new_n354), .ZN(new_n355));
  XNOR2_X1  g154(.A(KEYINPUT82), .B(G22gat), .ZN(new_n356));
  NAND2_X1  g155(.A1(G228gat), .A2(G233gat), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  XNOR2_X1  g157(.A(G78gat), .B(G106gat), .ZN(new_n359));
  AND2_X1   g158(.A1(G155gat), .A2(G162gat), .ZN(new_n360));
  NOR2_X1   g159(.A1(G155gat), .A2(G162gat), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  XNOR2_X1  g161(.A(G141gat), .B(G148gat), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT2), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n364), .B1(G155gat), .B2(G162gat), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n362), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(G141gat), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(G148gat), .ZN(new_n368));
  INV_X1    g167(.A(G148gat), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(G141gat), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  XNOR2_X1  g170(.A(G155gat), .B(G162gat), .ZN(new_n372));
  INV_X1    g171(.A(G155gat), .ZN(new_n373));
  INV_X1    g172(.A(G162gat), .ZN(new_n374));
  OAI21_X1  g173(.A(KEYINPUT2), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n371), .A2(new_n372), .A3(new_n375), .ZN(new_n376));
  AND2_X1   g175(.A1(new_n366), .A2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT29), .ZN(new_n378));
  AND2_X1   g177(.A1(G211gat), .A2(G218gat), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n379), .A2(KEYINPUT22), .ZN(new_n380));
  NOR2_X1   g179(.A1(G211gat), .A2(G218gat), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(G204gat), .ZN(new_n383));
  AND2_X1   g182(.A1(KEYINPUT74), .A2(G197gat), .ZN(new_n384));
  NOR2_X1   g183(.A1(KEYINPUT74), .A2(G197gat), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n383), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT74), .ZN(new_n387));
  INV_X1    g186(.A(G197gat), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(KEYINPUT74), .A2(G197gat), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n389), .A2(G204gat), .A3(new_n390), .ZN(new_n391));
  AOI211_X1 g190(.A(new_n380), .B(new_n382), .C1(new_n386), .C2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(new_n382), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n386), .A2(new_n391), .ZN(new_n394));
  INV_X1    g193(.A(new_n380), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n393), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n378), .B1(new_n392), .B2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT3), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n377), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n366), .A2(new_n376), .A3(new_n398), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(new_n378), .ZN(new_n401));
  NOR3_X1   g200(.A1(new_n384), .A2(new_n385), .A3(new_n383), .ZN(new_n402));
  AOI21_X1  g201(.A(G204gat), .B1(new_n389), .B2(new_n390), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n395), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(new_n382), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n394), .A2(new_n393), .A3(new_n395), .ZN(new_n406));
  AND3_X1   g205(.A1(new_n401), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n359), .B1(new_n399), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n366), .A2(new_n376), .ZN(new_n409));
  AOI21_X1  g208(.A(KEYINPUT29), .B1(new_n405), .B2(new_n406), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n409), .B1(new_n410), .B2(KEYINPUT3), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n392), .A2(new_n396), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(new_n401), .ZN(new_n413));
  INV_X1    g212(.A(new_n359), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n411), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  XNOR2_X1  g214(.A(KEYINPUT31), .B(G50gat), .ZN(new_n416));
  AND3_X1   g215(.A1(new_n408), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n416), .B1(new_n408), .B2(new_n415), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n358), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(new_n416), .ZN(new_n420));
  NOR3_X1   g219(.A1(new_n399), .A2(new_n407), .A3(new_n359), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n414), .B1(new_n411), .B2(new_n413), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n420), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n408), .A2(new_n415), .A3(new_n416), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n423), .A2(new_n357), .A3(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n356), .B1(new_n419), .B2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n419), .A2(new_n425), .A3(new_n356), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(G227gat), .A2(G233gat), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT27), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(G183gat), .ZN(new_n433));
  INV_X1    g232(.A(G183gat), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(KEYINPUT27), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT69), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n433), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n436), .B1(new_n433), .B2(new_n435), .ZN(new_n439));
  INV_X1    g238(.A(G190gat), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(KEYINPUT28), .ZN(new_n441));
  NOR3_X1   g240(.A1(new_n438), .A2(new_n439), .A3(new_n441), .ZN(new_n442));
  XNOR2_X1  g241(.A(KEYINPUT68), .B(KEYINPUT28), .ZN(new_n443));
  INV_X1    g242(.A(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n433), .A2(new_n435), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(KEYINPUT67), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT67), .ZN(new_n447));
  AOI21_X1  g246(.A(G190gat), .B1(new_n433), .B2(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n444), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  OAI21_X1  g248(.A(KEYINPUT70), .B1(new_n442), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n445), .A2(KEYINPUT69), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n451), .A2(new_n437), .A3(KEYINPUT28), .A4(new_n440), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n433), .A2(new_n447), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(new_n440), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n447), .B1(new_n433), .B2(new_n435), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n443), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT70), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n452), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(G169gat), .A2(G176gat), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT26), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NOR2_X1   g260(.A1(G169gat), .A2(G176gat), .ZN(new_n462));
  OR2_X1    g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  AOI22_X1  g262(.A1(new_n462), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n450), .A2(new_n458), .A3(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(G120gat), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(G113gat), .ZN(new_n469));
  INV_X1    g268(.A(G113gat), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(G120gat), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT1), .ZN(new_n473));
  INV_X1    g272(.A(G134gat), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(G127gat), .ZN(new_n475));
  INV_X1    g274(.A(G127gat), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(G134gat), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n472), .A2(new_n473), .A3(new_n475), .A4(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n475), .A2(new_n477), .ZN(new_n479));
  XNOR2_X1  g278(.A(G113gat), .B(G120gat), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n479), .B1(new_n480), .B2(KEYINPUT1), .ZN(new_n481));
  AND2_X1   g280(.A1(new_n478), .A2(new_n481), .ZN(new_n482));
  XNOR2_X1  g281(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n483));
  OAI21_X1  g282(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n484), .B1(new_n434), .B2(new_n440), .ZN(new_n485));
  NAND3_X1  g284(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n486));
  AND2_X1   g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n462), .A2(KEYINPUT23), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT23), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n489), .B1(G169gat), .B2(G176gat), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n488), .A2(new_n459), .A3(new_n490), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n483), .B1(new_n487), .B2(new_n491), .ZN(new_n492));
  NAND4_X1  g291(.A1(KEYINPUT65), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT65), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n486), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n485), .A2(new_n493), .A3(new_n495), .ZN(new_n496));
  AND3_X1   g295(.A1(new_n488), .A2(new_n459), .A3(new_n490), .ZN(new_n497));
  AND4_X1   g296(.A1(KEYINPUT66), .A2(new_n496), .A3(new_n497), .A4(KEYINPUT25), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT25), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n491), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g299(.A(KEYINPUT66), .B1(new_n500), .B2(new_n496), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n492), .B1(new_n498), .B2(new_n501), .ZN(new_n502));
  AND3_X1   g301(.A1(new_n467), .A2(new_n482), .A3(new_n502), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n482), .B1(new_n467), .B2(new_n502), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n431), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(KEYINPUT32), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT33), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  XNOR2_X1  g307(.A(KEYINPUT71), .B(G71gat), .ZN(new_n509));
  XNOR2_X1  g308(.A(new_n509), .B(G99gat), .ZN(new_n510));
  XOR2_X1   g309(.A(G15gat), .B(G43gat), .Z(new_n511));
  XOR2_X1   g310(.A(new_n510), .B(new_n511), .Z(new_n512));
  NAND3_X1  g311(.A1(new_n506), .A2(new_n508), .A3(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(new_n512), .ZN(new_n514));
  OAI211_X1 g313(.A(new_n505), .B(KEYINPUT32), .C1(new_n507), .C2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n467), .A2(new_n502), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n478), .A2(new_n481), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n467), .A2(new_n502), .A3(new_n482), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n518), .A2(new_n430), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(KEYINPUT34), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT34), .ZN(new_n522));
  NAND4_X1  g321(.A1(new_n518), .A2(new_n522), .A3(new_n430), .A4(new_n519), .ZN(new_n523));
  NAND4_X1  g322(.A1(new_n513), .A2(new_n515), .A3(new_n521), .A4(new_n523), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n503), .A2(new_n504), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n522), .B1(new_n525), .B2(new_n430), .ZN(new_n526));
  INV_X1    g325(.A(new_n523), .ZN(new_n527));
  OAI21_X1  g326(.A(KEYINPUT72), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT72), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n521), .A2(new_n529), .A3(new_n523), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n513), .A2(new_n515), .ZN(new_n532));
  AND3_X1   g331(.A1(new_n531), .A2(KEYINPUT73), .A3(new_n532), .ZN(new_n533));
  AOI21_X1  g332(.A(KEYINPUT73), .B1(new_n531), .B2(new_n532), .ZN(new_n534));
  OAI211_X1 g333(.A(new_n429), .B(new_n524), .C1(new_n533), .C2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n409), .A2(KEYINPUT3), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n536), .A2(new_n517), .A3(new_n400), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT76), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  AOI22_X1  g338(.A1(new_n409), .A2(KEYINPUT3), .B1(new_n478), .B2(new_n481), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n540), .A2(KEYINPUT76), .A3(new_n400), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT5), .ZN(new_n543));
  NAND2_X1  g342(.A1(G225gat), .A2(G233gat), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n542), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT77), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n482), .A2(new_n377), .A3(new_n547), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n478), .A2(new_n481), .A3(new_n366), .A4(new_n376), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(KEYINPUT77), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n548), .A2(new_n550), .A3(KEYINPUT4), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT79), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n552), .B1(new_n549), .B2(KEYINPUT4), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  NAND4_X1  g353(.A1(new_n548), .A2(new_n550), .A3(new_n552), .A4(KEYINPUT4), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(KEYINPUT80), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT80), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n554), .A2(new_n558), .A3(new_n555), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n546), .A2(new_n557), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n517), .A2(new_n409), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n548), .A2(new_n550), .A3(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n544), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n564), .A2(KEYINPUT5), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(KEYINPUT78), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT78), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n564), .A2(new_n567), .A3(KEYINPUT5), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n482), .A2(new_n377), .A3(KEYINPUT4), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT4), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n548), .A2(new_n550), .A3(new_n570), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n542), .A2(new_n544), .A3(new_n569), .A4(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n566), .A2(new_n568), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n560), .A2(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(G1gat), .B(G29gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n575), .B(KEYINPUT0), .ZN(new_n576));
  XNOR2_X1  g375(.A(G57gat), .B(G85gat), .ZN(new_n577));
  XOR2_X1   g376(.A(new_n576), .B(new_n577), .Z(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n574), .A2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT6), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n560), .A2(new_n573), .A3(new_n578), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  AND4_X1   g382(.A1(KEYINPUT81), .A2(new_n574), .A3(KEYINPUT6), .A4(new_n579), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n578), .B1(new_n560), .B2(new_n573), .ZN(new_n585));
  AOI21_X1  g384(.A(KEYINPUT81), .B1(new_n585), .B2(KEYINPUT6), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n583), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(G226gat), .ZN(new_n588));
  INV_X1    g387(.A(G233gat), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n452), .A2(new_n456), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n465), .B1(new_n592), .B2(KEYINPUT70), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n496), .A2(new_n497), .A3(KEYINPUT25), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT66), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n500), .A2(KEYINPUT66), .A3(new_n496), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  AOI22_X1  g397(.A1(new_n593), .A2(new_n458), .B1(new_n598), .B2(new_n492), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n591), .B1(new_n599), .B2(KEYINPUT29), .ZN(new_n600));
  INV_X1    g399(.A(new_n412), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n516), .A2(new_n590), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n600), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n590), .B1(new_n516), .B2(new_n378), .ZN(new_n604));
  OAI21_X1  g403(.A(KEYINPUT75), .B1(new_n599), .B2(new_n591), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT75), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n516), .A2(new_n606), .A3(new_n590), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n604), .B1(new_n605), .B2(new_n607), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n603), .B1(new_n608), .B2(new_n601), .ZN(new_n609));
  XNOR2_X1  g408(.A(G8gat), .B(G36gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(G64gat), .B(G92gat), .ZN(new_n611));
  XOR2_X1   g410(.A(new_n610), .B(new_n611), .Z(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n609), .A2(new_n613), .ZN(new_n614));
  OAI211_X1 g413(.A(new_n603), .B(new_n612), .C1(new_n608), .C2(new_n601), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n614), .A2(KEYINPUT30), .A3(new_n615), .ZN(new_n616));
  OR3_X1    g415(.A1(new_n609), .A2(KEYINPUT30), .A3(new_n613), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n587), .A2(new_n618), .ZN(new_n619));
  OAI21_X1  g418(.A(KEYINPUT35), .B1(new_n535), .B2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT86), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  OAI211_X1 g421(.A(KEYINPUT86), .B(KEYINPUT35), .C1(new_n535), .C2(new_n619), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n537), .A2(new_n538), .ZN(new_n624));
  AOI21_X1  g423(.A(KEYINPUT76), .B1(new_n540), .B2(new_n400), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n544), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n571), .A2(new_n569), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  AOI211_X1 g427(.A(KEYINPUT78), .B(new_n543), .C1(new_n562), .C2(new_n563), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n567), .B1(new_n564), .B2(KEYINPUT5), .ZN(new_n630));
  NOR3_X1   g429(.A1(new_n628), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  AND3_X1   g430(.A1(new_n554), .A2(new_n558), .A3(new_n555), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n558), .B1(new_n554), .B2(new_n555), .ZN(new_n633));
  NOR3_X1   g432(.A1(new_n632), .A2(new_n633), .A3(new_n545), .ZN(new_n634));
  OAI211_X1 g433(.A(KEYINPUT6), .B(new_n579), .C1(new_n631), .C2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT81), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n585), .A2(KEYINPUT81), .A3(KEYINPUT6), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  AOI22_X1  g438(.A1(new_n639), .A2(new_n583), .B1(new_n617), .B2(new_n616), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT35), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n521), .A2(new_n523), .ZN(new_n642));
  XOR2_X1   g441(.A(new_n532), .B(new_n642), .Z(new_n643));
  NAND4_X1  g442(.A1(new_n640), .A2(new_n641), .A3(new_n429), .A4(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n622), .A2(new_n623), .A3(new_n644), .ZN(new_n645));
  OAI211_X1 g444(.A(KEYINPUT36), .B(new_n524), .C1(new_n533), .C2(new_n534), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n646), .B1(new_n643), .B2(KEYINPUT36), .ZN(new_n647));
  INV_X1    g446(.A(new_n429), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n619), .A2(new_n648), .ZN(new_n649));
  AND2_X1   g448(.A1(new_n609), .A2(KEYINPUT37), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n613), .B1(new_n609), .B2(KEYINPUT37), .ZN(new_n651));
  OAI21_X1  g450(.A(KEYINPUT38), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n605), .A2(new_n607), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n653), .A2(new_n601), .A3(new_n600), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT84), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n600), .A2(new_n602), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n657), .A2(new_n412), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n658), .A2(KEYINPUT85), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n608), .A2(KEYINPUT84), .A3(new_n601), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT85), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n657), .A2(new_n661), .A3(new_n412), .ZN(new_n662));
  NAND4_X1  g461(.A1(new_n656), .A2(new_n659), .A3(new_n660), .A4(new_n662), .ZN(new_n663));
  AND2_X1   g462(.A1(new_n663), .A2(KEYINPUT37), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT38), .ZN(new_n665));
  OAI211_X1 g464(.A(new_n665), .B(new_n613), .C1(new_n609), .C2(KEYINPUT37), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n652), .B1(new_n664), .B2(new_n666), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n639), .A2(new_n583), .A3(new_n615), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT40), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n557), .A2(new_n559), .A3(new_n542), .ZN(new_n671));
  XOR2_X1   g470(.A(KEYINPUT83), .B(KEYINPUT39), .Z(new_n672));
  NAND3_X1  g471(.A1(new_n671), .A2(new_n563), .A3(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n673), .A2(new_n578), .ZN(new_n674));
  OR2_X1    g473(.A1(new_n562), .A2(new_n563), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(KEYINPUT39), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n676), .B1(new_n671), .B2(new_n563), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n670), .B1(new_n674), .B2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n677), .ZN(new_n679));
  NAND4_X1  g478(.A1(new_n679), .A2(KEYINPUT40), .A3(new_n578), .A4(new_n673), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n678), .A2(new_n680), .A3(new_n580), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n429), .B1(new_n681), .B2(new_n618), .ZN(new_n682));
  OAI211_X1 g481(.A(new_n647), .B(new_n649), .C1(new_n669), .C2(new_n682), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n355), .B1(new_n645), .B2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n587), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n686), .B(G1gat), .ZN(G1324gat));
  INV_X1    g486(.A(new_n618), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n684), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(G8gat), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT42), .ZN(new_n691));
  NAND2_X1  g490(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n692));
  OR2_X1    g491(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n693));
  NAND4_X1  g492(.A1(new_n684), .A2(new_n688), .A3(new_n692), .A4(new_n693), .ZN(new_n694));
  AND3_X1   g493(.A1(new_n694), .A2(KEYINPUT99), .A3(new_n691), .ZN(new_n695));
  AOI21_X1  g494(.A(KEYINPUT99), .B1(new_n694), .B2(new_n691), .ZN(new_n696));
  OAI221_X1 g495(.A(new_n690), .B1(new_n691), .B2(new_n694), .C1(new_n695), .C2(new_n696), .ZN(G1325gat));
  AOI21_X1  g496(.A(G15gat), .B1(new_n684), .B2(new_n643), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(KEYINPUT100), .ZN(new_n699));
  INV_X1    g498(.A(new_n647), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n684), .A2(G15gat), .A3(new_n700), .ZN(new_n701));
  AND2_X1   g500(.A1(new_n699), .A2(new_n701), .ZN(G1326gat));
  XNOR2_X1  g501(.A(KEYINPUT43), .B(G22gat), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n684), .A2(new_n648), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT101), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n705), .B(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT102), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n707), .A2(new_n708), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n704), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  OR2_X1    g511(.A1(new_n707), .A2(new_n708), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n713), .A2(new_n709), .A3(new_n703), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n712), .A2(new_n714), .ZN(G1327gat));
  NOR2_X1   g514(.A1(new_n291), .A2(new_n294), .ZN(new_n716));
  INV_X1    g515(.A(new_n716), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n717), .B1(new_n645), .B2(new_n683), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n344), .A2(new_n342), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n343), .B1(new_n336), .B2(new_n337), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n346), .B(KEYINPUT90), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n327), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(new_n353), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NOR3_X1   g524(.A1(new_n725), .A2(new_n243), .A3(new_n321), .ZN(new_n726));
  AND2_X1   g525(.A1(new_n718), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n727), .A2(new_n265), .A3(new_n685), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(KEYINPUT45), .ZN(new_n729));
  AND3_X1   g528(.A1(new_n419), .A2(new_n356), .A3(new_n425), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n524), .B1(new_n730), .B2(new_n426), .ZN(new_n731));
  AND3_X1   g530(.A1(new_n506), .A2(new_n508), .A3(new_n512), .ZN(new_n732));
  INV_X1    g531(.A(new_n515), .ZN(new_n733));
  AND3_X1   g532(.A1(new_n521), .A2(new_n529), .A3(new_n523), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n529), .B1(new_n521), .B2(new_n523), .ZN(new_n735));
  OAI22_X1  g534(.A1(new_n732), .A2(new_n733), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT73), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n531), .A2(KEYINPUT73), .A3(new_n532), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n731), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n641), .B1(new_n740), .B2(new_n640), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n644), .B1(new_n741), .B2(KEYINPUT86), .ZN(new_n742));
  INV_X1    g541(.A(new_n623), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n683), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT103), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n744), .A2(new_n745), .A3(new_n716), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT44), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND4_X1  g547(.A1(new_n744), .A2(new_n745), .A3(KEYINPUT44), .A4(new_n716), .ZN(new_n749));
  AND2_X1   g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n750), .A2(new_n685), .A3(new_n726), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(KEYINPUT104), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(G29gat), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n751), .A2(KEYINPUT104), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n729), .B1(new_n753), .B2(new_n754), .ZN(G1328gat));
  NAND4_X1  g554(.A1(new_n748), .A2(new_n688), .A3(new_n749), .A4(new_n726), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(G36gat), .ZN(new_n757));
  AOI211_X1 g556(.A(G36gat), .B(new_n618), .C1(KEYINPUT105), .C2(KEYINPUT46), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n718), .A2(new_n726), .A3(new_n758), .ZN(new_n759));
  NOR2_X1   g558(.A1(KEYINPUT105), .A2(KEYINPUT46), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n759), .B(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n757), .A2(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT106), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n762), .B(new_n763), .ZN(G1329gat));
  INV_X1    g563(.A(G43gat), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n647), .A2(new_n765), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n748), .A2(new_n749), .A3(new_n726), .A4(new_n766), .ZN(new_n767));
  AND2_X1   g566(.A1(new_n727), .A2(new_n643), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n767), .B1(new_n768), .B2(G43gat), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n769), .B(KEYINPUT47), .ZN(G1330gat));
  AND2_X1   g569(.A1(new_n648), .A2(G50gat), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n748), .A2(new_n749), .A3(new_n726), .A4(new_n771), .ZN(new_n772));
  AND2_X1   g571(.A1(new_n727), .A2(new_n648), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n772), .B1(new_n773), .B2(G50gat), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n774), .B(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g574(.A(new_n321), .ZN(new_n776));
  NOR3_X1   g575(.A1(new_n354), .A2(new_n776), .A3(new_n295), .ZN(new_n777));
  AND2_X1   g576(.A1(new_n744), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(new_n685), .ZN(new_n779));
  XOR2_X1   g578(.A(KEYINPUT107), .B(G57gat), .Z(new_n780));
  XNOR2_X1  g579(.A(new_n779), .B(new_n780), .ZN(G1332gat));
  XNOR2_X1  g580(.A(new_n618), .B(KEYINPUT108), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n782), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n778), .A2(new_n783), .ZN(new_n784));
  NOR2_X1   g583(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n785));
  XOR2_X1   g584(.A(new_n784), .B(new_n785), .Z(G1333gat));
  NAND3_X1  g585(.A1(new_n778), .A2(G71gat), .A3(new_n700), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n787), .B(KEYINPUT109), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n778), .A2(new_n643), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(new_n211), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(KEYINPUT50), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT50), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n788), .A2(new_n793), .A3(new_n790), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n792), .A2(new_n794), .ZN(G1334gat));
  NAND2_X1  g594(.A1(new_n778), .A2(new_n648), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g596(.A1(new_n354), .A2(new_n243), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n718), .A2(new_n798), .ZN(new_n799));
  XNOR2_X1  g598(.A(new_n799), .B(KEYINPUT51), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n800), .A2(new_n776), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n801), .A2(new_n246), .A3(new_n685), .ZN(new_n802));
  NOR3_X1   g601(.A1(new_n354), .A2(new_n243), .A3(new_n776), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n750), .A2(new_n803), .ZN(new_n804));
  OAI21_X1  g603(.A(G85gat), .B1(new_n804), .B2(new_n587), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n802), .A2(new_n805), .ZN(G1336gat));
  INV_X1    g605(.A(new_n782), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n748), .A2(new_n749), .A3(new_n807), .A4(new_n803), .ZN(new_n808));
  INV_X1    g607(.A(new_n245), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT52), .ZN(new_n811));
  NOR3_X1   g610(.A1(new_n782), .A2(G92gat), .A3(new_n776), .ZN(new_n812));
  INV_X1    g611(.A(new_n812), .ZN(new_n813));
  OAI211_X1 g612(.A(new_n810), .B(new_n811), .C1(new_n800), .C2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT51), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(KEYINPUT110), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n816), .B1(new_n718), .B2(new_n798), .ZN(new_n817));
  AND4_X1   g616(.A1(new_n744), .A2(new_n716), .A3(new_n798), .A4(new_n816), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n812), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(KEYINPUT111), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n748), .A2(new_n688), .A3(new_n749), .A4(new_n803), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(new_n809), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT111), .ZN(new_n823));
  OAI211_X1 g622(.A(new_n823), .B(new_n812), .C1(new_n817), .C2(new_n818), .ZN(new_n824));
  AND3_X1   g623(.A1(new_n820), .A2(new_n822), .A3(new_n824), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n814), .B1(new_n825), .B2(new_n811), .ZN(G1337gat));
  INV_X1    g625(.A(G99gat), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n801), .A2(new_n827), .A3(new_n643), .ZN(new_n828));
  OAI21_X1  g627(.A(G99gat), .B1(new_n804), .B2(new_n647), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(G1338gat));
  NAND4_X1  g629(.A1(new_n748), .A2(new_n648), .A3(new_n749), .A4(new_n803), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT113), .ZN(new_n832));
  XOR2_X1   g631(.A(KEYINPUT112), .B(G106gat), .Z(new_n833));
  NAND3_X1  g632(.A1(new_n831), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  NOR3_X1   g633(.A1(new_n776), .A2(new_n429), .A3(G106gat), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n835), .B1(new_n817), .B2(new_n818), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(KEYINPUT114), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT114), .ZN(new_n838));
  OAI211_X1 g637(.A(new_n838), .B(new_n835), .C1(new_n817), .C2(new_n818), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n834), .A2(new_n837), .A3(new_n839), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n832), .B1(new_n831), .B2(new_n833), .ZN(new_n841));
  OAI21_X1  g640(.A(KEYINPUT53), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n831), .A2(new_n833), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT53), .ZN(new_n844));
  INV_X1    g643(.A(new_n835), .ZN(new_n845));
  OAI211_X1 g644(.A(new_n843), .B(new_n844), .C1(new_n800), .C2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n842), .A2(new_n846), .ZN(G1339gat));
  NOR4_X1   g646(.A1(new_n354), .A2(new_n295), .A3(KEYINPUT115), .A4(new_n321), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT115), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n849), .B1(new_n322), .B2(new_n725), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT118), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n301), .A2(new_n303), .A3(new_n308), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n306), .A2(KEYINPUT54), .A3(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT54), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n304), .A2(new_n855), .A3(new_n305), .ZN(new_n856));
  AND3_X1   g655(.A1(new_n856), .A2(KEYINPUT116), .A3(new_n319), .ZN(new_n857));
  AOI21_X1  g656(.A(KEYINPUT116), .B1(new_n856), .B2(new_n319), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n854), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT55), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  OAI211_X1 g660(.A(KEYINPUT55), .B(new_n854), .C1(new_n857), .C2(new_n858), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n861), .A2(new_n317), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n284), .A2(new_n290), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n292), .B1(new_n282), .B2(new_n283), .ZN(new_n865));
  INV_X1    g664(.A(new_n288), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n864), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(new_n341), .ZN(new_n868));
  INV_X1    g667(.A(new_n340), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n868), .A2(new_n335), .A3(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT117), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND4_X1  g671(.A1(new_n868), .A2(KEYINPUT117), .A3(new_n335), .A4(new_n869), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n333), .B1(new_n331), .B2(new_n335), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n326), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND4_X1  g675(.A1(new_n867), .A2(new_n353), .A3(new_n876), .A4(new_n293), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n852), .B1(new_n863), .B2(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(new_n877), .ZN(new_n879));
  AND2_X1   g678(.A1(new_n317), .A2(new_n862), .ZN(new_n880));
  NAND4_X1  g679(.A1(new_n879), .A2(new_n880), .A3(KEYINPUT118), .A4(new_n861), .ZN(new_n881));
  INV_X1    g680(.A(new_n863), .ZN(new_n882));
  AND2_X1   g681(.A1(new_n353), .A2(new_n876), .ZN(new_n883));
  AOI22_X1  g682(.A1(new_n882), .A2(new_n354), .B1(new_n321), .B2(new_n883), .ZN(new_n884));
  OAI211_X1 g683(.A(new_n878), .B(new_n881), .C1(new_n884), .C2(new_n716), .ZN(new_n885));
  INV_X1    g684(.A(new_n243), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n851), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n887), .A2(new_n587), .A3(new_n535), .ZN(new_n888));
  AND2_X1   g687(.A1(new_n888), .A2(new_n782), .ZN(new_n889));
  AOI21_X1  g688(.A(G113gat), .B1(new_n889), .B2(new_n354), .ZN(new_n890));
  OAI21_X1  g689(.A(KEYINPUT119), .B1(new_n887), .B2(new_n648), .ZN(new_n891));
  OAI211_X1 g690(.A(new_n880), .B(new_n861), .C1(new_n723), .C2(new_n724), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n883), .A2(new_n321), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n716), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n881), .A2(new_n878), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n886), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  OR2_X1    g695(.A1(new_n848), .A2(new_n850), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT119), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n898), .A2(new_n899), .A3(new_n429), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n891), .A2(new_n900), .ZN(new_n901));
  AND4_X1   g700(.A1(new_n685), .A2(new_n901), .A3(new_n643), .A4(new_n782), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n725), .A2(new_n470), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n890), .B1(new_n902), .B2(new_n903), .ZN(G1340gat));
  AOI21_X1  g703(.A(G120gat), .B1(new_n889), .B2(new_n321), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n776), .A2(new_n468), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n905), .B1(new_n902), .B2(new_n906), .ZN(G1341gat));
  NAND3_X1  g706(.A1(new_n889), .A2(new_n476), .A3(new_n243), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n902), .A2(new_n243), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n908), .B1(new_n909), .B2(new_n476), .ZN(G1342gat));
  AOI21_X1  g709(.A(new_n474), .B1(new_n902), .B2(new_n716), .ZN(new_n911));
  NAND4_X1  g710(.A1(new_n888), .A2(new_n474), .A3(new_n618), .A4(new_n716), .ZN(new_n912));
  XNOR2_X1  g711(.A(new_n912), .B(KEYINPUT56), .ZN(new_n913));
  OR2_X1    g712(.A1(new_n911), .A2(new_n913), .ZN(G1343gat));
  NAND3_X1  g713(.A1(new_n782), .A2(new_n647), .A3(new_n685), .ZN(new_n915));
  XNOR2_X1  g714(.A(new_n915), .B(KEYINPUT120), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT57), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n917), .B1(new_n887), .B2(new_n429), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n898), .A2(KEYINPUT57), .A3(new_n648), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n916), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n367), .B1(new_n920), .B2(new_n354), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n700), .A2(new_n429), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n898), .A2(new_n685), .A3(new_n922), .ZN(new_n923));
  NOR4_X1   g722(.A1(new_n923), .A2(G141gat), .A3(new_n725), .A4(new_n807), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n921), .A2(new_n924), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT58), .ZN(new_n926));
  XNOR2_X1  g725(.A(new_n925), .B(new_n926), .ZN(G1344gat));
  NOR2_X1   g726(.A1(new_n923), .A2(new_n807), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n928), .A2(new_n369), .A3(new_n321), .ZN(new_n929));
  AOI211_X1 g728(.A(KEYINPUT59), .B(new_n369), .C1(new_n920), .C2(new_n321), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT59), .ZN(new_n931));
  OAI22_X1  g730(.A1(new_n884), .A2(new_n716), .B1(new_n863), .B2(new_n877), .ZN(new_n932));
  AOI22_X1  g731(.A1(new_n932), .A2(new_n886), .B1(new_n725), .B2(new_n322), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n917), .B1(new_n933), .B2(new_n429), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n934), .A2(new_n919), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n916), .A2(new_n776), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n931), .B1(new_n937), .B2(G148gat), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n929), .B1(new_n930), .B2(new_n938), .ZN(G1345gat));
  NAND3_X1  g738(.A1(new_n928), .A2(new_n373), .A3(new_n243), .ZN(new_n940));
  AND2_X1   g739(.A1(new_n920), .A2(new_n243), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n940), .B1(new_n941), .B2(new_n373), .ZN(G1346gat));
  AND2_X1   g741(.A1(new_n920), .A2(new_n716), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n618), .A2(new_n374), .A3(new_n716), .ZN(new_n944));
  OAI22_X1  g743(.A1(new_n943), .A2(new_n374), .B1(new_n923), .B2(new_n944), .ZN(G1347gat));
  INV_X1    g744(.A(KEYINPUT121), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n946), .B1(new_n887), .B2(new_n685), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n898), .A2(KEYINPUT121), .A3(new_n587), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n782), .A2(new_n535), .ZN(new_n950));
  AND2_X1   g749(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  AOI21_X1  g750(.A(G169gat), .B1(new_n951), .B2(new_n354), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n685), .A2(new_n618), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(new_n643), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n954), .B1(new_n891), .B2(new_n900), .ZN(new_n955));
  AND2_X1   g754(.A1(new_n354), .A2(G169gat), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n952), .B1(new_n955), .B2(new_n956), .ZN(G1348gat));
  INV_X1    g756(.A(G176gat), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n951), .A2(new_n958), .A3(new_n321), .ZN(new_n959));
  AND2_X1   g758(.A1(new_n955), .A2(new_n321), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n959), .B1(new_n960), .B2(new_n958), .ZN(G1349gat));
  INV_X1    g760(.A(new_n954), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n899), .B1(new_n898), .B2(new_n429), .ZN(new_n963));
  AOI211_X1 g762(.A(KEYINPUT119), .B(new_n648), .C1(new_n896), .C2(new_n897), .ZN(new_n964));
  OAI211_X1 g763(.A(new_n243), .B(new_n962), .C1(new_n963), .C2(new_n964), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT123), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND4_X1  g766(.A1(new_n901), .A2(KEYINPUT123), .A3(new_n243), .A4(new_n962), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n967), .A2(new_n968), .A3(G183gat), .ZN(new_n969));
  NOR3_X1   g768(.A1(new_n886), .A2(new_n439), .A3(new_n438), .ZN(new_n970));
  AOI21_X1  g769(.A(KEYINPUT121), .B1(new_n898), .B2(new_n587), .ZN(new_n971));
  AOI211_X1 g770(.A(new_n946), .B(new_n685), .C1(new_n896), .C2(new_n897), .ZN(new_n972));
  OAI211_X1 g771(.A(new_n950), .B(new_n970), .C1(new_n971), .C2(new_n972), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n973), .A2(KEYINPUT122), .ZN(new_n974));
  INV_X1    g773(.A(KEYINPUT122), .ZN(new_n975));
  NAND4_X1  g774(.A1(new_n949), .A2(new_n975), .A3(new_n950), .A4(new_n970), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n969), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n978), .A2(KEYINPUT60), .ZN(new_n979));
  INV_X1    g778(.A(KEYINPUT60), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n969), .A2(new_n977), .A3(new_n980), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n979), .A2(new_n981), .ZN(G1350gat));
  NAND3_X1  g781(.A1(new_n951), .A2(new_n440), .A3(new_n716), .ZN(new_n983));
  INV_X1    g782(.A(KEYINPUT61), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n955), .A2(new_n716), .ZN(new_n985));
  AOI21_X1  g784(.A(new_n984), .B1(new_n985), .B2(G190gat), .ZN(new_n986));
  AOI211_X1 g785(.A(KEYINPUT61), .B(new_n440), .C1(new_n955), .C2(new_n716), .ZN(new_n987));
  OAI21_X1  g786(.A(new_n983), .B1(new_n986), .B2(new_n987), .ZN(G1351gat));
  NAND2_X1  g787(.A1(new_n922), .A2(new_n807), .ZN(new_n989));
  AOI21_X1  g788(.A(new_n989), .B1(new_n947), .B2(new_n948), .ZN(new_n990));
  XOR2_X1   g789(.A(KEYINPUT124), .B(G197gat), .Z(new_n991));
  NAND3_X1  g790(.A1(new_n990), .A2(new_n354), .A3(new_n991), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n647), .A2(new_n953), .ZN(new_n993));
  INV_X1    g792(.A(new_n993), .ZN(new_n994));
  OR2_X1    g793(.A1(new_n994), .A2(KEYINPUT125), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n994), .A2(KEYINPUT125), .ZN(new_n996));
  AND3_X1   g795(.A1(new_n935), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  AND2_X1   g796(.A1(new_n997), .A2(new_n354), .ZN(new_n998));
  OAI21_X1  g797(.A(new_n992), .B1(new_n998), .B2(new_n991), .ZN(G1352gat));
  NAND4_X1  g798(.A1(new_n935), .A2(new_n321), .A3(new_n995), .A4(new_n996), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n1000), .A2(G204gat), .ZN(new_n1001));
  NOR2_X1   g800(.A1(new_n776), .A2(G204gat), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n990), .A2(new_n1002), .ZN(new_n1003));
  AND3_X1   g802(.A1(new_n1003), .A2(KEYINPUT126), .A3(KEYINPUT62), .ZN(new_n1004));
  AOI21_X1  g803(.A(KEYINPUT126), .B1(new_n1003), .B2(KEYINPUT62), .ZN(new_n1005));
  OAI221_X1 g804(.A(new_n1001), .B1(KEYINPUT62), .B2(new_n1003), .C1(new_n1004), .C2(new_n1005), .ZN(G1353gat));
  INV_X1    g805(.A(G211gat), .ZN(new_n1007));
  NAND3_X1  g806(.A1(new_n990), .A2(new_n1007), .A3(new_n243), .ZN(new_n1008));
  NAND2_X1  g807(.A1(new_n994), .A2(new_n243), .ZN(new_n1009));
  AOI21_X1  g808(.A(new_n1009), .B1(new_n934), .B2(new_n919), .ZN(new_n1010));
  INV_X1    g809(.A(KEYINPUT127), .ZN(new_n1011));
  OR2_X1    g810(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g811(.A(new_n1007), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1013));
  AND3_X1   g812(.A1(new_n1012), .A2(KEYINPUT63), .A3(new_n1013), .ZN(new_n1014));
  AOI21_X1  g813(.A(KEYINPUT63), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1015));
  OAI21_X1  g814(.A(new_n1008), .B1(new_n1014), .B2(new_n1015), .ZN(G1354gat));
  AOI21_X1  g815(.A(G218gat), .B1(new_n990), .B2(new_n716), .ZN(new_n1017));
  AND2_X1   g816(.A1(new_n716), .A2(G218gat), .ZN(new_n1018));
  AOI21_X1  g817(.A(new_n1017), .B1(new_n997), .B2(new_n1018), .ZN(G1355gat));
endmodule


