//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 0 1 1 1 1 0 1 0 1 0 0 0 1 0 0 0 0 0 1 1 1 1 0 0 1 0 0 1 1 1 1 0 1 0 1 1 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 1 1 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:53 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n448, new_n450, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n529, new_n530, new_n531, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n551, new_n552,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n596, new_n597, new_n598, new_n601, new_n602, new_n604, new_n605,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT65), .B(G69), .Z(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g021(.A(KEYINPUT66), .B(G452), .ZN(G391));
  NAND2_X1  g022(.A1(G94), .A2(G452), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT67), .Z(G173));
  NAND2_X1  g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g026(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g027(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT2), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR4_X1   g031(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n456), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  AOI22_X1  g035(.A1(new_n456), .A2(G2106), .B1(G567), .B2(new_n458), .ZN(G319));
  AND2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  INV_X1    g042(.A(new_n467), .ZN(new_n468));
  AOI22_X1  g043(.A1(new_n465), .A2(G137), .B1(G101), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  INV_X1    g045(.A(G125), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n470), .B1(new_n464), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n469), .A2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(G160));
  NAND2_X1  g050(.A1(new_n465), .A2(G136), .ZN(new_n476));
  INV_X1    g051(.A(new_n463), .ZN(new_n477));
  NAND2_X1  g052(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n466), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  OR2_X1    g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n481), .B(G2104), .C1(G112), .C2(new_n466), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n476), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G162));
  XNOR2_X1  g059(.A(KEYINPUT3), .B(G2104), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G2105), .ZN(new_n486));
  INV_X1    g061(.A(G126), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n466), .A2(G114), .ZN(new_n488));
  OAI21_X1  g063(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n489));
  OAI22_X1  g064(.A1(new_n486), .A2(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n491), .A2(new_n466), .A3(G138), .ZN(new_n492));
  NOR3_X1   g067(.A1(new_n464), .A2(KEYINPUT68), .A3(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT68), .ZN(new_n494));
  AND3_X1   g069(.A1(new_n491), .A2(new_n466), .A3(G138), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n494), .B1(new_n485), .B2(new_n495), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n493), .A2(new_n496), .ZN(new_n497));
  OAI211_X1 g072(.A(G138), .B(new_n466), .C1(new_n462), .C2(new_n463), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT4), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n490), .B1(new_n497), .B2(new_n499), .ZN(G164));
  NAND2_X1  g075(.A1(G75), .A2(G543), .ZN(new_n501));
  AND2_X1   g076(.A1(KEYINPUT5), .A2(G543), .ZN(new_n502));
  NOR2_X1   g077(.A1(KEYINPUT5), .A2(G543), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(G62), .ZN(new_n505));
  OAI21_X1  g080(.A(new_n501), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  AND2_X1   g081(.A1(KEYINPUT6), .A2(G651), .ZN(new_n507));
  NOR2_X1   g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  OAI21_X1  g083(.A(G543), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n506), .A2(G651), .B1(new_n510), .B2(G50), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT69), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n507), .A2(new_n508), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n512), .B1(new_n513), .B2(new_n504), .ZN(new_n514));
  XNOR2_X1  g089(.A(KEYINPUT5), .B(G543), .ZN(new_n515));
  OAI211_X1 g090(.A(new_n515), .B(KEYINPUT69), .C1(new_n508), .C2(new_n507), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(G88), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n511), .B1(new_n517), .B2(new_n518), .ZN(G303));
  INV_X1    g094(.A(G303), .ZN(G166));
  AND3_X1   g095(.A1(new_n515), .A2(G63), .A3(G651), .ZN(new_n521));
  NAND3_X1  g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  XOR2_X1   g097(.A(new_n522), .B(KEYINPUT7), .Z(new_n523));
  AOI211_X1 g098(.A(new_n521), .B(new_n523), .C1(G51), .C2(new_n510), .ZN(new_n524));
  AND2_X1   g099(.A1(new_n514), .A2(new_n516), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(G89), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n524), .A2(new_n526), .ZN(G286));
  INV_X1    g102(.A(G286), .ZN(G168));
  NAND2_X1  g103(.A1(new_n510), .A2(G52), .ZN(new_n529));
  INV_X1    g104(.A(G90), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n529), .B1(new_n517), .B2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT70), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n531), .B(new_n532), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n515), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n534));
  INV_X1    g109(.A(G651), .ZN(new_n535));
  OR2_X1    g110(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n533), .A2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT71), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n533), .A2(KEYINPUT71), .A3(new_n536), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n539), .A2(new_n540), .ZN(G171));
  NAND2_X1  g116(.A1(new_n525), .A2(G81), .ZN(new_n542));
  NAND2_X1  g117(.A1(G68), .A2(G543), .ZN(new_n543));
  INV_X1    g118(.A(G56), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n543), .B1(new_n504), .B2(new_n544), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n545), .A2(G651), .B1(new_n510), .B2(G43), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n542), .A2(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  NAND4_X1  g124(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT8), .ZN(new_n552));
  NAND4_X1  g127(.A1(G319), .A2(G483), .A3(G661), .A4(new_n552), .ZN(G188));
  NAND2_X1  g128(.A1(new_n525), .A2(G91), .ZN(new_n554));
  NAND2_X1  g129(.A1(KEYINPUT72), .A2(G53), .ZN(new_n555));
  OR3_X1    g130(.A1(new_n509), .A2(KEYINPUT9), .A3(new_n555), .ZN(new_n556));
  OAI21_X1  g131(.A(KEYINPUT9), .B1(new_n509), .B2(new_n555), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n515), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n559));
  OR2_X1    g134(.A1(new_n559), .A2(new_n535), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n554), .A2(new_n558), .A3(new_n560), .ZN(G299));
  INV_X1    g136(.A(G171), .ZN(G301));
  NAND3_X1  g137(.A1(new_n514), .A2(new_n516), .A3(G87), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(KEYINPUT73), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT73), .ZN(new_n565));
  NAND4_X1  g140(.A1(new_n514), .A2(new_n516), .A3(new_n565), .A4(G87), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n510), .A2(G49), .ZN(new_n568));
  OAI21_X1  g143(.A(G651), .B1(new_n515), .B2(G74), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n567), .A2(new_n571), .ZN(G288));
  NAND2_X1  g147(.A1(G73), .A2(G543), .ZN(new_n573));
  INV_X1    g148(.A(G61), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n573), .B1(new_n504), .B2(new_n574), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n575), .A2(G651), .B1(new_n510), .B2(G48), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n514), .A2(new_n516), .A3(G86), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(G305));
  AOI22_X1  g153(.A1(new_n515), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n579), .A2(new_n535), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT74), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n580), .A2(new_n581), .B1(G47), .B2(new_n510), .ZN(new_n582));
  XOR2_X1   g157(.A(KEYINPUT75), .B(G85), .Z(new_n583));
  OAI221_X1 g158(.A(new_n582), .B1(new_n581), .B2(new_n580), .C1(new_n517), .C2(new_n583), .ZN(G290));
  INV_X1    g159(.A(G92), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n517), .A2(new_n585), .ZN(new_n586));
  XNOR2_X1  g161(.A(new_n586), .B(KEYINPUT10), .ZN(new_n587));
  NAND2_X1  g162(.A1(G79), .A2(G543), .ZN(new_n588));
  INV_X1    g163(.A(G66), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n504), .B2(new_n589), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n590), .A2(G651), .B1(new_n510), .B2(G54), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n587), .A2(new_n591), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n592), .A2(G868), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n593), .B1(G171), .B2(G868), .ZN(G284));
  AOI21_X1  g169(.A(new_n593), .B1(G171), .B2(G868), .ZN(G321));
  INV_X1    g170(.A(G868), .ZN(new_n596));
  NOR2_X1   g171(.A1(G286), .A2(new_n596), .ZN(new_n597));
  XNOR2_X1  g172(.A(G299), .B(KEYINPUT76), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n597), .B1(new_n598), .B2(new_n596), .ZN(G280));
  XNOR2_X1  g174(.A(G280), .B(KEYINPUT77), .ZN(G297));
  INV_X1    g175(.A(new_n592), .ZN(new_n601));
  INV_X1    g176(.A(G559), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n602), .B2(G860), .ZN(G148));
  NAND2_X1  g178(.A1(new_n547), .A2(new_n596), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n592), .A2(G559), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n605), .B2(new_n596), .ZN(G323));
  XNOR2_X1  g181(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g182(.A1(new_n485), .A2(new_n468), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(KEYINPUT12), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT13), .ZN(new_n610));
  INV_X1    g185(.A(new_n610), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n611), .A2(G2100), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT78), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n465), .A2(G135), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n479), .A2(G123), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n466), .A2(G111), .ZN(new_n616));
  OAI21_X1  g191(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n617));
  OAI211_X1 g192(.A(new_n614), .B(new_n615), .C1(new_n616), .C2(new_n617), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(G2096), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n619), .B1(new_n611), .B2(G2100), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n613), .A2(new_n620), .ZN(G156));
  XNOR2_X1  g196(.A(KEYINPUT15), .B(G2435), .ZN(new_n622));
  XNOR2_X1  g197(.A(KEYINPUT80), .B(G2438), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  XOR2_X1   g199(.A(G2427), .B(G2430), .Z(new_n625));
  OR2_X1    g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  XOR2_X1   g201(.A(KEYINPUT79), .B(KEYINPUT14), .Z(new_n627));
  NAND2_X1  g202(.A1(new_n624), .A2(new_n625), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n626), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(G2451), .B(G2454), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT16), .ZN(new_n631));
  XNOR2_X1  g206(.A(G1341), .B(G1348), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n629), .B(new_n633), .Z(new_n634));
  XNOR2_X1  g209(.A(G2443), .B(G2446), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n634), .A2(new_n635), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n636), .A2(new_n637), .A3(G14), .ZN(new_n638));
  INV_X1    g213(.A(new_n638), .ZN(G401));
  XOR2_X1   g214(.A(G2067), .B(G2678), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT81), .ZN(new_n641));
  XOR2_X1   g216(.A(G2072), .B(G2078), .Z(new_n642));
  XOR2_X1   g217(.A(G2084), .B(G2090), .Z(new_n643));
  INV_X1    g218(.A(new_n643), .ZN(new_n644));
  NOR3_X1   g219(.A1(new_n641), .A2(new_n642), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT18), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n641), .A2(new_n642), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n642), .B(KEYINPUT17), .ZN(new_n648));
  OAI211_X1 g223(.A(new_n647), .B(new_n644), .C1(new_n641), .C2(new_n648), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n648), .A2(new_n641), .A3(new_n643), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n646), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2096), .B(G2100), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT82), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n651), .B(new_n653), .ZN(G227));
  XNOR2_X1  g229(.A(G1971), .B(G1976), .ZN(new_n655));
  XNOR2_X1  g230(.A(KEYINPUT83), .B(KEYINPUT19), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G1956), .B(G2474), .ZN(new_n658));
  XNOR2_X1  g233(.A(G1961), .B(G1966), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(KEYINPUT84), .B(KEYINPUT20), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(new_n660), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n658), .A2(new_n659), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  MUX2_X1   g241(.A(new_n666), .B(new_n665), .S(new_n657), .Z(new_n667));
  NAND2_X1  g242(.A1(new_n663), .A2(new_n667), .ZN(new_n668));
  INV_X1    g243(.A(G1981), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(G1986), .ZN(new_n671));
  XOR2_X1   g246(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT85), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n671), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1991), .B(G1996), .ZN(new_n675));
  OR2_X1    g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n674), .A2(new_n675), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(G229));
  INV_X1    g254(.A(G16), .ZN(new_n680));
  NOR2_X1   g255(.A1(G168), .A2(new_n680), .ZN(new_n681));
  AOI21_X1  g256(.A(new_n681), .B1(new_n680), .B2(G21), .ZN(new_n682));
  INV_X1    g257(.A(G1966), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(G164), .A2(G29), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n685), .B1(G27), .B2(G29), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n686), .A2(new_n443), .ZN(new_n687));
  INV_X1    g262(.A(G29), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n688), .A2(G26), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT28), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n465), .A2(G140), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n479), .A2(G128), .ZN(new_n692));
  OR2_X1    g267(.A1(G104), .A2(G2105), .ZN(new_n693));
  OAI211_X1 g268(.A(new_n693), .B(G2104), .C1(G116), .C2(new_n466), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n691), .A2(new_n692), .A3(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n690), .B1(new_n696), .B2(new_n688), .ZN(new_n697));
  INV_X1    g272(.A(G2067), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n682), .A2(new_n683), .ZN(new_n700));
  NAND4_X1  g275(.A1(new_n684), .A2(new_n687), .A3(new_n699), .A4(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n680), .A2(G19), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n702), .B1(new_n548), .B2(new_n680), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(G1341), .Z(new_n704));
  NAND2_X1  g279(.A1(new_n688), .A2(G32), .ZN(new_n705));
  AOI22_X1  g280(.A1(new_n465), .A2(G141), .B1(G105), .B2(new_n468), .ZN(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(new_n707));
  NAND3_X1  g282(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n708));
  XOR2_X1   g283(.A(new_n708), .B(KEYINPUT26), .Z(new_n709));
  INV_X1    g284(.A(G129), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n709), .B1(new_n486), .B2(new_n710), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n707), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n705), .B1(new_n712), .B2(new_n688), .ZN(new_n713));
  XNOR2_X1  g288(.A(KEYINPUT27), .B(G1996), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  OAI211_X1 g290(.A(new_n704), .B(new_n715), .C1(new_n443), .C2(new_n686), .ZN(new_n716));
  XNOR2_X1  g291(.A(KEYINPUT30), .B(G28), .ZN(new_n717));
  OR2_X1    g292(.A1(KEYINPUT31), .A2(G11), .ZN(new_n718));
  NAND2_X1  g293(.A1(KEYINPUT31), .A2(G11), .ZN(new_n719));
  AOI22_X1  g294(.A1(new_n717), .A2(new_n688), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(new_n618), .B2(new_n688), .ZN(new_n721));
  INV_X1    g296(.A(KEYINPUT24), .ZN(new_n722));
  INV_X1    g297(.A(G34), .ZN(new_n723));
  AOI21_X1  g298(.A(G29), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(new_n722), .B2(new_n723), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(G160), .B2(new_n688), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n721), .B1(new_n726), .B2(G2084), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n688), .A2(G35), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(G162), .B2(new_n688), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n729), .B(KEYINPUT29), .Z(new_n730));
  INV_X1    g305(.A(G2090), .ZN(new_n731));
  OAI221_X1 g306(.A(new_n727), .B1(G2084), .B2(new_n726), .C1(new_n730), .C2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n730), .A2(new_n731), .ZN(new_n733));
  AND2_X1   g308(.A1(new_n688), .A2(G33), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n735));
  INV_X1    g310(.A(KEYINPUT25), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(G139), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n485), .A2(new_n466), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n737), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(G115), .A2(G2104), .ZN(new_n741));
  INV_X1    g316(.A(G127), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n741), .B1(new_n464), .B2(new_n742), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n740), .B1(G2105), .B2(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(KEYINPUT90), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n744), .B(new_n745), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n734), .B1(new_n746), .B2(G29), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n747), .A2(new_n442), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n733), .A2(new_n748), .ZN(new_n749));
  NOR4_X1   g324(.A1(new_n701), .A2(new_n716), .A3(new_n732), .A4(new_n749), .ZN(new_n750));
  NOR2_X1   g325(.A1(G5), .A2(G16), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(G171), .B2(G16), .ZN(new_n752));
  INV_X1    g327(.A(G1961), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n752), .B(new_n753), .ZN(new_n754));
  NOR2_X1   g329(.A1(G4), .A2(G16), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(new_n601), .B2(G16), .ZN(new_n756));
  AND2_X1   g331(.A1(new_n756), .A2(G1348), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n756), .A2(G1348), .ZN(new_n758));
  XOR2_X1   g333(.A(KEYINPUT92), .B(KEYINPUT23), .Z(new_n759));
  NAND2_X1  g334(.A1(new_n680), .A2(G20), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n759), .B(new_n760), .ZN(new_n761));
  AND3_X1   g336(.A1(new_n554), .A2(new_n558), .A3(new_n560), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n761), .B1(new_n762), .B2(new_n680), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(G1956), .ZN(new_n764));
  NOR3_X1   g339(.A1(new_n757), .A2(new_n758), .A3(new_n764), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n747), .A2(new_n442), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT91), .ZN(new_n767));
  NAND4_X1  g342(.A1(new_n750), .A2(new_n754), .A3(new_n765), .A4(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n680), .A2(G22), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(G166), .B2(new_n680), .ZN(new_n770));
  INV_X1    g345(.A(G1971), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT89), .ZN(new_n773));
  INV_X1    g348(.A(KEYINPUT88), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(new_n567), .B2(new_n571), .ZN(new_n775));
  AOI211_X1 g350(.A(KEYINPUT88), .B(new_n570), .C1(new_n564), .C2(new_n566), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n777), .A2(G16), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G16), .B2(G23), .ZN(new_n779));
  XOR2_X1   g354(.A(KEYINPUT33), .B(G1976), .Z(new_n780));
  INV_X1    g355(.A(new_n780), .ZN(new_n781));
  OR2_X1    g356(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n779), .A2(new_n781), .ZN(new_n783));
  MUX2_X1   g358(.A(G6), .B(G305), .S(G16), .Z(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT32), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(new_n669), .ZN(new_n786));
  NAND4_X1  g361(.A1(new_n773), .A2(new_n782), .A3(new_n783), .A4(new_n786), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n787), .A2(KEYINPUT34), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n787), .A2(KEYINPUT34), .ZN(new_n789));
  MUX2_X1   g364(.A(G24), .B(G290), .S(G16), .Z(new_n790));
  XNOR2_X1  g365(.A(KEYINPUT87), .B(G1986), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n688), .A2(G25), .ZN(new_n793));
  INV_X1    g368(.A(G119), .ZN(new_n794));
  INV_X1    g369(.A(G131), .ZN(new_n795));
  OAI22_X1  g370(.A1(new_n794), .A2(new_n486), .B1(new_n739), .B2(new_n795), .ZN(new_n796));
  NOR2_X1   g371(.A1(G95), .A2(G2105), .ZN(new_n797));
  INV_X1    g372(.A(KEYINPUT86), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  OAI21_X1  g374(.A(G2104), .B1(new_n466), .B2(G107), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n796), .A2(new_n801), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n793), .B1(new_n802), .B2(new_n688), .ZN(new_n803));
  XOR2_X1   g378(.A(KEYINPUT35), .B(G1991), .Z(new_n804));
  INV_X1    g379(.A(new_n804), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n803), .B(new_n805), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n792), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n788), .A2(new_n789), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n808), .A2(KEYINPUT36), .ZN(new_n809));
  INV_X1    g384(.A(KEYINPUT36), .ZN(new_n810));
  NAND4_X1  g385(.A1(new_n788), .A2(new_n810), .A3(new_n789), .A4(new_n807), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n768), .B1(new_n809), .B2(new_n811), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT93), .ZN(G311));
  INV_X1    g388(.A(new_n812), .ZN(G150));
  NOR2_X1   g389(.A1(new_n592), .A2(new_n602), .ZN(new_n815));
  XOR2_X1   g390(.A(KEYINPUT94), .B(KEYINPUT38), .Z(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n510), .A2(G55), .ZN(new_n818));
  AOI22_X1  g393(.A1(new_n515), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n819));
  XNOR2_X1  g394(.A(KEYINPUT95), .B(G93), .ZN(new_n820));
  OAI221_X1 g395(.A(new_n818), .B1(new_n535), .B2(new_n819), .C1(new_n517), .C2(new_n820), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n547), .B(new_n821), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n817), .B(new_n822), .ZN(new_n823));
  AND2_X1   g398(.A1(new_n823), .A2(KEYINPUT39), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n823), .A2(KEYINPUT39), .ZN(new_n825));
  NOR3_X1   g400(.A1(new_n824), .A2(new_n825), .A3(G860), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n821), .A2(G860), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT37), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  XOR2_X1   g404(.A(new_n829), .B(KEYINPUT96), .Z(G145));
  XOR2_X1   g405(.A(KEYINPUT99), .B(G37), .Z(new_n831));
  INV_X1    g406(.A(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT98), .ZN(new_n833));
  OAI21_X1  g408(.A(KEYINPUT68), .B1(new_n464), .B2(new_n492), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n485), .A2(new_n495), .A3(new_n494), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n499), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n488), .A2(new_n489), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n837), .B1(new_n479), .B2(G126), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n696), .B(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n746), .B(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(new_n712), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  OR2_X1    g418(.A1(new_n746), .A2(new_n840), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n746), .A2(new_n840), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n844), .A2(new_n712), .A3(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n843), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n802), .A2(KEYINPUT97), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT97), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n849), .B1(new_n796), .B2(new_n801), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(new_n609), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n848), .A2(new_n609), .A3(new_n850), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n465), .A2(G142), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n479), .A2(G130), .ZN(new_n857));
  OR2_X1    g432(.A1(G106), .A2(G2105), .ZN(new_n858));
  OAI211_X1 g433(.A(new_n858), .B(G2104), .C1(G118), .C2(new_n466), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n856), .A2(new_n857), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n855), .A2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(new_n860), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n853), .A2(new_n862), .A3(new_n854), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n833), .B1(new_n847), .B2(new_n865), .ZN(new_n866));
  AOI211_X1 g441(.A(KEYINPUT98), .B(new_n864), .C1(new_n843), .C2(new_n846), .ZN(new_n867));
  OAI22_X1  g442(.A1(new_n866), .A2(new_n867), .B1(new_n847), .B2(new_n865), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n618), .B(new_n474), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(new_n483), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n832), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT100), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n865), .B1(new_n847), .B2(new_n872), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n873), .B1(new_n872), .B2(new_n847), .ZN(new_n874));
  INV_X1    g449(.A(new_n870), .ZN(new_n875));
  OAI211_X1 g450(.A(new_n874), .B(new_n875), .C1(new_n866), .C2(new_n867), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n871), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n877), .A2(KEYINPUT101), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT101), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n871), .A2(new_n876), .A3(new_n879), .ZN(new_n880));
  AND3_X1   g455(.A1(new_n878), .A2(KEYINPUT40), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(KEYINPUT40), .B1(new_n878), .B2(new_n880), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n881), .A2(new_n882), .ZN(G395));
  XNOR2_X1  g458(.A(new_n605), .B(new_n822), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n592), .B(new_n762), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT41), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n592), .B(G299), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n889), .A2(KEYINPUT41), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT102), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n888), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n885), .A2(KEYINPUT102), .A3(new_n887), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n886), .B1(new_n894), .B2(new_n884), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT42), .ZN(new_n896));
  OR2_X1    g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n777), .B(G166), .ZN(new_n898));
  XNOR2_X1  g473(.A(G290), .B(G305), .ZN(new_n899));
  OR2_X1    g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n898), .A2(new_n899), .ZN(new_n901));
  AND3_X1   g476(.A1(new_n900), .A2(KEYINPUT103), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n895), .A2(new_n896), .ZN(new_n903));
  AND3_X1   g478(.A1(new_n897), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n902), .B1(new_n897), .B2(new_n903), .ZN(new_n905));
  OAI21_X1  g480(.A(G868), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n821), .A2(new_n596), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(G295));
  NAND2_X1  g483(.A1(new_n906), .A2(new_n907), .ZN(G331));
  AOI21_X1  g484(.A(new_n822), .B1(new_n539), .B2(new_n540), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n539), .A2(new_n540), .A3(new_n822), .ZN(new_n912));
  AOI21_X1  g487(.A(G168), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(new_n912), .ZN(new_n914));
  NOR3_X1   g489(.A1(new_n914), .A2(G286), .A3(new_n910), .ZN(new_n915));
  OAI211_X1 g490(.A(new_n893), .B(new_n892), .C1(new_n913), .C2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n900), .A2(new_n901), .ZN(new_n917));
  OAI21_X1  g492(.A(G286), .B1(new_n914), .B2(new_n910), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n911), .A2(G168), .A3(new_n912), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n918), .A2(new_n919), .A3(new_n885), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n916), .A2(new_n917), .A3(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(G37), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT104), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n917), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n900), .A2(KEYINPUT104), .A3(new_n901), .ZN(new_n926));
  AOI22_X1  g501(.A1(new_n916), .A2(new_n920), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  OAI21_X1  g502(.A(KEYINPUT43), .B1(new_n923), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n925), .A2(new_n926), .ZN(new_n929));
  NAND4_X1  g504(.A1(new_n918), .A2(new_n919), .A3(KEYINPUT105), .A4(new_n885), .ZN(new_n930));
  AOI22_X1  g505(.A1(new_n918), .A2(new_n919), .B1(new_n888), .B2(new_n890), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT105), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n920), .A2(new_n932), .ZN(new_n933));
  OAI211_X1 g508(.A(new_n929), .B(new_n930), .C1(new_n931), .C2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT43), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n934), .A2(new_n935), .A3(new_n831), .A4(new_n921), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n928), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n935), .B1(new_n923), .B2(new_n927), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n934), .A2(KEYINPUT43), .A3(new_n831), .A4(new_n921), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  MUX2_X1   g515(.A(new_n937), .B(new_n940), .S(KEYINPUT44), .Z(G397));
  NAND2_X1  g516(.A1(G290), .A2(G1986), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  NOR2_X1   g518(.A1(G290), .A2(G1986), .ZN(new_n944));
  OR3_X1    g519(.A1(new_n943), .A2(KEYINPUT106), .A3(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(G1384), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n839), .A2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT45), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n469), .A2(new_n473), .A3(G40), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n952), .B1(new_n943), .B2(KEYINPUT106), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n712), .B(G1996), .ZN(new_n954));
  INV_X1    g529(.A(new_n802), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n955), .A2(new_n805), .ZN(new_n956));
  INV_X1    g531(.A(new_n956), .ZN(new_n957));
  XNOR2_X1  g532(.A(new_n695), .B(new_n698), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n955), .A2(new_n805), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n954), .A2(new_n957), .A3(new_n958), .A4(new_n959), .ZN(new_n960));
  AOI22_X1  g535(.A1(new_n945), .A2(new_n953), .B1(new_n960), .B2(new_n951), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n777), .A2(G1976), .ZN(new_n962));
  INV_X1    g537(.A(G1976), .ZN(new_n963));
  AOI21_X1  g538(.A(KEYINPUT52), .B1(G288), .B2(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(KEYINPUT107), .B1(new_n839), .B2(new_n946), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT107), .ZN(new_n966));
  AOI211_X1 g541(.A(new_n966), .B(G1384), .C1(new_n836), .C2(new_n838), .ZN(new_n967));
  NOR3_X1   g542(.A1(new_n965), .A2(new_n967), .A3(new_n950), .ZN(new_n968));
  INV_X1    g543(.A(G8), .ZN(new_n969));
  NOR3_X1   g544(.A1(new_n968), .A2(KEYINPUT109), .A3(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT109), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n966), .B1(G164), .B2(G1384), .ZN(new_n972));
  INV_X1    g547(.A(new_n950), .ZN(new_n973));
  AOI21_X1  g548(.A(G1384), .B1(new_n836), .B2(new_n838), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(KEYINPUT107), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n972), .A2(new_n973), .A3(new_n975), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n971), .B1(new_n976), .B2(G8), .ZN(new_n977));
  OAI211_X1 g552(.A(new_n962), .B(new_n964), .C1(new_n970), .C2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(KEYINPUT110), .ZN(new_n979));
  OAI21_X1  g554(.A(KEYINPUT109), .B1(new_n968), .B2(new_n969), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n976), .A2(new_n971), .A3(G8), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT110), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n982), .A2(new_n983), .A3(new_n962), .A4(new_n964), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n979), .A2(new_n984), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n950), .B1(new_n974), .B2(KEYINPUT45), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n949), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(new_n771), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT50), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n973), .B1(new_n974), .B2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n972), .A2(new_n975), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n991), .B1(new_n992), .B2(KEYINPUT50), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n988), .B1(new_n993), .B2(G2090), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT55), .ZN(new_n995));
  NOR3_X1   g570(.A1(G166), .A2(new_n995), .A3(new_n969), .ZN(new_n996));
  AOI21_X1  g571(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  OR2_X1    g573(.A1(new_n998), .A2(KEYINPUT108), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(KEYINPUT108), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n994), .A2(new_n999), .A3(G8), .A4(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(G305), .A2(G1981), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n576), .A2(new_n577), .A3(new_n669), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(KEYINPUT49), .ZN(new_n1005));
  OR2_X1    g580(.A1(new_n1004), .A2(KEYINPUT49), .ZN(new_n1006));
  AOI22_X1  g581(.A1(new_n980), .A2(new_n981), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n962), .B1(new_n970), .B2(new_n977), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1007), .B1(new_n1008), .B2(KEYINPUT52), .ZN(new_n1009));
  AND3_X1   g584(.A1(new_n985), .A2(new_n1001), .A3(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT113), .ZN(new_n1011));
  OAI21_X1  g586(.A(KEYINPUT50), .B1(new_n965), .B2(new_n967), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n950), .B1(new_n974), .B2(new_n989), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(KEYINPUT112), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT112), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1012), .A2(new_n1016), .A3(new_n1013), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1015), .A2(new_n731), .A3(new_n1017), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n969), .B1(new_n1018), .B2(new_n988), .ZN(new_n1019));
  INV_X1    g594(.A(new_n998), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1011), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(G2090), .B1(new_n1014), .B2(KEYINPUT112), .ZN(new_n1022));
  AOI22_X1  g597(.A1(new_n1022), .A2(new_n1017), .B1(new_n771), .B2(new_n987), .ZN(new_n1023));
  OAI211_X1 g598(.A(KEYINPUT113), .B(new_n998), .C1(new_n1023), .C2(new_n969), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1021), .A2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n948), .B1(new_n965), .B2(new_n967), .ZN(new_n1026));
  AOI21_X1  g601(.A(G1966), .B1(new_n1026), .B2(new_n986), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT114), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n965), .A2(new_n967), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n990), .B1(new_n1029), .B2(new_n989), .ZN(new_n1030));
  INV_X1    g605(.A(G2084), .ZN(new_n1031));
  AOI22_X1  g606(.A1(new_n1027), .A2(new_n1028), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(KEYINPUT45), .B1(new_n972), .B2(new_n975), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n974), .A2(KEYINPUT45), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(new_n973), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1033), .A2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g611(.A(KEYINPUT114), .B1(new_n1036), .B2(G1966), .ZN(new_n1037));
  AOI211_X1 g612(.A(new_n969), .B(G286), .C1(new_n1032), .C2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1010), .A2(new_n1025), .A3(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT116), .ZN(new_n1040));
  XOR2_X1   g615(.A(KEYINPUT115), .B(KEYINPUT63), .Z(new_n1041));
  AND3_X1   g616(.A1(new_n1039), .A2(new_n1040), .A3(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1040), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1043));
  AND2_X1   g618(.A1(new_n994), .A2(G8), .ZN(new_n1044));
  OR2_X1    g619(.A1(new_n1044), .A2(new_n1020), .ZN(new_n1045));
  AND4_X1   g620(.A1(KEYINPUT63), .A2(new_n1010), .A3(new_n1038), .A4(new_n1045), .ZN(new_n1046));
  NOR3_X1   g621(.A1(new_n1042), .A2(new_n1043), .A3(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(KEYINPUT121), .A2(KEYINPUT51), .ZN(new_n1048));
  OAI211_X1 g623(.A(new_n1028), .B(new_n683), .C1(new_n1033), .C2(new_n1035), .ZN(new_n1049));
  OAI211_X1 g624(.A(new_n991), .B(new_n1031), .C1(new_n992), .C2(KEYINPUT50), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1026), .A2(new_n986), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1028), .B1(new_n1052), .B2(new_n683), .ZN(new_n1053));
  NOR3_X1   g628(.A1(new_n1051), .A2(G286), .A3(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(G8), .B1(KEYINPUT121), .B2(KEYINPUT51), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1048), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1055), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1048), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1032), .A2(new_n1037), .ZN(new_n1059));
  OAI211_X1 g634(.A(new_n1057), .B(new_n1058), .C1(new_n1059), .C2(G286), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1056), .A2(new_n1060), .ZN(new_n1061));
  OAI211_X1 g636(.A(G8), .B(G286), .C1(new_n1051), .C2(new_n1053), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(KEYINPUT120), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT120), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1059), .A2(new_n1064), .A3(G8), .A4(G286), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1061), .A2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT124), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1067), .A2(new_n1068), .A3(KEYINPUT62), .ZN(new_n1069));
  AOI22_X1  g644(.A1(new_n1056), .A2(new_n1060), .B1(new_n1063), .B2(new_n1065), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT62), .ZN(new_n1071));
  OAI21_X1  g646(.A(KEYINPUT124), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  AND2_X1   g647(.A1(new_n949), .A2(new_n986), .ZN(new_n1073));
  AOI21_X1  g648(.A(KEYINPUT53), .B1(new_n1073), .B2(new_n443), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1074), .B1(new_n753), .B2(new_n993), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1036), .A2(KEYINPUT53), .A3(new_n443), .ZN(new_n1076));
  AOI21_X1  g651(.A(G301), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  AND3_X1   g652(.A1(new_n1010), .A2(new_n1025), .A3(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1069), .A2(new_n1072), .A3(new_n1078), .A4(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT54), .ZN(new_n1081));
  NAND2_X1  g656(.A1(G171), .A2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n468), .A2(G101), .ZN(new_n1083));
  INV_X1    g658(.A(G137), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1083), .B1(new_n739), .B2(new_n1084), .ZN(new_n1085));
  OAI211_X1 g660(.A(new_n473), .B(G40), .C1(new_n1085), .C2(KEYINPUT122), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1086), .B1(KEYINPUT122), .B2(new_n1085), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT123), .ZN(new_n1088));
  OR2_X1    g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  AND3_X1   g664(.A1(new_n949), .A2(KEYINPUT53), .A3(new_n443), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1089), .A2(new_n1090), .A3(new_n1034), .A4(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n539), .A2(KEYINPUT54), .A3(new_n540), .ZN(new_n1093));
  AND3_X1   g668(.A1(new_n1082), .A2(new_n1092), .A3(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1082), .A2(new_n1093), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1096));
  AOI22_X1  g671(.A1(new_n1094), .A2(new_n1075), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  AND3_X1   g672(.A1(new_n1010), .A2(new_n1025), .A3(new_n1097), .ZN(new_n1098));
  XNOR2_X1  g673(.A(KEYINPUT58), .B(G1341), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1099), .B1(new_n1029), .B2(new_n973), .ZN(new_n1100));
  INV_X1    g675(.A(G1996), .ZN(new_n1101));
  AND3_X1   g676(.A1(new_n949), .A2(new_n986), .A3(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n548), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1103));
  XOR2_X1   g678(.A(KEYINPUT118), .B(KEYINPUT59), .Z(new_n1104));
  INV_X1    g679(.A(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(G1348), .ZN(new_n1107));
  NOR3_X1   g682(.A1(new_n965), .A2(new_n967), .A3(KEYINPUT50), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1107), .B1(new_n1108), .B2(new_n990), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n968), .A2(new_n698), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1109), .A2(KEYINPUT60), .A3(new_n592), .A4(new_n1110), .ZN(new_n1111));
  OAI211_X1 g686(.A(new_n548), .B(new_n1104), .C1(new_n1100), .C2(new_n1102), .ZN(new_n1112));
  AND3_X1   g687(.A1(new_n1106), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT60), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1109), .A2(KEYINPUT60), .A3(new_n1110), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1116), .A2(new_n601), .A3(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(G1956), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1014), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT119), .ZN(new_n1121));
  AOI21_X1  g696(.A(KEYINPUT57), .B1(new_n558), .B2(KEYINPUT117), .ZN(new_n1122));
  XNOR2_X1  g697(.A(G299), .B(new_n1122), .ZN(new_n1123));
  XNOR2_X1  g698(.A(KEYINPUT56), .B(G2072), .ZN(new_n1124));
  AND3_X1   g699(.A1(new_n949), .A2(new_n986), .A3(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1125), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1120), .A2(new_n1121), .A3(new_n1123), .A4(new_n1126), .ZN(new_n1127));
  XNOR2_X1  g702(.A(new_n762), .B(new_n1122), .ZN(new_n1128));
  AOI21_X1  g703(.A(G1956), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1129));
  OAI211_X1 g704(.A(new_n1128), .B(new_n1121), .C1(new_n1129), .C2(new_n1125), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT61), .ZN(new_n1131));
  AND3_X1   g706(.A1(new_n1127), .A2(new_n1130), .A3(new_n1131), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1131), .B1(new_n1127), .B2(new_n1130), .ZN(new_n1133));
  OAI211_X1 g708(.A(new_n1113), .B(new_n1118), .C1(new_n1132), .C2(new_n1133), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1129), .A2(new_n1125), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1135), .A2(new_n1123), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1135), .A2(new_n1123), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n592), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1136), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  AOI22_X1  g714(.A1(new_n1066), .A2(new_n1061), .B1(new_n1134), .B2(new_n1139), .ZN(new_n1140));
  AND4_X1   g715(.A1(G8), .A2(new_n994), .A3(new_n999), .A4(new_n1000), .ZN(new_n1141));
  INV_X1    g716(.A(new_n984), .ZN(new_n1142));
  AOI22_X1  g717(.A1(new_n980), .A2(new_n981), .B1(G1976), .B2(new_n777), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n983), .B1(new_n1143), .B2(new_n964), .ZN(new_n1144));
  OAI211_X1 g719(.A(new_n1141), .B(new_n1009), .C1(new_n1142), .C2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n567), .A2(new_n963), .A3(new_n571), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1003), .B1(new_n1007), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1147), .A2(new_n982), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1145), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT111), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1145), .A2(KEYINPUT111), .A3(new_n1148), .ZN(new_n1152));
  AOI22_X1  g727(.A1(new_n1098), .A2(new_n1140), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1080), .A2(new_n1153), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n961), .B1(new_n1047), .B2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g730(.A(KEYINPUT46), .B1(new_n951), .B2(new_n1101), .ZN(new_n1156));
  OR2_X1    g731(.A1(new_n1156), .A2(KEYINPUT126), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1156), .A2(KEYINPUT126), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1101), .A2(KEYINPUT46), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n958), .A2(new_n712), .A3(new_n1159), .ZN(new_n1160));
  AOI22_X1  g735(.A1(new_n1157), .A2(new_n1158), .B1(new_n951), .B2(new_n1160), .ZN(new_n1161));
  XOR2_X1   g736(.A(new_n1161), .B(KEYINPUT47), .Z(new_n1162));
  NAND2_X1  g737(.A1(new_n944), .A2(new_n951), .ZN(new_n1163));
  XOR2_X1   g738(.A(new_n1163), .B(KEYINPUT127), .Z(new_n1164));
  OR2_X1    g739(.A1(new_n1164), .A2(KEYINPUT48), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n960), .A2(new_n951), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1164), .A2(KEYINPUT48), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1165), .A2(new_n1166), .A3(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n954), .A2(new_n958), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n957), .B1(new_n1169), .B2(new_n951), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1170), .B1(new_n698), .B2(new_n696), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n952), .B1(new_n1171), .B2(KEYINPUT125), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1172), .B1(KEYINPUT125), .B2(new_n1171), .ZN(new_n1173));
  AND3_X1   g748(.A1(new_n1162), .A2(new_n1168), .A3(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1155), .A2(new_n1174), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g750(.A(G319), .ZN(new_n1177));
  OR3_X1    g751(.A1(G401), .A2(new_n1177), .A3(G227), .ZN(new_n1178));
  AOI21_X1  g752(.A(new_n1178), .B1(new_n676), .B2(new_n677), .ZN(new_n1179));
  AOI21_X1  g753(.A(new_n879), .B1(new_n871), .B2(new_n876), .ZN(new_n1180));
  AND3_X1   g754(.A1(new_n871), .A2(new_n879), .A3(new_n876), .ZN(new_n1181));
  OAI211_X1 g755(.A(new_n937), .B(new_n1179), .C1(new_n1180), .C2(new_n1181), .ZN(G225));
  INV_X1    g756(.A(G225), .ZN(G308));
endmodule


