//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 0 0 1 0 0 1 0 0 1 1 0 0 1 0 0 0 1 1 1 0 1 0 0 1 1 0 1 1 1 0 0 1 0 0 1 1 1 0 0 0 1 0 1 0 0 0 0 0 1 0 0 1 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:42 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n740, new_n742,
    new_n743, new_n744, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n756, new_n757, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n835, new_n836, new_n837, new_n839, new_n840, new_n841, new_n843,
    new_n844, new_n845, new_n846, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n905, new_n906, new_n907, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n979, new_n980,
    new_n981, new_n982, new_n984, new_n985;
  XNOR2_X1  g000(.A(KEYINPUT69), .B(G71gat), .ZN(new_n202));
  INV_X1    g001(.A(G99gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XOR2_X1   g003(.A(G15gat), .B(G43gat), .Z(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(G227gat), .A2(G233gat), .ZN(new_n207));
  INV_X1    g006(.A(G169gat), .ZN(new_n208));
  INV_X1    g007(.A(G176gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  OR3_X1    g009(.A1(new_n210), .A2(KEYINPUT66), .A3(KEYINPUT26), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(KEYINPUT26), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n210), .A2(KEYINPUT26), .ZN(new_n213));
  AOI21_X1  g012(.A(KEYINPUT66), .B1(G169gat), .B2(G176gat), .ZN(new_n214));
  OAI211_X1 g013(.A(new_n211), .B(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(G183gat), .A2(G190gat), .ZN(new_n216));
  XNOR2_X1  g015(.A(KEYINPUT27), .B(G183gat), .ZN(new_n217));
  INV_X1    g016(.A(G190gat), .ZN(new_n218));
  AOI21_X1  g017(.A(KEYINPUT28), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n217), .A2(KEYINPUT28), .A3(new_n218), .ZN(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  OAI211_X1 g020(.A(new_n215), .B(new_n216), .C1(new_n219), .C2(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(KEYINPUT64), .B(KEYINPUT23), .ZN(new_n223));
  OAI21_X1  g022(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n224));
  INV_X1    g023(.A(new_n224), .ZN(new_n225));
  AOI22_X1  g024(.A1(new_n223), .A2(new_n210), .B1(new_n225), .B2(new_n216), .ZN(new_n226));
  NOR2_X1   g025(.A1(KEYINPUT65), .A2(KEYINPUT25), .ZN(new_n227));
  INV_X1    g026(.A(new_n227), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n208), .A2(new_n209), .A3(KEYINPUT23), .ZN(new_n229));
  AND2_X1   g028(.A1(G183gat), .A2(G190gat), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT24), .ZN(new_n231));
  AOI22_X1  g030(.A1(new_n230), .A2(new_n231), .B1(G169gat), .B2(G176gat), .ZN(new_n232));
  NAND4_X1  g031(.A1(new_n226), .A2(new_n228), .A3(new_n229), .A4(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT23), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(KEYINPUT64), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT64), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(KEYINPUT23), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n210), .A2(new_n235), .A3(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(G183gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(new_n218), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n240), .A2(KEYINPUT24), .A3(new_n216), .ZN(new_n241));
  NAND4_X1  g040(.A1(new_n232), .A2(new_n238), .A3(new_n241), .A4(new_n229), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(new_n227), .ZN(new_n243));
  NAND2_X1  g042(.A1(KEYINPUT65), .A2(KEYINPUT25), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n233), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n222), .A2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(G120gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(G113gat), .ZN(new_n248));
  INV_X1    g047(.A(G113gat), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(G120gat), .ZN(new_n250));
  AOI21_X1  g049(.A(KEYINPUT1), .B1(new_n248), .B2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT67), .ZN(new_n252));
  XNOR2_X1  g051(.A(G127gat), .B(G134gat), .ZN(new_n253));
  OR3_X1    g052(.A1(new_n251), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n252), .B1(new_n251), .B2(new_n253), .ZN(new_n255));
  AND2_X1   g054(.A1(KEYINPUT68), .A2(G113gat), .ZN(new_n256));
  NOR2_X1   g055(.A1(KEYINPUT68), .A2(G113gat), .ZN(new_n257));
  OAI21_X1  g056(.A(G120gat), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(KEYINPUT1), .B1(new_n258), .B2(new_n248), .ZN(new_n259));
  AOI22_X1  g058(.A1(new_n254), .A2(new_n255), .B1(new_n259), .B2(new_n253), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n246), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n222), .A2(new_n245), .A3(new_n260), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n207), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n206), .B1(new_n264), .B2(KEYINPUT33), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT32), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n262), .A2(new_n207), .A3(new_n263), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT34), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n271), .B1(new_n207), .B2(KEYINPUT70), .ZN(new_n272));
  OR2_X1    g071(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n270), .A2(new_n272), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n265), .A2(new_n267), .ZN(new_n275));
  NAND4_X1  g074(.A1(new_n269), .A2(new_n273), .A3(new_n274), .A4(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n273), .A2(new_n274), .ZN(new_n277));
  INV_X1    g076(.A(new_n275), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n277), .B1(new_n278), .B2(new_n268), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n276), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT88), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n276), .A2(new_n279), .A3(KEYINPUT88), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT84), .ZN(new_n286));
  XNOR2_X1  g085(.A(G197gat), .B(G204gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(KEYINPUT22), .ZN(new_n288));
  AND2_X1   g087(.A1(G211gat), .A2(G218gat), .ZN(new_n289));
  NOR2_X1   g088(.A1(G211gat), .A2(G218gat), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n288), .A2(new_n291), .ZN(new_n292));
  AND2_X1   g091(.A1(new_n290), .A2(KEYINPUT22), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n287), .B1(new_n293), .B2(new_n289), .ZN(new_n294));
  AND2_X1   g093(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(G226gat), .ZN(new_n296));
  INV_X1    g095(.A(G233gat), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT29), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n298), .B1(new_n246), .B2(new_n299), .ZN(new_n300));
  AOI211_X1 g099(.A(new_n296), .B(new_n297), .C1(new_n222), .C2(new_n245), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n295), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n246), .A2(new_n298), .ZN(new_n303));
  INV_X1    g102(.A(new_n295), .ZN(new_n304));
  AOI21_X1  g103(.A(KEYINPUT29), .B1(new_n222), .B2(new_n245), .ZN(new_n305));
  OAI211_X1 g104(.A(new_n303), .B(new_n304), .C1(new_n298), .C2(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n302), .A2(KEYINPUT71), .A3(new_n306), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n300), .A2(new_n301), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT71), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n308), .A2(new_n309), .A3(new_n304), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n307), .A2(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(G64gat), .B(G92gat), .ZN(new_n312));
  XNOR2_X1  g111(.A(new_n312), .B(G36gat), .ZN(new_n313));
  XNOR2_X1  g112(.A(new_n313), .B(KEYINPUT72), .ZN(new_n314));
  INV_X1    g113(.A(G8gat), .ZN(new_n315));
  XNOR2_X1  g114(.A(new_n314), .B(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n311), .A2(KEYINPUT30), .A3(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n307), .A2(new_n310), .A3(new_n316), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  AOI21_X1  g119(.A(KEYINPUT30), .B1(new_n311), .B2(new_n317), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n286), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  XNOR2_X1  g121(.A(KEYINPUT80), .B(KEYINPUT31), .ZN(new_n323));
  INV_X1    g122(.A(G50gat), .ZN(new_n324));
  XNOR2_X1  g123(.A(new_n323), .B(new_n324), .ZN(new_n325));
  XOR2_X1   g124(.A(G78gat), .B(G106gat), .Z(new_n326));
  XNOR2_X1  g125(.A(new_n325), .B(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(G22gat), .ZN(new_n328));
  NOR3_X1   g127(.A1(new_n327), .A2(KEYINPUT82), .A3(new_n328), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n329), .B1(new_n328), .B2(new_n327), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(G228gat), .ZN(new_n332));
  XNOR2_X1  g131(.A(G141gat), .B(G148gat), .ZN(new_n333));
  INV_X1    g132(.A(G162gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(KEYINPUT77), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT77), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(G162gat), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n335), .A2(new_n337), .A3(G155gat), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n333), .B1(new_n338), .B2(KEYINPUT2), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT78), .ZN(new_n340));
  XNOR2_X1  g139(.A(G155gat), .B(G162gat), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n339), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n340), .B1(new_n339), .B2(new_n341), .ZN(new_n344));
  XOR2_X1   g143(.A(KEYINPUT75), .B(KEYINPUT2), .Z(new_n345));
  NOR2_X1   g144(.A1(new_n345), .A2(new_n333), .ZN(new_n346));
  OAI21_X1  g145(.A(KEYINPUT74), .B1(G155gat), .B2(G162gat), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  NOR3_X1   g147(.A1(KEYINPUT74), .A2(G155gat), .A3(G162gat), .ZN(new_n349));
  INV_X1    g148(.A(G155gat), .ZN(new_n350));
  OAI22_X1  g149(.A1(new_n348), .A2(new_n349), .B1(new_n350), .B2(new_n334), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT76), .ZN(new_n352));
  NOR3_X1   g151(.A1(new_n346), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n333), .ZN(new_n354));
  XNOR2_X1  g153(.A(KEYINPUT75), .B(KEYINPUT2), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  OR3_X1    g155(.A1(KEYINPUT74), .A2(G155gat), .A3(G162gat), .ZN(new_n357));
  AOI22_X1  g156(.A1(new_n357), .A2(new_n347), .B1(G155gat), .B2(G162gat), .ZN(new_n358));
  AOI21_X1  g157(.A(KEYINPUT76), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  OAI22_X1  g158(.A1(new_n343), .A2(new_n344), .B1(new_n353), .B2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  AOI21_X1  g160(.A(KEYINPUT3), .B1(new_n304), .B2(new_n299), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n338), .A2(KEYINPUT2), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n364), .A2(new_n354), .A3(new_n341), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(KEYINPUT78), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(new_n342), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT3), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n352), .B1(new_n346), .B2(new_n351), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n356), .A2(new_n358), .A3(KEYINPUT76), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n367), .A2(new_n368), .A3(new_n371), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n304), .B1(new_n372), .B2(new_n299), .ZN(new_n373));
  OR4_X1    g172(.A1(new_n332), .A2(new_n363), .A3(new_n373), .A4(new_n297), .ZN(new_n374));
  AOI21_X1  g173(.A(KEYINPUT29), .B1(new_n295), .B2(KEYINPUT81), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n375), .B1(KEYINPUT81), .B2(new_n292), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n361), .B1(new_n376), .B2(new_n368), .ZN(new_n377));
  OAI22_X1  g176(.A1(new_n377), .A2(new_n373), .B1(new_n332), .B2(new_n297), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n331), .B1(new_n374), .B2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n374), .A2(new_n378), .A3(new_n331), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n311), .A2(new_n317), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT30), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND4_X1  g184(.A1(new_n385), .A2(KEYINPUT84), .A3(new_n319), .A4(new_n318), .ZN(new_n386));
  AND3_X1   g185(.A1(new_n322), .A2(new_n382), .A3(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT35), .ZN(new_n388));
  XNOR2_X1  g187(.A(KEYINPUT0), .B(G57gat), .ZN(new_n389));
  XNOR2_X1  g188(.A(new_n389), .B(G85gat), .ZN(new_n390));
  XNOR2_X1  g189(.A(G1gat), .B(G29gat), .ZN(new_n391));
  XOR2_X1   g190(.A(new_n390), .B(new_n391), .Z(new_n392));
  XNOR2_X1  g191(.A(new_n392), .B(KEYINPUT85), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n367), .A2(new_n260), .A3(new_n371), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(KEYINPUT4), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT4), .ZN(new_n397));
  NAND4_X1  g196(.A1(new_n367), .A2(new_n260), .A3(new_n397), .A4(new_n371), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n360), .A2(KEYINPUT3), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n400), .A2(new_n261), .A3(new_n372), .ZN(new_n401));
  NAND2_X1  g200(.A1(G225gat), .A2(G233gat), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n395), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n399), .A2(new_n401), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n360), .A2(new_n261), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT79), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n406), .A2(new_n407), .A3(new_n395), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n360), .A2(new_n261), .A3(KEYINPUT79), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n408), .A2(new_n403), .A3(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n405), .A2(new_n410), .A3(KEYINPUT5), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT86), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n403), .A2(KEYINPUT5), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n399), .A2(new_n401), .A3(new_n413), .ZN(new_n414));
  AND3_X1   g213(.A1(new_n411), .A2(new_n412), .A3(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n412), .B1(new_n411), .B2(new_n414), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n394), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n411), .A2(new_n414), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(KEYINPUT6), .B1(new_n419), .B2(new_n392), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n417), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n392), .B1(new_n411), .B2(new_n414), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(KEYINPUT6), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  NAND4_X1  g223(.A1(new_n285), .A2(new_n387), .A3(new_n388), .A4(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT73), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n321), .B1(new_n320), .B2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT6), .ZN(new_n428));
  INV_X1    g227(.A(new_n392), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n428), .B1(new_n418), .B2(new_n429), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n423), .B1(new_n430), .B2(new_n422), .ZN(new_n431));
  OAI211_X1 g230(.A(new_n427), .B(new_n431), .C1(new_n426), .C2(new_n320), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n382), .A2(new_n279), .A3(new_n276), .ZN(new_n433));
  OAI21_X1  g232(.A(KEYINPUT35), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n425), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n322), .A2(new_n386), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n418), .A2(KEYINPUT86), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n411), .A2(new_n412), .A3(new_n414), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n393), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n399), .A2(new_n401), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(new_n403), .ZN(new_n441));
  OR2_X1    g240(.A1(new_n441), .A2(KEYINPUT39), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n408), .A2(new_n409), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(new_n402), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n441), .A2(new_n444), .A3(KEYINPUT39), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n442), .A2(new_n393), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(KEYINPUT40), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT40), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n442), .A2(new_n445), .A3(new_n448), .A4(new_n393), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n439), .B1(new_n447), .B2(new_n449), .ZN(new_n450));
  AND3_X1   g249(.A1(new_n436), .A2(KEYINPUT87), .A3(new_n450), .ZN(new_n451));
  AOI21_X1  g250(.A(KEYINPUT87), .B1(new_n436), .B2(new_n450), .ZN(new_n452));
  AOI21_X1  g251(.A(KEYINPUT37), .B1(new_n307), .B2(new_n310), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n453), .A2(new_n317), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n302), .A2(new_n306), .ZN(new_n455));
  AOI21_X1  g254(.A(KEYINPUT38), .B1(new_n455), .B2(KEYINPUT37), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  OAI211_X1 g256(.A(new_n423), .B(new_n457), .C1(new_n439), .C2(new_n430), .ZN(new_n458));
  AND3_X1   g257(.A1(new_n307), .A2(KEYINPUT37), .A3(new_n310), .ZN(new_n459));
  NOR3_X1   g258(.A1(new_n459), .A2(new_n453), .A3(new_n317), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT38), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n383), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n382), .B1(new_n458), .B2(new_n462), .ZN(new_n463));
  NOR3_X1   g262(.A1(new_n451), .A2(new_n452), .A3(new_n463), .ZN(new_n464));
  AND3_X1   g263(.A1(new_n276), .A2(KEYINPUT36), .A3(new_n279), .ZN(new_n465));
  AOI21_X1  g264(.A(KEYINPUT36), .B1(new_n276), .B2(new_n279), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT83), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n382), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n380), .A2(KEYINPUT83), .A3(new_n381), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n467), .B1(new_n472), .B2(new_n432), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n435), .B1(new_n464), .B2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT96), .ZN(new_n476));
  INV_X1    g275(.A(G1gat), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(KEYINPUT16), .ZN(new_n478));
  AND2_X1   g277(.A1(G15gat), .A2(G22gat), .ZN(new_n479));
  NOR2_X1   g278(.A1(G15gat), .A2(G22gat), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n478), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(G15gat), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(new_n328), .ZN(new_n483));
  NAND2_X1  g282(.A1(G15gat), .A2(G22gat), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n483), .A2(new_n477), .A3(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n481), .A2(new_n485), .A3(KEYINPUT92), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT92), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n483), .A2(new_n487), .A3(new_n477), .A4(new_n484), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n486), .A2(G8gat), .A3(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT93), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n481), .A2(new_n490), .ZN(new_n491));
  XNOR2_X1  g290(.A(KEYINPUT94), .B(G8gat), .ZN(new_n492));
  OAI211_X1 g291(.A(new_n478), .B(KEYINPUT93), .C1(new_n479), .C2(new_n480), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n491), .A2(new_n485), .A3(new_n492), .A4(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n489), .A2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  OAI21_X1  g295(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n497));
  INV_X1    g296(.A(new_n497), .ZN(new_n498));
  NOR3_X1   g297(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n499));
  AND3_X1   g298(.A1(KEYINPUT90), .A2(G29gat), .A3(G36gat), .ZN(new_n500));
  AOI21_X1  g299(.A(KEYINPUT90), .B1(G29gat), .B2(G36gat), .ZN(new_n501));
  OAI22_X1  g300(.A1(new_n498), .A2(new_n499), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(G43gat), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n503), .A2(G50gat), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n324), .A2(G43gat), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n502), .A2(KEYINPUT15), .A3(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT15), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n508), .B1(new_n504), .B2(new_n505), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n324), .A2(G43gat), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n503), .A2(G50gat), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n510), .A2(new_n511), .A3(KEYINPUT15), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT14), .ZN(new_n513));
  INV_X1    g312(.A(G29gat), .ZN(new_n514));
  INV_X1    g313(.A(G36gat), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n513), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(new_n497), .ZN(new_n517));
  NAND2_X1  g316(.A1(G29gat), .A2(G36gat), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT90), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g319(.A1(KEYINPUT90), .A2(G29gat), .A3(G36gat), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND4_X1  g321(.A1(new_n509), .A2(new_n512), .A3(new_n517), .A4(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT91), .ZN(new_n525));
  AOI21_X1  g324(.A(KEYINPUT17), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT17), .ZN(new_n527));
  AOI211_X1 g326(.A(KEYINPUT91), .B(new_n527), .C1(new_n507), .C2(new_n523), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n496), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n495), .A2(new_n524), .ZN(new_n530));
  NAND2_X1  g329(.A1(G229gat), .A2(G233gat), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n529), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(KEYINPUT18), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT18), .ZN(new_n534));
  NAND4_X1  g333(.A1(new_n529), .A2(new_n534), .A3(new_n530), .A4(new_n531), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n531), .B(KEYINPUT13), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(new_n530), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n495), .A2(new_n524), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n537), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(KEYINPUT95), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT95), .ZN(new_n542));
  OAI211_X1 g341(.A(new_n542), .B(new_n537), .C1(new_n538), .C2(new_n539), .ZN(new_n543));
  AOI22_X1  g342(.A1(new_n533), .A2(new_n535), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(G113gat), .B(G141gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(G169gat), .B(G197gat), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n545), .B(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(KEYINPUT89), .B(KEYINPUT11), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n547), .B(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n549), .B(KEYINPUT12), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n476), .B1(new_n544), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n533), .A2(new_n535), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n541), .A2(new_n543), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n555), .A2(new_n550), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n552), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n555), .A2(new_n476), .A3(new_n550), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  XOR2_X1   g358(.A(G57gat), .B(G64gat), .Z(new_n560));
  OR2_X1    g359(.A1(G71gat), .A2(G78gat), .ZN(new_n561));
  NAND2_X1  g360(.A1(G71gat), .A2(G78gat), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT9), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n560), .A2(new_n563), .A3(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(G57gat), .B(G64gat), .ZN(new_n567));
  OAI211_X1 g366(.A(new_n562), .B(new_n561), .C1(new_n567), .C2(new_n564), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  XOR2_X1   g368(.A(G99gat), .B(G106gat), .Z(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT100), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT8), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n573), .B1(G99gat), .B2(G106gat), .ZN(new_n574));
  NOR2_X1   g373(.A1(G85gat), .A2(G92gat), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n572), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(G99gat), .A2(G106gat), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n577), .A2(KEYINPUT8), .ZN(new_n578));
  INV_X1    g377(.A(G85gat), .ZN(new_n579));
  INV_X1    g378(.A(G92gat), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n578), .A2(KEYINPUT100), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n576), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(G85gat), .A2(G92gat), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT7), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n571), .B1(new_n583), .B2(new_n589), .ZN(new_n590));
  AOI211_X1 g389(.A(new_n570), .B(new_n588), .C1(new_n576), .C2(new_n582), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n569), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  AND3_X1   g391(.A1(new_n578), .A2(KEYINPUT100), .A3(new_n581), .ZN(new_n593));
  AOI21_X1  g392(.A(KEYINPUT100), .B1(new_n578), .B2(new_n581), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n589), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n595), .A2(new_n570), .ZN(new_n596));
  INV_X1    g395(.A(new_n569), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n583), .A2(new_n571), .A3(new_n589), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(KEYINPUT102), .B(KEYINPUT10), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n592), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  NAND4_X1  g400(.A1(new_n596), .A2(new_n597), .A3(new_n598), .A4(KEYINPUT10), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(G230gat), .A2(G233gat), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(G120gat), .B(G148gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(new_n209), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(G204gat), .ZN(new_n608));
  AND2_X1   g407(.A1(new_n592), .A2(new_n599), .ZN(new_n609));
  OAI211_X1 g408(.A(new_n605), .B(new_n608), .C1(new_n604), .C2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n608), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n609), .A2(new_n604), .ZN(new_n612));
  INV_X1    g411(.A(new_n604), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n613), .B1(new_n601), .B2(new_n602), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n611), .B1(new_n612), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n610), .A2(new_n615), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n559), .A2(new_n616), .ZN(new_n617));
  AND2_X1   g416(.A1(new_n475), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT21), .ZN(new_n619));
  OAI211_X1 g418(.A(new_n489), .B(new_n494), .C1(new_n569), .C2(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n620), .B(G183gat), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n597), .A2(KEYINPUT21), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n620), .B(new_n239), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n625), .A2(new_n622), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n628));
  XOR2_X1   g427(.A(new_n628), .B(KEYINPUT99), .Z(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n627), .A2(new_n630), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n629), .B1(new_n624), .B2(new_n626), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(KEYINPUT97), .B(KEYINPUT98), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(G211gat), .ZN(new_n635));
  XOR2_X1   g434(.A(G127gat), .B(G155gat), .Z(new_n636));
  XOR2_X1   g435(.A(new_n635), .B(new_n636), .Z(new_n637));
  NAND2_X1  g436(.A1(G231gat), .A2(G233gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n637), .B(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n633), .A2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n639), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n631), .A2(new_n641), .A3(new_n632), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(G134gat), .B(G162gat), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  OAI22_X1  g445(.A1(new_n526), .A2(new_n528), .B1(new_n591), .B2(new_n590), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n596), .A2(new_n524), .A3(new_n598), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT101), .ZN(new_n649));
  NAND3_X1  g448(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n650));
  AND3_X1   g449(.A1(new_n648), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n649), .B1(new_n648), .B2(new_n650), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n647), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  AOI21_X1  g452(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(G190gat), .B(G218gat), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n654), .ZN(new_n658));
  OAI211_X1 g457(.A(new_n658), .B(new_n647), .C1(new_n651), .C2(new_n652), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n655), .A2(new_n657), .A3(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n657), .B1(new_n655), .B2(new_n659), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n646), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n662), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n664), .A2(new_n645), .A3(new_n660), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n644), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n618), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n668), .A2(new_n431), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(new_n477), .ZN(G1324gat));
  INV_X1    g469(.A(new_n436), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n673));
  OR2_X1    g472(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n672), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT42), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND4_X1  g476(.A1(new_n672), .A2(KEYINPUT42), .A3(new_n673), .A4(new_n674), .ZN(new_n678));
  OAI211_X1 g477(.A(new_n677), .B(new_n678), .C1(new_n315), .C2(new_n672), .ZN(G1325gat));
  INV_X1    g478(.A(KEYINPUT103), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n467), .B(new_n680), .ZN(new_n681));
  NOR3_X1   g480(.A1(new_n668), .A2(new_n482), .A3(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n668), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(new_n285), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n682), .B1(new_n482), .B2(new_n684), .ZN(G1326gat));
  NOR2_X1   g484(.A1(new_n668), .A2(new_n471), .ZN(new_n686));
  XOR2_X1   g485(.A(KEYINPUT43), .B(G22gat), .Z(new_n687));
  XNOR2_X1  g486(.A(new_n686), .B(new_n687), .ZN(G1327gat));
  NAND2_X1  g487(.A1(new_n475), .A2(new_n666), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n617), .A2(new_n644), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n431), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n691), .A2(new_n514), .A3(new_n692), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(KEYINPUT45), .ZN(new_n694));
  XOR2_X1   g493(.A(KEYINPUT104), .B(KEYINPUT44), .Z(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n689), .A2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT104), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT44), .ZN(new_n699));
  OAI211_X1 g498(.A(new_n475), .B(new_n666), .C1(new_n698), .C2(new_n699), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n690), .B1(new_n697), .B2(new_n700), .ZN(new_n701));
  AND2_X1   g500(.A1(new_n701), .A2(new_n692), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n694), .B1(new_n514), .B2(new_n702), .ZN(G1328gat));
  INV_X1    g502(.A(new_n689), .ZN(new_n704));
  INV_X1    g503(.A(new_n690), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NOR3_X1   g505(.A1(new_n706), .A2(G36gat), .A3(new_n671), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT46), .ZN(new_n708));
  OR2_X1    g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n707), .A2(new_n708), .ZN(new_n710));
  AND2_X1   g509(.A1(new_n701), .A2(new_n436), .ZN(new_n711));
  OAI211_X1 g510(.A(new_n709), .B(new_n710), .C1(new_n711), .C2(new_n515), .ZN(G1329gat));
  XOR2_X1   g511(.A(KEYINPUT105), .B(KEYINPUT47), .Z(new_n713));
  NOR2_X1   g512(.A1(new_n284), .A2(G43gat), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n704), .A2(new_n705), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(KEYINPUT106), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT106), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n691), .A2(new_n717), .A3(new_n714), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(new_n681), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n503), .B1(new_n701), .B2(new_n720), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n713), .B1(new_n719), .B2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(new_n467), .ZN(new_n723));
  AOI211_X1 g522(.A(new_n723), .B(new_n690), .C1(new_n697), .C2(new_n700), .ZN(new_n724));
  OAI211_X1 g523(.A(KEYINPUT47), .B(new_n715), .C1(new_n724), .C2(new_n503), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n722), .A2(new_n725), .ZN(G1330gat));
  INV_X1    g525(.A(KEYINPUT48), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n324), .B1(new_n701), .B2(new_n472), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n471), .A2(G50gat), .ZN(new_n729));
  INV_X1    g528(.A(new_n729), .ZN(new_n730));
  NOR3_X1   g529(.A1(new_n706), .A2(KEYINPUT107), .A3(new_n730), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n727), .B1(new_n728), .B2(new_n731), .ZN(new_n732));
  OAI22_X1  g531(.A1(new_n706), .A2(new_n730), .B1(KEYINPUT107), .B2(KEYINPUT48), .ZN(new_n733));
  INV_X1    g532(.A(new_n382), .ZN(new_n734));
  AOI211_X1 g533(.A(new_n727), .B(new_n324), .C1(new_n701), .C2(new_n734), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n732), .B1(new_n733), .B2(new_n735), .ZN(G1331gat));
  INV_X1    g535(.A(new_n559), .ZN(new_n737));
  NOR3_X1   g536(.A1(new_n737), .A2(new_n644), .A3(new_n666), .ZN(new_n738));
  AND3_X1   g537(.A1(new_n475), .A2(new_n616), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(new_n692), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g540(.A1(new_n739), .A2(new_n436), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n742), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n743));
  XOR2_X1   g542(.A(KEYINPUT49), .B(G64gat), .Z(new_n744));
  OAI21_X1  g543(.A(new_n743), .B1(new_n742), .B2(new_n744), .ZN(G1333gat));
  NAND4_X1  g544(.A1(new_n475), .A2(new_n616), .A3(new_n285), .A4(new_n738), .ZN(new_n746));
  OR2_X1    g545(.A1(new_n746), .A2(KEYINPUT108), .ZN(new_n747));
  INV_X1    g546(.A(G71gat), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n746), .A2(KEYINPUT108), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n747), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n739), .A2(G71gat), .A3(new_n720), .ZN(new_n751));
  XNOR2_X1  g550(.A(KEYINPUT109), .B(KEYINPUT50), .ZN(new_n752));
  AND3_X1   g551(.A1(new_n750), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n752), .B1(new_n750), .B2(new_n751), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n753), .A2(new_n754), .ZN(G1334gat));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n472), .ZN(new_n756));
  XOR2_X1   g555(.A(KEYINPUT110), .B(G78gat), .Z(new_n757));
  XNOR2_X1  g556(.A(new_n756), .B(new_n757), .ZN(G1335gat));
  NOR2_X1   g557(.A1(new_n737), .A2(new_n643), .ZN(new_n759));
  INV_X1    g558(.A(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(new_n616), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  AND2_X1   g561(.A1(new_n663), .A2(new_n665), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n698), .A2(new_n699), .ZN(new_n764));
  INV_X1    g563(.A(new_n463), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n436), .A2(new_n450), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT87), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n436), .A2(new_n450), .A3(KEYINPUT87), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n765), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(new_n473), .ZN(new_n771));
  AOI211_X1 g570(.A(new_n763), .B(new_n764), .C1(new_n771), .C2(new_n435), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n695), .B1(new_n475), .B2(new_n666), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n762), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NOR3_X1   g573(.A1(new_n774), .A2(new_n579), .A3(new_n431), .ZN(new_n775));
  OAI21_X1  g574(.A(KEYINPUT51), .B1(new_n689), .B2(new_n760), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT51), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n475), .A2(new_n777), .A3(new_n666), .A4(new_n759), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n776), .A2(new_n692), .A3(new_n616), .A4(new_n778), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n775), .B1(new_n579), .B2(new_n779), .ZN(G1336gat));
  NAND4_X1  g579(.A1(new_n776), .A2(new_n580), .A3(new_n616), .A4(new_n778), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n781), .A2(new_n671), .ZN(new_n782));
  INV_X1    g581(.A(new_n762), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n783), .B1(new_n697), .B2(new_n700), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n580), .B1(new_n784), .B2(new_n436), .ZN(new_n785));
  OAI21_X1  g584(.A(KEYINPUT52), .B1(new_n782), .B2(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(G92gat), .B1(new_n774), .B2(new_n671), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT52), .ZN(new_n788));
  OAI211_X1 g587(.A(new_n787), .B(new_n788), .C1(new_n671), .C2(new_n781), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n786), .A2(new_n789), .ZN(G1337gat));
  OAI21_X1  g589(.A(G99gat), .B1(new_n774), .B2(new_n681), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n776), .A2(new_n203), .A3(new_n616), .A4(new_n778), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n791), .B1(new_n284), .B2(new_n792), .ZN(G1338gat));
  OAI21_X1  g592(.A(G106gat), .B1(new_n774), .B2(new_n382), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT53), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n382), .A2(G106gat), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n776), .A2(new_n616), .A3(new_n778), .A4(new_n796), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n794), .A2(new_n795), .A3(new_n797), .ZN(new_n798));
  OAI211_X1 g597(.A(new_n472), .B(new_n762), .C1(new_n772), .C2(new_n773), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(G106gat), .ZN(new_n800));
  AND3_X1   g599(.A1(new_n800), .A2(KEYINPUT111), .A3(new_n797), .ZN(new_n801));
  OAI21_X1  g600(.A(KEYINPUT53), .B1(new_n800), .B2(KEYINPUT111), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n798), .B1(new_n801), .B2(new_n802), .ZN(G1339gat));
  NAND2_X1  g602(.A1(new_n738), .A2(new_n761), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n601), .A2(new_n602), .A3(new_n613), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n605), .A2(KEYINPUT54), .A3(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT54), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n608), .B1(new_n614), .B2(new_n807), .ZN(new_n808));
  AND3_X1   g607(.A1(new_n806), .A2(KEYINPUT55), .A3(new_n808), .ZN(new_n809));
  AOI21_X1  g608(.A(KEYINPUT55), .B1(new_n806), .B2(new_n808), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND4_X1  g610(.A1(new_n557), .A2(new_n811), .A3(new_n610), .A4(new_n558), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n544), .A2(new_n551), .ZN(new_n813));
  INV_X1    g612(.A(new_n549), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n531), .B1(new_n529), .B2(new_n530), .ZN(new_n815));
  NOR3_X1   g614(.A1(new_n538), .A2(new_n539), .A3(new_n537), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n814), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n813), .A2(new_n616), .A3(new_n817), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n666), .B1(new_n812), .B2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(new_n610), .ZN(new_n820));
  NOR3_X1   g619(.A1(new_n809), .A2(new_n810), .A3(new_n820), .ZN(new_n821));
  AND2_X1   g620(.A1(new_n813), .A2(new_n817), .ZN(new_n822));
  AND3_X1   g621(.A1(new_n666), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n644), .B1(new_n819), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n804), .A2(new_n824), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n436), .A2(new_n431), .ZN(new_n826));
  AND2_X1   g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(new_n433), .ZN(new_n828));
  AND2_X1   g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  OAI211_X1 g628(.A(new_n829), .B(new_n737), .C1(new_n257), .C2(new_n256), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n472), .A2(new_n284), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n827), .A2(new_n831), .ZN(new_n832));
  OAI21_X1  g631(.A(G113gat), .B1(new_n832), .B2(new_n559), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n830), .A2(new_n833), .ZN(G1340gat));
  OAI21_X1  g633(.A(G120gat), .B1(new_n832), .B2(new_n761), .ZN(new_n835));
  XOR2_X1   g634(.A(new_n835), .B(KEYINPUT112), .Z(new_n836));
  NAND3_X1  g635(.A1(new_n829), .A2(new_n247), .A3(new_n616), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(G1341gat));
  AOI21_X1  g637(.A(G127gat), .B1(new_n829), .B2(new_n643), .ZN(new_n839));
  INV_X1    g638(.A(G127gat), .ZN(new_n840));
  NOR3_X1   g639(.A1(new_n832), .A2(new_n840), .A3(new_n644), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n839), .A2(new_n841), .ZN(G1342gat));
  INV_X1    g641(.A(G134gat), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n829), .A2(new_n843), .A3(new_n666), .ZN(new_n844));
  XOR2_X1   g643(.A(new_n844), .B(KEYINPUT56), .Z(new_n845));
  OAI21_X1  g644(.A(G134gat), .B1(new_n832), .B2(new_n763), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(G1343gat));
  INV_X1    g646(.A(KEYINPUT57), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n825), .A2(new_n848), .A3(new_n734), .ZN(new_n849));
  NOR3_X1   g648(.A1(new_n467), .A2(new_n436), .A3(new_n431), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT115), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT113), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n818), .A2(new_n853), .ZN(new_n854));
  NAND4_X1  g653(.A1(new_n813), .A2(new_n616), .A3(KEYINPUT113), .A4(new_n817), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  AND2_X1   g655(.A1(new_n806), .A2(new_n808), .ZN(new_n857));
  OAI21_X1  g656(.A(KEYINPUT55), .B1(new_n857), .B2(KEYINPUT114), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT114), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n820), .B1(new_n810), .B2(new_n859), .ZN(new_n860));
  NAND4_X1  g659(.A1(new_n557), .A2(new_n858), .A3(new_n860), .A4(new_n558), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n852), .B1(new_n856), .B2(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(new_n862), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n856), .A2(new_n861), .A3(new_n852), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n863), .A2(new_n763), .A3(new_n864), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n666), .A2(new_n821), .A3(new_n822), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n643), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NOR4_X1   g666(.A1(new_n737), .A2(new_n644), .A3(new_n666), .A4(new_n616), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n472), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n851), .B1(new_n869), .B2(KEYINPUT57), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n870), .A2(G141gat), .A3(new_n737), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT58), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(KEYINPUT116), .ZN(new_n873));
  INV_X1    g672(.A(G141gat), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n720), .A2(new_n382), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(new_n827), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n874), .B1(new_n876), .B2(new_n559), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n871), .A2(new_n873), .A3(new_n877), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n872), .A2(KEYINPUT116), .ZN(new_n879));
  XOR2_X1   g678(.A(new_n878), .B(new_n879), .Z(G1344gat));
  INV_X1    g679(.A(KEYINPUT119), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT118), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n825), .A2(KEYINPUT57), .A3(new_n734), .ZN(new_n883));
  AND3_X1   g682(.A1(new_n856), .A2(new_n861), .A3(new_n852), .ZN(new_n884));
  NOR3_X1   g683(.A1(new_n884), .A2(new_n862), .A3(new_n666), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n644), .B1(new_n885), .B2(new_n823), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n471), .B1(new_n886), .B2(new_n804), .ZN(new_n887));
  OAI211_X1 g686(.A(new_n882), .B(new_n883), .C1(new_n887), .C2(KEYINPUT57), .ZN(new_n888));
  OR2_X1    g687(.A1(new_n883), .A2(new_n882), .ZN(new_n889));
  XNOR2_X1  g688(.A(new_n850), .B(KEYINPUT117), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n888), .A2(new_n616), .A3(new_n889), .A4(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT59), .ZN(new_n892));
  INV_X1    g691(.A(G148gat), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  AND2_X1   g693(.A1(new_n891), .A2(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(new_n876), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n896), .A2(new_n893), .A3(new_n616), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n893), .B1(new_n870), .B2(new_n616), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n897), .B1(new_n898), .B2(KEYINPUT59), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n881), .B1(new_n895), .B2(new_n899), .ZN(new_n900));
  OR2_X1    g699(.A1(new_n898), .A2(KEYINPUT59), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n891), .A2(new_n894), .ZN(new_n902));
  NAND4_X1  g701(.A1(new_n901), .A2(new_n902), .A3(KEYINPUT119), .A4(new_n897), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n900), .A2(new_n903), .ZN(G1345gat));
  INV_X1    g703(.A(new_n870), .ZN(new_n905));
  NOR3_X1   g704(.A1(new_n905), .A2(new_n350), .A3(new_n644), .ZN(new_n906));
  AOI21_X1  g705(.A(G155gat), .B1(new_n896), .B2(new_n643), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n906), .A2(new_n907), .ZN(G1346gat));
  NAND2_X1  g707(.A1(new_n335), .A2(new_n337), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n896), .A2(new_n909), .A3(new_n666), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n870), .A2(new_n666), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT120), .ZN(new_n912));
  XNOR2_X1  g711(.A(new_n911), .B(new_n912), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n910), .B1(new_n913), .B2(new_n909), .ZN(G1347gat));
  NOR2_X1   g713(.A1(new_n671), .A2(new_n692), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n812), .A2(new_n818), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(new_n763), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n643), .B1(new_n917), .B2(new_n866), .ZN(new_n918));
  OAI211_X1 g717(.A(new_n831), .B(new_n915), .C1(new_n918), .C2(new_n868), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT122), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND4_X1  g720(.A1(new_n825), .A2(KEYINPUT122), .A3(new_n831), .A4(new_n915), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  OAI21_X1  g722(.A(G169gat), .B1(new_n923), .B2(new_n559), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n828), .A2(new_n436), .ZN(new_n925));
  XOR2_X1   g724(.A(new_n925), .B(KEYINPUT121), .Z(new_n926));
  AOI21_X1  g725(.A(new_n692), .B1(new_n804), .B2(new_n824), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  INV_X1    g727(.A(new_n928), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n929), .A2(new_n208), .A3(new_n737), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n924), .A2(new_n930), .ZN(G1348gat));
  NOR3_X1   g730(.A1(new_n923), .A2(new_n209), .A3(new_n761), .ZN(new_n932));
  AOI21_X1  g731(.A(G176gat), .B1(new_n929), .B2(new_n616), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n932), .A2(new_n933), .ZN(G1349gat));
  INV_X1    g733(.A(KEYINPUT60), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n921), .A2(new_n643), .A3(new_n922), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n936), .A2(KEYINPUT123), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT123), .ZN(new_n938));
  NAND4_X1  g737(.A1(new_n921), .A2(new_n922), .A3(new_n938), .A4(new_n643), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n937), .A2(G183gat), .A3(new_n939), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT124), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n929), .A2(new_n643), .A3(new_n217), .ZN(new_n942));
  AND3_X1   g741(.A1(new_n940), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n941), .B1(new_n940), .B2(new_n942), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n935), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n940), .A2(new_n942), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n946), .A2(KEYINPUT124), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n940), .A2(new_n941), .A3(new_n942), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n947), .A2(KEYINPUT60), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n945), .A2(new_n949), .ZN(G1350gat));
  NAND3_X1  g749(.A1(new_n929), .A2(new_n218), .A3(new_n666), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT61), .ZN(new_n952));
  INV_X1    g751(.A(new_n923), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(new_n666), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n952), .B1(new_n954), .B2(G190gat), .ZN(new_n955));
  AOI211_X1 g754(.A(KEYINPUT61), .B(new_n218), .C1(new_n953), .C2(new_n666), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n951), .B1(new_n955), .B2(new_n956), .ZN(G1351gat));
  AND2_X1   g756(.A1(new_n681), .A2(new_n915), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n888), .A2(new_n889), .A3(new_n958), .ZN(new_n959));
  OAI21_X1  g758(.A(G197gat), .B1(new_n959), .B2(new_n559), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n681), .A2(new_n734), .A3(new_n436), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT125), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND4_X1  g762(.A1(new_n681), .A2(KEYINPUT125), .A3(new_n734), .A4(new_n436), .ZN(new_n964));
  AND3_X1   g763(.A1(new_n963), .A2(new_n927), .A3(new_n964), .ZN(new_n965));
  INV_X1    g764(.A(new_n965), .ZN(new_n966));
  OR2_X1    g765(.A1(new_n966), .A2(G197gat), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n960), .B1(new_n559), .B2(new_n967), .ZN(G1352gat));
  INV_X1    g767(.A(G204gat), .ZN(new_n969));
  NAND4_X1  g768(.A1(new_n963), .A2(new_n969), .A3(new_n927), .A4(new_n964), .ZN(new_n970));
  OR3_X1    g769(.A1(new_n970), .A2(KEYINPUT126), .A3(new_n761), .ZN(new_n971));
  OAI21_X1  g770(.A(KEYINPUT126), .B1(new_n970), .B2(new_n761), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n973), .B1(KEYINPUT127), .B2(KEYINPUT62), .ZN(new_n974));
  NAND4_X1  g773(.A1(new_n888), .A2(new_n616), .A3(new_n889), .A4(new_n958), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n975), .A2(G204gat), .ZN(new_n976));
  XOR2_X1   g775(.A(KEYINPUT127), .B(KEYINPUT62), .Z(new_n977));
  OAI211_X1 g776(.A(new_n974), .B(new_n976), .C1(new_n973), .C2(new_n977), .ZN(G1353gat));
  NAND4_X1  g777(.A1(new_n888), .A2(new_n643), .A3(new_n889), .A4(new_n958), .ZN(new_n979));
  AND3_X1   g778(.A1(new_n979), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n980));
  AOI21_X1  g779(.A(KEYINPUT63), .B1(new_n979), .B2(G211gat), .ZN(new_n981));
  OR2_X1    g780(.A1(new_n644), .A2(G211gat), .ZN(new_n982));
  OAI22_X1  g781(.A1(new_n980), .A2(new_n981), .B1(new_n966), .B2(new_n982), .ZN(G1354gat));
  OAI21_X1  g782(.A(G218gat), .B1(new_n959), .B2(new_n763), .ZN(new_n984));
  OR2_X1    g783(.A1(new_n763), .A2(G218gat), .ZN(new_n985));
  OAI21_X1  g784(.A(new_n984), .B1(new_n966), .B2(new_n985), .ZN(G1355gat));
endmodule


