

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808;

  NOR2_X1 U375 ( .A1(n517), .A2(n515), .ZN(n514) );
  XNOR2_X1 U376 ( .A(n682), .B(KEYINPUT75), .ZN(n517) );
  XNOR2_X1 U377 ( .A(n372), .B(KEYINPUT106), .ZN(n804) );
  XNOR2_X1 U378 ( .A(n434), .B(n433), .ZN(n371) );
  XNOR2_X1 U379 ( .A(n380), .B(KEYINPUT109), .ZN(n494) );
  NAND2_X1 U380 ( .A1(n444), .A2(n464), .ZN(n380) );
  XNOR2_X1 U381 ( .A(n643), .B(n592), .ZN(n686) );
  BUF_X1 U382 ( .A(n622), .Z(n643) );
  XNOR2_X1 U383 ( .A(KEYINPUT65), .B(KEYINPUT22), .ZN(n364) );
  NAND2_X1 U384 ( .A1(n622), .A2(n687), .ZN(n636) );
  NAND2_X1 U385 ( .A1(n739), .A2(n728), .ZN(n591) );
  XOR2_X1 U386 ( .A(KEYINPUT10), .B(n576), .Z(n793) );
  NAND2_X2 U387 ( .A1(n443), .A2(n732), .ZN(n441) );
  NAND2_X1 U388 ( .A1(n354), .A2(n371), .ZN(n678) );
  NAND2_X1 U389 ( .A1(n487), .A2(n490), .ZN(n354) );
  NOR2_X2 U390 ( .A1(n502), .A2(n501), .ZN(n524) );
  XNOR2_X2 U391 ( .A(n586), .B(n782), .ZN(n739) );
  OR2_X4 U392 ( .A1(n788), .A2(n499), .ZN(n730) );
  XNOR2_X2 U393 ( .A(n469), .B(KEYINPUT41), .ZN(n697) );
  OR2_X2 U394 ( .A1(n769), .A2(G902), .ZN(n551) );
  AND2_X2 U395 ( .A1(n732), .A2(n731), .ZN(n776) );
  NOR2_X1 U396 ( .A1(G953), .A2(G237), .ZN(n604) );
  NOR2_X1 U397 ( .A1(n672), .A2(n718), .ZN(n436) );
  NOR2_X1 U398 ( .A1(n421), .A2(n671), .ZN(n448) );
  AND2_X1 U399 ( .A1(n662), .A2(n670), .ZN(n667) );
  XNOR2_X1 U400 ( .A(n671), .B(n522), .ZN(n662) );
  INV_X2 U401 ( .A(G953), .ZN(n722) );
  AND2_X1 U402 ( .A1(n431), .A2(n373), .ZN(n503) );
  AND2_X1 U403 ( .A1(n489), .A2(n488), .ZN(n487) );
  NAND2_X1 U404 ( .A1(n435), .A2(n357), .ZN(n434) );
  XNOR2_X1 U405 ( .A(n663), .B(KEYINPUT33), .ZN(n718) );
  NOR2_X1 U406 ( .A1(n617), .A2(n449), .ZN(n618) );
  XNOR2_X1 U407 ( .A(n612), .B(KEYINPUT102), .ZN(n633) );
  XNOR2_X1 U408 ( .A(n600), .B(n386), .ZN(n628) );
  NOR2_X1 U409 ( .A1(n777), .A2(G902), .ZN(n566) );
  OR2_X1 U410 ( .A1(n401), .A2(n518), .ZN(n404) );
  XNOR2_X1 U411 ( .A(n537), .B(n476), .ZN(n475) );
  XNOR2_X1 U412 ( .A(n377), .B(n535), .ZN(n476) );
  XNOR2_X1 U413 ( .A(n378), .B(n536), .ZN(n377) );
  AND2_X1 U414 ( .A1(n722), .A2(G224), .ZN(n423) );
  XNOR2_X1 U415 ( .A(KEYINPUT76), .B(KEYINPUT2), .ZN(n680) );
  AND2_X2 U416 ( .A1(n699), .A2(n698), .ZN(n670) );
  XNOR2_X2 U417 ( .A(n486), .B(n555), .ZN(n795) );
  NAND2_X1 U418 ( .A1(n529), .A2(n765), .ZN(n394) );
  AND2_X1 U419 ( .A1(n804), .A2(KEYINPUT81), .ZN(n373) );
  INV_X1 U420 ( .A(G237), .ZN(n538) );
  NAND2_X1 U421 ( .A1(n684), .A2(n736), .ZN(n650) );
  NAND2_X1 U422 ( .A1(n587), .A2(G214), .ZN(n687) );
  XNOR2_X1 U423 ( .A(n385), .B(n384), .ZN(n689) );
  INV_X1 U424 ( .A(KEYINPUT105), .ZN(n384) );
  XNOR2_X1 U425 ( .A(n564), .B(KEYINPUT25), .ZN(n565) );
  XNOR2_X1 U426 ( .A(G134), .B(G131), .ZN(n532) );
  NAND2_X1 U427 ( .A1(n721), .A2(n516), .ZN(n515) );
  INV_X1 U428 ( .A(KEYINPUT82), .ZN(n493) );
  NOR2_X1 U429 ( .A1(n631), .A2(KEYINPUT69), .ZN(n624) );
  INV_X1 U430 ( .A(KEYINPUT47), .ZN(n396) );
  INV_X1 U431 ( .A(KEYINPUT0), .ZN(n466) );
  XNOR2_X1 U432 ( .A(KEYINPUT96), .B(KEYINPUT12), .ZN(n390) );
  XNOR2_X1 U433 ( .A(G143), .B(G140), .ZN(n605) );
  XNOR2_X1 U434 ( .A(G104), .B(G113), .ZN(n601) );
  XOR2_X1 U435 ( .A(G131), .B(G122), .Z(n602) );
  XNOR2_X1 U436 ( .A(n388), .B(KEYINPUT11), .ZN(n387) );
  NAND2_X1 U437 ( .A1(n604), .A2(G214), .ZN(n388) );
  XNOR2_X1 U438 ( .A(n504), .B(n645), .ZN(n684) );
  XNOR2_X1 U439 ( .A(n589), .B(n588), .ZN(n590) );
  XNOR2_X1 U440 ( .A(n399), .B(n616), .ZN(n617) );
  NAND2_X1 U441 ( .A1(n409), .A2(n361), .ZN(n399) );
  XNOR2_X1 U442 ( .A(n477), .B(n534), .ZN(n537) );
  XNOR2_X1 U443 ( .A(n533), .B(G119), .ZN(n477) );
  XNOR2_X1 U444 ( .A(G116), .B(G113), .ZN(n533) );
  XOR2_X1 U445 ( .A(G137), .B(G140), .Z(n555) );
  XNOR2_X1 U446 ( .A(n560), .B(n498), .ZN(n497) );
  INV_X1 U447 ( .A(KEYINPUT24), .ZN(n498) );
  XNOR2_X1 U448 ( .A(KEYINPUT9), .B(KEYINPUT7), .ZN(n595) );
  XNOR2_X1 U449 ( .A(G107), .B(G116), .ZN(n593) );
  XNOR2_X1 U450 ( .A(n594), .B(n596), .ZN(n481) );
  INV_X1 U451 ( .A(G128), .ZN(n530) );
  OR2_X1 U452 ( .A1(n450), .A2(n642), .ZN(n383) );
  XNOR2_X1 U453 ( .A(n436), .B(n664), .ZN(n435) );
  XNOR2_X1 U454 ( .A(n376), .B(KEYINPUT107), .ZN(n375) );
  INV_X1 U455 ( .A(KEYINPUT101), .ZN(n386) );
  XNOR2_X1 U456 ( .A(n610), .B(n355), .ZN(n627) );
  NOR2_X1 U457 ( .A1(n773), .A2(G902), .ZN(n610) );
  XOR2_X1 U458 ( .A(G104), .B(G110), .Z(n545) );
  NAND2_X1 U459 ( .A1(n510), .A2(KEYINPUT123), .ZN(n509) );
  NAND2_X1 U460 ( .A1(n513), .A2(n512), .ZN(n511) );
  NOR2_X1 U461 ( .A1(n641), .A2(n483), .ZN(n638) );
  AND2_X1 U462 ( .A1(n362), .A2(n493), .ZN(n492) );
  INV_X1 U463 ( .A(KEYINPUT84), .ZN(n571) );
  XNOR2_X1 U464 ( .A(n624), .B(n396), .ZN(n395) );
  INV_X1 U465 ( .A(KEYINPUT48), .ZN(n391) );
  XNOR2_X1 U466 ( .A(KEYINPUT85), .B(KEYINPUT18), .ZN(n574) );
  NAND2_X1 U467 ( .A1(G234), .A2(G237), .ZN(n540) );
  AND2_X1 U468 ( .A1(n356), .A2(n698), .ZN(n473) );
  NAND2_X1 U469 ( .A1(n519), .A2(n539), .ZN(n518) );
  INV_X1 U470 ( .A(G472), .ZN(n519) );
  AND2_X1 U471 ( .A1(n521), .A2(n520), .ZN(n403) );
  NAND2_X1 U472 ( .A1(G902), .A2(G472), .ZN(n520) );
  XNOR2_X1 U473 ( .A(KEYINPUT94), .B(KEYINPUT5), .ZN(n536) );
  OR2_X1 U474 ( .A1(n678), .A2(KEYINPUT44), .ZN(n360) );
  XNOR2_X1 U475 ( .A(G128), .B(G110), .ZN(n553) );
  INV_X1 U476 ( .A(KEYINPUT70), .ZN(n472) );
  AND2_X1 U477 ( .A1(n667), .A2(n438), .ZN(n663) );
  INV_X1 U478 ( .A(n698), .ZN(n657) );
  XNOR2_X1 U479 ( .A(n668), .B(KEYINPUT95), .ZN(n709) );
  INV_X1 U480 ( .A(KEYINPUT30), .ZN(n470) );
  INV_X1 U481 ( .A(KEYINPUT90), .ZN(n465) );
  NAND2_X1 U482 ( .A1(n403), .A2(n404), .ZN(n402) );
  XNOR2_X1 U483 ( .A(n607), .B(n606), .ZN(n773) );
  XNOR2_X1 U484 ( .A(n389), .B(n387), .ZN(n606) );
  XNOR2_X1 U485 ( .A(n605), .B(n390), .ZN(n389) );
  NAND2_X1 U486 ( .A1(n467), .A2(n686), .ZN(n469) );
  NOR2_X1 U487 ( .A1(n689), .A2(n468), .ZN(n467) );
  NAND2_X1 U488 ( .A1(n640), .A2(n484), .ZN(n483) );
  XNOR2_X1 U489 ( .A(n669), .B(KEYINPUT31), .ZN(n430) );
  AND2_X1 U490 ( .A1(n709), .A2(n400), .ZN(n669) );
  INV_X1 U491 ( .A(KEYINPUT114), .ZN(n406) );
  XNOR2_X1 U492 ( .A(n537), .B(n411), .ZN(n782) );
  XNOR2_X1 U493 ( .A(n585), .B(n506), .ZN(n411) );
  INV_X1 U494 ( .A(G122), .ZN(n506) );
  XNOR2_X1 U495 ( .A(n495), .B(n561), .ZN(n777) );
  XNOR2_X1 U496 ( .A(n593), .B(n595), .ZN(n479) );
  NAND2_X1 U497 ( .A1(n426), .A2(n732), .ZN(n424) );
  XOR2_X1 U498 ( .A(G101), .B(G146), .Z(n547) );
  AND2_X1 U499 ( .A1(n453), .A2(n460), .ZN(n452) );
  NAND2_X1 U500 ( .A1(G953), .A2(n723), .ZN(n460) );
  NOR2_X1 U501 ( .A1(n507), .A2(n454), .ZN(n455) );
  XNOR2_X1 U502 ( .A(n644), .B(KEYINPUT111), .ZN(n803) );
  XNOR2_X1 U503 ( .A(n382), .B(KEYINPUT43), .ZN(n381) );
  INV_X1 U504 ( .A(KEYINPUT35), .ZN(n433) );
  INV_X1 U505 ( .A(KEYINPUT32), .ZN(n446) );
  AND2_X1 U506 ( .A1(n375), .A2(n661), .ZN(n463) );
  INV_X1 U507 ( .A(n430), .ZN(n760) );
  INV_X1 U508 ( .A(KEYINPUT110), .ZN(n485) );
  NAND2_X1 U509 ( .A1(n379), .A2(n677), .ZN(n372) );
  INV_X1 U510 ( .A(n380), .ZN(n379) );
  XNOR2_X1 U511 ( .A(n416), .B(n415), .ZN(G60) );
  INV_X1 U512 ( .A(KEYINPUT60), .ZN(n415) );
  NAND2_X1 U513 ( .A1(n418), .A2(n417), .ZN(n416) );
  XNOR2_X1 U514 ( .A(n424), .B(n366), .ZN(n418) );
  INV_X1 U515 ( .A(KEYINPUT56), .ZN(n412) );
  NAND2_X1 U516 ( .A1(n414), .A2(n417), .ZN(n413) );
  XNOR2_X1 U517 ( .A(n742), .B(n367), .ZN(n414) );
  XOR2_X1 U518 ( .A(n609), .B(n608), .Z(n355) );
  OR2_X1 U519 ( .A1(n653), .A2(n544), .ZN(n356) );
  XNOR2_X1 U520 ( .A(KEYINPUT72), .B(n665), .ZN(n357) );
  INV_X1 U521 ( .A(n450), .ZN(n464) );
  NOR2_X1 U522 ( .A1(n689), .A2(n657), .ZN(n358) );
  XOR2_X1 U523 ( .A(n683), .B(KEYINPUT74), .Z(n359) );
  INV_X1 U524 ( .A(n676), .ZN(n437) );
  INV_X1 U525 ( .A(n699), .ZN(n676) );
  AND2_X1 U526 ( .A1(n676), .A2(n473), .ZN(n361) );
  NOR2_X1 U527 ( .A1(n409), .A2(n699), .ZN(n362) );
  AND2_X1 U528 ( .A1(n730), .A2(KEYINPUT123), .ZN(n363) );
  XNOR2_X1 U529 ( .A(n633), .B(n485), .ZN(n757) );
  XOR2_X1 U530 ( .A(n679), .B(KEYINPUT45), .Z(n365) );
  XNOR2_X1 U531 ( .A(n773), .B(KEYINPUT59), .ZN(n366) );
  XOR2_X1 U532 ( .A(n741), .B(n740), .Z(n367) );
  XOR2_X1 U533 ( .A(n401), .B(KEYINPUT62), .Z(n368) );
  AND2_X1 U534 ( .A1(n729), .A2(G475), .ZN(n369) );
  AND2_X1 U535 ( .A1(n729), .A2(G210), .ZN(n370) );
  INV_X1 U536 ( .A(KEYINPUT81), .ZN(n527) );
  AND2_X1 U537 ( .A1(KEYINPUT53), .A2(n722), .ZN(n461) );
  INV_X1 U538 ( .A(n461), .ZN(n454) );
  INV_X1 U539 ( .A(n780), .ZN(n417) );
  XNOR2_X1 U540 ( .A(n371), .B(G122), .ZN(G24) );
  XNOR2_X2 U541 ( .A(n551), .B(n550), .ZN(n671) );
  NAND2_X1 U542 ( .A1(n431), .A2(n804), .ZN(n374) );
  NAND2_X1 U543 ( .A1(n374), .A2(n527), .ZN(n525) );
  NAND2_X1 U544 ( .A1(n662), .A2(n676), .ZN(n376) );
  NAND2_X1 U545 ( .A1(n604), .A2(G210), .ZN(n378) );
  NOR2_X1 U546 ( .A1(n381), .A2(n643), .ZN(n644) );
  NOR2_X1 U547 ( .A1(n641), .A2(n383), .ZN(n382) );
  NAND2_X1 U548 ( .A1(n627), .A2(n628), .ZN(n385) );
  XNOR2_X1 U549 ( .A(n392), .B(n391), .ZN(n505) );
  NAND2_X1 U550 ( .A1(n397), .A2(n393), .ZN(n392) );
  NOR2_X1 U551 ( .A1(n395), .A2(n394), .ZN(n393) );
  XNOR2_X1 U552 ( .A(n398), .B(KEYINPUT46), .ZN(n397) );
  NOR2_X2 U553 ( .A1(n737), .A2(n806), .ZN(n398) );
  XNOR2_X1 U554 ( .A(n656), .B(n466), .ZN(n400) );
  XNOR2_X1 U555 ( .A(n656), .B(n466), .ZN(n658) );
  XNOR2_X1 U556 ( .A(n480), .B(n478), .ZN(n775) );
  XNOR2_X1 U557 ( .A(n482), .B(n481), .ZN(n480) );
  XNOR2_X1 U558 ( .A(n774), .B(n775), .ZN(n419) );
  NOR2_X1 U559 ( .A1(n775), .A2(G902), .ZN(n599) );
  XNOR2_X1 U560 ( .A(n486), .B(n475), .ZN(n401) );
  XNOR2_X1 U561 ( .A(n486), .B(n475), .ZN(n733) );
  NAND2_X1 U562 ( .A1(n403), .A2(n404), .ZN(n634) );
  NAND2_X1 U563 ( .A1(n618), .A2(KEYINPUT114), .ZN(n407) );
  NAND2_X1 U564 ( .A1(n405), .A2(n406), .ZN(n408) );
  NAND2_X1 U565 ( .A1(n407), .A2(n408), .ZN(n750) );
  INV_X1 U566 ( .A(n618), .ZN(n405) );
  AND2_X1 U567 ( .A1(n730), .A2(n369), .ZN(n426) );
  AND2_X1 U568 ( .A1(n730), .A2(n370), .ZN(n442) );
  AND2_X2 U569 ( .A1(n730), .A2(n729), .ZN(n731) );
  INV_X1 U570 ( .A(n636), .ZN(n484) );
  XNOR2_X1 U571 ( .A(n402), .B(KEYINPUT108), .ZN(n409) );
  XNOR2_X1 U572 ( .A(n634), .B(KEYINPUT108), .ZN(n660) );
  BUF_X1 U573 ( .A(n662), .Z(n450) );
  BUF_X1 U574 ( .A(n724), .Z(n410) );
  BUF_X1 U575 ( .A(n402), .Z(n706) );
  BUF_X1 U576 ( .A(n671), .Z(n449) );
  NAND2_X1 U577 ( .A1(n733), .A2(G472), .ZN(n521) );
  XNOR2_X1 U578 ( .A(n569), .B(KEYINPUT71), .ZN(n625) );
  AND2_X2 U579 ( .A1(n731), .A2(G472), .ZN(n443) );
  INV_X2 U580 ( .A(G125), .ZN(n420) );
  NAND2_X1 U581 ( .A1(n625), .A2(n686), .ZN(n445) );
  NAND2_X1 U582 ( .A1(n552), .A2(n448), .ZN(n569) );
  NAND2_X2 U583 ( .A1(n425), .A2(n727), .ZN(n732) );
  NAND2_X1 U584 ( .A1(n732), .A2(n442), .ZN(n742) );
  XNOR2_X1 U585 ( .A(n413), .B(n412), .ZN(G51) );
  XNOR2_X1 U586 ( .A(n422), .B(n523), .ZN(n578) );
  XNOR2_X1 U587 ( .A(n441), .B(n368), .ZN(n440) );
  XNOR2_X1 U588 ( .A(n471), .B(n470), .ZN(n552) );
  NAND2_X1 U589 ( .A1(n451), .A2(n452), .ZN(n457) );
  NOR2_X1 U590 ( .A1(n457), .A2(n455), .ZN(n456) );
  NAND2_X1 U591 ( .A1(n511), .A2(n509), .ZN(n508) );
  NOR2_X1 U592 ( .A1(n419), .A2(n780), .ZN(G63) );
  NAND2_X1 U593 ( .A1(n440), .A2(n417), .ZN(n439) );
  NAND2_X1 U594 ( .A1(n685), .A2(n359), .ZN(n499) );
  XNOR2_X2 U595 ( .A(n420), .B(G146), .ZN(n576) );
  NAND2_X1 U596 ( .A1(n678), .A2(KEYINPUT44), .ZN(n432) );
  NAND2_X1 U597 ( .A1(n670), .A2(n356), .ZN(n421) );
  NAND2_X1 U598 ( .A1(n514), .A2(n461), .ZN(n451) );
  XNOR2_X1 U599 ( .A(n576), .B(n423), .ZN(n422) );
  NAND2_X1 U600 ( .A1(n726), .A2(n725), .ZN(n425) );
  AND2_X1 U601 ( .A1(n427), .A2(n690), .ZN(n428) );
  NAND2_X1 U602 ( .A1(n430), .A2(n706), .ZN(n427) );
  NOR2_X1 U603 ( .A1(n675), .A2(n706), .ZN(n744) );
  NAND2_X1 U604 ( .A1(n429), .A2(n428), .ZN(n431) );
  NAND2_X1 U605 ( .A1(n675), .A2(n430), .ZN(n429) );
  NOR2_X1 U606 ( .A1(n432), .A2(KEYINPUT81), .ZN(n501) );
  NAND2_X1 U607 ( .A1(n432), .A2(n503), .ZN(n474) );
  AND2_X1 U608 ( .A1(n661), .A2(n437), .ZN(n677) );
  NAND2_X1 U609 ( .A1(n757), .A2(n438), .ZN(n641) );
  INV_X1 U610 ( .A(n661), .ZN(n438) );
  XNOR2_X1 U611 ( .A(n439), .B(KEYINPUT63), .ZN(G57) );
  AND2_X1 U612 ( .A1(n776), .A2(G469), .ZN(n771) );
  NAND2_X1 U613 ( .A1(n444), .A2(n463), .ZN(n447) );
  XNOR2_X2 U614 ( .A(n659), .B(n364), .ZN(n444) );
  XNOR2_X2 U615 ( .A(n445), .B(KEYINPUT39), .ZN(n646) );
  XNOR2_X2 U616 ( .A(n526), .B(n365), .ZN(n788) );
  XNOR2_X2 U617 ( .A(n447), .B(n446), .ZN(n805) );
  XNOR2_X1 U618 ( .A(n578), .B(n577), .ZN(n582) );
  NAND2_X1 U619 ( .A1(n508), .A2(n461), .ZN(n453) );
  NAND2_X1 U620 ( .A1(n456), .A2(n458), .ZN(G75) );
  NOR2_X1 U621 ( .A1(n514), .A2(n508), .ZN(n462) );
  NAND2_X1 U622 ( .A1(n462), .A2(n459), .ZN(n458) );
  AND2_X1 U623 ( .A1(n507), .A2(n723), .ZN(n459) );
  XNOR2_X1 U624 ( .A(n400), .B(n465), .ZN(n672) );
  NAND2_X1 U625 ( .A1(n686), .A2(n687), .ZN(n692) );
  INV_X1 U626 ( .A(n687), .ZN(n468) );
  NAND2_X1 U627 ( .A1(n697), .A2(n750), .ZN(n620) );
  NAND2_X1 U628 ( .A1(n660), .A2(n687), .ZN(n471) );
  NAND2_X1 U629 ( .A1(n494), .A2(n492), .ZN(n488) );
  NOR2_X1 U630 ( .A1(n672), .A2(n673), .ZN(n674) );
  XNOR2_X1 U631 ( .A(n724), .B(n472), .ZN(n726) );
  NAND2_X1 U632 ( .A1(n494), .A2(n362), .ZN(n500) );
  NAND2_X1 U633 ( .A1(n500), .A2(n491), .ZN(n490) );
  NAND2_X1 U634 ( .A1(n474), .A2(n525), .ZN(n502) );
  XNOR2_X2 U635 ( .A(n577), .B(n532), .ZN(n486) );
  XNOR2_X2 U636 ( .A(n598), .B(KEYINPUT4), .ZN(n577) );
  XNOR2_X2 U637 ( .A(n531), .B(n530), .ZN(n598) );
  XNOR2_X1 U638 ( .A(n598), .B(n479), .ZN(n478) );
  NAND2_X1 U639 ( .A1(n597), .A2(G217), .ZN(n482) );
  NAND2_X1 U640 ( .A1(n805), .A2(n493), .ZN(n489) );
  NOR2_X1 U641 ( .A1(n805), .A2(n493), .ZN(n491) );
  XNOR2_X1 U642 ( .A(n793), .B(n496), .ZN(n495) );
  XNOR2_X1 U643 ( .A(n562), .B(n497), .ZN(n496) );
  XNOR2_X1 U644 ( .A(n500), .B(G110), .ZN(G12) );
  NAND2_X1 U645 ( .A1(n505), .A2(n803), .ZN(n504) );
  NAND2_X1 U646 ( .A1(n517), .A2(n363), .ZN(n507) );
  INV_X1 U647 ( .A(n721), .ZN(n510) );
  INV_X1 U648 ( .A(n515), .ZN(n512) );
  INV_X1 U649 ( .A(n730), .ZN(n513) );
  INV_X1 U650 ( .A(KEYINPUT123), .ZN(n516) );
  INV_X1 U651 ( .A(KEYINPUT1), .ZN(n522) );
  XNOR2_X1 U652 ( .A(n575), .B(n574), .ZN(n523) );
  NAND2_X1 U653 ( .A1(n749), .A2(n655), .ZN(n656) );
  XNOR2_X2 U654 ( .A(n636), .B(KEYINPUT19), .ZN(n749) );
  XNOR2_X2 U655 ( .A(n591), .B(n590), .ZN(n622) );
  NAND2_X1 U656 ( .A1(n524), .A2(n360), .ZN(n526) );
  XOR2_X1 U657 ( .A(KEYINPUT36), .B(KEYINPUT83), .Z(n528) );
  AND2_X1 U658 ( .A1(n754), .A2(n632), .ZN(n529) );
  XNOR2_X2 U659 ( .A(G143), .B(KEYINPUT64), .ZN(n531) );
  XOR2_X1 U660 ( .A(KEYINPUT3), .B(G101), .Z(n534) );
  XNOR2_X1 U661 ( .A(G146), .B(G137), .ZN(n535) );
  INV_X1 U662 ( .A(G902), .ZN(n539) );
  NAND2_X1 U663 ( .A1(n539), .A2(n538), .ZN(n587) );
  XOR2_X1 U664 ( .A(KEYINPUT14), .B(KEYINPUT87), .Z(n541) );
  XNOR2_X1 U665 ( .A(n541), .B(n540), .ZN(n542) );
  NAND2_X1 U666 ( .A1(n542), .A2(G952), .ZN(n716) );
  NOR2_X1 U667 ( .A1(n716), .A2(G953), .ZN(n653) );
  NAND2_X1 U668 ( .A1(G902), .A2(n542), .ZN(n651) );
  OR2_X1 U669 ( .A1(n722), .A2(n651), .ZN(n543) );
  NOR2_X1 U670 ( .A1(n543), .A2(G900), .ZN(n544) );
  XNOR2_X1 U671 ( .A(G107), .B(n545), .ZN(n781) );
  XNOR2_X1 U672 ( .A(KEYINPUT67), .B(n781), .ZN(n580) );
  NAND2_X1 U673 ( .A1(G227), .A2(n722), .ZN(n546) );
  XNOR2_X1 U674 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U675 ( .A(n580), .B(n548), .ZN(n549) );
  XNOR2_X1 U676 ( .A(n795), .B(n549), .ZN(n769) );
  XOR2_X1 U677 ( .A(KEYINPUT66), .B(G469), .Z(n550) );
  XOR2_X1 U678 ( .A(KEYINPUT23), .B(G119), .Z(n554) );
  XNOR2_X1 U679 ( .A(n554), .B(n553), .ZN(n562) );
  XOR2_X1 U680 ( .A(n555), .B(KEYINPUT91), .Z(n559) );
  NAND2_X1 U681 ( .A1(n722), .A2(G234), .ZN(n557) );
  XNOR2_X1 U682 ( .A(KEYINPUT77), .B(KEYINPUT8), .ZN(n556) );
  XNOR2_X1 U683 ( .A(n557), .B(n556), .ZN(n597) );
  NAND2_X1 U684 ( .A1(G221), .A2(n597), .ZN(n558) );
  XNOR2_X1 U685 ( .A(n559), .B(n558), .ZN(n561) );
  INV_X1 U686 ( .A(KEYINPUT92), .ZN(n560) );
  XNOR2_X1 U687 ( .A(G902), .B(KEYINPUT15), .ZN(n728) );
  NAND2_X1 U688 ( .A1(G234), .A2(n728), .ZN(n563) );
  XNOR2_X1 U689 ( .A(KEYINPUT20), .B(n563), .ZN(n567) );
  NAND2_X1 U690 ( .A1(G217), .A2(n567), .ZN(n564) );
  XNOR2_X2 U691 ( .A(n566), .B(n565), .ZN(n699) );
  NAND2_X1 U692 ( .A1(n567), .A2(G221), .ZN(n568) );
  XOR2_X1 U693 ( .A(n568), .B(KEYINPUT21), .Z(n698) );
  INV_X1 U694 ( .A(KEYINPUT17), .ZN(n570) );
  NAND2_X1 U695 ( .A1(n570), .A2(KEYINPUT84), .ZN(n573) );
  NAND2_X1 U696 ( .A1(n571), .A2(KEYINPUT17), .ZN(n572) );
  NAND2_X1 U697 ( .A1(n573), .A2(n572), .ZN(n575) );
  INV_X1 U698 ( .A(n582), .ZN(n579) );
  NAND2_X1 U699 ( .A1(n579), .A2(n580), .ZN(n584) );
  INV_X1 U700 ( .A(n580), .ZN(n581) );
  NAND2_X1 U701 ( .A1(n582), .A2(n581), .ZN(n583) );
  NAND2_X1 U702 ( .A1(n584), .A2(n583), .ZN(n586) );
  XOR2_X1 U703 ( .A(KEYINPUT16), .B(KEYINPUT68), .Z(n585) );
  NAND2_X1 U704 ( .A1(n587), .A2(G210), .ZN(n589) );
  INV_X1 U705 ( .A(KEYINPUT86), .ZN(n588) );
  INV_X1 U706 ( .A(KEYINPUT38), .ZN(n592) );
  XOR2_X1 U707 ( .A(G134), .B(G122), .Z(n594) );
  XOR2_X1 U708 ( .A(KEYINPUT99), .B(KEYINPUT100), .Z(n596) );
  XNOR2_X1 U709 ( .A(n599), .B(G478), .ZN(n600) );
  XNOR2_X1 U710 ( .A(n602), .B(n601), .ZN(n603) );
  XNOR2_X1 U711 ( .A(n793), .B(n603), .ZN(n607) );
  XOR2_X1 U712 ( .A(KEYINPUT98), .B(KEYINPUT13), .Z(n609) );
  XNOR2_X1 U713 ( .A(KEYINPUT97), .B(G475), .ZN(n608) );
  INV_X1 U714 ( .A(n627), .ZN(n611) );
  NAND2_X1 U715 ( .A1(n628), .A2(n611), .ZN(n612) );
  INV_X1 U716 ( .A(n633), .ZN(n613) );
  NAND2_X1 U717 ( .A1(n646), .A2(n613), .ZN(n615) );
  INV_X1 U718 ( .A(KEYINPUT40), .ZN(n614) );
  XNOR2_X1 U719 ( .A(n615), .B(n614), .ZN(n737) );
  XOR2_X1 U720 ( .A(KEYINPUT113), .B(KEYINPUT28), .Z(n616) );
  XNOR2_X1 U721 ( .A(KEYINPUT115), .B(KEYINPUT42), .ZN(n619) );
  XNOR2_X1 U722 ( .A(n620), .B(n619), .ZN(n806) );
  INV_X1 U723 ( .A(n628), .ZN(n621) );
  AND2_X1 U724 ( .A1(n621), .A2(n627), .ZN(n759) );
  XNOR2_X1 U725 ( .A(KEYINPUT103), .B(n759), .ZN(n647) );
  NAND2_X1 U726 ( .A1(n647), .A2(n633), .ZN(n690) );
  AND2_X1 U727 ( .A1(n749), .A2(n690), .ZN(n623) );
  NAND2_X1 U728 ( .A1(n623), .A2(n750), .ZN(n631) );
  NAND2_X1 U729 ( .A1(n625), .A2(n643), .ZN(n626) );
  XNOR2_X1 U730 ( .A(n626), .B(KEYINPUT112), .ZN(n630) );
  NOR2_X1 U731 ( .A1(n628), .A2(n627), .ZN(n665) );
  INV_X1 U732 ( .A(n665), .ZN(n629) );
  OR2_X1 U733 ( .A1(n630), .A2(n629), .ZN(n754) );
  NAND2_X1 U734 ( .A1(n631), .A2(KEYINPUT69), .ZN(n632) );
  XNOR2_X1 U735 ( .A(KEYINPUT104), .B(KEYINPUT6), .ZN(n635) );
  XNOR2_X1 U736 ( .A(n706), .B(n635), .ZN(n661) );
  AND2_X1 U737 ( .A1(n676), .A2(n698), .ZN(n637) );
  AND2_X1 U738 ( .A1(n637), .A2(n356), .ZN(n640) );
  XNOR2_X1 U739 ( .A(n638), .B(n528), .ZN(n639) );
  NAND2_X1 U740 ( .A1(n639), .A2(n450), .ZN(n765) );
  NAND2_X1 U741 ( .A1(n640), .A2(n687), .ZN(n642) );
  INV_X1 U742 ( .A(KEYINPUT80), .ZN(n645) );
  BUF_X1 U743 ( .A(n646), .Z(n649) );
  INV_X1 U744 ( .A(n647), .ZN(n648) );
  NAND2_X1 U745 ( .A1(n649), .A2(n648), .ZN(n736) );
  XNOR2_X2 U746 ( .A(n650), .B(KEYINPUT78), .ZN(n724) );
  XOR2_X1 U747 ( .A(G898), .B(KEYINPUT88), .Z(n787) );
  NAND2_X1 U748 ( .A1(G953), .A2(n787), .ZN(n784) );
  NOR2_X1 U749 ( .A1(n651), .A2(n784), .ZN(n652) );
  NOR2_X1 U750 ( .A1(n653), .A2(n652), .ZN(n654) );
  XNOR2_X1 U751 ( .A(KEYINPUT89), .B(n654), .ZN(n655) );
  NAND2_X1 U752 ( .A1(n658), .A2(n358), .ZN(n659) );
  XOR2_X1 U753 ( .A(KEYINPUT34), .B(KEYINPUT73), .Z(n664) );
  NAND2_X1 U754 ( .A1(n667), .A2(n706), .ZN(n668) );
  INV_X1 U755 ( .A(n670), .ZN(n701) );
  OR2_X1 U756 ( .A1(n701), .A2(n449), .ZN(n673) );
  XNOR2_X1 U757 ( .A(n674), .B(KEYINPUT93), .ZN(n675) );
  INV_X1 U758 ( .A(KEYINPUT79), .ZN(n679) );
  NOR2_X1 U759 ( .A1(n724), .A2(n788), .ZN(n681) );
  NOR2_X2 U760 ( .A1(n681), .A2(n680), .ZN(n682) );
  NAND2_X1 U761 ( .A1(n736), .A2(KEYINPUT2), .ZN(n683) );
  BUF_X1 U762 ( .A(n684), .Z(n685) );
  NOR2_X1 U763 ( .A1(n687), .A2(n686), .ZN(n688) );
  NOR2_X1 U764 ( .A1(n689), .A2(n688), .ZN(n694) );
  INV_X1 U765 ( .A(n690), .ZN(n691) );
  NOR2_X1 U766 ( .A1(n692), .A2(n691), .ZN(n693) );
  NOR2_X1 U767 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U768 ( .A(n695), .B(KEYINPUT122), .ZN(n696) );
  NOR2_X1 U769 ( .A1(n718), .A2(n696), .ZN(n713) );
  INV_X1 U770 ( .A(n697), .ZN(n717) );
  NOR2_X1 U771 ( .A1(n437), .A2(n698), .ZN(n700) );
  XNOR2_X1 U772 ( .A(KEYINPUT49), .B(n700), .ZN(n705) );
  XOR2_X1 U773 ( .A(KEYINPUT50), .B(KEYINPUT121), .Z(n703) );
  NAND2_X1 U774 ( .A1(n701), .A2(n464), .ZN(n702) );
  XNOR2_X1 U775 ( .A(n703), .B(n702), .ZN(n704) );
  NAND2_X1 U776 ( .A1(n705), .A2(n704), .ZN(n707) );
  NOR2_X1 U777 ( .A1(n707), .A2(n706), .ZN(n708) );
  NOR2_X1 U778 ( .A1(n709), .A2(n708), .ZN(n710) );
  XOR2_X1 U779 ( .A(KEYINPUT51), .B(n710), .Z(n711) );
  NOR2_X1 U780 ( .A1(n717), .A2(n711), .ZN(n712) );
  NOR2_X1 U781 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U782 ( .A(n714), .B(KEYINPUT52), .ZN(n715) );
  NOR2_X1 U783 ( .A1(n716), .A2(n715), .ZN(n720) );
  NOR2_X1 U784 ( .A1(n718), .A2(n717), .ZN(n719) );
  NOR2_X1 U785 ( .A1(n720), .A2(n719), .ZN(n721) );
  INV_X1 U786 ( .A(KEYINPUT53), .ZN(n723) );
  INV_X1 U787 ( .A(n788), .ZN(n725) );
  INV_X1 U788 ( .A(KEYINPUT2), .ZN(n727) );
  INV_X1 U789 ( .A(n728), .ZN(n729) );
  INV_X1 U790 ( .A(G952), .ZN(n734) );
  AND2_X1 U791 ( .A1(n734), .A2(G953), .ZN(n780) );
  XNOR2_X1 U792 ( .A(G134), .B(KEYINPUT120), .ZN(n735) );
  XNOR2_X1 U793 ( .A(n736), .B(n735), .ZN(G36) );
  BUF_X1 U794 ( .A(n737), .Z(n738) );
  XOR2_X1 U795 ( .A(G131), .B(n738), .Z(G33) );
  BUF_X1 U796 ( .A(n739), .Z(n741) );
  XNOR2_X1 U797 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n740) );
  NAND2_X1 U798 ( .A1(n744), .A2(n757), .ZN(n743) );
  XNOR2_X1 U799 ( .A(n743), .B(G104), .ZN(G6) );
  NAND2_X1 U800 ( .A1(n744), .A2(n759), .ZN(n745) );
  XNOR2_X1 U801 ( .A(n745), .B(KEYINPUT27), .ZN(n746) );
  XOR2_X1 U802 ( .A(n746), .B(KEYINPUT26), .Z(n748) );
  XNOR2_X1 U803 ( .A(G107), .B(KEYINPUT116), .ZN(n747) );
  XNOR2_X1 U804 ( .A(n748), .B(n747), .ZN(G9) );
  XOR2_X1 U805 ( .A(KEYINPUT29), .B(KEYINPUT117), .Z(n752) );
  AND2_X1 U806 ( .A1(n749), .A2(n750), .ZN(n755) );
  NAND2_X1 U807 ( .A1(n755), .A2(n759), .ZN(n751) );
  XNOR2_X1 U808 ( .A(n752), .B(n751), .ZN(n753) );
  XOR2_X1 U809 ( .A(G128), .B(n753), .Z(G30) );
  XNOR2_X1 U810 ( .A(G143), .B(n754), .ZN(G45) );
  NAND2_X1 U811 ( .A1(n755), .A2(n757), .ZN(n756) );
  XNOR2_X1 U812 ( .A(n756), .B(G146), .ZN(G48) );
  NAND2_X1 U813 ( .A1(n760), .A2(n757), .ZN(n758) );
  XNOR2_X1 U814 ( .A(n758), .B(G113), .ZN(G15) );
  XOR2_X1 U815 ( .A(KEYINPUT118), .B(KEYINPUT119), .Z(n762) );
  NAND2_X1 U816 ( .A1(n760), .A2(n759), .ZN(n761) );
  XNOR2_X1 U817 ( .A(n762), .B(n761), .ZN(n763) );
  XNOR2_X1 U818 ( .A(G116), .B(n763), .ZN(G18) );
  XOR2_X1 U819 ( .A(G125), .B(KEYINPUT37), .Z(n764) );
  XNOR2_X1 U820 ( .A(n765), .B(n764), .ZN(G27) );
  XOR2_X1 U821 ( .A(KEYINPUT124), .B(KEYINPUT125), .Z(n767) );
  XNOR2_X1 U822 ( .A(KEYINPUT58), .B(KEYINPUT57), .ZN(n766) );
  XNOR2_X1 U823 ( .A(n767), .B(n766), .ZN(n768) );
  XNOR2_X1 U824 ( .A(n769), .B(n768), .ZN(n770) );
  XNOR2_X1 U825 ( .A(n771), .B(n770), .ZN(n772) );
  NOR2_X1 U826 ( .A1(n780), .A2(n772), .ZN(G54) );
  NAND2_X1 U827 ( .A1(n776), .A2(G478), .ZN(n774) );
  NAND2_X1 U828 ( .A1(n776), .A2(G217), .ZN(n778) );
  XNOR2_X1 U829 ( .A(n778), .B(n777), .ZN(n779) );
  NOR2_X1 U830 ( .A1(n780), .A2(n779), .ZN(G66) );
  XOR2_X1 U831 ( .A(n782), .B(n781), .Z(n783) );
  NAND2_X1 U832 ( .A1(n784), .A2(n783), .ZN(n792) );
  NAND2_X1 U833 ( .A1(G953), .A2(G224), .ZN(n785) );
  XOR2_X1 U834 ( .A(KEYINPUT61), .B(n785), .Z(n786) );
  NOR2_X1 U835 ( .A1(n787), .A2(n786), .ZN(n790) );
  NOR2_X1 U836 ( .A1(G953), .A2(n788), .ZN(n789) );
  NOR2_X1 U837 ( .A1(n790), .A2(n789), .ZN(n791) );
  XNOR2_X1 U838 ( .A(n792), .B(n791), .ZN(G69) );
  XOR2_X1 U839 ( .A(n793), .B(KEYINPUT126), .Z(n794) );
  XNOR2_X1 U840 ( .A(n795), .B(n794), .ZN(n798) );
  XNOR2_X1 U841 ( .A(n410), .B(n798), .ZN(n797) );
  NAND2_X1 U842 ( .A1(n797), .A2(n722), .ZN(n802) );
  XNOR2_X1 U843 ( .A(G227), .B(n798), .ZN(n799) );
  NAND2_X1 U844 ( .A1(n799), .A2(G900), .ZN(n800) );
  NAND2_X1 U845 ( .A1(n800), .A2(G953), .ZN(n801) );
  NAND2_X1 U846 ( .A1(n802), .A2(n801), .ZN(G72) );
  XNOR2_X1 U847 ( .A(G140), .B(n803), .ZN(G42) );
  XNOR2_X1 U848 ( .A(n804), .B(G101), .ZN(G3) );
  XOR2_X1 U849 ( .A(n805), .B(G119), .Z(G21) );
  XNOR2_X1 U850 ( .A(G137), .B(KEYINPUT127), .ZN(n808) );
  BUF_X1 U851 ( .A(n806), .Z(n807) );
  XNOR2_X1 U852 ( .A(n808), .B(n807), .ZN(G39) );
endmodule

