//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 0 0 1 0 0 1 1 1 1 0 1 1 1 1 0 1 0 0 0 0 1 1 0 1 1 1 0 0 0 0 0 1 0 1 1 0 1 0 0 0 0 1 1 0 0 0 1 0 0 0 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:31 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n716, new_n717,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n754, new_n755, new_n756, new_n757,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n792, new_n793, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT82), .ZN(new_n189));
  INV_X1    g003(.A(G146), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G143), .ZN(new_n191));
  INV_X1    g005(.A(G143), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G146), .ZN(new_n193));
  OR2_X1    g007(.A1(KEYINPUT0), .A2(G128), .ZN(new_n194));
  NAND2_X1  g008(.A1(KEYINPUT0), .A2(G128), .ZN(new_n195));
  AOI22_X1  g009(.A1(new_n191), .A2(new_n193), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n191), .A2(new_n193), .A3(new_n195), .ZN(new_n197));
  INV_X1    g011(.A(new_n197), .ZN(new_n198));
  OAI21_X1  g012(.A(G125), .B1(new_n196), .B2(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n191), .A2(new_n193), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n191), .A2(KEYINPUT1), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n200), .A2(new_n201), .A3(G128), .ZN(new_n202));
  INV_X1    g016(.A(G125), .ZN(new_n203));
  INV_X1    g017(.A(G128), .ZN(new_n204));
  OAI211_X1 g018(.A(new_n191), .B(new_n193), .C1(KEYINPUT1), .C2(new_n204), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n202), .A2(new_n203), .A3(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n199), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G953), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G224), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(KEYINPUT7), .ZN(new_n210));
  INV_X1    g024(.A(new_n210), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n189), .B1(new_n207), .B2(new_n211), .ZN(new_n212));
  AOI211_X1 g026(.A(KEYINPUT82), .B(new_n210), .C1(new_n199), .C2(new_n206), .ZN(new_n213));
  OAI22_X1  g027(.A1(new_n212), .A2(new_n213), .B1(new_n207), .B2(new_n211), .ZN(new_n214));
  INV_X1    g028(.A(G116), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n215), .A2(G119), .ZN(new_n216));
  XNOR2_X1  g030(.A(KEYINPUT65), .B(G116), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n216), .B1(new_n217), .B2(G119), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(KEYINPUT5), .ZN(new_n219));
  INV_X1    g033(.A(new_n216), .ZN(new_n220));
  OAI211_X1 g034(.A(new_n219), .B(G113), .C1(KEYINPUT5), .C2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT66), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n215), .A2(KEYINPUT65), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT65), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(G116), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n223), .A2(new_n225), .A3(G119), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(new_n220), .ZN(new_n227));
  OAI21_X1  g041(.A(KEYINPUT64), .B1(KEYINPUT2), .B2(G113), .ZN(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  NOR3_X1   g043(.A1(KEYINPUT64), .A2(KEYINPUT2), .A3(G113), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT2), .ZN(new_n231));
  INV_X1    g045(.A(G113), .ZN(new_n232));
  OAI22_X1  g046(.A1(new_n229), .A2(new_n230), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n222), .B1(new_n227), .B2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT64), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n235), .A2(new_n231), .A3(new_n232), .ZN(new_n236));
  AOI22_X1  g050(.A1(new_n236), .A2(new_n228), .B1(KEYINPUT2), .B2(G113), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n218), .A2(KEYINPUT66), .A3(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n234), .A2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT77), .ZN(new_n240));
  INV_X1    g054(.A(G107), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n240), .B1(new_n241), .B2(G104), .ZN(new_n242));
  INV_X1    g056(.A(G104), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n243), .A2(KEYINPUT77), .A3(G107), .ZN(new_n244));
  AND2_X1   g058(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  OAI21_X1  g059(.A(KEYINPUT3), .B1(new_n243), .B2(G107), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT3), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n247), .A2(new_n241), .A3(G104), .ZN(new_n248));
  AND2_X1   g062(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(G101), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n245), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n243), .A2(G107), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT78), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n253), .B1(G104), .B2(new_n241), .ZN(new_n254));
  NOR3_X1   g068(.A1(new_n243), .A2(KEYINPUT78), .A3(G107), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n252), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G101), .ZN(new_n257));
  AND2_X1   g071(.A1(new_n251), .A2(new_n257), .ZN(new_n258));
  AND3_X1   g072(.A1(new_n221), .A2(new_n239), .A3(new_n258), .ZN(new_n259));
  AOI22_X1  g073(.A1(new_n234), .A2(new_n238), .B1(new_n233), .B2(new_n227), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n242), .A2(new_n246), .A3(new_n248), .A4(new_n244), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n261), .A2(new_n262), .A3(G101), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n250), .B1(new_n245), .B2(new_n249), .ZN(new_n264));
  OAI21_X1  g078(.A(KEYINPUT4), .B1(new_n261), .B2(G101), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n263), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n260), .A2(new_n266), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n259), .A2(new_n267), .ZN(new_n268));
  XNOR2_X1  g082(.A(G110), .B(G122), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n214), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  XNOR2_X1  g084(.A(new_n269), .B(KEYINPUT8), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n258), .B1(new_n221), .B2(new_n239), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n271), .B1(new_n259), .B2(new_n272), .ZN(new_n273));
  AOI21_X1  g087(.A(G902), .B1(new_n270), .B2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(new_n269), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n275), .B1(new_n259), .B2(new_n267), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n221), .A2(new_n239), .A3(new_n258), .ZN(new_n277));
  OAI211_X1 g091(.A(new_n277), .B(new_n269), .C1(new_n260), .C2(new_n266), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n276), .A2(KEYINPUT6), .A3(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT6), .ZN(new_n280));
  OAI211_X1 g094(.A(new_n280), .B(new_n275), .C1(new_n259), .C2(new_n267), .ZN(new_n281));
  XNOR2_X1  g095(.A(new_n207), .B(new_n209), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n279), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n274), .A2(new_n283), .ZN(new_n284));
  OAI21_X1  g098(.A(G210), .B1(G237), .B2(G902), .ZN(new_n285));
  XOR2_X1   g099(.A(new_n285), .B(KEYINPUT83), .Z(new_n286));
  NAND2_X1  g100(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(new_n286), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n274), .A2(new_n283), .A3(new_n288), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n188), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT84), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  AND3_X1   g106(.A1(new_n274), .A2(new_n283), .A3(new_n288), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n288), .B1(new_n274), .B2(new_n283), .ZN(new_n294));
  OAI211_X1 g108(.A(new_n291), .B(new_n187), .C1(new_n293), .C2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  XNOR2_X1  g110(.A(G125), .B(G140), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT87), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(KEYINPUT19), .ZN(new_n299));
  OR2_X1    g113(.A1(new_n298), .A2(KEYINPUT19), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n297), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n301), .B1(new_n297), .B2(new_n300), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(new_n190), .ZN(new_n303));
  INV_X1    g117(.A(G140), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(G125), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n305), .A2(KEYINPUT16), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n306), .B1(new_n297), .B2(KEYINPUT16), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(G146), .ZN(new_n308));
  INV_X1    g122(.A(G237), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n309), .A2(new_n208), .A3(G214), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(new_n192), .ZN(new_n311));
  NOR2_X1   g125(.A1(G237), .A2(G953), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n312), .A2(G143), .A3(G214), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(G131), .ZN(new_n315));
  INV_X1    g129(.A(G131), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n311), .A2(new_n316), .A3(new_n313), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n303), .A2(new_n308), .A3(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(new_n313), .ZN(new_n321));
  AOI21_X1  g135(.A(G143), .B1(new_n312), .B2(G214), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(KEYINPUT18), .A2(G131), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n297), .A2(new_n190), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n203), .A2(G140), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n305), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(G146), .ZN(new_n328));
  AOI22_X1  g142(.A1(new_n323), .A2(new_n324), .B1(new_n325), .B2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT85), .ZN(new_n330));
  INV_X1    g144(.A(new_n324), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n330), .B1(new_n314), .B2(new_n331), .ZN(new_n332));
  AOI211_X1 g146(.A(KEYINPUT85), .B(new_n324), .C1(new_n311), .C2(new_n313), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n329), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT86), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  OAI211_X1 g150(.A(new_n329), .B(KEYINPUT86), .C1(new_n332), .C2(new_n333), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n320), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  XNOR2_X1  g152(.A(G113), .B(G122), .ZN(new_n339));
  XNOR2_X1  g153(.A(new_n339), .B(new_n243), .ZN(new_n340));
  OAI21_X1  g154(.A(KEYINPUT88), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n337), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n331), .B1(new_n321), .B2(new_n322), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(KEYINPUT85), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n314), .A2(new_n330), .A3(new_n331), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  AOI21_X1  g160(.A(KEYINPUT86), .B1(new_n346), .B2(new_n329), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n319), .B1(new_n342), .B2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT88), .ZN(new_n349));
  INV_X1    g163(.A(new_n340), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n348), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  AND2_X1   g165(.A1(new_n297), .A2(KEYINPUT16), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n190), .B1(new_n352), .B2(new_n306), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n314), .A2(KEYINPUT17), .A3(G131), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n353), .A2(new_n308), .A3(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT89), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND4_X1  g171(.A1(new_n353), .A2(new_n308), .A3(KEYINPUT89), .A4(new_n354), .ZN(new_n358));
  OAI211_X1 g172(.A(new_n357), .B(new_n358), .C1(KEYINPUT17), .C2(new_n318), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n336), .A2(new_n337), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n359), .A2(new_n360), .A3(new_n340), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n341), .A2(new_n351), .A3(new_n361), .ZN(new_n362));
  NOR2_X1   g176(.A1(G475), .A2(G902), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(KEYINPUT20), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT20), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n362), .A2(new_n366), .A3(new_n363), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(G952), .ZN(new_n369));
  AOI211_X1 g183(.A(G953), .B(new_n369), .C1(G234), .C2(G237), .ZN(new_n370));
  INV_X1    g184(.A(G902), .ZN(new_n371));
  AOI211_X1 g185(.A(new_n371), .B(new_n208), .C1(G234), .C2(G237), .ZN(new_n372));
  XNOR2_X1  g186(.A(KEYINPUT21), .B(G898), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n370), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  XNOR2_X1  g189(.A(KEYINPUT9), .B(G234), .ZN(new_n376));
  INV_X1    g190(.A(G217), .ZN(new_n377));
  NOR3_X1   g191(.A1(new_n376), .A2(new_n377), .A3(G953), .ZN(new_n378));
  XOR2_X1   g192(.A(new_n378), .B(KEYINPUT92), .Z(new_n379));
  NAND3_X1  g193(.A1(new_n223), .A2(new_n225), .A3(G122), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT90), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n217), .A2(KEYINPUT90), .A3(G122), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(G122), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(G116), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n384), .A2(new_n241), .A3(new_n386), .ZN(new_n387));
  XNOR2_X1  g201(.A(G128), .B(G143), .ZN(new_n388));
  INV_X1    g202(.A(G134), .ZN(new_n389));
  XNOR2_X1  g203(.A(new_n388), .B(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n387), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n384), .A2(KEYINPUT14), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT14), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n382), .A2(new_n383), .A3(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n392), .A2(new_n386), .A3(new_n394), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n391), .B1(G107), .B2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT91), .ZN(new_n397));
  OAI22_X1  g211(.A1(new_n397), .A2(KEYINPUT13), .B1(new_n192), .B2(G128), .ZN(new_n398));
  AND2_X1   g212(.A1(new_n397), .A2(KEYINPUT13), .ZN(new_n399));
  OAI21_X1  g213(.A(G134), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  XNOR2_X1  g214(.A(new_n400), .B(new_n388), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n380), .A2(new_n381), .ZN(new_n402));
  AOI21_X1  g216(.A(KEYINPUT90), .B1(new_n217), .B2(G122), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(new_n386), .ZN(new_n405));
  OAI21_X1  g219(.A(G107), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n401), .B1(new_n406), .B2(new_n387), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n379), .B1(new_n396), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n395), .A2(G107), .ZN(new_n409));
  INV_X1    g223(.A(new_n391), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(new_n379), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n406), .A2(new_n387), .ZN(new_n413));
  INV_X1    g227(.A(new_n401), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n411), .A2(new_n412), .A3(new_n415), .ZN(new_n416));
  AOI21_X1  g230(.A(G902), .B1(new_n408), .B2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT15), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n417), .A2(KEYINPUT93), .A3(new_n418), .A4(G478), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n408), .A2(new_n416), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n420), .A2(KEYINPUT93), .A3(new_n371), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n418), .A2(G478), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n417), .A2(KEYINPUT93), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n419), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(new_n361), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n340), .B1(new_n359), .B2(new_n360), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n371), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(G475), .ZN(new_n429));
  NAND4_X1  g243(.A1(new_n368), .A2(new_n375), .A3(new_n425), .A4(new_n429), .ZN(new_n430));
  NOR3_X1   g244(.A1(new_n292), .A2(new_n296), .A3(new_n430), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n377), .B1(G234), .B2(new_n371), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT23), .ZN(new_n433));
  INV_X1    g247(.A(G119), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n433), .B1(new_n434), .B2(G128), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(G128), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n204), .A2(KEYINPUT23), .A3(G119), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n435), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(G110), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n439), .B(KEYINPUT71), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n353), .A2(new_n308), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT70), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n442), .B1(new_n434), .B2(G128), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n204), .A2(KEYINPUT70), .A3(G119), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n443), .A2(new_n444), .A3(new_n436), .ZN(new_n445));
  XNOR2_X1  g259(.A(KEYINPUT24), .B(G110), .ZN(new_n446));
  OAI211_X1 g260(.A(new_n440), .B(new_n441), .C1(new_n445), .C2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n445), .A2(new_n446), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(KEYINPUT72), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT72), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n445), .A2(new_n450), .A3(new_n446), .ZN(new_n451));
  OR2_X1    g265(.A1(new_n438), .A2(G110), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n449), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(new_n325), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n454), .B1(new_n307), .B2(G146), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n453), .A2(KEYINPUT73), .A3(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  AOI21_X1  g271(.A(KEYINPUT73), .B1(new_n453), .B2(new_n455), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n447), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  XNOR2_X1  g273(.A(KEYINPUT22), .B(G137), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n208), .A2(G221), .A3(G234), .ZN(new_n461));
  XNOR2_X1  g275(.A(new_n460), .B(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n459), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n453), .A2(new_n455), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT73), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(new_n456), .ZN(new_n467));
  INV_X1    g281(.A(new_n462), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n467), .A2(new_n447), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n463), .A2(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(KEYINPUT25), .B1(new_n470), .B2(new_n371), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT25), .ZN(new_n472));
  AOI211_X1 g286(.A(new_n472), .B(G902), .C1(new_n463), .C2(new_n469), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n432), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n432), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n459), .A2(new_n462), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n468), .B1(new_n467), .B2(new_n447), .ZN(new_n477));
  OAI211_X1 g291(.A(new_n371), .B(new_n475), .C1(new_n476), .C2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(KEYINPUT74), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT74), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n470), .A2(new_n480), .A3(new_n371), .A4(new_n475), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n474), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n227), .A2(new_n233), .ZN(new_n484));
  NOR3_X1   g298(.A1(new_n227), .A2(new_n233), .A3(new_n222), .ZN(new_n485));
  AOI21_X1  g299(.A(KEYINPUT66), .B1(new_n218), .B2(new_n237), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT11), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n488), .B1(new_n389), .B2(G137), .ZN(new_n489));
  INV_X1    g303(.A(G137), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n490), .A2(KEYINPUT11), .A3(G134), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n389), .A2(G137), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n489), .A2(new_n491), .A3(new_n316), .A4(new_n492), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n389), .A2(G137), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n490), .A2(G134), .ZN(new_n495));
  OAI21_X1  g309(.A(G131), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n202), .A2(new_n493), .A3(new_n205), .A4(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n489), .A2(new_n491), .A3(new_n492), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(G131), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n194), .A2(new_n195), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(new_n200), .ZN(new_n502));
  AOI22_X1  g316(.A1(new_n500), .A2(new_n493), .B1(new_n502), .B2(new_n197), .ZN(new_n503));
  NOR3_X1   g317(.A1(new_n498), .A2(new_n503), .A3(KEYINPUT30), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT30), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n500), .A2(new_n493), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n502), .A2(new_n197), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n505), .B1(new_n508), .B2(new_n497), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n487), .B1(new_n504), .B2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT31), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n312), .A2(G210), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n512), .B(KEYINPUT27), .ZN(new_n513));
  XNOR2_X1  g327(.A(KEYINPUT26), .B(G101), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n513), .B(new_n514), .ZN(new_n515));
  NAND4_X1  g329(.A1(new_n239), .A2(new_n508), .A3(new_n484), .A4(new_n497), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n510), .A2(new_n511), .A3(new_n515), .A4(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT67), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  OAI21_X1  g333(.A(KEYINPUT30), .B1(new_n498), .B2(new_n503), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n508), .A2(new_n505), .A3(new_n497), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n260), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(new_n516), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n524), .A2(KEYINPUT67), .A3(new_n511), .A4(new_n515), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n519), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n510), .A2(new_n515), .A3(new_n516), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(KEYINPUT31), .ZN(new_n528));
  INV_X1    g342(.A(new_n515), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT28), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n508), .A2(new_n497), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n487), .A2(new_n531), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n530), .B1(new_n532), .B2(new_n516), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT68), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n534), .B1(new_n516), .B2(new_n530), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  AOI211_X1 g350(.A(new_n534), .B(new_n530), .C1(new_n532), .C2(new_n516), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n529), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n526), .A2(new_n528), .A3(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(G472), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n539), .A2(new_n540), .A3(new_n371), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(KEYINPUT32), .ZN(new_n542));
  AOI22_X1  g356(.A1(new_n239), .A2(new_n484), .B1(new_n508), .B2(new_n497), .ZN(new_n543));
  OAI211_X1 g357(.A(KEYINPUT68), .B(KEYINPUT28), .C1(new_n523), .C2(new_n543), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n544), .B1(new_n533), .B2(new_n535), .ZN(new_n545));
  AOI22_X1  g359(.A1(new_n545), .A2(new_n529), .B1(KEYINPUT31), .B2(new_n527), .ZN(new_n546));
  AOI21_X1  g360(.A(G902), .B1(new_n546), .B2(new_n526), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT32), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n547), .A2(new_n548), .A3(new_n540), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n542), .A2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT29), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n510), .A2(new_n516), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(new_n529), .ZN(new_n553));
  OAI211_X1 g367(.A(new_n551), .B(new_n553), .C1(new_n545), .C2(new_n529), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(KEYINPUT69), .ZN(new_n555));
  OAI21_X1  g369(.A(KEYINPUT28), .B1(new_n523), .B2(new_n543), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n516), .A2(new_n530), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NOR3_X1   g372(.A1(new_n558), .A2(new_n551), .A3(new_n529), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n559), .A2(G902), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n555), .A2(new_n560), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n554), .A2(KEYINPUT69), .ZN(new_n562));
  OAI21_X1  g376(.A(G472), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n483), .B1(new_n550), .B2(new_n563), .ZN(new_n564));
  OAI21_X1  g378(.A(G221), .B1(new_n376), .B2(G902), .ZN(new_n565));
  XNOR2_X1  g379(.A(new_n565), .B(KEYINPUT75), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT80), .ZN(new_n567));
  XOR2_X1   g381(.A(G110), .B(G140), .Z(new_n568));
  XNOR2_X1  g382(.A(new_n568), .B(KEYINPUT76), .ZN(new_n569));
  AND2_X1   g383(.A1(new_n208), .A2(G227), .ZN(new_n570));
  XOR2_X1   g384(.A(new_n569), .B(new_n570), .Z(new_n571));
  INV_X1    g385(.A(KEYINPUT79), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n251), .A2(new_n257), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n202), .A2(new_n205), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n572), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n574), .ZN(new_n576));
  NAND4_X1  g390(.A1(new_n576), .A2(KEYINPUT79), .A3(new_n251), .A4(new_n257), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n573), .A2(new_n574), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n575), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(new_n506), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT12), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n579), .A2(KEYINPUT12), .A3(new_n506), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT10), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n575), .A2(new_n585), .A3(new_n577), .ZN(new_n586));
  OAI211_X1 g400(.A(new_n507), .B(new_n263), .C1(new_n264), .C2(new_n265), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n576), .A2(KEYINPUT10), .A3(new_n251), .A4(new_n257), .ZN(new_n588));
  AND2_X1   g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n506), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n586), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n571), .B1(new_n584), .B2(new_n591), .ZN(new_n592));
  AND3_X1   g406(.A1(new_n586), .A2(new_n589), .A3(new_n590), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n590), .B1(new_n586), .B2(new_n589), .ZN(new_n594));
  INV_X1    g408(.A(new_n571), .ZN(new_n595));
  NOR3_X1   g409(.A1(new_n593), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n567), .B1(new_n592), .B2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n594), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n598), .A2(new_n591), .A3(new_n571), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n593), .B1(new_n583), .B2(new_n582), .ZN(new_n600));
  OAI211_X1 g414(.A(KEYINPUT80), .B(new_n599), .C1(new_n600), .C2(new_n571), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n597), .A2(new_n371), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(G469), .ZN(new_n603));
  NOR3_X1   g417(.A1(new_n593), .A2(new_n594), .A3(new_n571), .ZN(new_n604));
  AND3_X1   g418(.A1(new_n579), .A2(KEYINPUT12), .A3(new_n506), .ZN(new_n605));
  AOI21_X1  g419(.A(KEYINPUT12), .B1(new_n579), .B2(new_n506), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n591), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n604), .B1(new_n607), .B2(new_n571), .ZN(new_n608));
  INV_X1    g422(.A(G469), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n608), .A2(KEYINPUT81), .A3(new_n609), .A4(new_n371), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n607), .A2(new_n571), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n598), .A2(new_n591), .A3(new_n595), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n611), .A2(new_n609), .A3(new_n371), .A4(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT81), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n610), .A2(new_n615), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n566), .B1(new_n603), .B2(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n431), .A2(new_n564), .A3(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(G101), .ZN(G3));
  AOI211_X1 g433(.A(new_n483), .B(new_n566), .C1(new_n603), .C2(new_n616), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n539), .A2(new_n371), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(G472), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT94), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n622), .A2(new_n623), .A3(new_n541), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n621), .A2(KEYINPUT94), .A3(G472), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n620), .A2(new_n626), .ZN(new_n627));
  XOR2_X1   g441(.A(new_n627), .B(KEYINPUT95), .Z(new_n628));
  NAND2_X1  g442(.A1(new_n290), .A2(new_n375), .ZN(new_n629));
  AND3_X1   g443(.A1(new_n362), .A2(new_n366), .A3(new_n363), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n366), .B1(new_n362), .B2(new_n363), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n429), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT33), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n412), .B1(new_n411), .B2(new_n415), .ZN(new_n634));
  NOR3_X1   g448(.A1(new_n396), .A2(new_n407), .A3(new_n379), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n633), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT96), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n634), .A2(KEYINPUT97), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT97), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n408), .A2(new_n640), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n639), .A2(new_n641), .A3(KEYINPUT33), .A4(new_n416), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n420), .A2(KEYINPUT96), .A3(new_n633), .ZN(new_n643));
  AND2_X1   g457(.A1(new_n371), .A2(G478), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n638), .A2(new_n642), .A3(new_n643), .A4(new_n644), .ZN(new_n645));
  OR2_X1    g459(.A1(new_n417), .A2(G478), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n632), .A2(new_n647), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n629), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n628), .A2(new_n649), .ZN(new_n650));
  XOR2_X1   g464(.A(KEYINPUT34), .B(G104), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G6));
  AOI22_X1  g466(.A1(new_n365), .A2(new_n367), .B1(G475), .B2(new_n428), .ZN(new_n653));
  INV_X1    g467(.A(new_n425), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n629), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n628), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g471(.A(KEYINPUT35), .B(G107), .Z(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G9));
  INV_X1    g473(.A(KEYINPUT99), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n371), .B1(new_n476), .B2(new_n477), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(new_n472), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n470), .A2(KEYINPUT25), .A3(new_n371), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n475), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n468), .A2(KEYINPUT36), .ZN(new_n665));
  XOR2_X1   g479(.A(new_n665), .B(KEYINPUT98), .Z(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(new_n459), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n667), .A2(new_n371), .A3(new_n475), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n660), .B1(new_n664), .B2(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n474), .A2(KEYINPUT99), .A3(new_n668), .ZN(new_n671));
  AOI22_X1  g485(.A1(new_n624), .A2(new_n625), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n431), .A2(new_n672), .A3(new_n617), .ZN(new_n673));
  XOR2_X1   g487(.A(KEYINPUT37), .B(G110), .Z(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(G12));
  NOR3_X1   g489(.A1(new_n664), .A2(new_n669), .A3(new_n660), .ZN(new_n676));
  AOI21_X1  g490(.A(KEYINPUT99), .B1(new_n474), .B2(new_n668), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(new_n370), .ZN(new_n679));
  INV_X1    g493(.A(new_n372), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n679), .B1(new_n680), .B2(G900), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(KEYINPUT100), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n653), .A2(new_n654), .A3(new_n683), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n678), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n550), .A2(new_n563), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n685), .A2(new_n686), .A3(new_n617), .A4(new_n290), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G128), .ZN(G30));
  XOR2_X1   g502(.A(new_n682), .B(KEYINPUT39), .Z(new_n689));
  NAND2_X1  g503(.A1(new_n617), .A2(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT40), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n690), .B(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(new_n527), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n515), .B1(new_n532), .B2(new_n516), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n371), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(G472), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n550), .A2(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT102), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n550), .A2(KEYINPUT102), .A3(new_n696), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT103), .ZN(new_n702));
  OAI211_X1 g516(.A(new_n419), .B(new_n187), .C1(new_n423), .C2(new_n424), .ZN(new_n703));
  INV_X1    g517(.A(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(new_n632), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n702), .B1(new_n678), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n670), .A2(new_n671), .ZN(new_n708));
  NOR3_X1   g522(.A1(new_n708), .A2(new_n705), .A3(KEYINPUT103), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n287), .A2(new_n289), .ZN(new_n710));
  XOR2_X1   g524(.A(KEYINPUT101), .B(KEYINPUT38), .Z(new_n711));
  XOR2_X1   g525(.A(new_n710), .B(new_n711), .Z(new_n712));
  NOR3_X1   g526(.A1(new_n707), .A2(new_n709), .A3(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n692), .A2(new_n701), .A3(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G143), .ZN(G45));
  NAND3_X1  g529(.A1(new_n632), .A2(new_n647), .A3(new_n683), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n678), .A2(new_n716), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n717), .A2(new_n686), .A3(new_n617), .A4(new_n290), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G146), .ZN(G48));
  INV_X1    g533(.A(new_n566), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n608), .A2(new_n371), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(G469), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n616), .A2(new_n720), .A3(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT104), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n616), .A2(KEYINPUT104), .A3(new_n720), .A4(new_n722), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n564), .A2(new_n725), .A3(new_n649), .A4(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(KEYINPUT41), .B(G113), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n727), .B(new_n728), .ZN(G15));
  NAND4_X1  g543(.A1(new_n564), .A2(new_n725), .A3(new_n656), .A4(new_n726), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G116), .ZN(G18));
  NOR2_X1   g545(.A1(new_n678), .A2(new_n430), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n187), .B1(new_n293), .B2(new_n294), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n723), .A2(new_n733), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n732), .A2(new_n734), .A3(new_n686), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G119), .ZN(G21));
  INV_X1    g550(.A(new_n483), .ZN(new_n737));
  AOI22_X1  g551(.A1(new_n558), .A2(new_n529), .B1(new_n527), .B2(KEYINPUT31), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n526), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g553(.A1(G472), .A2(G902), .ZN(new_n740));
  AOI21_X1  g554(.A(KEYINPUT105), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT105), .ZN(new_n742));
  INV_X1    g556(.A(new_n740), .ZN(new_n743));
  AOI211_X1 g557(.A(new_n742), .B(new_n743), .C1(new_n526), .C2(new_n738), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n741), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n621), .A2(KEYINPUT106), .A3(G472), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT106), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n747), .B1(new_n547), .B2(new_n540), .ZN(new_n748));
  AND4_X1   g562(.A1(new_n737), .A2(new_n745), .A3(new_n746), .A4(new_n748), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n704), .A2(new_n632), .A3(new_n710), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n750), .A2(new_n374), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n749), .A2(new_n725), .A3(new_n726), .A4(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G122), .ZN(G24));
  XNOR2_X1  g567(.A(new_n716), .B(KEYINPUT107), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n745), .A2(new_n746), .A3(new_n748), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n755), .A2(new_n678), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n754), .A2(new_n756), .A3(new_n734), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G125), .ZN(G27));
  INV_X1    g572(.A(KEYINPUT111), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n542), .A2(new_n549), .A3(new_n759), .ZN(new_n760));
  AND2_X1   g574(.A1(new_n760), .A2(new_n563), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n550), .A2(KEYINPUT111), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n483), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n287), .A2(new_n720), .A3(new_n187), .A4(new_n289), .ZN(new_n764));
  INV_X1    g578(.A(new_n764), .ZN(new_n765));
  AND2_X1   g579(.A1(new_n610), .A2(new_n615), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT108), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n767), .B1(new_n600), .B2(new_n571), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n607), .A2(KEYINPUT108), .A3(new_n595), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n768), .A2(G469), .A3(new_n599), .A4(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(G469), .A2(G902), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n765), .B1(new_n766), .B2(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(KEYINPUT109), .ZN(new_n774));
  AND2_X1   g588(.A1(new_n770), .A2(new_n771), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(new_n616), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT109), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n776), .A2(new_n777), .A3(new_n765), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n774), .A2(new_n778), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n763), .A2(new_n779), .A3(KEYINPUT42), .A4(new_n754), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT42), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n777), .B1(new_n776), .B2(new_n765), .ZN(new_n782));
  AOI211_X1 g596(.A(KEYINPUT109), .B(new_n764), .C1(new_n775), .C2(new_n616), .ZN(new_n783));
  OAI211_X1 g597(.A(new_n754), .B(new_n564), .C1(new_n782), .C2(new_n783), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n781), .B1(new_n784), .B2(KEYINPUT110), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT110), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n686), .A2(new_n737), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n787), .B1(new_n774), .B2(new_n778), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n786), .B1(new_n788), .B2(new_n754), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n780), .B1(new_n785), .B2(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G131), .ZN(G33));
  INV_X1    g605(.A(new_n684), .ZN(new_n792));
  OAI211_X1 g606(.A(new_n564), .B(new_n792), .C1(new_n782), .C2(new_n783), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(G134), .ZN(G36));
  INV_X1    g608(.A(KEYINPUT112), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT45), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n597), .A2(new_n796), .A3(new_n601), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n768), .A2(KEYINPUT45), .A3(new_n599), .A4(new_n769), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n797), .A2(G469), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(new_n771), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT46), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n795), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n800), .A2(new_n795), .A3(new_n801), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n799), .A2(KEYINPUT46), .A3(new_n771), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n803), .A2(new_n616), .A3(new_n804), .A4(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n806), .A2(new_n720), .A3(new_n689), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n653), .A2(new_n647), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n809), .A2(KEYINPUT43), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT43), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n653), .A2(new_n811), .A3(new_n647), .ZN(new_n812));
  AND2_X1   g626(.A1(new_n810), .A2(new_n812), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n626), .A2(new_n678), .ZN(new_n814));
  AND3_X1   g628(.A1(new_n813), .A2(new_n814), .A3(KEYINPUT44), .ZN(new_n815));
  AOI21_X1  g629(.A(KEYINPUT44), .B1(new_n813), .B2(new_n814), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n710), .A2(new_n188), .ZN(new_n817));
  INV_X1    g631(.A(new_n817), .ZN(new_n818));
  NOR3_X1   g632(.A1(new_n815), .A2(new_n816), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n808), .A2(new_n819), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n820), .B(G137), .ZN(G39));
  NOR4_X1   g635(.A1(new_n686), .A2(new_n818), .A3(new_n737), .A4(new_n716), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n806), .A2(KEYINPUT47), .A3(new_n720), .ZN(new_n823));
  INV_X1    g637(.A(new_n823), .ZN(new_n824));
  AOI21_X1  g638(.A(KEYINPUT47), .B1(new_n806), .B2(new_n720), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n822), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n826), .B(G140), .ZN(G42));
  INV_X1    g641(.A(KEYINPUT51), .ZN(new_n828));
  INV_X1    g642(.A(new_n825), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n616), .A2(new_n722), .ZN(new_n830));
  INV_X1    g644(.A(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n831), .A2(new_n566), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n829), .A2(new_n823), .A3(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n810), .A2(new_n812), .A3(new_n370), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n745), .A2(new_n737), .A3(new_n748), .A4(new_n746), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(new_n817), .ZN(new_n837));
  XNOR2_X1  g651(.A(new_n837), .B(KEYINPUT115), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n828), .B1(new_n833), .B2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(new_n723), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n712), .A2(new_n840), .A3(new_n188), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n841), .A2(new_n836), .A3(KEYINPUT50), .ZN(new_n842));
  AOI21_X1  g656(.A(KEYINPUT50), .B1(new_n841), .B2(new_n836), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(new_n701), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n831), .A2(new_n765), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n846), .A2(new_n483), .A3(new_n679), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n632), .A2(new_n647), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n845), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n834), .A2(new_n846), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n850), .A2(KEYINPUT117), .A3(new_n756), .ZN(new_n851));
  AOI21_X1  g665(.A(KEYINPUT117), .B1(new_n850), .B2(new_n756), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n849), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n844), .B1(new_n853), .B2(KEYINPUT118), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT119), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT118), .ZN(new_n856));
  OAI211_X1 g670(.A(new_n856), .B(new_n849), .C1(new_n851), .C2(new_n852), .ZN(new_n857));
  AND3_X1   g671(.A1(new_n854), .A2(new_n855), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n855), .B1(new_n854), .B2(new_n857), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n839), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n850), .A2(new_n763), .ZN(new_n861));
  XOR2_X1   g675(.A(new_n861), .B(KEYINPUT48), .Z(new_n862));
  NAND2_X1  g676(.A1(new_n845), .A2(new_n847), .ZN(new_n863));
  OAI211_X1 g677(.A(G952), .B(new_n208), .C1(new_n863), .C2(new_n648), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n836), .A2(new_n734), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n865), .B(KEYINPUT120), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n862), .A2(new_n864), .A3(new_n866), .ZN(new_n867));
  OR2_X1    g681(.A1(new_n853), .A2(new_n844), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT116), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n869), .B1(new_n829), .B2(new_n823), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n824), .A2(new_n825), .A3(KEYINPUT116), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n832), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n868), .B1(new_n872), .B2(new_n838), .ZN(new_n873));
  OAI211_X1 g687(.A(new_n860), .B(new_n867), .C1(new_n873), .C2(KEYINPUT51), .ZN(new_n874));
  OAI211_X1 g688(.A(new_n754), .B(new_n756), .C1(new_n782), .C2(new_n783), .ZN(new_n875));
  AND2_X1   g689(.A1(new_n617), .A2(new_n686), .ZN(new_n876));
  NOR4_X1   g690(.A1(new_n818), .A2(new_n632), .A3(new_n654), .A4(new_n682), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n876), .A2(new_n877), .A3(new_n708), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n875), .A2(new_n878), .A3(new_n793), .ZN(new_n879));
  OAI211_X1 g693(.A(new_n431), .B(new_n617), .C1(new_n672), .C2(new_n564), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n655), .A2(new_n648), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n733), .A2(KEYINPUT84), .ZN(new_n882));
  AND3_X1   g696(.A1(new_n882), .A2(new_n375), .A3(new_n295), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n620), .A2(new_n626), .A3(new_n881), .A4(new_n883), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n880), .A2(new_n884), .A3(new_n735), .A4(new_n752), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n730), .A2(new_n727), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n879), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  AND2_X1   g701(.A1(new_n887), .A2(new_n790), .ZN(new_n888));
  INV_X1    g702(.A(new_n750), .ZN(new_n889));
  NOR4_X1   g703(.A1(new_n664), .A2(new_n669), .A3(new_n566), .A4(new_n682), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n697), .A2(new_n889), .A3(new_n776), .A4(new_n890), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n757), .A2(new_n687), .A3(new_n718), .A4(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(KEYINPUT52), .ZN(new_n893));
  OAI211_X1 g707(.A(new_n876), .B(new_n290), .C1(new_n685), .C2(new_n717), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT52), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n894), .A2(new_n895), .A3(new_n757), .A4(new_n891), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n893), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(KEYINPUT114), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n687), .A2(new_n718), .ZN(new_n899));
  AOI21_X1  g713(.A(KEYINPUT114), .B1(new_n899), .B2(KEYINPUT52), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n893), .A2(new_n900), .A3(new_n896), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n888), .A2(KEYINPUT53), .A3(new_n898), .A4(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT54), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n887), .A2(new_n790), .A3(new_n893), .A4(new_n896), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT53), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n902), .A2(new_n903), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n904), .A2(KEYINPUT53), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n898), .A2(new_n790), .A3(new_n887), .A4(new_n901), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n908), .B1(new_n909), .B2(KEYINPUT53), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n907), .B1(new_n910), .B2(new_n903), .ZN(new_n911));
  OAI22_X1  g725(.A1(new_n874), .A2(new_n911), .B1(G952), .B2(G953), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n737), .A2(new_n720), .A3(new_n187), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(KEYINPUT113), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n830), .A2(KEYINPUT49), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n712), .A2(new_n653), .A3(new_n915), .A4(new_n647), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n830), .A2(KEYINPUT49), .ZN(new_n917));
  OR4_X1    g731(.A1(new_n701), .A2(new_n914), .A3(new_n916), .A4(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n912), .A2(new_n918), .ZN(G75));
  NAND2_X1  g733(.A1(new_n902), .A2(new_n906), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n920), .A2(G902), .A3(new_n286), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT56), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n279), .A2(new_n281), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(new_n282), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(KEYINPUT55), .ZN(new_n925));
  AND3_X1   g739(.A1(new_n921), .A2(new_n922), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n925), .B1(new_n921), .B2(new_n922), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n369), .A2(G953), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n928), .B(KEYINPUT121), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n929), .B(KEYINPUT122), .Z(new_n930));
  INV_X1    g744(.A(new_n930), .ZN(new_n931));
  NOR3_X1   g745(.A1(new_n926), .A2(new_n927), .A3(new_n931), .ZN(G51));
  XOR2_X1   g746(.A(new_n771), .B(KEYINPUT57), .Z(new_n933));
  AND3_X1   g747(.A1(new_n902), .A2(new_n903), .A3(new_n906), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n903), .B1(new_n902), .B2(new_n906), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n933), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(new_n608), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n920), .A2(G902), .ZN(new_n938));
  OR2_X1    g752(.A1(new_n938), .A2(new_n799), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n929), .B1(new_n937), .B2(new_n939), .ZN(G54));
  NAND2_X1  g754(.A1(KEYINPUT58), .A2(G475), .ZN(new_n941));
  OR3_X1    g755(.A1(new_n938), .A2(new_n362), .A3(new_n941), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n362), .B1(new_n938), .B2(new_n941), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n929), .B1(new_n942), .B2(new_n943), .ZN(G60));
  AND3_X1   g758(.A1(new_n638), .A2(new_n643), .A3(new_n642), .ZN(new_n945));
  NAND2_X1  g759(.A1(G478), .A2(G902), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n946), .B(KEYINPUT59), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n945), .B1(new_n911), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n945), .A2(new_n947), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n920), .A2(KEYINPUT54), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n949), .B1(new_n950), .B2(new_n907), .ZN(new_n951));
  NOR3_X1   g765(.A1(new_n948), .A2(new_n931), .A3(new_n951), .ZN(G63));
  INV_X1    g766(.A(KEYINPUT61), .ZN(new_n953));
  NAND2_X1  g767(.A1(G217), .A2(G902), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n954), .B(KEYINPUT60), .Z(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n956), .B1(new_n902), .B2(new_n906), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n957), .A2(new_n667), .ZN(new_n958));
  INV_X1    g772(.A(new_n958), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n930), .B1(new_n957), .B2(new_n470), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n953), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n920), .A2(new_n955), .ZN(new_n962));
  INV_X1    g776(.A(new_n470), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n964), .A2(KEYINPUT61), .A3(new_n930), .A4(new_n958), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n961), .A2(new_n965), .ZN(G66));
  NOR2_X1   g780(.A1(new_n885), .A2(new_n886), .ZN(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(G224), .A2(G953), .ZN(new_n969));
  OAI22_X1  g783(.A1(new_n968), .A2(G953), .B1(new_n373), .B2(new_n969), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n970), .B(KEYINPUT123), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n923), .B1(G898), .B2(new_n208), .ZN(new_n972));
  XOR2_X1   g786(.A(new_n971), .B(new_n972), .Z(G69));
  NOR2_X1   g787(.A1(new_n504), .A2(new_n509), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n974), .B(new_n302), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n975), .B1(G900), .B2(G953), .ZN(new_n976));
  AND2_X1   g790(.A1(new_n894), .A2(new_n757), .ZN(new_n977));
  AND3_X1   g791(.A1(new_n820), .A2(new_n793), .A3(new_n977), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n808), .A2(new_n889), .A3(new_n763), .ZN(new_n979));
  NAND4_X1  g793(.A1(new_n978), .A2(new_n790), .A3(new_n826), .A4(new_n979), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n976), .B1(new_n980), .B2(G953), .ZN(new_n981));
  INV_X1    g795(.A(KEYINPUT125), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n564), .A2(new_n817), .A3(new_n881), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n983), .A2(new_n690), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n984), .B1(new_n808), .B2(new_n819), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n826), .A2(new_n985), .ZN(new_n986));
  AND3_X1   g800(.A1(new_n977), .A2(new_n714), .A3(KEYINPUT62), .ZN(new_n987));
  AOI21_X1  g801(.A(KEYINPUT62), .B1(new_n977), .B2(new_n714), .ZN(new_n988));
  NOR2_X1   g802(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n982), .B1(new_n986), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n977), .A2(new_n714), .ZN(new_n991));
  INV_X1    g805(.A(KEYINPUT62), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n977), .A2(new_n714), .A3(KEYINPUT62), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n995), .A2(KEYINPUT125), .A3(new_n826), .A4(new_n985), .ZN(new_n996));
  AOI21_X1  g810(.A(G953), .B1(new_n990), .B2(new_n996), .ZN(new_n997));
  XOR2_X1   g811(.A(new_n975), .B(KEYINPUT124), .Z(new_n998));
  OAI21_X1  g812(.A(new_n981), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n208), .B1(G227), .B2(G900), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g815(.A(new_n1000), .ZN(new_n1002));
  OAI211_X1 g816(.A(new_n981), .B(new_n1002), .C1(new_n997), .C2(new_n998), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1001), .A2(new_n1003), .ZN(G72));
  NOR2_X1   g818(.A1(new_n524), .A2(new_n529), .ZN(new_n1005));
  AND3_X1   g819(.A1(new_n990), .A2(new_n967), .A3(new_n996), .ZN(new_n1006));
  XNOR2_X1  g820(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1007));
  NOR2_X1   g821(.A1(new_n540), .A2(new_n371), .ZN(new_n1008));
  XOR2_X1   g822(.A(new_n1007), .B(new_n1008), .Z(new_n1009));
  INV_X1    g823(.A(new_n1009), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n1005), .B1(new_n1006), .B2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n1010), .B1(new_n553), .B2(new_n527), .ZN(new_n1012));
  OAI211_X1 g826(.A(new_n908), .B(new_n1012), .C1(new_n909), .C2(KEYINPUT53), .ZN(new_n1013));
  INV_X1    g827(.A(KEYINPUT127), .ZN(new_n1014));
  XNOR2_X1  g828(.A(new_n1013), .B(new_n1014), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n1009), .B1(new_n980), .B2(new_n968), .ZN(new_n1016));
  NOR2_X1   g830(.A1(new_n552), .A2(new_n515), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n929), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  AND3_X1   g832(.A1(new_n1011), .A2(new_n1015), .A3(new_n1018), .ZN(G57));
endmodule


