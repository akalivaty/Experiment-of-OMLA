

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U550 ( .A1(n719), .A2(G8), .ZN(n720) );
  NAND2_X1 U551 ( .A1(G160), .A2(G40), .ZN(n810) );
  XNOR2_X1 U552 ( .A(n547), .B(KEYINPUT17), .ZN(n903) );
  NAND2_X1 U553 ( .A1(n587), .A2(n583), .ZN(n547) );
  INV_X4 U554 ( .A(G2105), .ZN(n583) );
  BUF_X1 U555 ( .A(n706), .Z(n907) );
  NOR2_X1 U556 ( .A1(n597), .A2(n596), .ZN(G164) );
  NOR2_X2 U557 ( .A1(n725), .A2(n724), .ZN(n727) );
  AND2_X1 U558 ( .A1(n536), .A2(n535), .ZN(n534) );
  NAND2_X1 U559 ( .A1(n517), .A2(n544), .ZN(n533) );
  AND2_X1 U560 ( .A1(n530), .A2(n527), .ZN(n526) );
  NOR2_X1 U561 ( .A1(n753), .A2(n752), .ZN(n735) );
  BUF_X2 U562 ( .A(n903), .Z(n514) );
  OR2_X2 U563 ( .A1(n784), .A2(G1966), .ZN(n772) );
  NOR2_X4 U564 ( .A1(n810), .A2(n716), .ZN(n736) );
  INV_X2 U565 ( .A(n736), .ZN(n719) );
  XNOR2_X2 U566 ( .A(n765), .B(KEYINPUT100), .ZN(n777) );
  OR2_X1 U567 ( .A1(G286), .A2(KEYINPUT102), .ZN(n529) );
  AND2_X1 U568 ( .A1(G286), .A2(KEYINPUT102), .ZN(n531) );
  AND2_X1 U569 ( .A1(n780), .A2(KEYINPUT103), .ZN(n542) );
  NAND2_X1 U570 ( .A1(n525), .A2(n523), .ZN(n522) );
  NOR2_X1 U571 ( .A1(n674), .A2(n559), .ZN(n657) );
  XNOR2_X1 U572 ( .A(n733), .B(n732), .ZN(n752) );
  XNOR2_X1 U573 ( .A(n729), .B(n728), .ZN(n731) );
  NOR2_X1 U574 ( .A1(G2084), .A2(n719), .ZN(n773) );
  NOR2_X1 U575 ( .A1(n524), .A2(KEYINPUT102), .ZN(n523) );
  INV_X1 U576 ( .A(n770), .ZN(n524) );
  NAND2_X1 U577 ( .A1(n518), .A2(n528), .ZN(n527) );
  AND2_X1 U578 ( .A1(n542), .A2(n544), .ZN(n537) );
  NOR2_X1 U579 ( .A1(n780), .A2(KEYINPUT103), .ZN(n539) );
  NOR2_X1 U580 ( .A1(n790), .A2(n541), .ZN(n540) );
  AND2_X1 U581 ( .A1(n790), .A2(n545), .ZN(n538) );
  INV_X1 U582 ( .A(n950), .ZN(n787) );
  AND2_X1 U583 ( .A1(n784), .A2(n553), .ZN(n552) );
  XOR2_X1 U584 ( .A(n616), .B(KEYINPUT15), .Z(n946) );
  NOR2_X1 U585 ( .A1(n609), .A2(n608), .ZN(n748) );
  NOR2_X1 U586 ( .A1(G651), .A2(G543), .ZN(n660) );
  NAND2_X1 U587 ( .A1(n713), .A2(n712), .ZN(n714) );
  OR2_X1 U588 ( .A1(n796), .A2(n795), .ZN(n515) );
  AND2_X1 U589 ( .A1(G8), .A2(n721), .ZN(n516) );
  AND2_X1 U590 ( .A1(n791), .A2(n538), .ZN(n517) );
  OR2_X1 U591 ( .A1(n770), .A2(KEYINPUT102), .ZN(n518) );
  OR2_X1 U592 ( .A1(n540), .A2(n539), .ZN(n519) );
  NAND2_X1 U593 ( .A1(n787), .A2(n786), .ZN(n520) );
  OR2_X1 U594 ( .A1(n520), .A2(n552), .ZN(n521) );
  INV_X1 U595 ( .A(KEYINPUT103), .ZN(n545) );
  NAND2_X1 U596 ( .A1(n777), .A2(n531), .ZN(n530) );
  NAND2_X1 U597 ( .A1(n526), .A2(n522), .ZN(n532) );
  INV_X1 U598 ( .A(n777), .ZN(n525) );
  NAND2_X1 U599 ( .A1(n770), .A2(n529), .ZN(n528) );
  NAND2_X1 U600 ( .A1(n532), .A2(G8), .ZN(n771) );
  NAND2_X1 U601 ( .A1(n534), .A2(n533), .ZN(n782) );
  NAND2_X1 U602 ( .A1(n519), .A2(n544), .ZN(n535) );
  NAND2_X1 U603 ( .A1(n543), .A2(n537), .ZN(n536) );
  INV_X1 U604 ( .A(n542), .ZN(n541) );
  INV_X1 U605 ( .A(n791), .ZN(n543) );
  INV_X1 U606 ( .A(n952), .ZN(n544) );
  NAND2_X1 U607 ( .A1(n707), .A2(n546), .ZN(n711) );
  NAND2_X1 U608 ( .A1(n514), .A2(G137), .ZN(n546) );
  NAND2_X1 U609 ( .A1(n548), .A2(n521), .ZN(n549) );
  INV_X1 U610 ( .A(n798), .ZN(n548) );
  NOR2_X1 U611 ( .A1(n798), .A2(KEYINPUT33), .ZN(n551) );
  NAND2_X1 U612 ( .A1(n550), .A2(n549), .ZN(n833) );
  NAND2_X1 U613 ( .A1(n783), .A2(n551), .ZN(n550) );
  INV_X1 U614 ( .A(KEYINPUT33), .ZN(n553) );
  INV_X1 U615 ( .A(G2104), .ZN(n587) );
  NOR2_X2 U616 ( .A1(G2104), .A2(n583), .ZN(n906) );
  XNOR2_X2 U617 ( .A(n771), .B(KEYINPUT32), .ZN(n791) );
  NOR2_X1 U618 ( .A1(G164), .A2(G1384), .ZN(n811) );
  XNOR2_X2 U619 ( .A(n714), .B(KEYINPUT65), .ZN(G160) );
  AND2_X1 U620 ( .A1(n841), .A2(n835), .ZN(n554) );
  INV_X1 U621 ( .A(KEYINPUT31), .ZN(n726) );
  AND2_X2 U622 ( .A1(n583), .A2(G2104), .ZN(n708) );
  NAND2_X1 U623 ( .A1(n554), .A2(n831), .ZN(n832) );
  INV_X1 U624 ( .A(n748), .ZN(n943) );
  NOR2_X1 U625 ( .A1(n577), .A2(n576), .ZN(G171) );
  NAND2_X1 U626 ( .A1(n660), .A2(G89), .ZN(n555) );
  XNOR2_X1 U627 ( .A(n555), .B(KEYINPUT4), .ZN(n557) );
  XOR2_X1 U628 ( .A(G543), .B(KEYINPUT0), .Z(n674) );
  INV_X1 U629 ( .A(G651), .ZN(n559) );
  NAND2_X1 U630 ( .A1(G76), .A2(n657), .ZN(n556) );
  NAND2_X1 U631 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U632 ( .A(n558), .B(KEYINPUT5), .ZN(n567) );
  NOR2_X1 U633 ( .A1(G543), .A2(n559), .ZN(n560) );
  XOR2_X1 U634 ( .A(KEYINPUT1), .B(n560), .Z(n672) );
  NAND2_X1 U635 ( .A1(n672), .A2(G63), .ZN(n561) );
  XNOR2_X1 U636 ( .A(n561), .B(KEYINPUT74), .ZN(n564) );
  NOR2_X1 U637 ( .A1(G651), .A2(n674), .ZN(n562) );
  XNOR2_X2 U638 ( .A(KEYINPUT64), .B(n562), .ZN(n668) );
  NAND2_X1 U639 ( .A1(G51), .A2(n668), .ZN(n563) );
  NAND2_X1 U640 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U641 ( .A(KEYINPUT6), .B(n565), .Z(n566) );
  NAND2_X1 U642 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U643 ( .A(n568), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U644 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U645 ( .A1(G64), .A2(n672), .ZN(n569) );
  XNOR2_X1 U646 ( .A(n569), .B(KEYINPUT68), .ZN(n572) );
  NAND2_X1 U647 ( .A1(n668), .A2(G52), .ZN(n570) );
  XOR2_X1 U648 ( .A(KEYINPUT69), .B(n570), .Z(n571) );
  NAND2_X1 U649 ( .A1(n572), .A2(n571), .ZN(n577) );
  NAND2_X1 U650 ( .A1(G90), .A2(n660), .ZN(n574) );
  NAND2_X1 U651 ( .A1(G77), .A2(n657), .ZN(n573) );
  NAND2_X1 U652 ( .A1(n574), .A2(n573), .ZN(n575) );
  XOR2_X1 U653 ( .A(KEYINPUT9), .B(n575), .Z(n576) );
  AND2_X1 U654 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U655 ( .A1(G2105), .A2(G2104), .ZN(n578) );
  XOR2_X1 U656 ( .A(KEYINPUT66), .B(n578), .Z(n706) );
  NAND2_X1 U657 ( .A1(G111), .A2(n907), .ZN(n579) );
  XOR2_X1 U658 ( .A(KEYINPUT75), .B(n579), .Z(n581) );
  NAND2_X1 U659 ( .A1(n708), .A2(G99), .ZN(n580) );
  NAND2_X1 U660 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U661 ( .A(KEYINPUT76), .B(n582), .ZN(n586) );
  NAND2_X1 U662 ( .A1(n906), .A2(G123), .ZN(n584) );
  XOR2_X1 U663 ( .A(KEYINPUT18), .B(n584), .Z(n585) );
  NOR2_X1 U664 ( .A1(n586), .A2(n585), .ZN(n589) );
  NAND2_X1 U665 ( .A1(n514), .A2(G135), .ZN(n588) );
  NAND2_X1 U666 ( .A1(n589), .A2(n588), .ZN(n1021) );
  XNOR2_X1 U667 ( .A(G2096), .B(n1021), .ZN(n590) );
  OR2_X1 U668 ( .A1(G2100), .A2(n590), .ZN(G156) );
  NAND2_X1 U669 ( .A1(n903), .A2(G138), .ZN(n591) );
  XNOR2_X1 U670 ( .A(KEYINPUT87), .B(n591), .ZN(n597) );
  NAND2_X1 U671 ( .A1(G114), .A2(n907), .ZN(n595) );
  NAND2_X1 U672 ( .A1(G102), .A2(n708), .ZN(n593) );
  NAND2_X1 U673 ( .A1(G126), .A2(n906), .ZN(n592) );
  AND2_X1 U674 ( .A1(n593), .A2(n592), .ZN(n594) );
  NAND2_X1 U675 ( .A1(n595), .A2(n594), .ZN(n596) );
  INV_X1 U676 ( .A(G132), .ZN(G219) );
  INV_X1 U677 ( .A(G82), .ZN(G220) );
  INV_X1 U678 ( .A(G120), .ZN(G236) );
  INV_X1 U679 ( .A(G69), .ZN(G235) );
  INV_X1 U680 ( .A(G108), .ZN(G238) );
  NAND2_X1 U681 ( .A1(G7), .A2(G661), .ZN(n598) );
  XOR2_X1 U682 ( .A(n598), .B(KEYINPUT10), .Z(n850) );
  NAND2_X1 U683 ( .A1(n850), .A2(G567), .ZN(n599) );
  XOR2_X1 U684 ( .A(KEYINPUT11), .B(n599), .Z(G234) );
  NAND2_X1 U685 ( .A1(n672), .A2(G56), .ZN(n600) );
  XNOR2_X1 U686 ( .A(n600), .B(KEYINPUT14), .ZN(n602) );
  NAND2_X1 U687 ( .A1(G43), .A2(n668), .ZN(n601) );
  NAND2_X1 U688 ( .A1(n602), .A2(n601), .ZN(n609) );
  NAND2_X1 U689 ( .A1(G68), .A2(n657), .ZN(n605) );
  NAND2_X1 U690 ( .A1(n660), .A2(G81), .ZN(n603) );
  XNOR2_X1 U691 ( .A(n603), .B(KEYINPUT12), .ZN(n604) );
  NAND2_X1 U692 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X1 U693 ( .A(n606), .B(KEYINPUT13), .ZN(n607) );
  XNOR2_X1 U694 ( .A(KEYINPUT71), .B(n607), .ZN(n608) );
  NAND2_X1 U695 ( .A1(n748), .A2(G860), .ZN(G153) );
  XOR2_X1 U696 ( .A(G171), .B(KEYINPUT72), .Z(G301) );
  NAND2_X1 U697 ( .A1(n672), .A2(G66), .ZN(n611) );
  NAND2_X1 U698 ( .A1(G54), .A2(n668), .ZN(n610) );
  NAND2_X1 U699 ( .A1(n611), .A2(n610), .ZN(n615) );
  NAND2_X1 U700 ( .A1(G92), .A2(n660), .ZN(n613) );
  NAND2_X1 U701 ( .A1(G79), .A2(n657), .ZN(n612) );
  NAND2_X1 U702 ( .A1(n613), .A2(n612), .ZN(n614) );
  NOR2_X1 U703 ( .A1(n615), .A2(n614), .ZN(n616) );
  NOR2_X1 U704 ( .A1(n946), .A2(G868), .ZN(n617) );
  XNOR2_X1 U705 ( .A(n617), .B(KEYINPUT73), .ZN(n619) );
  NAND2_X1 U706 ( .A1(G301), .A2(G868), .ZN(n618) );
  NAND2_X1 U707 ( .A1(n619), .A2(n618), .ZN(G284) );
  NAND2_X1 U708 ( .A1(G91), .A2(n660), .ZN(n621) );
  NAND2_X1 U709 ( .A1(G78), .A2(n657), .ZN(n620) );
  NAND2_X1 U710 ( .A1(n621), .A2(n620), .ZN(n624) );
  NAND2_X1 U711 ( .A1(n672), .A2(G65), .ZN(n622) );
  XOR2_X1 U712 ( .A(KEYINPUT70), .B(n622), .Z(n623) );
  NOR2_X1 U713 ( .A1(n624), .A2(n623), .ZN(n626) );
  NAND2_X1 U714 ( .A1(G53), .A2(n668), .ZN(n625) );
  NAND2_X1 U715 ( .A1(n626), .A2(n625), .ZN(G299) );
  INV_X1 U716 ( .A(G868), .ZN(n678) );
  NOR2_X1 U717 ( .A1(G286), .A2(n678), .ZN(n628) );
  NOR2_X1 U718 ( .A1(G868), .A2(G299), .ZN(n627) );
  NOR2_X1 U719 ( .A1(n628), .A2(n627), .ZN(G297) );
  INV_X1 U720 ( .A(G860), .ZN(n629) );
  NAND2_X1 U721 ( .A1(n629), .A2(G559), .ZN(n630) );
  NAND2_X1 U722 ( .A1(n630), .A2(n946), .ZN(n631) );
  XNOR2_X1 U723 ( .A(n631), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U724 ( .A1(G868), .A2(n943), .ZN(n634) );
  NAND2_X1 U725 ( .A1(G868), .A2(n946), .ZN(n632) );
  NOR2_X1 U726 ( .A1(G559), .A2(n632), .ZN(n633) );
  NOR2_X1 U727 ( .A1(n634), .A2(n633), .ZN(G282) );
  NAND2_X1 U728 ( .A1(G559), .A2(n946), .ZN(n635) );
  XNOR2_X1 U729 ( .A(n635), .B(KEYINPUT77), .ZN(n636) );
  XOR2_X1 U730 ( .A(n943), .B(n636), .Z(n686) );
  NOR2_X1 U731 ( .A1(n686), .A2(G860), .ZN(n643) );
  NAND2_X1 U732 ( .A1(n672), .A2(G67), .ZN(n638) );
  NAND2_X1 U733 ( .A1(G55), .A2(n668), .ZN(n637) );
  NAND2_X1 U734 ( .A1(n638), .A2(n637), .ZN(n642) );
  NAND2_X1 U735 ( .A1(G93), .A2(n660), .ZN(n640) );
  NAND2_X1 U736 ( .A1(G80), .A2(n657), .ZN(n639) );
  NAND2_X1 U737 ( .A1(n640), .A2(n639), .ZN(n641) );
  NOR2_X1 U738 ( .A1(n642), .A2(n641), .ZN(n682) );
  XNOR2_X1 U739 ( .A(n643), .B(n682), .ZN(G145) );
  NAND2_X1 U740 ( .A1(G85), .A2(n660), .ZN(n645) );
  NAND2_X1 U741 ( .A1(G72), .A2(n657), .ZN(n644) );
  NAND2_X1 U742 ( .A1(n645), .A2(n644), .ZN(n648) );
  NAND2_X1 U743 ( .A1(G47), .A2(n668), .ZN(n646) );
  XNOR2_X1 U744 ( .A(KEYINPUT67), .B(n646), .ZN(n647) );
  NOR2_X1 U745 ( .A1(n648), .A2(n647), .ZN(n650) );
  NAND2_X1 U746 ( .A1(n672), .A2(G60), .ZN(n649) );
  NAND2_X1 U747 ( .A1(n650), .A2(n649), .ZN(G290) );
  NAND2_X1 U748 ( .A1(G88), .A2(n660), .ZN(n652) );
  NAND2_X1 U749 ( .A1(G75), .A2(n657), .ZN(n651) );
  NAND2_X1 U750 ( .A1(n652), .A2(n651), .ZN(n656) );
  NAND2_X1 U751 ( .A1(n672), .A2(G62), .ZN(n654) );
  NAND2_X1 U752 ( .A1(G50), .A2(n668), .ZN(n653) );
  NAND2_X1 U753 ( .A1(n654), .A2(n653), .ZN(n655) );
  NOR2_X1 U754 ( .A1(n656), .A2(n655), .ZN(G166) );
  INV_X1 U755 ( .A(G166), .ZN(G303) );
  NAND2_X1 U756 ( .A1(G73), .A2(n657), .ZN(n658) );
  XOR2_X1 U757 ( .A(KEYINPUT2), .B(n658), .Z(n665) );
  NAND2_X1 U758 ( .A1(n672), .A2(G61), .ZN(n659) );
  XNOR2_X1 U759 ( .A(n659), .B(KEYINPUT80), .ZN(n662) );
  NAND2_X1 U760 ( .A1(G86), .A2(n660), .ZN(n661) );
  NAND2_X1 U761 ( .A1(n662), .A2(n661), .ZN(n663) );
  XOR2_X1 U762 ( .A(KEYINPUT81), .B(n663), .Z(n664) );
  NOR2_X1 U763 ( .A1(n665), .A2(n664), .ZN(n667) );
  NAND2_X1 U764 ( .A1(G48), .A2(n668), .ZN(n666) );
  NAND2_X1 U765 ( .A1(n667), .A2(n666), .ZN(G305) );
  NAND2_X1 U766 ( .A1(G651), .A2(G74), .ZN(n670) );
  NAND2_X1 U767 ( .A1(G49), .A2(n668), .ZN(n669) );
  NAND2_X1 U768 ( .A1(n670), .A2(n669), .ZN(n671) );
  NOR2_X1 U769 ( .A1(n672), .A2(n671), .ZN(n673) );
  XNOR2_X1 U770 ( .A(KEYINPUT78), .B(n673), .ZN(n677) );
  NAND2_X1 U771 ( .A1(n674), .A2(G87), .ZN(n675) );
  XOR2_X1 U772 ( .A(KEYINPUT79), .B(n675), .Z(n676) );
  NAND2_X1 U773 ( .A1(n677), .A2(n676), .ZN(G288) );
  NAND2_X1 U774 ( .A1(n678), .A2(n682), .ZN(n689) );
  XNOR2_X1 U775 ( .A(KEYINPUT19), .B(KEYINPUT82), .ZN(n680) );
  XOR2_X1 U776 ( .A(G290), .B(G303), .Z(n679) );
  XNOR2_X1 U777 ( .A(n680), .B(n679), .ZN(n681) );
  XNOR2_X1 U778 ( .A(n682), .B(n681), .ZN(n684) );
  XOR2_X1 U779 ( .A(G305), .B(G299), .Z(n683) );
  XNOR2_X1 U780 ( .A(n684), .B(n683), .ZN(n685) );
  XOR2_X1 U781 ( .A(n685), .B(G288), .Z(n920) );
  XNOR2_X1 U782 ( .A(n920), .B(n686), .ZN(n687) );
  NAND2_X1 U783 ( .A1(n687), .A2(G868), .ZN(n688) );
  NAND2_X1 U784 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U785 ( .A(n690), .B(KEYINPUT83), .ZN(G295) );
  NAND2_X1 U786 ( .A1(G2078), .A2(G2084), .ZN(n691) );
  XOR2_X1 U787 ( .A(KEYINPUT20), .B(n691), .Z(n692) );
  NAND2_X1 U788 ( .A1(G2090), .A2(n692), .ZN(n693) );
  XNOR2_X1 U789 ( .A(KEYINPUT21), .B(n693), .ZN(n694) );
  NAND2_X1 U790 ( .A1(n694), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U791 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U792 ( .A1(G483), .A2(G661), .ZN(n704) );
  NOR2_X1 U793 ( .A1(G235), .A2(G236), .ZN(n695) );
  XNOR2_X1 U794 ( .A(n695), .B(KEYINPUT85), .ZN(n696) );
  NOR2_X1 U795 ( .A1(G238), .A2(n696), .ZN(n697) );
  NAND2_X1 U796 ( .A1(G57), .A2(n697), .ZN(n854) );
  NAND2_X1 U797 ( .A1(n854), .A2(G567), .ZN(n703) );
  NOR2_X1 U798 ( .A1(G220), .A2(G219), .ZN(n698) );
  XOR2_X1 U799 ( .A(KEYINPUT22), .B(n698), .Z(n699) );
  NOR2_X1 U800 ( .A1(G218), .A2(n699), .ZN(n700) );
  XNOR2_X1 U801 ( .A(KEYINPUT84), .B(n700), .ZN(n701) );
  NAND2_X1 U802 ( .A1(n701), .A2(G96), .ZN(n855) );
  NAND2_X1 U803 ( .A1(n855), .A2(G2106), .ZN(n702) );
  NAND2_X1 U804 ( .A1(n703), .A2(n702), .ZN(n856) );
  NOR2_X1 U805 ( .A1(n704), .A2(n856), .ZN(n705) );
  XNOR2_X1 U806 ( .A(n705), .B(KEYINPUT86), .ZN(n853) );
  NAND2_X1 U807 ( .A1(G36), .A2(n853), .ZN(G176) );
  NAND2_X1 U808 ( .A1(G125), .A2(n906), .ZN(n713) );
  NAND2_X1 U809 ( .A1(G113), .A2(n706), .ZN(n707) );
  NAND2_X1 U810 ( .A1(G101), .A2(n708), .ZN(n709) );
  XNOR2_X1 U811 ( .A(KEYINPUT23), .B(n709), .ZN(n710) );
  NOR2_X1 U812 ( .A1(n711), .A2(n710), .ZN(n712) );
  INV_X1 U813 ( .A(n811), .ZN(n716) );
  XNOR2_X1 U814 ( .A(G2078), .B(KEYINPUT25), .ZN(n1003) );
  NOR2_X1 U815 ( .A1(n719), .A2(n1003), .ZN(n718) );
  INV_X1 U816 ( .A(G1961), .ZN(n942) );
  NOR2_X1 U817 ( .A1(n736), .A2(n942), .ZN(n717) );
  NOR2_X1 U818 ( .A1(n718), .A2(n717), .ZN(n760) );
  NOR2_X1 U819 ( .A1(G171), .A2(n760), .ZN(n725) );
  XNOR2_X2 U820 ( .A(n720), .B(KEYINPUT94), .ZN(n784) );
  INV_X1 U821 ( .A(n773), .ZN(n721) );
  NAND2_X1 U822 ( .A1(n772), .A2(n516), .ZN(n722) );
  XNOR2_X1 U823 ( .A(n722), .B(KEYINPUT30), .ZN(n723) );
  NOR2_X1 U824 ( .A1(n723), .A2(G168), .ZN(n724) );
  XNOR2_X1 U825 ( .A(n727), .B(n726), .ZN(n764) );
  INV_X1 U826 ( .A(G299), .ZN(n753) );
  INV_X1 U827 ( .A(KEYINPUT96), .ZN(n733) );
  NAND2_X1 U828 ( .A1(n736), .A2(G2072), .ZN(n729) );
  INV_X1 U829 ( .A(KEYINPUT27), .ZN(n728) );
  NAND2_X1 U830 ( .A1(G1956), .A2(n719), .ZN(n730) );
  NAND2_X1 U831 ( .A1(n731), .A2(n730), .ZN(n732) );
  INV_X1 U832 ( .A(KEYINPUT28), .ZN(n734) );
  XNOR2_X1 U833 ( .A(n735), .B(n734), .ZN(n757) );
  INV_X1 U834 ( .A(n946), .ZN(n919) );
  NOR2_X1 U835 ( .A1(n943), .A2(n919), .ZN(n741) );
  NAND2_X1 U836 ( .A1(n736), .A2(G1996), .ZN(n737) );
  XNOR2_X1 U837 ( .A(n737), .B(KEYINPUT26), .ZN(n739) );
  NAND2_X1 U838 ( .A1(G1341), .A2(n719), .ZN(n738) );
  NAND2_X1 U839 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U840 ( .A(KEYINPUT97), .B(n740), .ZN(n747) );
  NAND2_X1 U841 ( .A1(n741), .A2(n747), .ZN(n746) );
  NAND2_X1 U842 ( .A1(n719), .A2(G1348), .ZN(n742) );
  XNOR2_X1 U843 ( .A(n742), .B(KEYINPUT98), .ZN(n744) );
  NAND2_X1 U844 ( .A1(n736), .A2(G2067), .ZN(n743) );
  NAND2_X1 U845 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U846 ( .A1(n746), .A2(n745), .ZN(n751) );
  NAND2_X1 U847 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U848 ( .A1(n749), .A2(n919), .ZN(n750) );
  NAND2_X1 U849 ( .A1(n751), .A2(n750), .ZN(n755) );
  NAND2_X1 U850 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U851 ( .A1(n755), .A2(n754), .ZN(n756) );
  NAND2_X1 U852 ( .A1(n757), .A2(n756), .ZN(n759) );
  XNOR2_X1 U853 ( .A(KEYINPUT99), .B(KEYINPUT29), .ZN(n758) );
  XNOR2_X1 U854 ( .A(n759), .B(n758), .ZN(n762) );
  NAND2_X1 U855 ( .A1(n760), .A2(G171), .ZN(n761) );
  NAND2_X1 U856 ( .A1(n762), .A2(n761), .ZN(n763) );
  NAND2_X1 U857 ( .A1(n764), .A2(n763), .ZN(n765) );
  NOR2_X1 U858 ( .A1(n784), .A2(G1971), .ZN(n766) );
  XOR2_X1 U859 ( .A(KEYINPUT101), .B(n766), .Z(n768) );
  NOR2_X1 U860 ( .A1(G2090), .A2(n719), .ZN(n767) );
  NOR2_X1 U861 ( .A1(n768), .A2(n767), .ZN(n769) );
  NAND2_X1 U862 ( .A1(n769), .A2(G303), .ZN(n770) );
  INV_X1 U863 ( .A(n772), .ZN(n776) );
  NAND2_X1 U864 ( .A1(n773), .A2(G8), .ZN(n774) );
  XNOR2_X1 U865 ( .A(KEYINPUT95), .B(n774), .ZN(n775) );
  NOR2_X1 U866 ( .A1(n776), .A2(n775), .ZN(n778) );
  NAND2_X1 U867 ( .A1(n778), .A2(n777), .ZN(n790) );
  NOR2_X1 U868 ( .A1(G1976), .A2(G288), .ZN(n953) );
  NOR2_X1 U869 ( .A1(G1971), .A2(G303), .ZN(n779) );
  NOR2_X1 U870 ( .A1(n953), .A2(n779), .ZN(n780) );
  NAND2_X1 U871 ( .A1(G288), .A2(G1976), .ZN(n781) );
  XOR2_X1 U872 ( .A(KEYINPUT104), .B(n781), .Z(n952) );
  XNOR2_X1 U873 ( .A(n782), .B(KEYINPUT105), .ZN(n783) );
  XNOR2_X1 U874 ( .A(G1981), .B(G305), .ZN(n950) );
  AND2_X1 U875 ( .A1(n953), .A2(KEYINPUT33), .ZN(n785) );
  INV_X1 U876 ( .A(n784), .ZN(n796) );
  NAND2_X1 U877 ( .A1(n785), .A2(n796), .ZN(n786) );
  NOR2_X1 U878 ( .A1(G1981), .A2(G305), .ZN(n788) );
  XNOR2_X1 U879 ( .A(n788), .B(KEYINPUT24), .ZN(n789) );
  NAND2_X1 U880 ( .A1(n789), .A2(n796), .ZN(n797) );
  AND2_X1 U881 ( .A1(n791), .A2(n790), .ZN(n794) );
  NAND2_X1 U882 ( .A1(G166), .A2(G8), .ZN(n792) );
  NOR2_X1 U883 ( .A1(G2090), .A2(n792), .ZN(n793) );
  NOR2_X1 U884 ( .A1(n794), .A2(n793), .ZN(n795) );
  NAND2_X1 U885 ( .A1(n797), .A2(n515), .ZN(n798) );
  NAND2_X1 U886 ( .A1(G140), .A2(n514), .ZN(n800) );
  NAND2_X1 U887 ( .A1(G104), .A2(n708), .ZN(n799) );
  NAND2_X1 U888 ( .A1(n800), .A2(n799), .ZN(n801) );
  XNOR2_X1 U889 ( .A(KEYINPUT34), .B(n801), .ZN(n807) );
  NAND2_X1 U890 ( .A1(G116), .A2(n907), .ZN(n802) );
  XOR2_X1 U891 ( .A(KEYINPUT89), .B(n802), .Z(n804) );
  NAND2_X1 U892 ( .A1(n906), .A2(G128), .ZN(n803) );
  NAND2_X1 U893 ( .A1(n804), .A2(n803), .ZN(n805) );
  XOR2_X1 U894 ( .A(n805), .B(KEYINPUT35), .Z(n806) );
  NOR2_X1 U895 ( .A1(n807), .A2(n806), .ZN(n808) );
  XOR2_X1 U896 ( .A(KEYINPUT36), .B(n808), .Z(n809) );
  XOR2_X1 U897 ( .A(KEYINPUT90), .B(n809), .Z(n913) );
  XNOR2_X1 U898 ( .A(KEYINPUT37), .B(G2067), .ZN(n843) );
  NOR2_X1 U899 ( .A1(n913), .A2(n843), .ZN(n1037) );
  NOR2_X1 U900 ( .A1(n810), .A2(n811), .ZN(n812) );
  XNOR2_X1 U901 ( .A(n812), .B(KEYINPUT88), .ZN(n845) );
  NAND2_X1 U902 ( .A1(n1037), .A2(n845), .ZN(n841) );
  NAND2_X1 U903 ( .A1(n906), .A2(G129), .ZN(n814) );
  NAND2_X1 U904 ( .A1(G117), .A2(n907), .ZN(n813) );
  NAND2_X1 U905 ( .A1(n814), .A2(n813), .ZN(n817) );
  NAND2_X1 U906 ( .A1(n708), .A2(G105), .ZN(n815) );
  XOR2_X1 U907 ( .A(KEYINPUT38), .B(n815), .Z(n816) );
  NOR2_X1 U908 ( .A1(n817), .A2(n816), .ZN(n819) );
  NAND2_X1 U909 ( .A1(n514), .A2(G141), .ZN(n818) );
  NAND2_X1 U910 ( .A1(n819), .A2(n818), .ZN(n885) );
  NAND2_X1 U911 ( .A1(G1996), .A2(n885), .ZN(n820) );
  XNOR2_X1 U912 ( .A(n820), .B(KEYINPUT92), .ZN(n829) );
  NAND2_X1 U913 ( .A1(n708), .A2(G95), .ZN(n822) );
  NAND2_X1 U914 ( .A1(G107), .A2(n907), .ZN(n821) );
  NAND2_X1 U915 ( .A1(n822), .A2(n821), .ZN(n825) );
  NAND2_X1 U916 ( .A1(G119), .A2(n906), .ZN(n823) );
  XNOR2_X1 U917 ( .A(KEYINPUT91), .B(n823), .ZN(n824) );
  NOR2_X1 U918 ( .A1(n825), .A2(n824), .ZN(n827) );
  NAND2_X1 U919 ( .A1(n514), .A2(G131), .ZN(n826) );
  NAND2_X1 U920 ( .A1(n827), .A2(n826), .ZN(n886) );
  NAND2_X1 U921 ( .A1(G1991), .A2(n886), .ZN(n828) );
  NAND2_X1 U922 ( .A1(n829), .A2(n828), .ZN(n1024) );
  NAND2_X1 U923 ( .A1(n1024), .A2(n845), .ZN(n830) );
  XOR2_X1 U924 ( .A(n830), .B(KEYINPUT93), .Z(n835) );
  XNOR2_X1 U925 ( .A(G1986), .B(G290), .ZN(n962) );
  NAND2_X1 U926 ( .A1(n962), .A2(n845), .ZN(n831) );
  OR2_X2 U927 ( .A1(n833), .A2(n832), .ZN(n848) );
  NOR2_X1 U928 ( .A1(n885), .A2(G1996), .ZN(n834) );
  XNOR2_X1 U929 ( .A(n834), .B(KEYINPUT106), .ZN(n1017) );
  INV_X1 U930 ( .A(n835), .ZN(n838) );
  NOR2_X1 U931 ( .A1(G1986), .A2(G290), .ZN(n836) );
  NOR2_X1 U932 ( .A1(G1991), .A2(n886), .ZN(n1020) );
  NOR2_X1 U933 ( .A1(n836), .A2(n1020), .ZN(n837) );
  NOR2_X1 U934 ( .A1(n838), .A2(n837), .ZN(n839) );
  NOR2_X1 U935 ( .A1(n1017), .A2(n839), .ZN(n840) );
  XNOR2_X1 U936 ( .A(n840), .B(KEYINPUT39), .ZN(n842) );
  NAND2_X1 U937 ( .A1(n842), .A2(n841), .ZN(n844) );
  NAND2_X1 U938 ( .A1(n913), .A2(n843), .ZN(n1034) );
  NAND2_X1 U939 ( .A1(n844), .A2(n1034), .ZN(n846) );
  NAND2_X1 U940 ( .A1(n846), .A2(n845), .ZN(n847) );
  NAND2_X1 U941 ( .A1(n848), .A2(n847), .ZN(n849) );
  XNOR2_X1 U942 ( .A(n849), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U943 ( .A1(G2106), .A2(n850), .ZN(G217) );
  INV_X1 U944 ( .A(n850), .ZN(G223) );
  AND2_X1 U945 ( .A1(G15), .A2(G2), .ZN(n851) );
  NAND2_X1 U946 ( .A1(G661), .A2(n851), .ZN(G259) );
  NAND2_X1 U947 ( .A1(G3), .A2(G1), .ZN(n852) );
  NAND2_X1 U948 ( .A1(n853), .A2(n852), .ZN(G188) );
  XNOR2_X1 U949 ( .A(G96), .B(KEYINPUT107), .ZN(G221) );
  NOR2_X1 U950 ( .A1(n855), .A2(n854), .ZN(G325) );
  XOR2_X1 U951 ( .A(KEYINPUT108), .B(G325), .Z(G261) );
  INV_X1 U953 ( .A(n856), .ZN(G319) );
  XNOR2_X1 U954 ( .A(G1956), .B(G2474), .ZN(n866) );
  XOR2_X1 U955 ( .A(G1976), .B(G1971), .Z(n858) );
  XOR2_X1 U956 ( .A(G1986), .B(n942), .Z(n857) );
  XNOR2_X1 U957 ( .A(n858), .B(n857), .ZN(n862) );
  XOR2_X1 U958 ( .A(G1966), .B(G1981), .Z(n860) );
  XNOR2_X1 U959 ( .A(G1996), .B(G1991), .ZN(n859) );
  XNOR2_X1 U960 ( .A(n860), .B(n859), .ZN(n861) );
  XOR2_X1 U961 ( .A(n862), .B(n861), .Z(n864) );
  XNOR2_X1 U962 ( .A(KEYINPUT112), .B(KEYINPUT41), .ZN(n863) );
  XNOR2_X1 U963 ( .A(n864), .B(n863), .ZN(n865) );
  XNOR2_X1 U964 ( .A(n866), .B(n865), .ZN(G229) );
  XNOR2_X1 U965 ( .A(G2072), .B(G2078), .ZN(n867) );
  XNOR2_X1 U966 ( .A(n867), .B(KEYINPUT42), .ZN(n877) );
  XOR2_X1 U967 ( .A(KEYINPUT43), .B(KEYINPUT110), .Z(n869) );
  XNOR2_X1 U968 ( .A(KEYINPUT109), .B(G2096), .ZN(n868) );
  XNOR2_X1 U969 ( .A(n869), .B(n868), .ZN(n873) );
  XOR2_X1 U970 ( .A(G2100), .B(G2090), .Z(n871) );
  XNOR2_X1 U971 ( .A(G2067), .B(G2084), .ZN(n870) );
  XNOR2_X1 U972 ( .A(n871), .B(n870), .ZN(n872) );
  XOR2_X1 U973 ( .A(n873), .B(n872), .Z(n875) );
  XNOR2_X1 U974 ( .A(KEYINPUT111), .B(G2678), .ZN(n874) );
  XNOR2_X1 U975 ( .A(n875), .B(n874), .ZN(n876) );
  XNOR2_X1 U976 ( .A(n877), .B(n876), .ZN(G227) );
  NAND2_X1 U977 ( .A1(G124), .A2(n906), .ZN(n878) );
  XNOR2_X1 U978 ( .A(n878), .B(KEYINPUT44), .ZN(n880) );
  NAND2_X1 U979 ( .A1(G112), .A2(n907), .ZN(n879) );
  NAND2_X1 U980 ( .A1(n880), .A2(n879), .ZN(n884) );
  NAND2_X1 U981 ( .A1(G136), .A2(n514), .ZN(n882) );
  NAND2_X1 U982 ( .A1(G100), .A2(n708), .ZN(n881) );
  NAND2_X1 U983 ( .A1(n882), .A2(n881), .ZN(n883) );
  NOR2_X1 U984 ( .A1(n884), .A2(n883), .ZN(G162) );
  XNOR2_X1 U985 ( .A(G160), .B(n885), .ZN(n887) );
  XNOR2_X1 U986 ( .A(n887), .B(n886), .ZN(n891) );
  XOR2_X1 U987 ( .A(KEYINPUT114), .B(KEYINPUT113), .Z(n889) );
  XNOR2_X1 U988 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n888) );
  XNOR2_X1 U989 ( .A(n889), .B(n888), .ZN(n890) );
  XOR2_X1 U990 ( .A(n891), .B(n890), .Z(n893) );
  XNOR2_X1 U991 ( .A(G164), .B(G162), .ZN(n892) );
  XNOR2_X1 U992 ( .A(n893), .B(n892), .ZN(n902) );
  NAND2_X1 U993 ( .A1(n906), .A2(G130), .ZN(n895) );
  NAND2_X1 U994 ( .A1(G118), .A2(n907), .ZN(n894) );
  NAND2_X1 U995 ( .A1(n895), .A2(n894), .ZN(n900) );
  NAND2_X1 U996 ( .A1(G142), .A2(n514), .ZN(n897) );
  NAND2_X1 U997 ( .A1(G106), .A2(n708), .ZN(n896) );
  NAND2_X1 U998 ( .A1(n897), .A2(n896), .ZN(n898) );
  XOR2_X1 U999 ( .A(KEYINPUT45), .B(n898), .Z(n899) );
  NOR2_X1 U1000 ( .A1(n900), .A2(n899), .ZN(n901) );
  XOR2_X1 U1001 ( .A(n902), .B(n901), .Z(n915) );
  NAND2_X1 U1002 ( .A1(G139), .A2(n514), .ZN(n905) );
  NAND2_X1 U1003 ( .A1(G103), .A2(n708), .ZN(n904) );
  NAND2_X1 U1004 ( .A1(n905), .A2(n904), .ZN(n912) );
  NAND2_X1 U1005 ( .A1(n906), .A2(G127), .ZN(n909) );
  NAND2_X1 U1006 ( .A1(G115), .A2(n907), .ZN(n908) );
  NAND2_X1 U1007 ( .A1(n909), .A2(n908), .ZN(n910) );
  XOR2_X1 U1008 ( .A(KEYINPUT47), .B(n910), .Z(n911) );
  NOR2_X1 U1009 ( .A1(n912), .A2(n911), .ZN(n1027) );
  XNOR2_X1 U1010 ( .A(n913), .B(n1027), .ZN(n914) );
  XNOR2_X1 U1011 ( .A(n915), .B(n914), .ZN(n916) );
  XOR2_X1 U1012 ( .A(n1021), .B(n916), .Z(n917) );
  NOR2_X1 U1013 ( .A1(G37), .A2(n917), .ZN(n918) );
  XOR2_X1 U1014 ( .A(KEYINPUT115), .B(n918), .Z(G395) );
  XOR2_X1 U1015 ( .A(n943), .B(n919), .Z(n921) );
  XNOR2_X1 U1016 ( .A(n921), .B(n920), .ZN(n923) );
  XNOR2_X1 U1017 ( .A(G286), .B(G171), .ZN(n922) );
  XNOR2_X1 U1018 ( .A(n923), .B(n922), .ZN(n924) );
  NOR2_X1 U1019 ( .A1(G37), .A2(n924), .ZN(n925) );
  XNOR2_X1 U1020 ( .A(KEYINPUT116), .B(n925), .ZN(G397) );
  XOR2_X1 U1021 ( .A(G2451), .B(G2430), .Z(n927) );
  XNOR2_X1 U1022 ( .A(G2438), .B(G2443), .ZN(n926) );
  XNOR2_X1 U1023 ( .A(n927), .B(n926), .ZN(n933) );
  XOR2_X1 U1024 ( .A(G2435), .B(G2454), .Z(n929) );
  XNOR2_X1 U1025 ( .A(G1348), .B(G1341), .ZN(n928) );
  XNOR2_X1 U1026 ( .A(n929), .B(n928), .ZN(n931) );
  XOR2_X1 U1027 ( .A(G2446), .B(G2427), .Z(n930) );
  XNOR2_X1 U1028 ( .A(n931), .B(n930), .ZN(n932) );
  XOR2_X1 U1029 ( .A(n933), .B(n932), .Z(n934) );
  NAND2_X1 U1030 ( .A1(G14), .A2(n934), .ZN(n941) );
  NAND2_X1 U1031 ( .A1(G319), .A2(n941), .ZN(n938) );
  NOR2_X1 U1032 ( .A1(G229), .A2(G227), .ZN(n935) );
  XOR2_X1 U1033 ( .A(KEYINPUT49), .B(n935), .Z(n936) );
  XNOR2_X1 U1034 ( .A(n936), .B(KEYINPUT117), .ZN(n937) );
  NOR2_X1 U1035 ( .A1(n938), .A2(n937), .ZN(n940) );
  NOR2_X1 U1036 ( .A1(G395), .A2(G397), .ZN(n939) );
  NAND2_X1 U1037 ( .A1(n940), .A2(n939), .ZN(G225) );
  INV_X1 U1038 ( .A(G225), .ZN(G308) );
  INV_X1 U1039 ( .A(G57), .ZN(G237) );
  INV_X1 U1040 ( .A(n941), .ZN(G401) );
  INV_X1 U1041 ( .A(G16), .ZN(n990) );
  XOR2_X1 U1042 ( .A(KEYINPUT56), .B(n990), .Z(n966) );
  XNOR2_X1 U1043 ( .A(G171), .B(n942), .ZN(n945) );
  XNOR2_X1 U1044 ( .A(n943), .B(G1341), .ZN(n944) );
  NOR2_X1 U1045 ( .A1(n945), .A2(n944), .ZN(n948) );
  XNOR2_X1 U1046 ( .A(G1348), .B(n946), .ZN(n947) );
  NAND2_X1 U1047 ( .A1(n948), .A2(n947), .ZN(n958) );
  XOR2_X1 U1048 ( .A(G168), .B(G1966), .Z(n949) );
  NOR2_X1 U1049 ( .A1(n950), .A2(n949), .ZN(n951) );
  XOR2_X1 U1050 ( .A(KEYINPUT57), .B(n951), .Z(n956) );
  NOR2_X1 U1051 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1052 ( .A(n954), .B(KEYINPUT124), .ZN(n955) );
  NAND2_X1 U1053 ( .A1(n956), .A2(n955), .ZN(n957) );
  NOR2_X1 U1054 ( .A1(n958), .A2(n957), .ZN(n964) );
  XOR2_X1 U1055 ( .A(G303), .B(G1971), .Z(n960) );
  XOR2_X1 U1056 ( .A(G299), .B(G1956), .Z(n959) );
  NAND2_X1 U1057 ( .A1(n960), .A2(n959), .ZN(n961) );
  NOR2_X1 U1058 ( .A1(n962), .A2(n961), .ZN(n963) );
  NAND2_X1 U1059 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1060 ( .A1(n966), .A2(n965), .ZN(n1047) );
  XOR2_X1 U1061 ( .A(G5), .B(G1961), .Z(n980) );
  XOR2_X1 U1062 ( .A(G1956), .B(G20), .Z(n972) );
  XOR2_X1 U1063 ( .A(G1981), .B(G6), .Z(n967) );
  XNOR2_X1 U1064 ( .A(KEYINPUT125), .B(n967), .ZN(n969) );
  XNOR2_X1 U1065 ( .A(G19), .B(G1341), .ZN(n968) );
  NOR2_X1 U1066 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1067 ( .A(KEYINPUT126), .B(n970), .ZN(n971) );
  NAND2_X1 U1068 ( .A1(n972), .A2(n971), .ZN(n975) );
  XOR2_X1 U1069 ( .A(KEYINPUT59), .B(G1348), .Z(n973) );
  XNOR2_X1 U1070 ( .A(G4), .B(n973), .ZN(n974) );
  NOR2_X1 U1071 ( .A1(n975), .A2(n974), .ZN(n976) );
  XOR2_X1 U1072 ( .A(KEYINPUT60), .B(n976), .Z(n978) );
  XNOR2_X1 U1073 ( .A(G1966), .B(G21), .ZN(n977) );
  NOR2_X1 U1074 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1075 ( .A1(n980), .A2(n979), .ZN(n988) );
  XNOR2_X1 U1076 ( .A(G1986), .B(G24), .ZN(n982) );
  XNOR2_X1 U1077 ( .A(G23), .B(G1976), .ZN(n981) );
  NOR2_X1 U1078 ( .A1(n982), .A2(n981), .ZN(n985) );
  XNOR2_X1 U1079 ( .A(G1971), .B(KEYINPUT127), .ZN(n983) );
  XNOR2_X1 U1080 ( .A(n983), .B(G22), .ZN(n984) );
  NAND2_X1 U1081 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1082 ( .A(KEYINPUT58), .B(n986), .ZN(n987) );
  NOR2_X1 U1083 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1084 ( .A(KEYINPUT61), .B(n989), .ZN(n991) );
  NAND2_X1 U1085 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1086 ( .A1(n992), .A2(G11), .ZN(n1045) );
  INV_X1 U1087 ( .A(KEYINPUT55), .ZN(n1039) );
  XNOR2_X1 U1088 ( .A(G2090), .B(G35), .ZN(n1009) );
  XOR2_X1 U1089 ( .A(G1991), .B(G25), .Z(n993) );
  NAND2_X1 U1090 ( .A1(G28), .A2(n993), .ZN(n994) );
  XNOR2_X1 U1091 ( .A(n994), .B(KEYINPUT119), .ZN(n1002) );
  XNOR2_X1 U1092 ( .A(G1996), .B(G32), .ZN(n1000) );
  XNOR2_X1 U1093 ( .A(G2067), .B(KEYINPUT120), .ZN(n995) );
  XNOR2_X1 U1094 ( .A(n995), .B(G26), .ZN(n997) );
  XNOR2_X1 U1095 ( .A(G33), .B(G2072), .ZN(n996) );
  NOR2_X1 U1096 ( .A1(n997), .A2(n996), .ZN(n998) );
  XNOR2_X1 U1097 ( .A(KEYINPUT121), .B(n998), .ZN(n999) );
  NOR2_X1 U1098 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1099 ( .A1(n1002), .A2(n1001), .ZN(n1006) );
  XOR2_X1 U1100 ( .A(G27), .B(n1003), .Z(n1004) );
  XNOR2_X1 U1101 ( .A(KEYINPUT122), .B(n1004), .ZN(n1005) );
  NOR2_X1 U1102 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1103 ( .A(KEYINPUT53), .B(n1007), .ZN(n1008) );
  NOR2_X1 U1104 ( .A1(n1009), .A2(n1008), .ZN(n1012) );
  XOR2_X1 U1105 ( .A(G2084), .B(G34), .Z(n1010) );
  XNOR2_X1 U1106 ( .A(KEYINPUT54), .B(n1010), .ZN(n1011) );
  NAND2_X1 U1107 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XOR2_X1 U1108 ( .A(n1039), .B(n1013), .Z(n1014) );
  NOR2_X1 U1109 ( .A1(G29), .A2(n1014), .ZN(n1015) );
  XNOR2_X1 U1110 ( .A(n1015), .B(KEYINPUT123), .ZN(n1043) );
  XOR2_X1 U1111 ( .A(G2090), .B(G162), .Z(n1016) );
  NOR2_X1 U1112 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XOR2_X1 U1113 ( .A(KEYINPUT51), .B(n1018), .Z(n1026) );
  XOR2_X1 U1114 ( .A(G160), .B(G2084), .Z(n1019) );
  NOR2_X1 U1115 ( .A1(n1020), .A2(n1019), .ZN(n1022) );
  NAND2_X1 U1116 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NOR2_X1 U1117 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1118 ( .A1(n1026), .A2(n1025), .ZN(n1033) );
  XOR2_X1 U1119 ( .A(G2072), .B(n1027), .Z(n1029) );
  XOR2_X1 U1120 ( .A(G164), .B(G2078), .Z(n1028) );
  NOR2_X1 U1121 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  XOR2_X1 U1122 ( .A(KEYINPUT118), .B(n1030), .Z(n1031) );
  XNOR2_X1 U1123 ( .A(KEYINPUT50), .B(n1031), .ZN(n1032) );
  NOR2_X1 U1124 ( .A1(n1033), .A2(n1032), .ZN(n1035) );
  NAND2_X1 U1125 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  NOR2_X1 U1126 ( .A1(n1037), .A2(n1036), .ZN(n1038) );
  XNOR2_X1 U1127 ( .A(n1038), .B(KEYINPUT52), .ZN(n1040) );
  NAND2_X1 U1128 ( .A1(n1040), .A2(n1039), .ZN(n1041) );
  NAND2_X1 U1129 ( .A1(G29), .A2(n1041), .ZN(n1042) );
  NAND2_X1 U1130 ( .A1(n1043), .A2(n1042), .ZN(n1044) );
  NOR2_X1 U1131 ( .A1(n1045), .A2(n1044), .ZN(n1046) );
  NAND2_X1 U1132 ( .A1(n1047), .A2(n1046), .ZN(n1048) );
  XNOR2_X1 U1133 ( .A(KEYINPUT62), .B(n1048), .ZN(G150) );
  INV_X1 U1134 ( .A(G150), .ZN(G311) );
endmodule

