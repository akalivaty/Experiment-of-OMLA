//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 0 0 0 1 0 0 0 0 1 0 0 0 0 0 0 1 1 1 1 1 0 1 0 1 0 0 1 1 1 1 1 0 1 1 1 1 0 1 1 1 1 1 1 1 0 1 0 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:37 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1274, new_n1275, new_n1276, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1350, new_n1351, new_n1352;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G13), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  OAI21_X1  g0007(.A(G250), .B1(G257), .B2(G264), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NOR2_X1   g0013(.A1(G58), .A2(G68), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(G50), .ZN(new_n216));
  OAI22_X1  g0016(.A1(new_n209), .A2(KEYINPUT0), .B1(new_n213), .B2(new_n216), .ZN(new_n217));
  AOI21_X1  g0017(.A(new_n217), .B1(KEYINPUT0), .B2(new_n209), .ZN(new_n218));
  XNOR2_X1  g0018(.A(new_n218), .B(KEYINPUT64), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n205), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT1), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n219), .A2(new_n227), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  INV_X1    g0029(.A(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(KEYINPUT2), .B(G226), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XNOR2_X1  g0037(.A(G50), .B(G68), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G58), .B(G77), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n238), .B(new_n239), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT65), .ZN(new_n241));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XOR2_X1   g0042(.A(G107), .B(G116), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  INV_X1    g0044(.A(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n241), .B(new_n245), .ZN(G351));
  INV_X1    g0046(.A(G1), .ZN(new_n247));
  OAI21_X1  g0047(.A(new_n247), .B1(G41), .B2(G45), .ZN(new_n248));
  INV_X1    g0048(.A(G274), .ZN(new_n249));
  NOR2_X1   g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  AND2_X1   g0050(.A1(G33), .A2(G41), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n248), .B1(new_n210), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(KEYINPUT66), .ZN(new_n253));
  INV_X1    g0053(.A(new_n210), .ZN(new_n254));
  NAND2_X1  g0054(.A1(G33), .A2(G41), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT66), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n256), .A2(new_n257), .A3(new_n248), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n253), .A2(new_n258), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n250), .B1(new_n259), .B2(G238), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT3), .ZN(new_n261));
  INV_X1    g0061(.A(G33), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  AOI21_X1  g0064(.A(G1698), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G226), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n263), .A2(new_n264), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n267), .A2(G232), .A3(G1698), .ZN(new_n268));
  NAND2_X1  g0068(.A1(G33), .A2(G97), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n266), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  OAI21_X1  g0070(.A(KEYINPUT68), .B1(new_n251), .B2(new_n210), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT68), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n254), .A2(new_n272), .A3(new_n255), .ZN(new_n273));
  AND2_X1   g0073(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n270), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n260), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(KEYINPUT13), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT13), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n260), .A2(new_n278), .A3(new_n275), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G169), .ZN(new_n281));
  AND2_X1   g0081(.A1(new_n277), .A2(new_n279), .ZN(new_n282));
  AOI22_X1  g0082(.A1(new_n281), .A2(KEYINPUT14), .B1(new_n282), .B2(G179), .ZN(new_n283));
  INV_X1    g0083(.A(G169), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n284), .B1(new_n277), .B2(new_n279), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT14), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n283), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n211), .A2(new_n262), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G68), .ZN(new_n291));
  AOI22_X1  g0091(.A1(new_n290), .A2(G50), .B1(G20), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n211), .A2(G33), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n292), .B1(new_n202), .B2(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(new_n210), .ZN(new_n296));
  AND3_X1   g0096(.A1(new_n294), .A2(KEYINPUT11), .A3(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(new_n296), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n211), .A2(G1), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n298), .A2(G68), .A3(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G13), .ZN(new_n302));
  NOR3_X1   g0102(.A1(new_n302), .A2(new_n211), .A3(G1), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  OAI21_X1  g0104(.A(KEYINPUT12), .B1(new_n304), .B2(G68), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  NOR3_X1   g0106(.A1(new_n304), .A2(KEYINPUT12), .A3(G68), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n301), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  AOI21_X1  g0108(.A(KEYINPUT11), .B1(new_n294), .B2(new_n296), .ZN(new_n309));
  NOR3_X1   g0109(.A1(new_n297), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n280), .A2(G200), .ZN(new_n312));
  INV_X1    g0112(.A(G190), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n310), .B1(new_n280), .B2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  AOI22_X1  g0115(.A1(new_n288), .A2(new_n311), .B1(new_n312), .B2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(G58), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n317), .A2(new_n291), .ZN(new_n318));
  OAI21_X1  g0118(.A(G20), .B1(new_n318), .B2(new_n214), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n290), .A2(G159), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  AND2_X1   g0122(.A1(KEYINPUT3), .A2(G33), .ZN(new_n323));
  NOR2_X1   g0123(.A1(KEYINPUT3), .A2(G33), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT7), .ZN(new_n325));
  NOR4_X1   g0125(.A1(new_n323), .A2(new_n324), .A3(new_n325), .A4(G20), .ZN(new_n326));
  OAI21_X1  g0126(.A(KEYINPUT71), .B1(new_n323), .B2(new_n324), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT71), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n263), .A2(new_n328), .A3(new_n264), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n327), .A2(new_n329), .A3(new_n211), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n326), .B1(new_n330), .B2(new_n325), .ZN(new_n331));
  OAI211_X1 g0131(.A(KEYINPUT16), .B(new_n322), .C1(new_n331), .C2(new_n291), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT16), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n325), .B1(new_n267), .B2(G20), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n323), .A2(new_n324), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n335), .A2(KEYINPUT7), .A3(new_n211), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n291), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n333), .B1(new_n337), .B2(new_n321), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n332), .A2(new_n296), .A3(new_n338), .ZN(new_n339));
  XNOR2_X1  g0139(.A(KEYINPUT8), .B(G58), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n340), .A2(new_n299), .ZN(new_n341));
  XNOR2_X1  g0141(.A(new_n341), .B(KEYINPUT72), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n303), .A2(new_n296), .ZN(new_n343));
  AOI22_X1  g0143(.A1(new_n342), .A2(new_n343), .B1(new_n340), .B2(new_n303), .ZN(new_n344));
  AND2_X1   g0144(.A1(new_n339), .A2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(new_n250), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n346), .B1(new_n252), .B2(new_n230), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(G226), .A2(G1698), .ZN(new_n349));
  NAND2_X1  g0149(.A1(KEYINPUT73), .A2(G223), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n349), .B1(new_n350), .B2(G1698), .ZN(new_n351));
  AOI22_X1  g0151(.A1(new_n267), .A2(new_n351), .B1(G33), .B2(G87), .ZN(new_n352));
  INV_X1    g0152(.A(G1698), .ZN(new_n353));
  OAI211_X1 g0153(.A(G223), .B(new_n353), .C1(new_n323), .C2(new_n324), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT73), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  AND2_X1   g0156(.A1(new_n352), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n271), .A2(new_n273), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n348), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  OAI21_X1  g0159(.A(KEYINPUT74), .B1(new_n359), .B2(G179), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n358), .B1(new_n352), .B2(new_n356), .ZN(new_n361));
  NOR4_X1   g0161(.A1(new_n361), .A2(new_n347), .A3(KEYINPUT74), .A4(G179), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n359), .A2(new_n284), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n360), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  OAI21_X1  g0165(.A(KEYINPUT18), .B1(new_n345), .B2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT74), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n361), .A2(new_n347), .ZN(new_n368));
  INV_X1    g0168(.A(G179), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n367), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n368), .A2(G169), .ZN(new_n371));
  NOR3_X1   g0171(.A1(new_n370), .A2(new_n371), .A3(new_n362), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT18), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n339), .A2(new_n344), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n372), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  XNOR2_X1  g0175(.A(KEYINPUT75), .B(G190), .ZN(new_n376));
  NOR3_X1   g0176(.A1(new_n361), .A2(new_n347), .A3(new_n376), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n377), .B1(G200), .B2(new_n359), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n378), .A2(new_n344), .A3(new_n339), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT17), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n378), .A2(KEYINPUT17), .A3(new_n344), .A4(new_n339), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n366), .A2(new_n375), .A3(new_n381), .A4(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(G50), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n299), .A2(new_n385), .ZN(new_n386));
  AOI22_X1  g0186(.A1(new_n343), .A2(new_n386), .B1(new_n385), .B2(new_n303), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n340), .A2(new_n293), .ZN(new_n388));
  INV_X1    g0188(.A(G150), .ZN(new_n389));
  OAI22_X1  g0189(.A1(new_n201), .A2(new_n211), .B1(new_n289), .B2(new_n389), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n296), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n387), .A2(new_n391), .ZN(new_n392));
  XNOR2_X1  g0192(.A(new_n392), .B(KEYINPUT9), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n259), .A2(G226), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n394), .A2(KEYINPUT67), .A3(new_n346), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT67), .ZN(new_n396));
  INV_X1    g0196(.A(G226), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n397), .B1(new_n253), .B2(new_n258), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n396), .B1(new_n398), .B2(new_n250), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n353), .B1(new_n263), .B2(new_n264), .ZN(new_n400));
  AOI22_X1  g0200(.A1(new_n400), .A2(G223), .B1(new_n335), .B2(G77), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n265), .A2(G222), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(new_n274), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n395), .A2(new_n399), .A3(G190), .A4(new_n404), .ZN(new_n405));
  AND2_X1   g0205(.A1(new_n393), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n395), .A2(new_n399), .A3(new_n404), .ZN(new_n407));
  AND3_X1   g0207(.A1(new_n407), .A2(KEYINPUT70), .A3(G200), .ZN(new_n408));
  AOI21_X1  g0208(.A(KEYINPUT70), .B1(new_n407), .B2(G200), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n406), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(KEYINPUT10), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT10), .ZN(new_n412));
  OAI211_X1 g0212(.A(new_n406), .B(new_n412), .C1(new_n408), .C2(new_n409), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  OR2_X1    g0214(.A1(new_n407), .A2(G179), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n407), .A2(new_n284), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n415), .A2(new_n392), .A3(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n267), .A2(G232), .A3(new_n353), .ZN(new_n419));
  OAI211_X1 g0219(.A(G238), .B(G1698), .C1(new_n323), .C2(new_n324), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n335), .A2(G107), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n419), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(new_n274), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n252), .A2(KEYINPUT66), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n257), .B1(new_n256), .B2(new_n248), .ZN(new_n425));
  OAI21_X1  g0225(.A(G244), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n423), .A2(new_n426), .A3(new_n346), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(new_n284), .ZN(new_n428));
  XNOR2_X1  g0228(.A(KEYINPUT15), .B(G87), .ZN(new_n429));
  OAI22_X1  g0229(.A1(new_n429), .A2(new_n293), .B1(new_n211), .B2(new_n202), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n340), .A2(new_n289), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n296), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n303), .A2(new_n202), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n298), .A2(G77), .A3(new_n300), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n432), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n423), .A2(new_n426), .A3(new_n369), .A4(new_n346), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n428), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n435), .B1(new_n427), .B2(G200), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT69), .ZN(new_n439));
  OAI22_X1  g0239(.A1(new_n438), .A2(new_n439), .B1(new_n313), .B2(new_n427), .ZN(new_n440));
  AOI211_X1 g0240(.A(KEYINPUT69), .B(new_n435), .C1(new_n427), .C2(G200), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n437), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n418), .A2(new_n442), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n316), .A2(new_n384), .A3(new_n414), .A4(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  OAI211_X1 g0245(.A(G244), .B(new_n353), .C1(new_n323), .C2(new_n324), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(KEYINPUT4), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT4), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n267), .A2(new_n448), .A3(G244), .A4(new_n353), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  OAI211_X1 g0250(.A(G250), .B(G1698), .C1(new_n323), .C2(new_n324), .ZN(new_n451));
  NAND2_X1  g0251(.A1(G33), .A2(G283), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n450), .A2(new_n454), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n358), .B1(new_n455), .B2(KEYINPUT76), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n453), .B1(new_n447), .B2(new_n449), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT76), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n456), .A2(new_n459), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n251), .A2(new_n210), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n461), .A2(new_n249), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT77), .ZN(new_n463));
  XNOR2_X1  g0263(.A(KEYINPUT5), .B(G41), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n247), .A2(G45), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n462), .A2(new_n463), .A3(new_n464), .A4(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n256), .A2(G274), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n464), .A2(new_n466), .ZN(new_n469));
  OAI21_X1  g0269(.A(KEYINPUT77), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n461), .B1(new_n466), .B2(new_n464), .ZN(new_n471));
  AOI22_X1  g0271(.A1(new_n467), .A2(new_n470), .B1(G257), .B2(new_n471), .ZN(new_n472));
  AOI21_X1  g0272(.A(KEYINPUT78), .B1(new_n460), .B2(new_n472), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n274), .B1(new_n457), .B2(new_n458), .ZN(new_n474));
  AND3_X1   g0274(.A1(new_n450), .A2(new_n458), .A3(new_n454), .ZN(new_n475));
  OAI211_X1 g0275(.A(KEYINPUT78), .B(new_n472), .C1(new_n474), .C2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n284), .B1(new_n473), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n467), .A2(new_n470), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n471), .A2(G257), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n481), .B1(new_n456), .B2(new_n459), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n482), .A2(KEYINPUT79), .A3(new_n369), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT79), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n472), .B1(new_n474), .B2(new_n475), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n484), .B1(new_n485), .B2(G179), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT6), .ZN(new_n488));
  INV_X1    g0288(.A(G97), .ZN(new_n489));
  INV_X1    g0289(.A(G107), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NOR2_X1   g0291(.A1(G97), .A2(G107), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n488), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n490), .A2(KEYINPUT6), .A3(G97), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  AOI22_X1  g0295(.A1(new_n495), .A2(G20), .B1(G77), .B2(new_n290), .ZN(new_n496));
  AND2_X1   g0296(.A1(new_n334), .A2(new_n336), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n496), .B1(new_n497), .B2(new_n490), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(new_n296), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n303), .A2(new_n489), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n343), .B1(G1), .B2(new_n262), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(G97), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n499), .A2(new_n500), .A3(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n478), .A2(new_n487), .A3(new_n504), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n504), .B1(G200), .B2(new_n485), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT78), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n485), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(new_n476), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n506), .B1(new_n313), .B2(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n505), .A2(KEYINPUT80), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n505), .A2(new_n510), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT80), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT81), .ZN(new_n515));
  XNOR2_X1  g0315(.A(new_n465), .B(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(G250), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n461), .A2(new_n517), .ZN(new_n518));
  AOI22_X1  g0318(.A1(new_n516), .A2(new_n518), .B1(G274), .B2(new_n466), .ZN(new_n519));
  OAI211_X1 g0319(.A(G244), .B(G1698), .C1(new_n323), .C2(new_n324), .ZN(new_n520));
  OAI211_X1 g0320(.A(G238), .B(new_n353), .C1(new_n323), .C2(new_n324), .ZN(new_n521));
  NAND2_X1  g0321(.A1(G33), .A2(G116), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n520), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(new_n274), .ZN(new_n524));
  AND3_X1   g0324(.A1(new_n519), .A2(new_n524), .A3(G179), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n284), .B1(new_n519), .B2(new_n524), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT19), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n211), .B1(new_n269), .B2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(G87), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n492), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n211), .B(G68), .C1(new_n323), .C2(new_n324), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n528), .B1(new_n293), .B2(new_n489), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n296), .ZN(new_n536));
  INV_X1    g0336(.A(new_n429), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n343), .B(new_n537), .C1(G1), .C2(new_n262), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n429), .A2(new_n303), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n536), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(KEYINPUT82), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT82), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n536), .A2(new_n538), .A3(new_n542), .A4(new_n539), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n527), .B1(new_n544), .B2(KEYINPUT83), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT83), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n541), .A2(new_n546), .A3(new_n543), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n519), .A2(new_n524), .A3(G190), .ZN(new_n548));
  INV_X1    g0348(.A(G200), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n549), .B1(new_n519), .B2(new_n524), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n536), .B(new_n539), .C1(new_n530), .C2(new_n501), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  AOI22_X1  g0352(.A1(new_n545), .A2(new_n547), .B1(new_n548), .B2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(new_n553), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n304), .A2(G116), .ZN(new_n555));
  INV_X1    g0355(.A(G116), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n501), .A2(new_n556), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n452), .B(new_n211), .C1(G33), .C2(new_n489), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n556), .A2(G20), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n558), .A2(new_n296), .A3(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT20), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n560), .A2(new_n561), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n562), .B1(KEYINPUT84), .B2(new_n563), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n563), .A2(KEYINPUT84), .ZN(new_n565));
  INV_X1    g0365(.A(new_n565), .ZN(new_n566));
  AOI211_X1 g0366(.A(new_n555), .B(new_n557), .C1(new_n564), .C2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n400), .A2(G264), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n265), .A2(G257), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n335), .A2(G303), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n274), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n471), .A2(G270), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n572), .A2(new_n479), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(G200), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n567), .B(new_n575), .C1(new_n376), .C2(new_n574), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n555), .B1(new_n502), .B2(G116), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n563), .A2(KEYINPUT84), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n578), .B1(new_n561), .B2(new_n560), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n577), .B1(new_n579), .B2(new_n565), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n580), .A2(G169), .A3(new_n574), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT21), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n580), .A2(KEYINPUT21), .A3(G169), .A4(new_n574), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n574), .A2(new_n369), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(new_n580), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n576), .A2(new_n583), .A3(new_n584), .A4(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n267), .A2(new_n211), .A3(G87), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(KEYINPUT22), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT22), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n267), .A2(new_n590), .A3(new_n211), .A4(G87), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n522), .A2(G20), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT23), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n594), .B1(new_n211), .B2(G107), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n490), .A2(KEYINPUT23), .A3(G20), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n593), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n592), .A2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT24), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n592), .A2(KEYINPUT24), .A3(new_n597), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n600), .A2(new_n296), .A3(new_n601), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n343), .B(G107), .C1(G1), .C2(new_n262), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT85), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n604), .B(KEYINPUT25), .C1(new_n304), .C2(G107), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT25), .ZN(new_n606));
  AOI21_X1  g0406(.A(G107), .B1(new_n606), .B2(KEYINPUT85), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n303), .B(new_n607), .C1(KEYINPUT85), .C2(new_n606), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n603), .A2(new_n605), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(KEYINPUT86), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT86), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n603), .A2(new_n611), .A3(new_n605), .A4(new_n608), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n602), .A2(new_n613), .ZN(new_n614));
  OAI211_X1 g0414(.A(G257), .B(G1698), .C1(new_n323), .C2(new_n324), .ZN(new_n615));
  NAND2_X1  g0415(.A1(G33), .A2(G294), .ZN(new_n616));
  OAI211_X1 g0416(.A(G250), .B(new_n353), .C1(new_n323), .C2(new_n324), .ZN(new_n617));
  OAI211_X1 g0417(.A(new_n615), .B(new_n616), .C1(new_n617), .C2(KEYINPUT87), .ZN(new_n618));
  AND2_X1   g0418(.A1(new_n617), .A2(KEYINPUT87), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n274), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n471), .A2(G264), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n620), .A2(new_n479), .A3(new_n621), .ZN(new_n622));
  OR2_X1    g0422(.A1(new_n622), .A2(G179), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n284), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n614), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n620), .A2(new_n479), .A3(G190), .A4(new_n621), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n622), .A2(G200), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n602), .A2(new_n626), .A3(new_n627), .A4(new_n613), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n625), .A2(new_n628), .ZN(new_n629));
  NOR3_X1   g0429(.A1(new_n554), .A2(new_n587), .A3(new_n629), .ZN(new_n630));
  AND4_X1   g0430(.A1(new_n445), .A2(new_n511), .A3(new_n514), .A4(new_n630), .ZN(G372));
  INV_X1    g0431(.A(KEYINPUT90), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT89), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n407), .A2(G200), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT70), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n407), .A2(KEYINPUT70), .A3(G200), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n412), .B1(new_n638), .B2(new_n406), .ZN(new_n639));
  INV_X1    g0439(.A(new_n413), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n633), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n411), .A2(KEYINPUT89), .A3(new_n413), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n310), .B1(new_n283), .B2(new_n287), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n437), .B1(new_n315), .B2(new_n312), .ZN(new_n645));
  OAI21_X1  g0445(.A(KEYINPUT88), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n381), .A2(new_n382), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n287), .ZN(new_n649));
  OAI22_X1  g0449(.A1(new_n285), .A2(new_n286), .B1(new_n280), .B2(new_n369), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n311), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT88), .ZN(new_n652));
  INV_X1    g0452(.A(new_n437), .ZN(new_n653));
  INV_X1    g0453(.A(new_n312), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n653), .B1(new_n654), .B2(new_n314), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n651), .A2(new_n652), .A3(new_n655), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n646), .A2(new_n648), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n366), .A2(new_n375), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n643), .B1(new_n657), .B2(new_n659), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n632), .B1(new_n660), .B2(new_n418), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n651), .A2(new_n655), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n647), .B1(new_n662), .B2(KEYINPUT88), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n658), .B1(new_n663), .B2(new_n656), .ZN(new_n664));
  OAI211_X1 g0464(.A(KEYINPUT90), .B(new_n417), .C1(new_n664), .C2(new_n643), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n661), .A2(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(KEYINPUT26), .B1(new_n505), .B2(new_n554), .ZN(new_n667));
  AOI22_X1  g0467(.A1(new_n581), .A2(new_n582), .B1(new_n580), .B2(new_n585), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n668), .A2(new_n625), .A3(new_n584), .ZN(new_n669));
  OR2_X1    g0469(.A1(new_n525), .A2(new_n526), .ZN(new_n670));
  AOI22_X1  g0470(.A1(new_n670), .A2(new_n544), .B1(new_n548), .B2(new_n552), .ZN(new_n671));
  AND2_X1   g0471(.A1(new_n671), .A2(new_n628), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n505), .A2(new_n669), .A3(new_n510), .A4(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n670), .A2(new_n544), .ZN(new_n674));
  INV_X1    g0474(.A(new_n504), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n675), .B1(new_n509), .B2(new_n284), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT26), .ZN(new_n677));
  NAND4_X1  g0477(.A1(new_n676), .A2(new_n677), .A3(new_n487), .A4(new_n671), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n667), .A2(new_n673), .A3(new_n674), .A4(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n445), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n666), .A2(new_n680), .ZN(G369));
  NOR2_X1   g0481(.A1(new_n302), .A2(G20), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n682), .A2(KEYINPUT91), .A3(new_n247), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n247), .A2(new_n211), .A3(G13), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT91), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT27), .ZN(new_n688));
  OAI21_X1  g0488(.A(G213), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT92), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n687), .A2(new_n691), .A3(new_n688), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n691), .B1(new_n687), .B2(new_n688), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n690), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(KEYINPUT93), .ZN(new_n696));
  AND2_X1   g0496(.A1(new_n683), .A2(new_n686), .ZN(new_n697));
  OAI21_X1  g0497(.A(KEYINPUT92), .B1(new_n697), .B2(KEYINPUT27), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(new_n692), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT93), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n699), .A2(new_n700), .A3(new_n690), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n696), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g0502(.A(KEYINPUT94), .B(G343), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(new_n567), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n668), .A2(new_n584), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n708), .B1(new_n587), .B2(new_n706), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(G330), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n704), .A2(new_n614), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(new_n628), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(new_n625), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n625), .A2(new_n704), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n710), .A2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n625), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n719), .B1(new_n711), .B2(new_n628), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n707), .A2(new_n705), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n715), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n718), .A2(new_n723), .ZN(G399));
  NOR2_X1   g0524(.A1(new_n207), .A2(G41), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n531), .A2(G116), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n726), .A2(G1), .A3(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n728), .B1(new_n216), .B2(new_n726), .ZN(new_n729));
  XNOR2_X1  g0529(.A(new_n729), .B(KEYINPUT28), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n679), .A2(new_n705), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n731), .A2(KEYINPUT29), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT29), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n478), .A2(new_n487), .A3(new_n504), .A4(new_n671), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(KEYINPUT26), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n676), .A2(new_n553), .A3(new_n677), .A4(new_n487), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n673), .A2(new_n735), .A3(new_n674), .A4(new_n736), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n733), .B1(new_n737), .B2(new_n705), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n732), .A2(new_n738), .ZN(new_n739));
  NAND4_X1  g0539(.A1(new_n514), .A2(new_n511), .A3(new_n630), .A4(new_n705), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT31), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n519), .A2(new_n524), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n574), .A2(new_n622), .A3(new_n369), .A4(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(new_n482), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n620), .A2(new_n621), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n519), .A2(new_n524), .A3(G179), .ZN(new_n746));
  NOR3_X1   g0546(.A1(new_n574), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n508), .A2(new_n476), .A3(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT30), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n744), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n508), .A2(KEYINPUT30), .A3(new_n476), .A4(new_n747), .ZN(new_n751));
  AOI211_X1 g0551(.A(new_n741), .B(new_n705), .C1(new_n750), .C2(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n748), .A2(new_n749), .ZN(new_n753));
  INV_X1    g0553(.A(new_n744), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n753), .A2(new_n751), .A3(new_n754), .ZN(new_n755));
  AOI21_X1  g0555(.A(KEYINPUT31), .B1(new_n755), .B2(new_n704), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n752), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n740), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(G330), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n739), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n730), .B1(new_n761), .B2(G1), .ZN(G364));
  INV_X1    g0562(.A(new_n710), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n247), .B1(new_n682), .B2(G45), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n725), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n763), .A2(new_n766), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n767), .B1(G330), .B2(new_n709), .ZN(new_n768));
  INV_X1    g0568(.A(KEYINPUT95), .ZN(new_n769));
  AND2_X1   g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(G13), .A2(G33), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(G20), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  OR2_X1    g0574(.A1(new_n709), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n267), .A2(new_n206), .ZN(new_n776));
  INV_X1    g0576(.A(G355), .ZN(new_n777));
  OAI22_X1  g0577(.A1(new_n776), .A2(new_n777), .B1(G116), .B2(new_n206), .ZN(new_n778));
  INV_X1    g0578(.A(G45), .ZN(new_n779));
  OR2_X1    g0579(.A1(new_n240), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n327), .A2(new_n329), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(new_n206), .ZN(new_n783));
  INV_X1    g0583(.A(new_n216), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n783), .B1(new_n779), .B2(new_n784), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n778), .B1(new_n780), .B2(new_n785), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n254), .B1(new_n211), .B2(G169), .ZN(new_n787));
  OR2_X1    g0587(.A1(new_n787), .A2(KEYINPUT96), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n787), .A2(KEYINPUT96), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(new_n773), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n766), .B1(new_n786), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n211), .A2(G190), .ZN(new_n794));
  NOR2_X1   g0594(.A1(G179), .A2(G200), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n267), .B1(new_n797), .B2(G329), .ZN(new_n798));
  INV_X1    g0598(.A(G294), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n795), .A2(G190), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(G20), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n798), .B1(new_n799), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n369), .A2(G200), .ZN(new_n804));
  INV_X1    g0604(.A(KEYINPUT98), .ZN(new_n805));
  XNOR2_X1  g0605(.A(new_n804), .B(new_n805), .ZN(new_n806));
  NOR3_X1   g0606(.A1(new_n806), .A2(new_n211), .A3(G190), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n803), .B1(G283), .B2(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n211), .A2(new_n369), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(G200), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n810), .A2(new_n376), .ZN(new_n811));
  AND2_X1   g0611(.A1(new_n811), .A2(G326), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n809), .A2(new_n313), .A3(G200), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  XNOR2_X1  g0614(.A(KEYINPUT33), .B(G317), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n812), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n809), .A2(new_n549), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n817), .A2(new_n376), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n817), .A2(G190), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n818), .A2(G322), .B1(new_n819), .B2(G311), .ZN(new_n820));
  NOR3_X1   g0620(.A1(new_n806), .A2(new_n211), .A3(new_n313), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n821), .A2(G303), .ZN(new_n822));
  NAND4_X1  g0622(.A1(new_n808), .A2(new_n816), .A3(new_n820), .A4(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n807), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n824), .A2(new_n490), .ZN(new_n825));
  INV_X1    g0625(.A(new_n821), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n826), .A2(new_n530), .ZN(new_n827));
  INV_X1    g0627(.A(G159), .ZN(new_n828));
  NOR3_X1   g0628(.A1(new_n796), .A2(KEYINPUT32), .A3(new_n828), .ZN(new_n829));
  NOR4_X1   g0629(.A1(new_n825), .A2(new_n827), .A3(new_n335), .A4(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n801), .A2(G97), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n814), .A2(G68), .ZN(new_n832));
  OAI21_X1  g0632(.A(KEYINPUT32), .B1(new_n796), .B2(new_n828), .ZN(new_n833));
  NAND4_X1  g0633(.A1(new_n830), .A2(new_n831), .A3(new_n832), .A4(new_n833), .ZN(new_n834));
  AOI22_X1  g0634(.A1(new_n818), .A2(G58), .B1(new_n819), .B2(G77), .ZN(new_n835));
  INV_X1    g0635(.A(new_n811), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n835), .B1(new_n385), .B2(new_n836), .ZN(new_n837));
  XNOR2_X1  g0637(.A(new_n837), .B(KEYINPUT97), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n823), .B1(new_n834), .B2(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n793), .B1(new_n839), .B2(new_n790), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n770), .B1(new_n775), .B2(new_n840), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n841), .B1(new_n769), .B2(new_n768), .ZN(G396));
  INV_X1    g0642(.A(KEYINPUT101), .ZN(new_n843));
  INV_X1    g0643(.A(new_n703), .ZN(new_n844));
  NAND4_X1  g0644(.A1(new_n696), .A2(new_n435), .A3(new_n701), .A4(new_n844), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n845), .B1(new_n440), .B2(new_n441), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n846), .A2(new_n437), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n700), .B1(new_n699), .B2(new_n690), .ZN(new_n848));
  AOI211_X1 g0648(.A(KEYINPUT93), .B(new_n689), .C1(new_n698), .C2(new_n692), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n437), .B1(new_n850), .B2(new_n844), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n843), .B1(new_n847), .B2(new_n852), .ZN(new_n853));
  AOI211_X1 g0653(.A(KEYINPUT101), .B(new_n851), .C1(new_n846), .C2(new_n437), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n731), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n679), .A2(new_n705), .A3(new_n855), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n766), .B1(new_n859), .B2(new_n759), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n860), .B1(new_n759), .B2(new_n859), .ZN(new_n861));
  INV_X1    g0661(.A(new_n790), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(new_n772), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n766), .B1(new_n863), .B2(G77), .ZN(new_n864));
  XNOR2_X1  g0664(.A(new_n864), .B(KEYINPUT99), .ZN(new_n865));
  AOI22_X1  g0665(.A1(new_n811), .A2(G303), .B1(new_n819), .B2(G116), .ZN(new_n866));
  INV_X1    g0666(.A(G283), .ZN(new_n867));
  INV_X1    g0667(.A(new_n818), .ZN(new_n868));
  OAI221_X1 g0668(.A(new_n866), .B1(new_n867), .B2(new_n813), .C1(new_n799), .C2(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n826), .A2(new_n490), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n824), .A2(new_n530), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n797), .A2(G311), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n872), .A2(new_n335), .A3(new_n831), .ZN(new_n873));
  NOR4_X1   g0673(.A1(new_n869), .A2(new_n870), .A3(new_n871), .A4(new_n873), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n824), .A2(new_n291), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n875), .B1(G50), .B2(new_n821), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n782), .B1(G132), .B2(new_n797), .ZN(new_n877));
  OAI211_X1 g0677(.A(new_n876), .B(new_n877), .C1(new_n317), .C2(new_n802), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT34), .ZN(new_n879));
  AOI22_X1  g0679(.A1(G137), .A2(new_n811), .B1(new_n814), .B2(G150), .ZN(new_n880));
  INV_X1    g0680(.A(new_n819), .ZN(new_n881));
  XOR2_X1   g0681(.A(KEYINPUT100), .B(G143), .Z(new_n882));
  OAI221_X1 g0682(.A(new_n880), .B1(new_n828), .B2(new_n881), .C1(new_n868), .C2(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n878), .B1(new_n879), .B2(new_n883), .ZN(new_n884));
  OR2_X1    g0684(.A1(new_n883), .A2(new_n879), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n874), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  OAI221_X1 g0686(.A(new_n865), .B1(new_n862), .B2(new_n886), .C1(new_n855), .C2(new_n772), .ZN(new_n887));
  AND2_X1   g0687(.A1(new_n861), .A2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(G384));
  AOI211_X1 g0689(.A(new_n556), .B(new_n213), .C1(new_n495), .C2(KEYINPUT35), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n890), .B1(KEYINPUT35), .B2(new_n495), .ZN(new_n891));
  XOR2_X1   g0691(.A(new_n891), .B(KEYINPUT36), .Z(new_n892));
  OR3_X1    g0692(.A1(new_n216), .A2(new_n202), .A3(new_n318), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n385), .A2(G68), .ZN(new_n894));
  AOI211_X1 g0694(.A(new_n247), .B(G13), .C1(new_n893), .C2(new_n894), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n892), .A2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(G330), .ZN(new_n897));
  INV_X1    g0697(.A(new_n344), .ZN(new_n898));
  AND2_X1   g0698(.A1(new_n332), .A2(new_n296), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n322), .B1(new_n331), .B2(new_n291), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(new_n333), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n898), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n379), .B1(new_n902), .B2(new_n702), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n902), .A2(new_n365), .ZN(new_n904));
  OAI21_X1  g0704(.A(KEYINPUT37), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n372), .A2(new_n374), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n850), .A2(new_n374), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT37), .ZN(new_n908));
  NAND4_X1  g0708(.A1(new_n906), .A2(new_n907), .A3(new_n908), .A4(new_n379), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n905), .A2(new_n909), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n902), .A2(new_n702), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n383), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n910), .A2(KEYINPUT38), .A3(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n906), .A2(new_n907), .A3(new_n379), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(KEYINPUT37), .ZN(new_n915));
  INV_X1    g0715(.A(new_n907), .ZN(new_n916));
  AOI22_X1  g0716(.A1(new_n909), .A2(new_n915), .B1(new_n383), .B2(new_n916), .ZN(new_n917));
  XOR2_X1   g0717(.A(KEYINPUT103), .B(KEYINPUT38), .Z(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n913), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n704), .A2(new_n311), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n316), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n921), .B1(new_n283), .B2(new_n287), .ZN(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  NAND4_X1  g0725(.A1(new_n758), .A2(new_n855), .A3(new_n920), .A4(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(KEYINPUT40), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n856), .B1(new_n740), .B2(new_n757), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n910), .A2(new_n912), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT38), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(KEYINPUT40), .B1(new_n931), .B2(new_n913), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n928), .A2(new_n925), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n927), .A2(new_n933), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n444), .B1(new_n740), .B2(new_n757), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n897), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n936), .B1(new_n935), .B2(new_n934), .ZN(new_n937));
  XOR2_X1   g0737(.A(new_n937), .B(KEYINPUT104), .Z(new_n938));
  AOI21_X1  g0738(.A(new_n923), .B1(new_n316), .B2(new_n921), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n939), .B1(new_n858), .B2(new_n852), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n931), .A2(new_n913), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT39), .ZN(new_n943));
  INV_X1    g0743(.A(new_n913), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n915), .A2(new_n909), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n383), .A2(new_n916), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n919), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n943), .B1(new_n944), .B2(new_n947), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n931), .A2(KEYINPUT39), .A3(new_n913), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n644), .A2(KEYINPUT102), .A3(new_n705), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT102), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n951), .B1(new_n651), .B2(new_n704), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n948), .A2(new_n949), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n658), .A2(new_n702), .ZN(new_n955));
  AND3_X1   g0755(.A1(new_n942), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n445), .B1(new_n732), .B2(new_n738), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n666), .A2(new_n957), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n956), .B(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n938), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n960), .B1(new_n247), .B2(new_n682), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT105), .ZN(new_n962));
  OAI22_X1  g0762(.A1(new_n961), .A2(new_n962), .B1(new_n938), .B2(new_n959), .ZN(new_n963));
  AND2_X1   g0763(.A1(new_n961), .A2(new_n962), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n896), .B1(new_n963), .B2(new_n964), .ZN(G367));
  NAND3_X1  g0765(.A1(new_n704), .A2(new_n551), .A3(new_n674), .ZN(new_n966));
  AND2_X1   g0766(.A1(new_n704), .A2(new_n551), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n966), .B1(new_n967), .B2(new_n671), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n968), .B(KEYINPUT106), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT43), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n971), .B(KEYINPUT107), .ZN(new_n972));
  INV_X1    g0772(.A(new_n969), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(KEYINPUT43), .ZN(new_n974));
  INV_X1    g0774(.A(new_n505), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(new_n704), .ZN(new_n976));
  OAI211_X1 g0776(.A(new_n505), .B(new_n510), .C1(new_n675), .C2(new_n705), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n721), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n713), .A2(new_n715), .A3(new_n980), .ZN(new_n981));
  OAI21_X1  g0781(.A(KEYINPUT42), .B1(new_n979), .B2(new_n981), .ZN(new_n982));
  AND2_X1   g0782(.A1(new_n510), .A2(new_n719), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n705), .B1(new_n983), .B2(new_n975), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  NOR3_X1   g0785(.A1(new_n979), .A2(KEYINPUT42), .A3(new_n981), .ZN(new_n986));
  OAI211_X1 g0786(.A(new_n972), .B(new_n974), .C1(new_n985), .C2(new_n986), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n971), .B(KEYINPUT107), .Z(new_n988));
  OAI21_X1  g0788(.A(new_n974), .B1(new_n985), .B2(new_n986), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n987), .A2(new_n990), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n718), .A2(new_n979), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n991), .B(new_n992), .ZN(new_n993));
  XOR2_X1   g0793(.A(new_n725), .B(KEYINPUT41), .Z(new_n994));
  INV_X1    g0794(.A(KEYINPUT45), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n995), .B1(new_n979), .B2(new_n722), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n723), .A2(KEYINPUT45), .A3(new_n978), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT44), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n999), .B1(new_n978), .B2(new_n723), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n979), .A2(KEYINPUT44), .A3(new_n722), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n998), .A2(new_n1002), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n1003), .A2(new_n717), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n718), .B1(new_n998), .B2(new_n1002), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n716), .A2(new_n721), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1007), .A2(new_n981), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n763), .B(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT108), .ZN(new_n1010));
  NAND4_X1  g0810(.A1(new_n1009), .A2(new_n739), .A3(new_n1010), .A4(new_n759), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1009), .A2(new_n739), .A3(new_n759), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1012), .A2(KEYINPUT108), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1006), .A2(new_n1011), .A3(new_n1013), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n994), .B1(new_n1014), .B2(new_n761), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n993), .B1(new_n1015), .B2(new_n765), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n791), .B1(new_n206), .B2(new_n429), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n783), .A2(new_n236), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n766), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT46), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1020), .B1(new_n826), .B2(new_n556), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n821), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n814), .A2(G294), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n811), .A2(G311), .B1(new_n819), .B2(G283), .ZN(new_n1024));
  NAND4_X1  g0824(.A1(new_n1021), .A2(new_n1022), .A3(new_n1023), .A4(new_n1024), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n818), .A2(G303), .B1(G107), .B2(new_n801), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n781), .B1(G317), .B2(new_n797), .ZN(new_n1027));
  OAI211_X1 g0827(.A(new_n1026), .B(new_n1027), .C1(new_n824), .C2(new_n489), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(G50), .A2(new_n819), .B1(new_n814), .B2(G159), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n1029), .B1(new_n836), .B2(new_n882), .C1(new_n389), .C2(new_n868), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n821), .A2(G58), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n807), .A2(G77), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n802), .A2(new_n291), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n335), .B1(new_n797), .B2(G137), .ZN(new_n1035));
  NAND4_X1  g0835(.A1(new_n1031), .A2(new_n1032), .A3(new_n1034), .A4(new_n1035), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n1025), .A2(new_n1028), .B1(new_n1030), .B2(new_n1036), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(KEYINPUT109), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT47), .ZN(new_n1039));
  OR2_X1    g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n862), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1019), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(new_n973), .B2(new_n774), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1016), .A2(new_n1043), .ZN(G387));
  OAI22_X1  g0844(.A1(new_n776), .A2(new_n727), .B1(G107), .B2(new_n206), .ZN(new_n1045));
  OR2_X1    g0845(.A1(new_n233), .A2(new_n779), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n727), .ZN(new_n1047));
  AOI211_X1 g0847(.A(G45), .B(new_n1047), .C1(G68), .C2(G77), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n340), .A2(G50), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT50), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n783), .B1(new_n1048), .B2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1045), .B1(new_n1046), .B2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n766), .B1(new_n1052), .B2(new_n792), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n818), .A2(G317), .B1(new_n819), .B2(G303), .ZN(new_n1054));
  OR2_X1    g0854(.A1(new_n1054), .A2(KEYINPUT110), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1054), .A2(KEYINPUT110), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(G322), .A2(new_n811), .B1(new_n814), .B2(G311), .ZN(new_n1057));
  AND3_X1   g0857(.A1(new_n1055), .A2(new_n1056), .A3(new_n1057), .ZN(new_n1058));
  OR2_X1    g0858(.A1(new_n1058), .A2(KEYINPUT48), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1058), .A2(KEYINPUT48), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n821), .A2(G294), .B1(G283), .B2(new_n801), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1059), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT49), .ZN(new_n1063));
  OR2_X1    g0863(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n824), .A2(new_n556), .ZN(new_n1066));
  AOI211_X1 g0866(.A(new_n781), .B(new_n1066), .C1(G326), .C2(new_n797), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1064), .A2(new_n1065), .A3(new_n1067), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n824), .A2(new_n489), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n811), .A2(G159), .B1(new_n819), .B2(G68), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n1070), .B(new_n781), .C1(new_n389), .C2(new_n796), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n826), .A2(new_n202), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n537), .A2(new_n801), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n1073), .B1(new_n340), .B2(new_n813), .C1(new_n868), .C2(new_n385), .ZN(new_n1074));
  OR4_X1    g0874(.A1(new_n1069), .A2(new_n1071), .A3(new_n1072), .A4(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1068), .A2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1053), .B1(new_n1076), .B2(new_n790), .ZN(new_n1077));
  INV_X1    g0877(.A(KEYINPUT111), .ZN(new_n1078));
  AND2_X1   g0878(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1079), .B1(new_n716), .B2(new_n773), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1080), .B1(new_n1078), .B2(new_n1077), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n1009), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n760), .A2(new_n1082), .A3(KEYINPUT112), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1083), .A2(new_n725), .A3(new_n1012), .ZN(new_n1084));
  AOI21_X1  g0884(.A(KEYINPUT112), .B1(new_n760), .B2(new_n1082), .ZN(new_n1085));
  OAI221_X1 g0885(.A(new_n1081), .B1(new_n764), .B2(new_n1082), .C1(new_n1084), .C2(new_n1085), .ZN(G393));
  NOR2_X1   g0886(.A1(new_n760), .A2(new_n1082), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n1014), .B(new_n725), .C1(new_n1087), .C2(new_n1006), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1006), .A2(new_n765), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n791), .B1(new_n489), .B2(new_n206), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n245), .A2(new_n783), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n766), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  AOI211_X1 g0892(.A(new_n267), .B(new_n825), .C1(G322), .C2(new_n797), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(G311), .A2(new_n818), .B1(new_n811), .B2(G317), .ZN(new_n1094));
  XOR2_X1   g0894(.A(new_n1094), .B(KEYINPUT52), .Z(new_n1095));
  OAI211_X1 g0895(.A(new_n1093), .B(new_n1095), .C1(new_n867), .C2(new_n826), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n814), .A2(G303), .B1(G116), .B2(new_n801), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1097), .B1(new_n799), .B2(new_n881), .ZN(new_n1098));
  XNOR2_X1  g0898(.A(new_n1098), .B(KEYINPUT113), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(G150), .A2(new_n811), .B1(new_n818), .B2(G159), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(new_n1100), .B(KEYINPUT51), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n871), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n881), .A2(new_n340), .B1(new_n385), .B2(new_n813), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1103), .B1(G77), .B2(new_n801), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n821), .A2(G68), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n882), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n782), .B1(new_n797), .B2(new_n1106), .ZN(new_n1107));
  NAND4_X1  g0907(.A1(new_n1102), .A2(new_n1104), .A3(new_n1105), .A4(new_n1107), .ZN(new_n1108));
  OAI22_X1  g0908(.A1(new_n1096), .A2(new_n1099), .B1(new_n1101), .B2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1092), .B1(new_n1109), .B2(new_n790), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1110), .B1(new_n978), .B2(new_n774), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1088), .A2(new_n1089), .A3(new_n1111), .ZN(G390));
  NAND2_X1  g0912(.A1(new_n948), .A2(new_n949), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1113), .A2(new_n771), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(G116), .A2(new_n818), .B1(new_n814), .B2(G107), .ZN(new_n1115));
  OAI221_X1 g0915(.A(new_n1115), .B1(new_n489), .B2(new_n881), .C1(new_n867), .C2(new_n836), .ZN(new_n1116));
  OAI221_X1 g0916(.A(new_n335), .B1(new_n796), .B2(new_n799), .C1(new_n802), .C2(new_n202), .ZN(new_n1117));
  NOR4_X1   g0917(.A1(new_n1116), .A2(new_n827), .A3(new_n875), .A4(new_n1117), .ZN(new_n1118));
  OR2_X1    g0918(.A1(new_n1118), .A2(KEYINPUT116), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1118), .A2(KEYINPUT116), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n821), .A2(G150), .ZN(new_n1121));
  XOR2_X1   g0921(.A(new_n1121), .B(KEYINPUT53), .Z(new_n1122));
  AOI22_X1  g0922(.A1(new_n814), .A2(G137), .B1(G159), .B2(new_n801), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(KEYINPUT54), .B(G143), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n818), .A2(G132), .B1(new_n819), .B2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n807), .A2(G50), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n811), .A2(G128), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n335), .B1(new_n797), .B2(G125), .ZN(new_n1129));
  AND3_X1   g0929(.A1(new_n1127), .A2(new_n1128), .A3(new_n1129), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n1122), .A2(new_n1123), .A3(new_n1126), .A4(new_n1130), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1119), .A2(new_n1120), .A3(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(new_n790), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n862), .A2(new_n340), .A3(new_n772), .ZN(new_n1134));
  NAND4_X1  g0934(.A1(new_n1114), .A2(new_n766), .A3(new_n1133), .A4(new_n1134), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(new_n1135), .B(KEYINPUT117), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1113), .B1(new_n940), .B2(new_n953), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n737), .A2(new_n855), .A3(new_n705), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1138), .A2(new_n852), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1139), .A2(new_n925), .ZN(new_n1140));
  AND3_X1   g0940(.A1(new_n920), .A2(new_n952), .A3(new_n950), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1137), .A2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n758), .A2(G330), .A3(new_n855), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n1144), .A2(new_n939), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1143), .A2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n928), .A2(G330), .A3(new_n925), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1137), .A2(new_n1142), .A3(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1136), .B1(new_n1149), .B2(new_n764), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n858), .A2(new_n852), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n925), .B1(new_n928), .B2(G330), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1151), .B1(new_n1145), .B2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n897), .B1(new_n740), .B2(new_n757), .ZN(new_n1154));
  INV_X1    g0954(.A(KEYINPUT114), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n856), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n759), .A2(KEYINPUT114), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n925), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1147), .A2(new_n852), .A3(new_n1138), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1153), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1154), .A2(new_n445), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n666), .A2(new_n1161), .A3(new_n957), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1160), .A2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(new_n1149), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1165), .A2(new_n725), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n1164), .A2(new_n1149), .ZN(new_n1167));
  OAI21_X1  g0967(.A(KEYINPUT115), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1167), .ZN(new_n1169));
  INV_X1    g0969(.A(KEYINPUT115), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n726), .B1(new_n1164), .B2(new_n1149), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1169), .A2(new_n1170), .A3(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1150), .B1(new_n1168), .B2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(G378));
  AOI211_X1 g0974(.A(new_n1033), .B(new_n1072), .C1(G283), .C2(new_n797), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n781), .A2(G41), .ZN(new_n1176));
  OAI211_X1 g0976(.A(new_n1175), .B(new_n1176), .C1(new_n317), .C2(new_n824), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n818), .A2(G107), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n814), .A2(G97), .ZN(new_n1179));
  AND2_X1   g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  OAI221_X1 g0980(.A(new_n1180), .B1(new_n556), .B2(new_n836), .C1(new_n429), .C2(new_n881), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n1177), .A2(new_n1181), .ZN(new_n1182));
  OR2_X1    g0982(.A1(new_n1182), .A2(KEYINPUT58), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1182), .A2(KEYINPUT58), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n385), .B1(G33), .B2(G41), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n1183), .B(new_n1184), .C1(new_n1176), .C2(new_n1185), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(G137), .A2(new_n819), .B1(new_n814), .B2(G132), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(new_n811), .A2(G125), .B1(G150), .B2(new_n801), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(new_n821), .A2(new_n1125), .B1(G128), .B2(new_n818), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT118), .ZN(new_n1190));
  AND2_X1   g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n1187), .B(new_n1188), .C1(new_n1191), .C2(new_n1192), .ZN(new_n1193));
  OR2_X1    g0993(.A1(new_n1193), .A2(KEYINPUT59), .ZN(new_n1194));
  AOI211_X1 g0994(.A(G33), .B(G41), .C1(new_n797), .C2(G124), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1195), .B1(new_n824), .B2(new_n828), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1196), .B1(new_n1193), .B2(KEYINPUT59), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1186), .B1(new_n1194), .B2(new_n1197), .ZN(new_n1198));
  OAI221_X1 g0998(.A(new_n766), .B1(G50), .B2(new_n863), .C1(new_n1198), .C2(new_n862), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n641), .A2(new_n417), .A3(new_n642), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n850), .A2(new_n392), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1200), .A2(new_n1202), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n641), .A2(new_n417), .A3(new_n642), .A4(new_n1201), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  XNOR2_X1  g1005(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(new_n1205), .B(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1199), .B1(new_n1207), .B2(new_n771), .ZN(new_n1208));
  AND3_X1   g1008(.A1(new_n758), .A2(new_n855), .A3(new_n925), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n1209), .A2(new_n932), .B1(new_n926), .B2(KEYINPUT40), .ZN(new_n1210));
  NOR3_X1   g1010(.A1(new_n1210), .A2(new_n1207), .A3(new_n897), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1206), .ZN(new_n1212));
  XNOR2_X1  g1012(.A(new_n1205), .B(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(new_n934), .B2(G330), .ZN(new_n1214));
  OAI21_X1  g1014(.A(KEYINPUT119), .B1(new_n1211), .B2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1215), .A2(new_n956), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1207), .B1(new_n1210), .B2(new_n897), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n934), .A2(G330), .A3(new_n1213), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n956), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1219), .A2(KEYINPUT119), .A3(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1216), .A2(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1208), .B1(new_n1222), .B2(new_n765), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n855), .B1(new_n759), .B2(KEYINPUT114), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n939), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1145), .A2(new_n1139), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1144), .A2(new_n939), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1228), .A2(new_n1147), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n1226), .A2(new_n1227), .B1(new_n1151), .B2(new_n1229), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1163), .B1(new_n1149), .B2(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(KEYINPUT57), .B1(new_n1222), .B2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1231), .A2(KEYINPUT57), .ZN(new_n1233));
  AND3_X1   g1033(.A1(new_n1217), .A2(new_n956), .A3(new_n1218), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n956), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n725), .B1(new_n1233), .B2(new_n1236), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1223), .B1(new_n1232), .B2(new_n1237), .ZN(G375));
  NOR2_X1   g1038(.A1(new_n1230), .A2(new_n1162), .ZN(new_n1239));
  OAI211_X1 g1039(.A(new_n1162), .B(new_n1153), .C1(new_n1158), .C2(new_n1159), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  NOR3_X1   g1041(.A1(new_n1239), .A2(new_n1241), .A3(new_n994), .ZN(new_n1242));
  XNOR2_X1  g1042(.A(new_n1242), .B(KEYINPUT120), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n766), .B1(new_n863), .B2(G68), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n819), .A2(G107), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n814), .A2(G116), .ZN(new_n1246));
  AND2_X1   g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  OAI221_X1 g1047(.A(new_n1247), .B1(new_n867), .B2(new_n868), .C1(new_n799), .C2(new_n836), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n267), .B1(new_n797), .B2(G303), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1032), .A2(new_n1073), .A3(new_n1249), .ZN(new_n1250));
  AOI211_X1 g1050(.A(new_n1248), .B(new_n1250), .C1(G97), .C2(new_n821), .ZN(new_n1251));
  OR2_X1    g1051(.A1(new_n1251), .A2(KEYINPUT121), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1251), .A2(KEYINPUT121), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n818), .A2(G137), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1254), .B1(new_n385), .B2(new_n802), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1255), .B1(G132), .B2(new_n811), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n782), .B1(G128), .B2(new_n797), .ZN(new_n1257));
  AOI22_X1  g1057(.A1(G150), .A2(new_n819), .B1(new_n814), .B2(new_n1125), .ZN(new_n1258));
  AOI22_X1  g1058(.A1(G58), .A2(new_n807), .B1(new_n821), .B2(G159), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1256), .A2(new_n1257), .A3(new_n1258), .A4(new_n1259), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1252), .A2(new_n1253), .A3(new_n1260), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1244), .B1(new_n1261), .B2(new_n790), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1262), .B1(new_n925), .B2(new_n772), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1263), .B1(new_n1230), .B2(new_n764), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1243), .A2(new_n1265), .ZN(G381));
  INV_X1    g1066(.A(G390), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1267), .A2(new_n888), .ZN(new_n1268));
  OR3_X1    g1068(.A1(new_n1268), .A2(G396), .A3(G393), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1150), .B1(new_n1169), .B2(new_n1171), .ZN(new_n1270));
  OAI211_X1 g1070(.A(new_n1223), .B(new_n1270), .C1(new_n1232), .C2(new_n1237), .ZN(new_n1271));
  NOR4_X1   g1071(.A1(new_n1269), .A2(G381), .A3(G387), .A4(new_n1271), .ZN(new_n1272));
  XOR2_X1   g1072(.A(new_n1272), .B(KEYINPUT122), .Z(G407));
  AND2_X1   g1073(.A1(new_n703), .A2(G213), .ZN(new_n1274));
  XNOR2_X1  g1074(.A(new_n1274), .B(KEYINPUT123), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1275), .ZN(new_n1276));
  OAI211_X1 g1076(.A(G407), .B(G213), .C1(new_n1271), .C2(new_n1276), .ZN(G409));
  XNOR2_X1  g1077(.A(G393), .B(G396), .ZN(new_n1278));
  AND3_X1   g1078(.A1(new_n1016), .A2(G390), .A3(new_n1043), .ZN(new_n1279));
  AOI21_X1  g1079(.A(G390), .B1(new_n1016), .B2(new_n1043), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1278), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(G387), .A2(new_n1267), .ZN(new_n1282));
  XOR2_X1   g1082(.A(G393), .B(G396), .Z(new_n1283));
  NAND3_X1  g1083(.A1(new_n1016), .A2(G390), .A3(new_n1043), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1282), .A2(new_n1283), .A3(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1281), .A2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1217), .A2(new_n956), .A3(new_n1218), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1208), .B1(new_n1289), .B2(new_n765), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1220), .B1(new_n1219), .B2(KEYINPUT119), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT119), .ZN(new_n1292));
  AOI211_X1 g1092(.A(new_n1292), .B(new_n956), .C1(new_n1217), .C2(new_n1218), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1231), .B1(new_n1291), .B2(new_n1293), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1290), .B1(new_n994), .B2(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1295), .A2(new_n1270), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1296), .B1(G375), .B2(new_n1173), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1297), .A2(new_n1276), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT125), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT60), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1301), .B1(new_n1160), .B2(new_n1163), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n725), .B1(new_n1302), .B2(new_n1241), .ZN(new_n1303));
  NOR3_X1   g1103(.A1(new_n1160), .A2(new_n1163), .A3(new_n1301), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1300), .B1(new_n1303), .B2(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1164), .A2(KEYINPUT60), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1306), .A2(new_n1240), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1304), .ZN(new_n1308));
  NAND4_X1  g1108(.A1(new_n1307), .A2(new_n1308), .A3(KEYINPUT125), .A4(new_n725), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1305), .A2(new_n1309), .ZN(new_n1310));
  AOI21_X1  g1110(.A(G384), .B1(new_n1310), .B2(new_n1265), .ZN(new_n1311));
  AOI211_X1 g1111(.A(new_n888), .B(new_n1264), .C1(new_n1305), .C2(new_n1309), .ZN(new_n1312));
  NOR2_X1   g1112(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT62), .ZN(new_n1315));
  NOR2_X1   g1115(.A1(new_n1314), .A2(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1297), .A2(KEYINPUT124), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT124), .ZN(new_n1318));
  OAI211_X1 g1118(.A(new_n1296), .B(new_n1318), .C1(G375), .C2(new_n1173), .ZN(new_n1319));
  NAND4_X1  g1119(.A1(new_n1317), .A2(new_n1276), .A3(new_n1313), .A4(new_n1319), .ZN(new_n1320));
  AOI22_X1  g1120(.A1(new_n1299), .A2(new_n1316), .B1(new_n1320), .B2(new_n1315), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n726), .B1(new_n1306), .B2(new_n1240), .ZN(new_n1322));
  AOI21_X1  g1122(.A(KEYINPUT125), .B1(new_n1322), .B2(new_n1308), .ZN(new_n1323));
  NOR3_X1   g1123(.A1(new_n1303), .A2(new_n1300), .A3(new_n1304), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n1265), .B1(new_n1323), .B2(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1325), .A2(new_n888), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1310), .A2(G384), .A3(new_n1265), .ZN(new_n1327));
  NAND4_X1  g1127(.A1(new_n1326), .A2(G2897), .A3(new_n1275), .A4(new_n1327), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1275), .A2(G2897), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n1329), .B1(new_n1311), .B2(new_n1312), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1328), .A2(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1331), .A2(new_n1298), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT61), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1332), .A2(new_n1333), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n1286), .B1(new_n1321), .B2(new_n1334), .ZN(new_n1335));
  AND3_X1   g1135(.A1(new_n1281), .A2(new_n1285), .A3(new_n1333), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1326), .A2(KEYINPUT63), .A3(new_n1327), .ZN(new_n1337));
  OAI21_X1  g1137(.A(new_n1336), .B1(new_n1298), .B2(new_n1337), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1317), .A2(new_n1276), .A3(new_n1319), .ZN(new_n1339));
  AOI21_X1  g1139(.A(new_n1338), .B1(new_n1339), .B2(new_n1331), .ZN(new_n1340));
  XOR2_X1   g1140(.A(KEYINPUT126), .B(KEYINPUT63), .Z(new_n1341));
  NAND2_X1  g1141(.A1(new_n1320), .A2(new_n1341), .ZN(new_n1342));
  AOI21_X1  g1142(.A(KEYINPUT127), .B1(new_n1340), .B2(new_n1342), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1339), .A2(new_n1331), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(new_n1281), .A2(new_n1285), .A3(new_n1333), .ZN(new_n1345));
  INV_X1    g1145(.A(new_n1337), .ZN(new_n1346));
  AOI21_X1  g1146(.A(new_n1345), .B1(new_n1299), .B2(new_n1346), .ZN(new_n1347));
  AND4_X1   g1147(.A1(KEYINPUT127), .A2(new_n1342), .A3(new_n1344), .A4(new_n1347), .ZN(new_n1348));
  OAI21_X1  g1148(.A(new_n1335), .B1(new_n1343), .B2(new_n1348), .ZN(G405));
  NOR2_X1   g1149(.A1(G375), .A2(new_n1173), .ZN(new_n1350));
  AOI21_X1  g1150(.A(new_n1350), .B1(G375), .B2(new_n1270), .ZN(new_n1351));
  XNOR2_X1  g1151(.A(new_n1351), .B(new_n1314), .ZN(new_n1352));
  XNOR2_X1  g1152(.A(new_n1352), .B(new_n1286), .ZN(G402));
endmodule


