//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 0 1 1 0 0 1 0 1 0 1 0 1 0 0 0 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 1 0 0 0 0 1 0 1 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:50 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n669, new_n670, new_n671, new_n672, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n684,
    new_n685, new_n686, new_n688, new_n689, new_n690, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n720, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979;
  INV_X1    g000(.A(KEYINPUT11), .ZN(new_n187));
  INV_X1    g001(.A(G134), .ZN(new_n188));
  OAI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G137), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(G137), .ZN(new_n190));
  INV_X1    g004(.A(G137), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n191), .A2(KEYINPUT11), .A3(G134), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n189), .A2(new_n190), .A3(new_n192), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n193), .A2(G131), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G131), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n191), .A2(G134), .ZN(new_n197));
  AOI21_X1  g011(.A(new_n196), .B1(new_n190), .B2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G143), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G146), .ZN(new_n201));
  OAI21_X1  g015(.A(KEYINPUT65), .B1(new_n200), .B2(G146), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT65), .ZN(new_n203));
  INV_X1    g017(.A(G146), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n203), .A2(new_n204), .A3(G143), .ZN(new_n205));
  AND2_X1   g019(.A1(new_n202), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G128), .ZN(new_n207));
  OAI21_X1  g021(.A(KEYINPUT1), .B1(new_n200), .B2(G146), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT68), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n207), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n204), .A2(G143), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n211), .A2(KEYINPUT68), .A3(KEYINPUT1), .ZN(new_n212));
  AOI22_X1  g026(.A1(new_n201), .A2(new_n206), .B1(new_n210), .B2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT1), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n201), .A2(new_n211), .A3(new_n214), .A4(G128), .ZN(new_n215));
  INV_X1    g029(.A(new_n215), .ZN(new_n216));
  OAI211_X1 g030(.A(new_n195), .B(new_n199), .C1(new_n213), .C2(new_n216), .ZN(new_n217));
  XOR2_X1   g031(.A(G116), .B(G119), .Z(new_n218));
  XNOR2_X1  g032(.A(KEYINPUT2), .B(G113), .ZN(new_n219));
  XNOR2_X1  g033(.A(new_n218), .B(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(KEYINPUT67), .A2(G131), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n193), .A2(new_n223), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n189), .A2(new_n192), .A3(new_n222), .A4(new_n190), .ZN(new_n225));
  AND3_X1   g039(.A1(new_n224), .A2(KEYINPUT69), .A3(new_n225), .ZN(new_n226));
  AOI21_X1  g040(.A(KEYINPUT69), .B1(new_n224), .B2(new_n225), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  AND2_X1   g042(.A1(KEYINPUT0), .A2(G128), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n201), .A2(new_n211), .A3(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(KEYINPUT66), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT66), .ZN(new_n232));
  NAND4_X1  g046(.A1(new_n201), .A2(new_n211), .A3(new_n229), .A4(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n202), .A2(new_n205), .A3(new_n201), .ZN(new_n235));
  OR3_X1    g049(.A1(KEYINPUT64), .A2(KEYINPUT0), .A3(G128), .ZN(new_n236));
  OAI21_X1  g050(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n237));
  INV_X1    g051(.A(new_n229), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n235), .A2(new_n236), .A3(new_n237), .A4(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n234), .A2(new_n239), .ZN(new_n240));
  OAI211_X1 g054(.A(new_n217), .B(new_n221), .C1(new_n228), .C2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT72), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT28), .ZN(new_n243));
  AND3_X1   g057(.A1(new_n241), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n242), .B1(new_n241), .B2(new_n243), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  XNOR2_X1  g060(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n247));
  XNOR2_X1  g061(.A(new_n247), .B(G101), .ZN(new_n248));
  NOR2_X1   g062(.A1(G237), .A2(G953), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G210), .ZN(new_n250));
  XNOR2_X1  g064(.A(new_n248), .B(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT71), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n208), .A2(new_n209), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n253), .A2(G128), .A3(new_n212), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n216), .B1(new_n254), .B2(new_n235), .ZN(new_n255));
  NOR3_X1   g069(.A1(new_n255), .A2(new_n194), .A3(new_n198), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n224), .A2(new_n225), .ZN(new_n257));
  AND3_X1   g071(.A1(new_n257), .A2(new_n239), .A3(new_n234), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n220), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n241), .A2(new_n259), .ZN(new_n260));
  XOR2_X1   g074(.A(KEYINPUT70), .B(KEYINPUT28), .Z(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n252), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  AOI211_X1 g077(.A(KEYINPUT71), .B(new_n261), .C1(new_n241), .C2(new_n259), .ZN(new_n264));
  OAI211_X1 g078(.A(new_n246), .B(new_n251), .C1(new_n263), .C2(new_n264), .ZN(new_n265));
  OAI211_X1 g079(.A(new_n217), .B(KEYINPUT30), .C1(new_n228), .C2(new_n240), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT30), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n267), .B1(new_n256), .B2(new_n258), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n266), .A2(new_n268), .A3(new_n220), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(new_n241), .ZN(new_n270));
  INV_X1    g084(.A(new_n251), .ZN(new_n271));
  AOI21_X1  g085(.A(KEYINPUT29), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n265), .A2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(G902), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT69), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n257), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n224), .A2(KEYINPUT69), .A3(new_n225), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n240), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n278), .A2(new_n256), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n279), .A2(new_n221), .ZN(new_n280));
  NOR3_X1   g094(.A1(new_n278), .A2(new_n256), .A3(new_n220), .ZN(new_n281));
  OR2_X1    g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(KEYINPUT28), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n283), .A2(KEYINPUT29), .A3(new_n251), .A4(new_n246), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n273), .A2(new_n274), .A3(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(G472), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n246), .B1(new_n263), .B2(new_n264), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n269), .A2(new_n251), .A3(new_n241), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT31), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND4_X1  g104(.A1(new_n269), .A2(KEYINPUT31), .A3(new_n251), .A4(new_n241), .ZN(new_n291));
  AOI22_X1  g105(.A1(new_n287), .A2(new_n271), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NOR2_X1   g106(.A1(G472), .A2(G902), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  NOR3_X1   g108(.A1(new_n292), .A2(KEYINPUT32), .A3(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT32), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n290), .A2(new_n291), .ZN(new_n297));
  OAI21_X1  g111(.A(KEYINPUT72), .B1(new_n281), .B2(KEYINPUT28), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n241), .A2(new_n242), .A3(new_n243), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n260), .A2(new_n262), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(KEYINPUT71), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n260), .A2(new_n252), .A3(new_n262), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n300), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n297), .B1(new_n304), .B2(new_n251), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n296), .B1(new_n305), .B2(new_n293), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n286), .B1(new_n295), .B2(new_n306), .ZN(new_n307));
  XOR2_X1   g121(.A(KEYINPUT24), .B(G110), .Z(new_n308));
  XNOR2_X1  g122(.A(G119), .B(G128), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT23), .ZN(new_n311));
  INV_X1    g125(.A(G119), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n311), .B1(new_n312), .B2(G128), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(G128), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n207), .A2(KEYINPUT23), .A3(G119), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n313), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(G110), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT73), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n316), .A2(KEYINPUT73), .A3(G110), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(G125), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(G140), .ZN(new_n323));
  INV_X1    g137(.A(G140), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G125), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n323), .A2(new_n325), .A3(KEYINPUT74), .ZN(new_n326));
  OR3_X1    g140(.A1(new_n324), .A2(KEYINPUT74), .A3(G125), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(KEYINPUT16), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n325), .A2(KEYINPUT16), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  AOI21_X1  g145(.A(G146), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT16), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n333), .B1(new_n326), .B2(new_n327), .ZN(new_n334));
  NOR3_X1   g148(.A1(new_n334), .A2(new_n204), .A3(new_n330), .ZN(new_n335));
  OAI211_X1 g149(.A(new_n310), .B(new_n321), .C1(new_n332), .C2(new_n335), .ZN(new_n336));
  NOR3_X1   g150(.A1(new_n324), .A2(KEYINPUT74), .A3(G125), .ZN(new_n337));
  XNOR2_X1  g151(.A(G125), .B(G140), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n337), .B1(new_n338), .B2(KEYINPUT74), .ZN(new_n339));
  OAI211_X1 g153(.A(G146), .B(new_n331), .C1(new_n339), .C2(new_n333), .ZN(new_n340));
  OAI22_X1  g154(.A1(new_n316), .A2(G110), .B1(new_n308), .B2(new_n309), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n338), .A2(new_n204), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n340), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n336), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(KEYINPUT76), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT76), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n336), .A2(new_n346), .A3(new_n343), .ZN(new_n347));
  XNOR2_X1  g161(.A(KEYINPUT75), .B(KEYINPUT22), .ZN(new_n348));
  XNOR2_X1  g162(.A(new_n348), .B(G137), .ZN(new_n349));
  INV_X1    g163(.A(G953), .ZN(new_n350));
  AND3_X1   g164(.A1(new_n350), .A2(G221), .A3(G234), .ZN(new_n351));
  XOR2_X1   g165(.A(new_n349), .B(new_n351), .Z(new_n352));
  NAND3_X1  g166(.A1(new_n345), .A2(new_n347), .A3(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(new_n352), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n344), .A2(new_n354), .A3(KEYINPUT76), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(new_n274), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(KEYINPUT25), .ZN(new_n358));
  INV_X1    g172(.A(G217), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n359), .B1(G234), .B2(new_n274), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT25), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n356), .A2(new_n361), .A3(new_n274), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n358), .A2(new_n360), .A3(new_n362), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n360), .A2(G902), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n356), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  OAI21_X1  g181(.A(G214), .B1(G237), .B2(G902), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n322), .B1(new_n234), .B2(new_n239), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(KEYINPUT81), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT81), .ZN(new_n373));
  AOI22_X1  g187(.A1(new_n370), .A2(new_n373), .B1(new_n322), .B2(new_n255), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT7), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n350), .A2(G224), .ZN(new_n376));
  XNOR2_X1  g190(.A(new_n376), .B(KEYINPUT82), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT83), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n375), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n377), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(KEYINPUT83), .ZN(new_n381));
  NAND4_X1  g195(.A1(new_n372), .A2(new_n374), .A3(new_n379), .A4(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT5), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n383), .A2(new_n312), .A3(G116), .ZN(new_n384));
  OAI211_X1 g198(.A(G113), .B(new_n384), .C1(new_n218), .C2(new_n383), .ZN(new_n385));
  OR2_X1    g199(.A1(new_n218), .A2(new_n219), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT77), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT3), .ZN(new_n389));
  INV_X1    g203(.A(G107), .ZN(new_n390));
  NAND4_X1  g204(.A1(new_n388), .A2(new_n389), .A3(new_n390), .A4(G104), .ZN(new_n391));
  INV_X1    g205(.A(G104), .ZN(new_n392));
  AOI22_X1  g206(.A1(new_n392), .A2(G107), .B1(KEYINPUT77), .B2(KEYINPUT3), .ZN(new_n393));
  OAI22_X1  g207(.A1(new_n392), .A2(G107), .B1(KEYINPUT77), .B2(KEYINPUT3), .ZN(new_n394));
  INV_X1    g208(.A(G101), .ZN(new_n395));
  NAND4_X1  g209(.A1(new_n391), .A2(new_n393), .A3(new_n394), .A4(new_n395), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n390), .A2(G104), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n392), .A2(G107), .ZN(new_n398));
  OAI21_X1  g212(.A(G101), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n396), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n387), .A2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(new_n400), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n402), .A2(new_n386), .A3(new_n385), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  XOR2_X1   g218(.A(G110), .B(G122), .Z(new_n405));
  XOR2_X1   g219(.A(new_n405), .B(KEYINPUT8), .Z(new_n406));
  NAND2_X1  g220(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  NOR3_X1   g221(.A1(new_n213), .A2(G125), .A3(new_n216), .ZN(new_n408));
  OAI22_X1  g222(.A1(new_n408), .A2(new_n370), .B1(new_n375), .B2(new_n377), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n391), .A2(new_n393), .A3(new_n394), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(G101), .ZN(new_n411));
  NAND4_X1  g225(.A1(new_n411), .A2(KEYINPUT78), .A3(KEYINPUT4), .A4(new_n396), .ZN(new_n412));
  NAND2_X1  g226(.A1(KEYINPUT78), .A2(KEYINPUT4), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n410), .A2(G101), .A3(new_n413), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n412), .A2(new_n220), .A3(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(new_n405), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n415), .A2(new_n403), .A3(new_n416), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n382), .A2(new_n407), .A3(new_n409), .A4(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n415), .A2(new_n403), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(new_n405), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n420), .A2(KEYINPUT6), .A3(new_n417), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT6), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n419), .A2(new_n422), .A3(new_n405), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  AND3_X1   g238(.A1(new_n372), .A2(new_n374), .A3(new_n380), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n380), .B1(new_n372), .B2(new_n374), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  OAI211_X1 g241(.A(new_n274), .B(new_n418), .C1(new_n424), .C2(new_n427), .ZN(new_n428));
  OAI21_X1  g242(.A(G210), .B1(G237), .B2(G902), .ZN(new_n429));
  XNOR2_X1  g243(.A(new_n429), .B(KEYINPUT84), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  OAI211_X1 g245(.A(new_n421), .B(new_n423), .C1(new_n425), .C2(new_n426), .ZN(new_n432));
  INV_X1    g246(.A(new_n430), .ZN(new_n433));
  NAND4_X1  g247(.A1(new_n432), .A2(new_n274), .A3(new_n433), .A4(new_n418), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n369), .B1(new_n431), .B2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(G469), .ZN(new_n436));
  XNOR2_X1  g250(.A(G110), .B(G140), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n350), .A2(G227), .ZN(new_n438));
  XNOR2_X1  g252(.A(new_n437), .B(new_n438), .ZN(new_n439));
  OAI21_X1  g253(.A(KEYINPUT79), .B1(new_n226), .B2(new_n227), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT79), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n276), .A2(new_n441), .A3(new_n277), .ZN(new_n442));
  AND2_X1   g256(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  OAI211_X1 g257(.A(new_n402), .B(KEYINPUT10), .C1(new_n213), .C2(new_n216), .ZN(new_n444));
  AOI22_X1  g258(.A1(new_n208), .A2(G128), .B1(new_n201), .B2(new_n211), .ZN(new_n445));
  OAI211_X1 g259(.A(new_n399), .B(new_n396), .C1(new_n216), .C2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT10), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n412), .A2(new_n414), .ZN(new_n449));
  OAI211_X1 g263(.A(new_n444), .B(new_n448), .C1(new_n449), .C2(new_n240), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n443), .A2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n276), .A2(new_n277), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n450), .A2(new_n453), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n439), .B1(new_n452), .B2(new_n454), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n439), .B1(new_n443), .B2(new_n450), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n255), .A2(new_n400), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(new_n446), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(new_n453), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT80), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT12), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n459), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  AOI22_X1  g276(.A1(new_n457), .A2(new_n446), .B1(new_n276), .B2(new_n277), .ZN(new_n463));
  OAI21_X1  g277(.A(KEYINPUT80), .B1(new_n463), .B2(KEYINPUT12), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n458), .A2(KEYINPUT12), .A3(new_n257), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n456), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  OAI211_X1 g281(.A(new_n436), .B(new_n274), .C1(new_n455), .C2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(new_n456), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(new_n454), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n451), .B1(new_n465), .B2(new_n466), .ZN(new_n471));
  OAI211_X1 g285(.A(new_n470), .B(G469), .C1(new_n471), .C2(new_n439), .ZN(new_n472));
  NAND2_X1  g286(.A1(G469), .A2(G902), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n468), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(G221), .ZN(new_n475));
  XNOR2_X1  g289(.A(KEYINPUT9), .B(G234), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n475), .B1(new_n477), .B2(new_n274), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n249), .A2(G143), .A3(G214), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(G143), .B1(new_n249), .B2(G214), .ZN(new_n482));
  OAI21_X1  g296(.A(G131), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT17), .ZN(new_n484));
  INV_X1    g298(.A(G237), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n485), .A2(new_n350), .A3(G214), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(new_n200), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n487), .A2(new_n196), .A3(new_n480), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n483), .A2(new_n484), .A3(new_n488), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n204), .B1(new_n334), .B2(new_n330), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n487), .A2(new_n480), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n491), .A2(KEYINPUT17), .A3(G131), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n489), .A2(new_n490), .A3(new_n340), .A4(new_n492), .ZN(new_n493));
  XNOR2_X1  g307(.A(G113), .B(G122), .ZN(new_n494));
  XNOR2_X1  g308(.A(new_n494), .B(new_n392), .ZN(new_n495));
  NAND2_X1  g309(.A1(KEYINPUT18), .A2(G131), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n491), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n487), .A2(KEYINPUT18), .A3(G131), .A4(new_n480), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  OAI211_X1 g313(.A(KEYINPUT85), .B(new_n342), .C1(new_n328), .C2(new_n204), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT85), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n339), .A2(new_n501), .A3(G146), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n499), .A2(new_n500), .A3(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n493), .A2(new_n495), .A3(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n495), .B1(new_n493), .B2(new_n503), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n274), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(G475), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT20), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n326), .A2(new_n327), .A3(KEYINPUT19), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT86), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n323), .A2(new_n325), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n511), .B1(new_n512), .B2(KEYINPUT19), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT19), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n338), .A2(KEYINPUT86), .A3(new_n514), .ZN(new_n515));
  NAND4_X1  g329(.A1(new_n510), .A2(new_n513), .A3(new_n204), .A4(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n483), .A2(new_n488), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n516), .A2(new_n340), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(new_n503), .ZN(new_n519));
  INV_X1    g333(.A(new_n495), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(new_n504), .ZN(new_n522));
  NOR2_X1   g336(.A1(G475), .A2(G902), .ZN(new_n523));
  XNOR2_X1  g337(.A(new_n523), .B(KEYINPUT87), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n509), .B1(new_n522), .B2(new_n525), .ZN(new_n526));
  AOI211_X1 g340(.A(KEYINPUT20), .B(new_n524), .C1(new_n521), .C2(new_n504), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n508), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(G234), .A2(G237), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n529), .A2(G952), .A3(new_n350), .ZN(new_n530));
  XOR2_X1   g344(.A(KEYINPUT21), .B(G898), .Z(new_n531));
  NAND3_X1  g345(.A1(new_n529), .A2(G902), .A3(G953), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(G116), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n535), .A2(KEYINPUT14), .A3(G122), .ZN(new_n536));
  XNOR2_X1  g350(.A(G116), .B(G122), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  OAI211_X1 g352(.A(G107), .B(new_n536), .C1(new_n538), .C2(KEYINPUT14), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n537), .A2(new_n390), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT88), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n541), .B1(new_n200), .B2(G128), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n207), .A2(KEYINPUT88), .A3(G143), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n200), .A2(G128), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n546), .A2(G134), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n188), .B1(new_n544), .B2(new_n545), .ZN(new_n548));
  OAI211_X1 g362(.A(new_n539), .B(new_n540), .C1(new_n547), .C2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT13), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n544), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n546), .A2(new_n551), .A3(G134), .ZN(new_n552));
  XNOR2_X1  g366(.A(new_n537), .B(new_n390), .ZN(new_n553));
  OAI211_X1 g367(.A(new_n544), .B(new_n545), .C1(new_n550), .C2(new_n188), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  NOR3_X1   g369(.A1(new_n476), .A2(new_n359), .A3(G953), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n549), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n556), .B1(new_n549), .B2(new_n555), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n274), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT89), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(KEYINPUT15), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n561), .A2(KEYINPUT15), .ZN(new_n564));
  OAI21_X1  g378(.A(G478), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n560), .A2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(new_n559), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(new_n557), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n569), .A2(new_n274), .A3(new_n565), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  NOR3_X1   g385(.A1(new_n528), .A2(new_n534), .A3(new_n571), .ZN(new_n572));
  AND4_X1   g386(.A1(new_n435), .A2(new_n474), .A3(new_n479), .A4(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n307), .A2(new_n367), .A3(new_n573), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n574), .B(G101), .ZN(G3));
  NAND2_X1  g389(.A1(new_n474), .A2(new_n479), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n576), .A2(new_n366), .ZN(new_n577));
  INV_X1    g391(.A(G472), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n578), .B1(new_n305), .B2(new_n274), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n292), .A2(new_n294), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AND2_X1   g395(.A1(new_n577), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n569), .A2(KEYINPUT33), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT33), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n568), .A2(new_n584), .A3(new_n557), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n583), .A2(new_n585), .A3(G478), .ZN(new_n586));
  OR2_X1    g400(.A1(new_n560), .A2(G478), .ZN(new_n587));
  NAND2_X1  g401(.A1(G478), .A2(G902), .ZN(new_n588));
  AND3_X1   g402(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  AND4_X1   g403(.A1(new_n435), .A2(new_n533), .A3(new_n528), .A4(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n582), .A2(new_n590), .ZN(new_n591));
  XNOR2_X1  g405(.A(KEYINPUT90), .B(KEYINPUT34), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n592), .B(new_n392), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n591), .B(new_n593), .ZN(G6));
  AOI211_X1 g408(.A(new_n369), .B(new_n534), .C1(new_n431), .C2(new_n434), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n522), .A2(new_n525), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(KEYINPUT20), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT91), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n522), .A2(new_n509), .A3(new_n525), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  OAI21_X1  g414(.A(KEYINPUT91), .B1(new_n526), .B2(new_n527), .ZN(new_n601));
  AND4_X1   g415(.A1(new_n571), .A2(new_n600), .A3(new_n508), .A4(new_n601), .ZN(new_n602));
  AOI21_X1  g416(.A(KEYINPUT92), .B1(new_n595), .B2(new_n602), .ZN(new_n603));
  AND4_X1   g417(.A1(KEYINPUT92), .A2(new_n435), .A3(new_n602), .A4(new_n533), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n582), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  XOR2_X1   g419(.A(KEYINPUT35), .B(G107), .Z(new_n606));
  XNOR2_X1  g420(.A(new_n605), .B(new_n606), .ZN(G9));
  AOI21_X1  g421(.A(new_n361), .B1(new_n356), .B2(new_n274), .ZN(new_n608));
  AOI211_X1 g422(.A(KEYINPUT25), .B(G902), .C1(new_n353), .C2(new_n355), .ZN(new_n609));
  INV_X1    g423(.A(new_n360), .ZN(new_n610));
  NOR3_X1   g424(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n352), .A2(KEYINPUT36), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n612), .B(new_n344), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(new_n364), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  OAI21_X1  g429(.A(KEYINPUT93), .B1(new_n611), .B2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT93), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n363), .A2(new_n617), .A3(new_n614), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n619), .A2(new_n573), .A3(new_n581), .ZN(new_n620));
  XOR2_X1   g434(.A(new_n620), .B(KEYINPUT37), .Z(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(G110), .ZN(G12));
  INV_X1    g436(.A(new_n435), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n576), .A2(new_n623), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n350), .A2(G900), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n625), .A2(G902), .A3(new_n529), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT94), .ZN(new_n627));
  OR2_X1    g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n626), .A2(new_n627), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n628), .A2(new_n530), .A3(new_n629), .ZN(new_n630));
  XOR2_X1   g444(.A(new_n630), .B(KEYINPUT95), .Z(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  AND2_X1   g446(.A1(new_n602), .A2(new_n632), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n307), .A2(new_n619), .A3(new_n624), .A4(new_n633), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(G128), .ZN(G30));
  INV_X1    g449(.A(new_n576), .ZN(new_n636));
  XOR2_X1   g450(.A(new_n631), .B(KEYINPUT39), .Z(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  XOR2_X1   g452(.A(new_n638), .B(KEYINPUT40), .Z(new_n639));
  NOR2_X1   g453(.A1(new_n611), .A2(new_n615), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n431), .A2(new_n434), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT96), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(KEYINPUT38), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n642), .B(KEYINPUT96), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT38), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n641), .B1(new_n645), .B2(new_n648), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n639), .A2(new_n368), .A3(new_n649), .ZN(new_n650));
  AOI22_X1  g464(.A1(new_n597), .A2(new_n599), .B1(G475), .B2(new_n507), .ZN(new_n651));
  INV_X1    g465(.A(new_n571), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n271), .B1(new_n280), .B2(new_n281), .ZN(new_n654));
  OR2_X1    g468(.A1(new_n654), .A2(KEYINPUT97), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n654), .A2(KEYINPUT97), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n655), .A2(new_n288), .A3(new_n656), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n578), .B1(new_n657), .B2(new_n274), .ZN(new_n658));
  OAI21_X1  g472(.A(KEYINPUT32), .B1(new_n292), .B2(new_n294), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n305), .A2(new_n296), .A3(new_n293), .ZN(new_n660));
  AOI211_X1 g474(.A(KEYINPUT98), .B(new_n658), .C1(new_n659), .C2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT98), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n659), .A2(new_n660), .ZN(new_n663));
  INV_X1    g477(.A(new_n658), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n662), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n653), .B1(new_n661), .B2(new_n665), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n650), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(new_n200), .ZN(G45));
  NAND3_X1  g482(.A1(new_n589), .A2(new_n528), .A3(new_n632), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n307), .A2(new_n619), .A3(new_n624), .A4(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(KEYINPUT99), .B(G146), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(G48));
  NAND2_X1  g487(.A1(new_n465), .A2(new_n466), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n454), .B1(new_n450), .B2(new_n443), .ZN(new_n675));
  INV_X1    g489(.A(new_n439), .ZN(new_n676));
  AOI22_X1  g490(.A1(new_n674), .A2(new_n469), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  OAI21_X1  g491(.A(G469), .B1(new_n677), .B2(G902), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n678), .A2(new_n479), .A3(new_n468), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n307), .A2(new_n367), .A3(new_n590), .A4(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(KEYINPUT41), .B(G113), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G15));
  NAND3_X1  g497(.A1(new_n307), .A2(new_n367), .A3(new_n680), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n603), .A2(new_n604), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(new_n535), .ZN(G18));
  NOR2_X1   g501(.A1(new_n623), .A2(new_n679), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n307), .A2(new_n619), .A3(new_n572), .A4(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(KEYINPUT100), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G119), .ZN(G21));
  NAND2_X1  g505(.A1(new_n653), .A2(KEYINPUT101), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT101), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n693), .B1(new_n651), .B2(new_n652), .ZN(new_n694));
  AND4_X1   g508(.A1(new_n435), .A2(new_n692), .A3(new_n533), .A4(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n283), .A2(new_n246), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(new_n271), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n294), .B1(new_n697), .B2(new_n297), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n579), .A2(new_n698), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n695), .A2(new_n367), .A3(new_n680), .A4(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G122), .ZN(G24));
  NOR3_X1   g515(.A1(new_n640), .A2(new_n579), .A3(new_n698), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT102), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n669), .B(new_n703), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n702), .A2(new_n688), .A3(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G125), .ZN(G27));
  NOR2_X1   g520(.A1(new_n478), .A2(new_n369), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n431), .A2(new_n434), .A3(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  XOR2_X1   g523(.A(new_n473), .B(KEYINPUT103), .Z(new_n710));
  NAND3_X1  g524(.A1(new_n468), .A2(new_n472), .A3(new_n710), .ZN(new_n711));
  AND2_X1   g525(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n307), .A2(new_n704), .A3(new_n712), .A4(new_n367), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT42), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n366), .B1(new_n663), .B2(new_n286), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n716), .A2(KEYINPUT42), .A3(new_n704), .A4(new_n712), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G131), .ZN(G33));
  AND4_X1   g533(.A1(new_n307), .A2(new_n367), .A3(new_n712), .A4(new_n633), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(new_n188), .ZN(G36));
  INV_X1    g535(.A(new_n581), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n723));
  NOR3_X1   g537(.A1(new_n723), .A2(new_n528), .A3(KEYINPUT43), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT104), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n528), .B(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(new_n589), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n724), .B1(new_n727), .B2(KEYINPUT43), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n722), .A2(new_n728), .A3(new_n641), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT44), .ZN(new_n730));
  OR2_X1    g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n642), .A2(new_n369), .ZN(new_n732));
  XOR2_X1   g546(.A(new_n732), .B(KEYINPUT105), .Z(new_n733));
  AND2_X1   g547(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n470), .B1(new_n471), .B2(new_n439), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT45), .ZN(new_n736));
  OR2_X1    g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n735), .A2(new_n736), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n737), .A2(G469), .A3(new_n738), .ZN(new_n739));
  AOI21_X1  g553(.A(KEYINPUT46), .B1(new_n739), .B2(new_n710), .ZN(new_n740));
  INV_X1    g554(.A(new_n468), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n739), .A2(KEYINPUT46), .A3(new_n710), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n478), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  AND2_X1   g558(.A1(new_n744), .A2(new_n637), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n729), .A2(new_n730), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n734), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G137), .ZN(G39));
  INV_X1    g562(.A(new_n732), .ZN(new_n749));
  NOR3_X1   g563(.A1(new_n307), .A2(new_n367), .A3(new_n749), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n744), .A2(KEYINPUT47), .ZN(new_n751));
  INV_X1    g565(.A(new_n743), .ZN(new_n752));
  NOR3_X1   g566(.A1(new_n752), .A2(new_n740), .A3(new_n741), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT47), .ZN(new_n754));
  NOR3_X1   g568(.A1(new_n753), .A2(new_n754), .A3(new_n478), .ZN(new_n755));
  OAI211_X1 g569(.A(new_n670), .B(new_n750), .C1(new_n751), .C2(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(KEYINPUT106), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n744), .A2(KEYINPUT47), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n754), .B1(new_n753), .B2(new_n478), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT106), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n760), .A2(new_n761), .A3(new_n670), .A4(new_n750), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n757), .A2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT107), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n763), .B(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(new_n324), .ZN(G42));
  OR2_X1    g580(.A1(G952), .A2(G953), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT54), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT53), .ZN(new_n769));
  AND3_X1   g583(.A1(new_n600), .A2(new_n601), .A3(new_n508), .ZN(new_n770));
  AND3_X1   g584(.A1(new_n307), .A2(new_n619), .A3(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT112), .ZN(new_n772));
  NOR3_X1   g586(.A1(new_n576), .A2(new_n571), .A3(new_n631), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n771), .A2(new_n772), .A3(new_n732), .A4(new_n773), .ZN(new_n774));
  OAI211_X1 g588(.A(new_n571), .B(new_n508), .C1(new_n526), .C2(new_n527), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n775), .B1(new_n651), .B2(new_n723), .ZN(new_n776));
  AND3_X1   g590(.A1(new_n435), .A2(new_n776), .A3(new_n533), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n577), .A2(new_n581), .A3(new_n777), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n574), .A2(new_n620), .A3(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n307), .A2(new_n619), .A3(new_n770), .A4(new_n732), .ZN(new_n781));
  INV_X1    g595(.A(new_n773), .ZN(new_n782));
  OAI21_X1  g596(.A(KEYINPUT112), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  AND4_X1   g597(.A1(new_n718), .A2(new_n774), .A3(new_n780), .A4(new_n783), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n689), .B1(new_n684), .B2(new_n685), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n681), .A2(new_n700), .ZN(new_n786));
  NOR3_X1   g600(.A1(new_n785), .A2(new_n786), .A3(new_n720), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n702), .A2(new_n704), .A3(new_n712), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT113), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT52), .ZN(new_n790));
  AND3_X1   g604(.A1(new_n692), .A2(new_n435), .A3(new_n694), .ZN(new_n791));
  AND4_X1   g605(.A1(new_n479), .A2(new_n640), .A3(new_n632), .A4(new_n711), .ZN(new_n792));
  OAI211_X1 g606(.A(new_n791), .B(new_n792), .C1(new_n661), .C2(new_n665), .ZN(new_n793));
  INV_X1    g607(.A(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n634), .A2(new_n705), .A3(new_n671), .ZN(new_n795));
  OAI211_X1 g609(.A(new_n789), .B(new_n790), .C1(new_n794), .C2(new_n795), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n784), .A2(new_n787), .A3(new_n788), .A4(new_n796), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n790), .B1(new_n794), .B2(new_n795), .ZN(new_n798));
  AND3_X1   g612(.A1(new_n634), .A2(new_n705), .A3(new_n671), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n799), .A2(KEYINPUT52), .A3(new_n793), .ZN(new_n800));
  AND3_X1   g614(.A1(new_n798), .A2(new_n800), .A3(KEYINPUT113), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n769), .B1(new_n797), .B2(new_n801), .ZN(new_n802));
  AOI22_X1  g616(.A1(new_n663), .A2(new_n286), .B1(new_n616), .B2(new_n618), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n803), .A2(new_n770), .A3(new_n732), .A4(new_n773), .ZN(new_n804));
  AOI22_X1  g618(.A1(new_n715), .A2(new_n717), .B1(new_n804), .B2(KEYINPUT112), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n781), .A2(new_n782), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n779), .B1(new_n806), .B2(new_n772), .ZN(new_n807));
  AND4_X1   g621(.A1(new_n787), .A2(new_n805), .A3(new_n807), .A4(new_n788), .ZN(new_n808));
  AOI21_X1  g622(.A(KEYINPUT52), .B1(new_n799), .B2(new_n793), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n803), .B(new_n624), .C1(new_n633), .C2(new_n670), .ZN(new_n810));
  AND4_X1   g624(.A1(KEYINPUT52), .A2(new_n793), .A3(new_n810), .A4(new_n705), .ZN(new_n811));
  OAI211_X1 g625(.A(new_n808), .B(KEYINPUT53), .C1(new_n809), .C2(new_n811), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n768), .B1(new_n802), .B2(new_n812), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n798), .A2(new_n800), .A3(KEYINPUT113), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n808), .A2(KEYINPUT53), .A3(new_n796), .A4(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT114), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n809), .A2(new_n811), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n787), .A2(new_n805), .A3(new_n807), .A4(new_n788), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n769), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n815), .A2(new_n816), .A3(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(new_n796), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n818), .A2(new_n821), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n822), .A2(KEYINPUT114), .A3(KEYINPUT53), .A4(new_n814), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n820), .A2(new_n823), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n813), .B1(new_n824), .B2(new_n768), .ZN(new_n825));
  INV_X1    g639(.A(new_n728), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n699), .A2(new_n367), .ZN(new_n827));
  NOR3_X1   g641(.A1(new_n826), .A2(new_n827), .A3(new_n530), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n678), .A2(new_n468), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n829), .B(KEYINPUT108), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n830), .A2(new_n478), .ZN(new_n831));
  OAI211_X1 g645(.A(new_n733), .B(new_n828), .C1(new_n760), .C2(new_n831), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n832), .B1(KEYINPUT115), .B2(KEYINPUT51), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n645), .A2(new_n648), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n827), .A2(new_n679), .ZN(new_n835));
  INV_X1    g649(.A(new_n530), .ZN(new_n836));
  AND3_X1   g650(.A1(new_n728), .A2(new_n369), .A3(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n834), .A2(new_n835), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n838), .A2(KEYINPUT50), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT50), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n834), .A2(new_n837), .A3(new_n840), .A4(new_n835), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n709), .A2(KEYINPUT116), .A3(new_n468), .A4(new_n678), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT116), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n843), .B1(new_n829), .B2(new_n708), .ZN(new_n844));
  AND3_X1   g658(.A1(new_n842), .A2(new_n836), .A3(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n845), .A2(new_n702), .A3(new_n728), .ZN(new_n846));
  AND3_X1   g660(.A1(new_n839), .A2(new_n841), .A3(new_n846), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n661), .A2(new_n665), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n848), .A2(new_n367), .A3(new_n845), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT117), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n848), .A2(KEYINPUT117), .A3(new_n367), .A4(new_n845), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n851), .A2(new_n651), .A3(new_n723), .A4(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n847), .A2(new_n853), .ZN(new_n854));
  OR2_X1    g668(.A1(new_n833), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n828), .A2(new_n688), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n851), .A2(new_n852), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n589), .A2(new_n528), .ZN(new_n858));
  OAI211_X1 g672(.A(G952), .B(new_n350), .C1(new_n857), .C2(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n854), .A2(KEYINPUT118), .ZN(new_n860));
  OR2_X1    g674(.A1(new_n760), .A2(new_n831), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT115), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n861), .A2(new_n862), .A3(new_n733), .A4(new_n828), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT118), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n847), .A2(new_n864), .A3(new_n853), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n860), .A2(new_n863), .A3(new_n833), .A4(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT51), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n859), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n825), .A2(new_n855), .A3(new_n856), .A4(new_n868), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n845), .A2(new_n716), .A3(new_n728), .ZN(new_n870));
  XNOR2_X1  g684(.A(KEYINPUT119), .B(KEYINPUT48), .ZN(new_n871));
  XNOR2_X1  g685(.A(new_n870), .B(new_n871), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n767), .B1(new_n869), .B2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT49), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n707), .B1(new_n830), .B2(new_n874), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n875), .A2(new_n366), .A3(new_n727), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n876), .B(KEYINPUT109), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n830), .A2(new_n874), .ZN(new_n878));
  XOR2_X1   g692(.A(new_n878), .B(KEYINPUT110), .Z(new_n879));
  NAND4_X1  g693(.A1(new_n877), .A2(new_n848), .A3(new_n834), .A4(new_n879), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n880), .B(KEYINPUT111), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n873), .A2(new_n881), .ZN(G75));
  NAND4_X1  g696(.A1(new_n820), .A2(G902), .A3(new_n430), .A4(new_n823), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT120), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n424), .A2(new_n427), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n886), .A2(new_n432), .ZN(new_n887));
  XOR2_X1   g701(.A(new_n887), .B(KEYINPUT55), .Z(new_n888));
  INV_X1    g702(.A(KEYINPUT56), .ZN(new_n889));
  AOI22_X1  g703(.A1(new_n885), .A2(new_n888), .B1(new_n889), .B2(new_n883), .ZN(new_n890));
  AND4_X1   g704(.A1(KEYINPUT120), .A2(new_n883), .A3(new_n889), .A4(new_n888), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n350), .A2(G952), .ZN(new_n892));
  NOR3_X1   g706(.A1(new_n890), .A2(new_n891), .A3(new_n892), .ZN(G51));
  XOR2_X1   g707(.A(KEYINPUT121), .B(KEYINPUT57), .Z(new_n894));
  INV_X1    g708(.A(new_n894), .ZN(new_n895));
  OR2_X1    g709(.A1(new_n710), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n710), .A2(new_n895), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n824), .A2(new_n768), .ZN(new_n898));
  AOI21_X1  g712(.A(KEYINPUT54), .B1(new_n820), .B2(new_n823), .ZN(new_n899));
  OAI211_X1 g713(.A(new_n896), .B(new_n897), .C1(new_n898), .C2(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(new_n677), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  XOR2_X1   g716(.A(new_n739), .B(KEYINPUT122), .Z(new_n903));
  NAND4_X1  g717(.A1(new_n820), .A2(G902), .A3(new_n823), .A4(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n892), .B1(new_n902), .B2(new_n904), .ZN(G54));
  INV_X1    g719(.A(new_n892), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n820), .A2(KEYINPUT58), .A3(G902), .A4(new_n823), .ZN(new_n907));
  INV_X1    g721(.A(G475), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n906), .B1(new_n909), .B2(new_n522), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n909), .A2(new_n522), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT123), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n909), .A2(KEYINPUT123), .A3(new_n522), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n910), .B1(new_n913), .B2(new_n914), .ZN(G60));
  AND2_X1   g729(.A1(new_n583), .A2(new_n585), .ZN(new_n916));
  XOR2_X1   g730(.A(new_n588), .B(KEYINPUT59), .Z(new_n917));
  OAI21_X1  g731(.A(new_n916), .B1(new_n825), .B2(new_n917), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n916), .A2(new_n917), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n919), .B1(new_n898), .B2(new_n899), .ZN(new_n920));
  AND3_X1   g734(.A1(new_n918), .A2(new_n906), .A3(new_n920), .ZN(G63));
  NAND2_X1  g735(.A1(G217), .A2(G902), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(KEYINPUT60), .ZN(new_n923));
  OAI211_X1 g737(.A(new_n355), .B(new_n353), .C1(new_n824), .C2(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(new_n923), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n820), .A2(new_n613), .A3(new_n823), .A4(new_n925), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n924), .A2(new_n906), .A3(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT61), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND4_X1  g743(.A1(new_n924), .A2(KEYINPUT61), .A3(new_n906), .A4(new_n926), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n929), .A2(new_n930), .ZN(G66));
  INV_X1    g745(.A(KEYINPUT124), .ZN(new_n932));
  NOR3_X1   g746(.A1(new_n785), .A2(new_n786), .A3(new_n779), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n933), .A2(G953), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n531), .A2(G224), .ZN(new_n935));
  AOI211_X1 g749(.A(new_n932), .B(new_n934), .C1(G953), .C2(new_n935), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n936), .B1(new_n932), .B2(new_n934), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n424), .B1(G898), .B2(new_n350), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n937), .B(new_n938), .ZN(G69));
  NAND2_X1  g753(.A1(new_n266), .A2(new_n268), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n510), .A2(new_n513), .A3(new_n515), .ZN(new_n941));
  XOR2_X1   g755(.A(new_n941), .B(KEYINPUT125), .Z(new_n942));
  XNOR2_X1  g756(.A(new_n940), .B(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(new_n747), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n944), .B1(new_n757), .B2(new_n762), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n638), .A2(new_n749), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n946), .A2(new_n716), .A3(new_n776), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n947), .B(KEYINPUT126), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT62), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n949), .B1(new_n667), .B2(new_n795), .ZN(new_n950));
  OAI211_X1 g764(.A(KEYINPUT62), .B(new_n799), .C1(new_n650), .C2(new_n666), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  AND3_X1   g766(.A1(new_n945), .A2(new_n948), .A3(new_n952), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n943), .B1(new_n953), .B2(G953), .ZN(new_n954));
  INV_X1    g768(.A(new_n720), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n745), .A2(new_n716), .A3(new_n791), .ZN(new_n956));
  AND3_X1   g770(.A1(new_n956), .A2(new_n718), .A3(new_n799), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n945), .A2(new_n955), .A3(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n625), .B1(new_n958), .B2(new_n350), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n954), .B1(new_n943), .B2(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n350), .B1(G227), .B2(G900), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n960), .B(new_n961), .ZN(G72));
  NAND4_X1  g776(.A1(new_n945), .A2(new_n955), .A3(new_n933), .A4(new_n957), .ZN(new_n963));
  NAND2_X1  g777(.A1(G472), .A2(G902), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n964), .B(KEYINPUT63), .Z(new_n965));
  NAND2_X1  g779(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n966), .A2(new_n271), .A3(new_n241), .A4(new_n269), .ZN(new_n967));
  INV_X1    g781(.A(new_n965), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n968), .B1(new_n802), .B2(new_n812), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n270), .A2(new_n271), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n970), .A2(new_n288), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n892), .B1(new_n969), .B2(new_n971), .ZN(new_n972));
  NAND4_X1  g786(.A1(new_n945), .A2(new_n933), .A3(new_n948), .A4(new_n952), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n973), .A2(new_n965), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n974), .A2(new_n251), .A3(new_n270), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n967), .A2(new_n972), .A3(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT127), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n967), .A2(new_n975), .A3(KEYINPUT127), .A4(new_n972), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n978), .A2(new_n979), .ZN(G57));
endmodule


