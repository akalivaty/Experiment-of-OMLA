//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 1 0 1 0 0 0 1 0 0 0 1 0 1 0 0 0 0 0 0 0 0 0 1 1 0 0 0 1 0 1 0 0 0 0 0 0 1 1 1 1 0 1 1 1 0 0 1 0 0 0 0 0 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n745, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n831, new_n832, new_n834, new_n835,
    new_n837, new_n838, new_n839, new_n840, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n899, new_n900, new_n901, new_n902,
    new_n904, new_n905, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n919,
    new_n921, new_n922, new_n923, new_n924, new_n926, new_n927, new_n928,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n939, new_n940, new_n941, new_n942, new_n943, new_n945,
    new_n946, new_n947, new_n948, new_n950, new_n951, new_n952, new_n953;
  INV_X1    g000(.A(KEYINPUT87), .ZN(new_n202));
  INV_X1    g001(.A(G43gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n203), .A2(G50gat), .ZN(new_n204));
  INV_X1    g003(.A(G50gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n205), .A2(G43gat), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n202), .B1(new_n204), .B2(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n205), .A2(G43gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n203), .A2(G50gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n208), .A2(new_n209), .A3(KEYINPUT87), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n207), .A2(KEYINPUT15), .A3(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT15), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n212), .B1(new_n204), .B2(new_n206), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(G29gat), .ZN(new_n215));
  INV_X1    g014(.A(G36gat), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n215), .A2(new_n216), .A3(KEYINPUT14), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT14), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n218), .B1(G29gat), .B2(G36gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(G29gat), .A2(G36gat), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n217), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n214), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT17), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n211), .A2(new_n221), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n221), .B1(new_n211), .B2(new_n213), .ZN(new_n227));
  AND3_X1   g026(.A1(new_n208), .A2(new_n209), .A3(KEYINPUT87), .ZN(new_n228));
  AOI21_X1  g027(.A(KEYINPUT87), .B1(new_n208), .B2(new_n209), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n222), .B1(new_n230), .B2(KEYINPUT15), .ZN(new_n231));
  OAI21_X1  g030(.A(KEYINPUT17), .B1(new_n227), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(KEYINPUT98), .A2(KEYINPUT7), .ZN(new_n233));
  INV_X1    g032(.A(G85gat), .ZN(new_n234));
  INV_X1    g033(.A(G92gat), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n233), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  NAND4_X1  g035(.A1(KEYINPUT98), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n237));
  AND2_X1   g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(G99gat), .A2(G106gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(KEYINPUT8), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT99), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n234), .A2(new_n235), .ZN(new_n242));
  AND3_X1   g041(.A1(new_n240), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n241), .B1(new_n240), .B2(new_n242), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n238), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  XOR2_X1   g044(.A(G99gat), .B(G106gat), .Z(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n246), .ZN(new_n248));
  OAI211_X1 g047(.A(new_n238), .B(new_n248), .C1(new_n243), .C2(new_n244), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n226), .A2(new_n232), .A3(new_n250), .ZN(new_n251));
  NAND3_X1  g050(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n227), .A2(new_n231), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n253), .A2(new_n249), .A3(new_n247), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n251), .A2(new_n252), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(G190gat), .ZN(new_n256));
  INV_X1    g055(.A(G190gat), .ZN(new_n257));
  NAND4_X1  g056(.A1(new_n251), .A2(new_n257), .A3(new_n252), .A4(new_n254), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(G218gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT97), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n256), .A2(G218gat), .A3(new_n258), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n261), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT100), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND4_X1  g065(.A1(new_n261), .A2(new_n262), .A3(KEYINPUT100), .A4(new_n263), .ZN(new_n267));
  XOR2_X1   g066(.A(G134gat), .B(G162gat), .Z(new_n268));
  XNOR2_X1  g067(.A(new_n268), .B(KEYINPUT96), .ZN(new_n269));
  NAND2_X1  g068(.A1(G232gat), .A2(G233gat), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT41), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  XOR2_X1   g071(.A(new_n269), .B(new_n272), .Z(new_n273));
  AND3_X1   g072(.A1(new_n266), .A2(new_n267), .A3(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(new_n273), .ZN(new_n275));
  AND2_X1   g074(.A1(new_n261), .A2(new_n263), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n266), .A2(new_n276), .A3(new_n267), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n274), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(G120gat), .B(G148gat), .ZN(new_n279));
  INV_X1    g078(.A(G176gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n279), .B(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(G204gat), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n281), .B(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  XNOR2_X1  g083(.A(G71gat), .B(G78gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(G71gat), .A2(G78gat), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT9), .ZN(new_n287));
  AND3_X1   g086(.A1(new_n286), .A2(KEYINPUT91), .A3(new_n287), .ZN(new_n288));
  AOI21_X1  g087(.A(KEYINPUT91), .B1(new_n286), .B2(new_n287), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  XNOR2_X1  g089(.A(G57gat), .B(G64gat), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n285), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT93), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n294), .B1(new_n288), .B2(new_n289), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n286), .A2(new_n287), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT91), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n286), .A2(KEYINPUT91), .A3(new_n287), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n298), .A2(KEYINPUT93), .A3(new_n299), .ZN(new_n300));
  AND2_X1   g099(.A1(new_n295), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n291), .A2(KEYINPUT92), .ZN(new_n302));
  INV_X1    g101(.A(G64gat), .ZN(new_n303));
  OR3_X1    g102(.A1(new_n303), .A2(KEYINPUT92), .A3(G57gat), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n302), .A2(new_n285), .A3(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n293), .B1(new_n301), .B2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT101), .ZN(new_n308));
  NAND4_X1  g107(.A1(new_n307), .A2(new_n308), .A3(new_n249), .A4(new_n247), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT10), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n295), .A2(new_n300), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n298), .A2(new_n299), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n312), .A2(new_n291), .ZN(new_n313));
  OAI22_X1  g112(.A1(new_n311), .A2(new_n305), .B1(new_n313), .B2(new_n285), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n236), .A2(new_n237), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT8), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n316), .B1(G99gat), .B2(G106gat), .ZN(new_n317));
  NOR2_X1   g116(.A1(G85gat), .A2(G92gat), .ZN(new_n318));
  OAI21_X1  g117(.A(KEYINPUT99), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n240), .A2(new_n241), .A3(new_n242), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n315), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n308), .B1(new_n321), .B2(new_n248), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n250), .B1(new_n314), .B2(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n309), .A2(new_n310), .A3(new_n323), .ZN(new_n324));
  NAND4_X1  g123(.A1(new_n307), .A2(KEYINPUT10), .A3(new_n249), .A4(new_n247), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(G230gat), .A2(G233gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n309), .A2(new_n323), .ZN(new_n329));
  INV_X1    g128(.A(new_n327), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n284), .B1(new_n328), .B2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT102), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n328), .A2(new_n333), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n330), .B1(new_n324), .B2(new_n325), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(KEYINPUT102), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n283), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT103), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n338), .B1(new_n329), .B2(new_n330), .ZN(new_n339));
  AOI211_X1 g138(.A(KEYINPUT103), .B(new_n327), .C1(new_n309), .C2(new_n323), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n337), .A2(KEYINPUT104), .A3(new_n341), .ZN(new_n342));
  AOI21_X1  g141(.A(KEYINPUT102), .B1(new_n326), .B2(new_n327), .ZN(new_n343));
  AOI211_X1 g142(.A(new_n333), .B(new_n330), .C1(new_n324), .C2(new_n325), .ZN(new_n344));
  OAI211_X1 g143(.A(new_n284), .B(new_n341), .C1(new_n343), .C2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT104), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n332), .B1(new_n342), .B2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  XNOR2_X1  g148(.A(G15gat), .B(G22gat), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT16), .ZN(new_n351));
  OR2_X1    g150(.A1(new_n351), .A2(G1gat), .ZN(new_n352));
  AND2_X1   g151(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n350), .A2(G1gat), .ZN(new_n354));
  OAI21_X1  g153(.A(G8gat), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n350), .A2(new_n352), .ZN(new_n356));
  INV_X1    g155(.A(G8gat), .ZN(new_n357));
  OAI211_X1 g156(.A(new_n356), .B(new_n357), .C1(G1gat), .C2(new_n350), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n355), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n226), .A2(new_n232), .A3(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(G229gat), .A2(G233gat), .ZN(new_n362));
  AOI21_X1  g161(.A(KEYINPUT88), .B1(new_n253), .B2(new_n359), .ZN(new_n363));
  AND4_X1   g162(.A1(KEYINPUT88), .A2(new_n223), .A3(new_n359), .A4(new_n225), .ZN(new_n364));
  OAI211_X1 g163(.A(new_n361), .B(new_n362), .C1(new_n363), .C2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(KEYINPUT89), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT18), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT88), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n223), .A2(new_n225), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n368), .B1(new_n369), .B2(new_n360), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n253), .A2(KEYINPUT88), .A3(new_n359), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT89), .ZN(new_n373));
  NAND4_X1  g172(.A1(new_n372), .A2(new_n373), .A3(new_n362), .A4(new_n361), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n366), .A2(new_n367), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(KEYINPUT90), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n369), .A2(new_n360), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n372), .A2(new_n377), .ZN(new_n378));
  XNOR2_X1  g177(.A(new_n362), .B(KEYINPUT13), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  NAND4_X1  g180(.A1(new_n372), .A2(KEYINPUT18), .A3(new_n362), .A4(new_n361), .ZN(new_n382));
  XNOR2_X1  g181(.A(G113gat), .B(G141gat), .ZN(new_n383));
  XNOR2_X1  g182(.A(G169gat), .B(G197gat), .ZN(new_n384));
  XNOR2_X1  g183(.A(new_n383), .B(new_n384), .ZN(new_n385));
  XNOR2_X1  g184(.A(KEYINPUT86), .B(KEYINPUT11), .ZN(new_n386));
  XNOR2_X1  g185(.A(new_n385), .B(new_n386), .ZN(new_n387));
  XNOR2_X1  g186(.A(new_n387), .B(KEYINPUT12), .ZN(new_n388));
  AND3_X1   g187(.A1(new_n381), .A2(new_n382), .A3(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT90), .ZN(new_n390));
  NAND4_X1  g189(.A1(new_n366), .A2(new_n374), .A3(new_n390), .A4(new_n367), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n376), .A2(new_n389), .A3(new_n391), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n375), .A2(new_n381), .A3(new_n382), .ZN(new_n393));
  INV_X1    g192(.A(new_n388), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n392), .A2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n349), .A2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT21), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n360), .B1(new_n314), .B2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(G183gat), .ZN(new_n401));
  XNOR2_X1  g200(.A(new_n400), .B(new_n401), .ZN(new_n402));
  AND2_X1   g201(.A1(G231gat), .A2(G233gat), .ZN(new_n403));
  OR2_X1    g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n402), .A2(new_n403), .ZN(new_n405));
  XNOR2_X1  g204(.A(KEYINPUT94), .B(KEYINPUT95), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  AND3_X1   g206(.A1(new_n404), .A2(new_n405), .A3(new_n407), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n407), .B1(new_n404), .B2(new_n405), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n314), .A2(new_n399), .ZN(new_n410));
  XNOR2_X1  g209(.A(G127gat), .B(G155gat), .ZN(new_n411));
  INV_X1    g210(.A(G211gat), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n411), .B(new_n412), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n410), .B(new_n413), .ZN(new_n414));
  XOR2_X1   g213(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n415));
  XNOR2_X1  g214(.A(new_n414), .B(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  OR3_X1    g216(.A1(new_n408), .A2(new_n409), .A3(new_n417), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n417), .B1(new_n408), .B2(new_n409), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n278), .A2(new_n398), .A3(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT77), .ZN(new_n422));
  NAND2_X1  g221(.A1(G225gat), .A2(G233gat), .ZN(new_n423));
  INV_X1    g222(.A(G134gat), .ZN(new_n424));
  AOI21_X1  g223(.A(KEYINPUT1), .B1(new_n424), .B2(G127gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(KEYINPUT68), .B(G120gat), .ZN(new_n426));
  INV_X1    g225(.A(G113gat), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  AND2_X1   g227(.A1(new_n427), .A2(G120gat), .ZN(new_n429));
  OAI221_X1 g228(.A(new_n425), .B1(G127gat), .B2(new_n424), .C1(new_n428), .C2(new_n429), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n424), .A2(G127gat), .ZN(new_n431));
  XNOR2_X1  g230(.A(new_n431), .B(KEYINPUT67), .ZN(new_n432));
  XNOR2_X1  g231(.A(KEYINPUT66), .B(G134gat), .ZN(new_n433));
  INV_X1    g232(.A(G127gat), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  XNOR2_X1  g234(.A(G113gat), .B(G120gat), .ZN(new_n436));
  OAI22_X1  g235(.A1(new_n432), .A2(new_n435), .B1(KEYINPUT1), .B2(new_n436), .ZN(new_n437));
  AND2_X1   g236(.A1(new_n430), .A2(new_n437), .ZN(new_n438));
  XNOR2_X1  g237(.A(G141gat), .B(G148gat), .ZN(new_n439));
  OR2_X1    g238(.A1(G155gat), .A2(G162gat), .ZN(new_n440));
  OR2_X1    g239(.A1(new_n440), .A2(KEYINPUT2), .ZN(new_n441));
  NAND2_X1  g240(.A1(G155gat), .A2(G162gat), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n439), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  OAI211_X1 g242(.A(new_n442), .B(new_n440), .C1(new_n439), .C2(KEYINPUT2), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT74), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  AND2_X1   g245(.A1(new_n440), .A2(new_n442), .ZN(new_n447));
  OAI211_X1 g246(.A(new_n447), .B(KEYINPUT74), .C1(KEYINPUT2), .C2(new_n439), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n443), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n438), .A2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n449), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n430), .A2(new_n437), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n423), .B1(new_n450), .B2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT5), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n422), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n451), .A2(KEYINPUT75), .A3(KEYINPUT3), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT3), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n449), .A2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT75), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n460), .B1(new_n449), .B2(new_n458), .ZN(new_n461));
  NAND4_X1  g260(.A1(new_n457), .A2(new_n452), .A3(new_n459), .A4(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(new_n423), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT4), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n463), .B1(new_n450), .B2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT76), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n449), .A2(new_n466), .ZN(new_n467));
  AOI211_X1 g266(.A(KEYINPUT76), .B(new_n443), .C1(new_n446), .C2(new_n448), .ZN(new_n468));
  OAI211_X1 g267(.A(KEYINPUT4), .B(new_n438), .C1(new_n467), .C2(new_n468), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n462), .A2(new_n465), .A3(new_n469), .ZN(new_n470));
  XNOR2_X1  g269(.A(new_n452), .B(new_n449), .ZN(new_n471));
  OAI211_X1 g270(.A(KEYINPUT77), .B(KEYINPUT5), .C1(new_n471), .C2(new_n423), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n456), .A2(new_n470), .A3(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n438), .B1(new_n467), .B2(new_n468), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(new_n464), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n438), .A2(KEYINPUT4), .A3(new_n449), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n476), .A2(new_n462), .A3(new_n455), .A4(new_n477), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n478), .A2(new_n463), .ZN(new_n479));
  OAI21_X1  g278(.A(KEYINPUT82), .B1(new_n474), .B2(new_n479), .ZN(new_n480));
  OR2_X1    g279(.A1(new_n478), .A2(new_n463), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT82), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n481), .A2(new_n482), .A3(new_n473), .ZN(new_n483));
  XNOR2_X1  g282(.A(KEYINPUT0), .B(G57gat), .ZN(new_n484));
  XNOR2_X1  g283(.A(new_n484), .B(G85gat), .ZN(new_n485));
  XNOR2_X1  g284(.A(G1gat), .B(G29gat), .ZN(new_n486));
  XOR2_X1   g285(.A(new_n485), .B(new_n486), .Z(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n480), .A2(new_n483), .A3(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT84), .ZN(new_n490));
  OAI211_X1 g289(.A(new_n473), .B(new_n487), .C1(new_n463), .C2(new_n478), .ZN(new_n491));
  XOR2_X1   g290(.A(KEYINPUT78), .B(KEYINPUT6), .Z(new_n492));
  INV_X1    g291(.A(new_n492), .ZN(new_n493));
  AND2_X1   g292(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  AND3_X1   g293(.A1(new_n489), .A2(new_n490), .A3(new_n494), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n490), .B1(new_n489), .B2(new_n494), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n487), .B1(new_n481), .B2(new_n473), .ZN(new_n497));
  INV_X1    g296(.A(new_n497), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n498), .A2(new_n493), .ZN(new_n499));
  NOR3_X1   g298(.A1(new_n495), .A2(new_n496), .A3(new_n499), .ZN(new_n500));
  XNOR2_X1  g299(.A(KEYINPUT27), .B(G183gat), .ZN(new_n501));
  XNOR2_X1  g300(.A(new_n501), .B(KEYINPUT65), .ZN(new_n502));
  OAI21_X1  g301(.A(KEYINPUT28), .B1(new_n502), .B2(G190gat), .ZN(new_n503));
  INV_X1    g302(.A(new_n501), .ZN(new_n504));
  AOI21_X1  g303(.A(G190gat), .B1(new_n504), .B2(KEYINPUT64), .ZN(new_n505));
  AOI21_X1  g304(.A(KEYINPUT64), .B1(new_n401), .B2(KEYINPUT27), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n506), .A2(KEYINPUT28), .ZN(new_n507));
  NAND2_X1  g306(.A1(G169gat), .A2(G176gat), .ZN(new_n508));
  NOR2_X1   g307(.A1(G169gat), .A2(G176gat), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n509), .A2(KEYINPUT26), .ZN(new_n510));
  AOI22_X1  g309(.A1(new_n505), .A2(new_n507), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n509), .A2(KEYINPUT26), .ZN(new_n512));
  NAND2_X1  g311(.A1(G183gat), .A2(G190gat), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n503), .A2(new_n511), .A3(new_n512), .A4(new_n513), .ZN(new_n514));
  AND2_X1   g313(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(new_n257), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n509), .A2(KEYINPUT23), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT23), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n518), .B1(G169gat), .B2(G176gat), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n516), .A2(new_n517), .A3(new_n519), .A4(new_n508), .ZN(new_n520));
  NOR2_X1   g319(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n521));
  NOR3_X1   g320(.A1(new_n515), .A2(new_n521), .A3(new_n257), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n523), .B(KEYINPUT25), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n514), .A2(new_n524), .ZN(new_n525));
  AND2_X1   g324(.A1(G226gat), .A2(G233gat), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT29), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n526), .B1(new_n525), .B2(new_n529), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(G197gat), .B(G204gat), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT22), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n533), .B1(new_n412), .B2(new_n260), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  XOR2_X1   g335(.A(G211gat), .B(G218gat), .Z(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(KEYINPUT71), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n536), .B(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n531), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n528), .A2(KEYINPUT72), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT72), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n543), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n530), .B1(new_n542), .B2(new_n544), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n541), .B1(new_n545), .B2(new_n540), .ZN(new_n546));
  XOR2_X1   g345(.A(G8gat), .B(G36gat), .Z(new_n547));
  XNOR2_X1  g346(.A(new_n547), .B(G64gat), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(new_n235), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n546), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT37), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n550), .B1(new_n546), .B2(new_n552), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n553), .B1(new_n552), .B2(new_n546), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(KEYINPUT38), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n552), .B1(new_n545), .B2(new_n540), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n556), .B1(new_n540), .B2(new_n531), .ZN(new_n557));
  OR2_X1    g356(.A1(new_n557), .A2(KEYINPUT85), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT38), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n557), .A2(KEYINPUT85), .ZN(new_n560));
  NAND4_X1  g359(.A1(new_n558), .A2(new_n559), .A3(new_n553), .A4(new_n560), .ZN(new_n561));
  NAND4_X1  g360(.A1(new_n500), .A2(new_n551), .A3(new_n555), .A4(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(G22gat), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n467), .A2(new_n468), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n536), .A2(new_n537), .ZN(new_n565));
  INV_X1    g364(.A(new_n537), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n529), .B1(new_n566), .B2(new_n535), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n458), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  AOI22_X1  g367(.A1(new_n564), .A2(new_n568), .B1(G228gat), .B2(G233gat), .ZN(new_n569));
  AOI21_X1  g368(.A(KEYINPUT29), .B1(new_n449), .B2(new_n458), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n569), .B1(new_n539), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n539), .A2(new_n529), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n449), .B1(new_n572), .B2(new_n458), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n539), .B1(new_n459), .B2(new_n529), .ZN(new_n574));
  OAI211_X1 g373(.A(G228gat), .B(G233gat), .C1(new_n573), .C2(new_n574), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n563), .B1(new_n571), .B2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n571), .A2(new_n563), .A3(new_n575), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n577), .A2(KEYINPUT79), .A3(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(G78gat), .B(G106gat), .ZN(new_n580));
  XNOR2_X1  g379(.A(KEYINPUT31), .B(G50gat), .ZN(new_n581));
  XOR2_X1   g380(.A(new_n580), .B(new_n581), .Z(new_n582));
  OR2_X1    g381(.A1(new_n579), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT79), .ZN(new_n584));
  INV_X1    g383(.A(new_n578), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n584), .B1(new_n585), .B2(new_n576), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n586), .A2(new_n579), .A3(new_n582), .ZN(new_n587));
  AND2_X1   g386(.A1(new_n583), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT30), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n551), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n590), .A2(KEYINPUT73), .ZN(new_n591));
  INV_X1    g390(.A(new_n551), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n592), .A2(KEYINPUT30), .ZN(new_n593));
  INV_X1    g392(.A(new_n546), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n594), .A2(new_n549), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT73), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n551), .A2(new_n596), .A3(new_n589), .ZN(new_n597));
  NAND4_X1  g396(.A1(new_n591), .A2(new_n593), .A3(new_n595), .A4(new_n597), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n476), .A2(new_n462), .A3(new_n477), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(new_n463), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n487), .B1(new_n600), .B2(KEYINPUT39), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT39), .ZN(new_n602));
  AND2_X1   g401(.A1(new_n471), .A2(new_n423), .ZN(new_n603));
  AOI211_X1 g402(.A(new_n602), .B(new_n603), .C1(new_n599), .C2(new_n463), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT40), .ZN(new_n605));
  NOR3_X1   g404(.A1(new_n601), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(KEYINPUT83), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n605), .B1(new_n601), .B2(new_n604), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(KEYINPUT81), .ZN(new_n609));
  NAND4_X1  g408(.A1(new_n598), .A2(new_n607), .A3(new_n489), .A4(new_n609), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n562), .A2(new_n588), .A3(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n598), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n499), .B1(new_n498), .B2(new_n494), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  AND2_X1   g414(.A1(new_n588), .A2(KEYINPUT80), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n588), .A2(KEYINPUT80), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n615), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT36), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n525), .B(new_n452), .ZN(new_n620));
  NAND2_X1  g419(.A1(G227gat), .A2(G233gat), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT34), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n624), .B1(new_n621), .B2(KEYINPUT70), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n620), .A2(new_n622), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n627), .A2(KEYINPUT32), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT69), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(G15gat), .B(G43gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n631), .B(G71gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(G99gat), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT33), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n633), .B1(new_n627), .B2(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n627), .A2(KEYINPUT69), .A3(KEYINPUT32), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n630), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  OAI211_X1 g436(.A(new_n627), .B(KEYINPUT32), .C1(new_n634), .C2(new_n633), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n626), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n637), .A2(new_n638), .A3(new_n626), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n623), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n641), .ZN(new_n643));
  INV_X1    g442(.A(new_n623), .ZN(new_n644));
  NOR3_X1   g443(.A1(new_n643), .A2(new_n639), .A3(new_n644), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n619), .B1(new_n642), .B2(new_n645), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n644), .B1(new_n643), .B2(new_n639), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n640), .A2(new_n623), .A3(new_n641), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n647), .A2(new_n648), .A3(KEYINPUT36), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n611), .A2(new_n618), .A3(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n647), .A2(new_n648), .A3(new_n588), .ZN(new_n652));
  OAI21_X1  g451(.A(KEYINPUT35), .B1(new_n615), .B2(new_n652), .ZN(new_n653));
  OR3_X1    g452(.A1(new_n500), .A2(KEYINPUT35), .A3(new_n598), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n653), .B1(new_n654), .B2(new_n652), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n421), .B1(new_n651), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n656), .A2(new_n613), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g457(.A1(new_n656), .A2(new_n598), .ZN(new_n659));
  NAND2_X1  g458(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n351), .A2(new_n357), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n659), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT42), .ZN(new_n663));
  OR2_X1    g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n662), .A2(new_n663), .ZN(new_n665));
  OAI211_X1 g464(.A(new_n664), .B(new_n665), .C1(new_n357), .C2(new_n659), .ZN(G1325gat));
  NOR2_X1   g465(.A1(new_n642), .A2(new_n645), .ZN(new_n667));
  AOI21_X1  g466(.A(G15gat), .B1(new_n656), .B2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n650), .ZN(new_n669));
  AND2_X1   g468(.A1(new_n656), .A2(G15gat), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n668), .B1(new_n669), .B2(new_n670), .ZN(G1326gat));
  NOR2_X1   g470(.A1(new_n616), .A2(new_n617), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n656), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g473(.A(KEYINPUT43), .B(G22gat), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n674), .B(new_n675), .ZN(G1327gat));
  AOI21_X1  g475(.A(new_n278), .B1(new_n651), .B2(new_n655), .ZN(new_n677));
  NOR3_X1   g476(.A1(new_n420), .A2(new_n349), .A3(new_n397), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n680), .A2(new_n215), .A3(new_n613), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n681), .B(KEYINPUT45), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n651), .A2(new_n655), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n277), .A2(new_n275), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n266), .A2(new_n267), .A3(new_n273), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  AOI21_X1  g485(.A(KEYINPUT44), .B1(new_n683), .B2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT44), .ZN(new_n688));
  AOI211_X1 g487(.A(new_n688), .B(new_n278), .C1(new_n651), .C2(new_n655), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  AND3_X1   g489(.A1(new_n690), .A2(new_n613), .A3(new_n678), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n682), .B1(new_n215), .B2(new_n691), .ZN(G1328gat));
  INV_X1    g491(.A(new_n687), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n677), .A2(KEYINPUT44), .ZN(new_n694));
  NAND4_X1  g493(.A1(new_n693), .A2(new_n598), .A3(new_n678), .A4(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT106), .ZN(new_n696));
  OR2_X1    g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n695), .A2(new_n696), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n697), .A2(G36gat), .A3(new_n698), .ZN(new_n699));
  NOR3_X1   g498(.A1(new_n679), .A2(G36gat), .A3(new_n612), .ZN(new_n700));
  XNOR2_X1  g499(.A(KEYINPUT105), .B(KEYINPUT46), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n700), .B(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n699), .A2(new_n702), .ZN(G1329gat));
  NAND4_X1  g502(.A1(new_n690), .A2(G43gat), .A3(new_n669), .A4(new_n678), .ZN(new_n704));
  INV_X1    g503(.A(new_n667), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n203), .B1(new_n679), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n707), .B(KEYINPUT47), .ZN(G1330gat));
  NOR2_X1   g507(.A1(new_n672), .A2(G50gat), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n680), .A2(KEYINPUT107), .A3(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(new_n588), .ZN(new_n711));
  AND3_X1   g510(.A1(new_n690), .A2(new_n711), .A3(new_n678), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n710), .B1(new_n712), .B2(new_n205), .ZN(new_n713));
  AOI22_X1  g512(.A1(new_n680), .A2(new_n709), .B1(KEYINPUT107), .B2(KEYINPUT48), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n690), .A2(new_n673), .A3(new_n678), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT48), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n715), .A2(new_n716), .A3(G50gat), .ZN(new_n717));
  AOI22_X1  g516(.A1(new_n713), .A2(KEYINPUT48), .B1(new_n714), .B2(new_n717), .ZN(G1331gat));
  NAND4_X1  g517(.A1(new_n684), .A2(new_n420), .A3(new_n685), .A4(new_n397), .ZN(new_n719));
  INV_X1    g518(.A(new_n719), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n683), .A2(new_n349), .A3(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT108), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n721), .B(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(new_n613), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n724), .B(G57gat), .ZN(G1332gat));
  OR2_X1    g524(.A1(new_n721), .A2(KEYINPUT108), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n721), .A2(KEYINPUT108), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n728), .A2(new_n612), .ZN(new_n729));
  NOR2_X1   g528(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n730));
  AND2_X1   g529(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n729), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n732), .B1(new_n729), .B2(new_n730), .ZN(G1333gat));
  XNOR2_X1  g532(.A(KEYINPUT109), .B(KEYINPUT50), .ZN(new_n734));
  INV_X1    g533(.A(new_n734), .ZN(new_n735));
  AOI21_X1  g534(.A(G71gat), .B1(new_n723), .B2(new_n667), .ZN(new_n736));
  INV_X1    g535(.A(G71gat), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n650), .A2(new_n737), .ZN(new_n738));
  AND3_X1   g537(.A1(new_n726), .A2(new_n727), .A3(new_n738), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n735), .B1(new_n736), .B2(new_n739), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n737), .B1(new_n728), .B2(new_n705), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n723), .A2(new_n738), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n741), .A2(new_n734), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n740), .A2(new_n743), .ZN(G1334gat));
  NAND2_X1  g543(.A1(new_n723), .A2(new_n673), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g545(.A1(new_n420), .A2(new_n396), .ZN(new_n747));
  NAND4_X1  g546(.A1(new_n693), .A2(new_n349), .A3(new_n694), .A4(new_n747), .ZN(new_n748));
  NOR3_X1   g547(.A1(new_n748), .A2(new_n234), .A3(new_n614), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n683), .A2(new_n686), .A3(new_n747), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT51), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n677), .A2(KEYINPUT51), .A3(new_n747), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n754), .A2(new_n613), .A3(new_n349), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n749), .B1(new_n234), .B2(new_n755), .ZN(G1336gat));
  NAND4_X1  g555(.A1(new_n690), .A2(new_n598), .A3(new_n349), .A4(new_n747), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(G92gat), .ZN(new_n758));
  NOR3_X1   g557(.A1(new_n612), .A2(G92gat), .A3(new_n348), .ZN(new_n759));
  AOI21_X1  g558(.A(KEYINPUT52), .B1(new_n754), .B2(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT110), .ZN(new_n762));
  AOI22_X1  g561(.A1(new_n752), .A2(new_n753), .B1(new_n762), .B2(new_n759), .ZN(new_n763));
  OR2_X1    g562(.A1(new_n759), .A2(new_n762), .ZN(new_n764));
  AOI22_X1  g563(.A1(new_n757), .A2(G92gat), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT52), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n761), .B1(new_n765), .B2(new_n766), .ZN(G1337gat));
  INV_X1    g566(.A(G99gat), .ZN(new_n768));
  NOR3_X1   g567(.A1(new_n748), .A2(new_n768), .A3(new_n650), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n754), .A2(new_n667), .A3(new_n349), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n769), .B1(new_n768), .B2(new_n770), .ZN(G1338gat));
  OAI21_X1  g570(.A(G106gat), .B1(new_n748), .B2(new_n588), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT53), .ZN(new_n773));
  INV_X1    g572(.A(G106gat), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n754), .A2(new_n774), .A3(new_n711), .A4(new_n349), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n772), .A2(new_n773), .A3(new_n775), .ZN(new_n776));
  AOI211_X1 g575(.A(G106gat), .B(new_n348), .C1(new_n752), .C2(new_n753), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n690), .A2(new_n673), .A3(new_n349), .A4(new_n747), .ZN(new_n778));
  AOI22_X1  g577(.A1(new_n777), .A2(new_n711), .B1(new_n778), .B2(G106gat), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n776), .B1(new_n779), .B2(new_n773), .ZN(G1339gat));
  INV_X1    g579(.A(KEYINPUT55), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n324), .A2(new_n330), .A3(new_n325), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(KEYINPUT54), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n783), .B1(new_n334), .B2(new_n336), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n283), .B1(new_n328), .B2(KEYINPUT54), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n781), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT111), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n342), .A2(new_n347), .ZN(new_n789));
  INV_X1    g588(.A(new_n785), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n343), .A2(new_n344), .ZN(new_n791));
  OAI211_X1 g590(.A(KEYINPUT55), .B(new_n790), .C1(new_n791), .C2(new_n783), .ZN(new_n792));
  OAI211_X1 g591(.A(KEYINPUT111), .B(new_n781), .C1(new_n784), .C2(new_n785), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n788), .A2(new_n789), .A3(new_n792), .A4(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n372), .A2(new_n361), .ZN(new_n795));
  INV_X1    g594(.A(new_n362), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n372), .A2(new_n377), .A3(new_n379), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  AOI21_X1  g598(.A(KEYINPUT112), .B1(new_n799), .B2(new_n387), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT112), .ZN(new_n801));
  INV_X1    g600(.A(new_n387), .ZN(new_n802));
  AOI211_X1 g601(.A(new_n801), .B(new_n802), .C1(new_n797), .C2(new_n798), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n800), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(new_n392), .ZN(new_n805));
  OAI22_X1  g604(.A1(new_n794), .A2(new_n397), .B1(new_n348), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(new_n278), .ZN(new_n807));
  INV_X1    g606(.A(new_n794), .ZN(new_n808));
  INV_X1    g607(.A(new_n805), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n808), .A2(new_n686), .A3(new_n809), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n420), .B1(new_n807), .B2(new_n810), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n719), .A2(new_n349), .ZN(new_n812));
  OAI211_X1 g611(.A(new_n667), .B(new_n672), .C1(new_n811), .C2(new_n812), .ZN(new_n813));
  AND2_X1   g612(.A1(new_n593), .A2(new_n595), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n814), .A2(new_n613), .A3(new_n591), .A4(new_n597), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  OAI21_X1  g616(.A(G113gat), .B1(new_n817), .B2(new_n397), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n807), .A2(new_n810), .ZN(new_n819));
  INV_X1    g618(.A(new_n420), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(new_n812), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n652), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  AND2_X1   g622(.A1(new_n823), .A2(new_n613), .ZN(new_n824));
  OR2_X1    g623(.A1(new_n824), .A2(KEYINPUT113), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(KEYINPUT113), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n825), .A2(new_n612), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n396), .A2(new_n427), .ZN(new_n828));
  XOR2_X1   g627(.A(new_n828), .B(KEYINPUT114), .Z(new_n829));
  OAI21_X1  g628(.A(new_n818), .B1(new_n827), .B2(new_n829), .ZN(G1340gat));
  OAI21_X1  g629(.A(G120gat), .B1(new_n817), .B2(new_n348), .ZN(new_n831));
  OR2_X1    g630(.A1(new_n348), .A2(new_n426), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n831), .B1(new_n827), .B2(new_n832), .ZN(G1341gat));
  NOR3_X1   g632(.A1(new_n817), .A2(new_n434), .A3(new_n820), .ZN(new_n834));
  OR2_X1    g633(.A1(new_n827), .A2(new_n820), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n834), .B1(new_n835), .B2(new_n434), .ZN(G1342gat));
  OR2_X1    g635(.A1(new_n278), .A2(new_n433), .ZN(new_n837));
  OR3_X1    g636(.A1(new_n827), .A2(KEYINPUT56), .A3(new_n837), .ZN(new_n838));
  OAI21_X1  g637(.A(G134gat), .B1(new_n817), .B2(new_n278), .ZN(new_n839));
  OAI21_X1  g638(.A(KEYINPUT56), .B1(new_n827), .B2(new_n837), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n838), .A2(new_n839), .A3(new_n840), .ZN(G1343gat));
  AOI21_X1  g640(.A(new_n588), .B1(new_n821), .B2(new_n822), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n669), .A2(new_n815), .ZN(new_n843));
  AND2_X1   g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(G141gat), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n844), .A2(new_n845), .A3(new_n396), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT58), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n396), .A2(new_n786), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n345), .A2(new_n346), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n345), .A2(new_n346), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n792), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  OAI22_X1  g650(.A1(new_n848), .A2(new_n851), .B1(new_n348), .B2(new_n805), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n278), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n810), .A2(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n812), .B1(new_n854), .B2(new_n820), .ZN(new_n855));
  OAI21_X1  g654(.A(KEYINPUT57), .B1(new_n855), .B2(new_n672), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT57), .ZN(new_n857));
  OAI211_X1 g656(.A(new_n857), .B(new_n711), .C1(new_n811), .C2(new_n812), .ZN(new_n858));
  NAND4_X1  g657(.A1(new_n856), .A2(new_n843), .A3(new_n858), .A4(new_n396), .ZN(new_n859));
  AND2_X1   g658(.A1(new_n859), .A2(KEYINPUT117), .ZN(new_n860));
  OAI21_X1  g659(.A(G141gat), .B1(new_n859), .B2(KEYINPUT117), .ZN(new_n861));
  OAI211_X1 g660(.A(new_n846), .B(new_n847), .C1(new_n860), .C2(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT115), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n846), .A2(new_n863), .ZN(new_n864));
  NAND4_X1  g663(.A1(new_n844), .A2(KEYINPUT115), .A3(new_n845), .A4(new_n396), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n859), .A2(G141gat), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  AND3_X1   g666(.A1(new_n867), .A2(KEYINPUT116), .A3(KEYINPUT58), .ZN(new_n868));
  AOI21_X1  g667(.A(KEYINPUT116), .B1(new_n867), .B2(KEYINPUT58), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n862), .B1(new_n868), .B2(new_n869), .ZN(G1344gat));
  INV_X1    g669(.A(KEYINPUT120), .ZN(new_n871));
  INV_X1    g670(.A(G148gat), .ZN(new_n872));
  AND3_X1   g671(.A1(new_n856), .A2(new_n843), .A3(new_n858), .ZN(new_n873));
  AOI211_X1 g672(.A(KEYINPUT59), .B(new_n872), .C1(new_n873), .C2(new_n349), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n857), .B1(new_n855), .B2(new_n672), .ZN(new_n875));
  OAI211_X1 g674(.A(KEYINPUT57), .B(new_n711), .C1(new_n811), .C2(new_n812), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(new_n815), .ZN(new_n878));
  AOI21_X1  g677(.A(KEYINPUT118), .B1(new_n650), .B2(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT118), .ZN(new_n880));
  AOI211_X1 g679(.A(new_n880), .B(new_n815), .C1(new_n646), .C2(new_n649), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n877), .A2(new_n349), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(KEYINPUT119), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT119), .ZN(new_n885));
  NAND4_X1  g684(.A1(new_n877), .A2(new_n885), .A3(new_n882), .A4(new_n349), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n884), .A2(G148gat), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n874), .B1(new_n887), .B2(KEYINPUT59), .ZN(new_n888));
  INV_X1    g687(.A(new_n844), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n349), .A2(new_n872), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n871), .B1(new_n888), .B2(new_n891), .ZN(new_n892));
  INV_X1    g691(.A(new_n891), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT59), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n872), .B1(new_n883), .B2(KEYINPUT119), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n894), .B1(new_n895), .B2(new_n886), .ZN(new_n896));
  OAI211_X1 g695(.A(KEYINPUT120), .B(new_n893), .C1(new_n896), .C2(new_n874), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n892), .A2(new_n897), .ZN(G1345gat));
  NAND2_X1  g697(.A1(new_n844), .A2(new_n420), .ZN(new_n899));
  XNOR2_X1  g698(.A(new_n899), .B(KEYINPUT121), .ZN(new_n900));
  INV_X1    g699(.A(G155gat), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n820), .A2(new_n901), .ZN(new_n902));
  AOI22_X1  g701(.A1(new_n900), .A2(new_n901), .B1(new_n873), .B2(new_n902), .ZN(G1346gat));
  AOI21_X1  g702(.A(G162gat), .B1(new_n844), .B2(new_n686), .ZN(new_n904));
  AND2_X1   g703(.A1(new_n873), .A2(new_n686), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n904), .B1(new_n905), .B2(G162gat), .ZN(G1347gat));
  NOR2_X1   g705(.A1(new_n612), .A2(new_n613), .ZN(new_n907));
  INV_X1    g706(.A(new_n907), .ZN(new_n908));
  OR2_X1    g707(.A1(new_n813), .A2(new_n908), .ZN(new_n909));
  OAI21_X1  g708(.A(G169gat), .B1(new_n909), .B2(new_n397), .ZN(new_n910));
  XNOR2_X1  g709(.A(new_n910), .B(KEYINPUT123), .ZN(new_n911));
  AND2_X1   g710(.A1(new_n823), .A2(new_n907), .ZN(new_n912));
  INV_X1    g711(.A(G169gat), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n912), .A2(new_n913), .A3(new_n396), .ZN(new_n914));
  XNOR2_X1  g713(.A(new_n914), .B(KEYINPUT122), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n911), .A2(new_n915), .ZN(G1348gat));
  OAI21_X1  g715(.A(G176gat), .B1(new_n909), .B2(new_n348), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n912), .A2(new_n280), .A3(new_n349), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  XNOR2_X1  g718(.A(new_n919), .B(KEYINPUT124), .ZN(G1349gat));
  OAI21_X1  g719(.A(G183gat), .B1(new_n909), .B2(new_n820), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n820), .A2(new_n502), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n912), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  XNOR2_X1  g723(.A(new_n924), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g724(.A(G190gat), .B1(new_n909), .B2(new_n278), .ZN(new_n926));
  XNOR2_X1  g725(.A(new_n926), .B(KEYINPUT61), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n912), .A2(new_n257), .A3(new_n686), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(G1351gat));
  NOR2_X1   g728(.A1(new_n669), .A2(new_n908), .ZN(new_n930));
  AND2_X1   g729(.A1(new_n842), .A2(new_n930), .ZN(new_n931));
  INV_X1    g730(.A(G197gat), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n931), .A2(new_n932), .A3(new_n396), .ZN(new_n933));
  AND2_X1   g732(.A1(new_n877), .A2(new_n930), .ZN(new_n934));
  AND2_X1   g733(.A1(new_n934), .A2(new_n396), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n933), .B1(new_n935), .B2(new_n932), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT125), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n936), .B(new_n937), .ZN(G1352gat));
  AND3_X1   g737(.A1(new_n931), .A2(new_n282), .A3(new_n349), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT62), .ZN(new_n940));
  OR2_X1    g739(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n939), .A2(new_n940), .ZN(new_n942));
  AND3_X1   g741(.A1(new_n877), .A2(new_n349), .A3(new_n930), .ZN(new_n943));
  OAI211_X1 g742(.A(new_n941), .B(new_n942), .C1(new_n282), .C2(new_n943), .ZN(G1353gat));
  AOI21_X1  g743(.A(new_n412), .B1(new_n934), .B2(new_n420), .ZN(new_n945));
  XNOR2_X1  g744(.A(new_n945), .B(KEYINPUT63), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n931), .A2(new_n412), .A3(new_n420), .ZN(new_n947));
  XOR2_X1   g746(.A(new_n947), .B(KEYINPUT126), .Z(new_n948));
  NAND2_X1  g747(.A1(new_n946), .A2(new_n948), .ZN(G1354gat));
  AOI21_X1  g748(.A(new_n260), .B1(new_n934), .B2(new_n686), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n278), .A2(G218gat), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n950), .B1(new_n931), .B2(new_n951), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT127), .ZN(new_n953));
  XNOR2_X1  g752(.A(new_n952), .B(new_n953), .ZN(G1355gat));
endmodule


