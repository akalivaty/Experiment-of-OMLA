

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765;

  BUF_X1 U374 ( .A(n677), .Z(n351) );
  AND2_X2 U375 ( .A1(n708), .A2(n542), .ZN(n530) );
  NOR2_X1 U376 ( .A1(G953), .A2(G237), .ZN(n495) );
  XNOR2_X1 U377 ( .A(n416), .B(n415), .ZN(n500) );
  INV_X1 U378 ( .A(G953), .ZN(n760) );
  XNOR2_X2 U379 ( .A(n369), .B(n386), .ZN(n464) );
  XNOR2_X2 U380 ( .A(n502), .B(n468), .ZN(n754) );
  XNOR2_X2 U381 ( .A(n591), .B(n478), .ZN(n542) );
  NAND2_X1 U382 ( .A1(n514), .A2(n537), .ZN(n729) );
  XNOR2_X1 U383 ( .A(n600), .B(KEYINPUT19), .ZN(n607) );
  INV_X1 U384 ( .A(n593), .ZN(n714) );
  NOR2_X1 U385 ( .A1(n545), .A2(n579), .ZN(n546) );
  BUF_X1 U386 ( .A(n541), .Z(n543) );
  XNOR2_X1 U387 ( .A(n381), .B(n380), .ZN(n765) );
  NAND2_X1 U388 ( .A1(n615), .A2(n614), .ZN(n688) );
  BUF_X1 U389 ( .A(n513), .Z(n723) );
  XNOR2_X1 U390 ( .A(n382), .B(n361), .ZN(n513) );
  NAND2_X1 U391 ( .A1(n607), .A2(n429), .ZN(n369) );
  NAND2_X2 U392 ( .A1(n365), .A2(n364), .ZN(n611) );
  XNOR2_X1 U393 ( .A(n611), .B(n392), .ZN(n727) );
  INV_X1 U394 ( .A(KEYINPUT38), .ZN(n392) );
  NAND2_X1 U395 ( .A1(n611), .A2(n726), .ZN(n600) );
  NOR2_X1 U396 ( .A1(n765), .A2(n764), .ZN(n598) );
  NAND2_X1 U397 ( .A1(n727), .A2(n726), .ZN(n383) );
  BUF_X1 U398 ( .A(n542), .Z(n707) );
  XNOR2_X1 U399 ( .A(G101), .B(KEYINPUT3), .ZN(n415) );
  XNOR2_X1 U400 ( .A(G116), .B(G113), .ZN(n414) );
  XNOR2_X1 U401 ( .A(G110), .B(G107), .ZN(n472) );
  XNOR2_X1 U402 ( .A(n597), .B(KEYINPUT39), .ZN(n629) );
  OR2_X1 U403 ( .A1(n671), .A2(n353), .ZN(n364) );
  AND2_X1 U404 ( .A1(n367), .A2(n366), .ZN(n365) );
  XNOR2_X1 U405 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U406 ( .A(n490), .B(KEYINPUT95), .ZN(n491) );
  XNOR2_X1 U407 ( .A(n466), .B(n363), .ZN(n506) );
  NOR2_X1 U408 ( .A1(n376), .A2(n544), .ZN(n375) );
  NOR2_X1 U409 ( .A1(n400), .A2(KEYINPUT85), .ZN(n376) );
  NAND2_X1 U410 ( .A1(n372), .A2(n355), .ZN(n371) );
  AND2_X1 U411 ( .A1(n388), .A2(KEYINPUT44), .ZN(n387) );
  NAND2_X1 U412 ( .A1(n391), .A2(n390), .ZN(n388) );
  XNOR2_X1 U413 ( .A(n422), .B(n421), .ZN(n564) );
  INV_X1 U414 ( .A(G237), .ZN(n418) );
  XNOR2_X1 U415 ( .A(n458), .B(n457), .ZN(n489) );
  XNOR2_X1 U416 ( .A(G143), .B(G113), .ZN(n433) );
  INV_X1 U417 ( .A(n383), .ZN(n724) );
  NAND2_X1 U418 ( .A1(n384), .A2(n352), .ZN(n366) );
  AND2_X1 U419 ( .A1(n708), .A2(n592), .ZN(n404) );
  INV_X1 U420 ( .A(KEYINPUT0), .ZN(n386) );
  NOR2_X1 U421 ( .A1(n729), .A2(n463), .ZN(n368) );
  XNOR2_X1 U422 ( .A(G128), .B(G110), .ZN(n479) );
  XNOR2_X1 U423 ( .A(G122), .B(G107), .ZN(n444) );
  XOR2_X1 U424 ( .A(G140), .B(G146), .Z(n470) );
  XNOR2_X1 U425 ( .A(G104), .B(G101), .ZN(n469) );
  INV_X1 U426 ( .A(KEYINPUT4), .ZN(n394) );
  XNOR2_X1 U427 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n406) );
  INV_X1 U428 ( .A(KEYINPUT41), .ZN(n582) );
  NOR2_X1 U429 ( .A1(n729), .A2(n383), .ZN(n583) );
  XNOR2_X1 U430 ( .A(n374), .B(n373), .ZN(n372) );
  INV_X1 U431 ( .A(KEYINPUT34), .ZN(n373) );
  NAND2_X1 U432 ( .A1(n513), .A2(n534), .ZN(n374) );
  XNOR2_X1 U433 ( .A(n417), .B(n500), .ZN(n560) );
  AND2_X1 U434 ( .A1(n647), .A2(G953), .ZN(n752) );
  NAND2_X1 U435 ( .A1(n577), .A2(n393), .ZN(n627) );
  XNOR2_X1 U436 ( .A(n379), .B(n377), .ZN(n764) );
  XNOR2_X1 U437 ( .A(n589), .B(n378), .ZN(n377) );
  NAND2_X1 U438 ( .A1(n740), .A2(n608), .ZN(n379) );
  INV_X1 U439 ( .A(KEYINPUT107), .ZN(n378) );
  INV_X1 U440 ( .A(KEYINPUT40), .ZN(n380) );
  NAND2_X1 U441 ( .A1(n541), .A2(n519), .ZN(n521) );
  NAND2_X1 U442 ( .A1(n396), .A2(n397), .ZN(n579) );
  NAND2_X1 U443 ( .A1(n543), .A2(n398), .ZN(n397) );
  NOR2_X1 U444 ( .A1(n359), .A2(n544), .ZN(n398) );
  AND2_X1 U445 ( .A1(n419), .A2(G210), .ZN(n352) );
  OR2_X1 U446 ( .A1(n384), .A2(n352), .ZN(n353) );
  XOR2_X1 U447 ( .A(G134), .B(G131), .Z(n354) );
  XOR2_X1 U448 ( .A(n614), .B(n516), .Z(n355) );
  XOR2_X1 U449 ( .A(KEYINPUT14), .B(KEYINPUT89), .Z(n356) );
  XOR2_X1 U450 ( .A(n566), .B(KEYINPUT103), .Z(n357) );
  AND2_X1 U451 ( .A1(n389), .A2(n387), .ZN(n358) );
  OR2_X1 U452 ( .A1(n707), .A2(KEYINPUT85), .ZN(n359) );
  INV_X1 U453 ( .A(n400), .ZN(n399) );
  AND2_X1 U454 ( .A1(n707), .A2(KEYINPUT85), .ZN(n400) );
  AND2_X1 U455 ( .A1(n627), .A2(n701), .ZN(n360) );
  XOR2_X1 U456 ( .A(n511), .B(KEYINPUT33), .Z(n361) );
  XNOR2_X1 U457 ( .A(n517), .B(KEYINPUT77), .ZN(n362) );
  XOR2_X1 U458 ( .A(n465), .B(KEYINPUT22), .Z(n363) );
  INV_X1 U459 ( .A(n632), .ZN(n384) );
  NAND2_X1 U460 ( .A1(n671), .A2(n352), .ZN(n367) );
  NAND2_X1 U461 ( .A1(n464), .A2(n368), .ZN(n466) );
  XNOR2_X2 U462 ( .A(n370), .B(n477), .ZN(n591) );
  OR2_X2 U463 ( .A1(n665), .A2(G902), .ZN(n370) );
  XNOR2_X2 U464 ( .A(n371), .B(n362), .ZN(n677) );
  NAND2_X1 U465 ( .A1(n395), .A2(n375), .ZN(n396) );
  NAND2_X1 U466 ( .A1(n629), .A2(n689), .ZN(n381) );
  NAND2_X1 U467 ( .A1(n530), .A2(n571), .ZN(n382) );
  NAND2_X1 U468 ( .A1(n628), .A2(n627), .ZN(n640) );
  NAND2_X1 U469 ( .A1(n628), .A2(n360), .ZN(n637) );
  XNOR2_X1 U470 ( .A(n560), .B(n385), .ZN(n671) );
  XNOR2_X1 U471 ( .A(n411), .B(n410), .ZN(n385) );
  INV_X1 U472 ( .A(n464), .ZN(n512) );
  NOR2_X1 U473 ( .A1(n563), .A2(n391), .ZN(n526) );
  NAND2_X1 U474 ( .A1(n563), .A2(n390), .ZN(n389) );
  INV_X1 U475 ( .A(KEYINPUT65), .ZN(n390) );
  INV_X1 U476 ( .A(n539), .ZN(n391) );
  INV_X2 U477 ( .A(KEYINPUT10), .ZN(n430) );
  NOR2_X2 U478 ( .A1(n596), .A2(n595), .ZN(n612) );
  XNOR2_X1 U479 ( .A(n583), .B(n582), .ZN(n740) );
  INV_X1 U480 ( .A(n611), .ZN(n393) );
  XNOR2_X2 U481 ( .A(n411), .B(n354), .ZN(n502) );
  XNOR2_X2 U482 ( .A(n447), .B(n394), .ZN(n411) );
  NOR2_X2 U483 ( .A1(n506), .A2(n571), .ZN(n541) );
  NAND2_X1 U484 ( .A1(n543), .A2(n399), .ZN(n395) );
  XNOR2_X2 U485 ( .A(n432), .B(n431), .ZN(n753) );
  XNOR2_X2 U486 ( .A(n430), .B(G140), .ZN(n431) );
  XNOR2_X2 U487 ( .A(n405), .B(G128), .ZN(n447) );
  XOR2_X1 U488 ( .A(KEYINPUT84), .B(KEYINPUT48), .Z(n401) );
  XNOR2_X1 U489 ( .A(KEYINPUT81), .B(KEYINPUT23), .ZN(n402) );
  XOR2_X1 U490 ( .A(n622), .B(KEYINPUT74), .Z(n403) );
  INV_X1 U491 ( .A(KEYINPUT93), .ZN(n421) );
  NOR2_X1 U492 ( .A1(n623), .A2(n403), .ZN(n624) );
  NOR2_X1 U493 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U494 ( .A(KEYINPUT94), .B(KEYINPUT20), .ZN(n457) );
  XNOR2_X1 U495 ( .A(n552), .B(KEYINPUT45), .ZN(n580) );
  XNOR2_X1 U496 ( .A(n482), .B(n402), .ZN(n488) );
  BUF_X1 U497 ( .A(n637), .Z(n759) );
  INV_X1 U498 ( .A(n553), .ZN(n703) );
  XNOR2_X2 U499 ( .A(G143), .B(KEYINPUT64), .ZN(n405) );
  XNOR2_X2 U500 ( .A(G146), .B(G125), .ZN(n432) );
  XNOR2_X1 U501 ( .A(n432), .B(n406), .ZN(n409) );
  NAND2_X1 U502 ( .A1(n760), .A2(G224), .ZN(n407) );
  XNOR2_X1 U503 ( .A(n407), .B(KEYINPUT88), .ZN(n408) );
  XNOR2_X1 U504 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X2 U505 ( .A(G122), .B(G104), .ZN(n439) );
  XNOR2_X1 U506 ( .A(KEYINPUT73), .B(KEYINPUT16), .ZN(n412) );
  XNOR2_X1 U507 ( .A(n439), .B(n412), .ZN(n413) );
  XNOR2_X1 U508 ( .A(n413), .B(n472), .ZN(n417) );
  XNOR2_X1 U509 ( .A(n414), .B(G119), .ZN(n416) );
  XNOR2_X1 U510 ( .A(G902), .B(KEYINPUT15), .ZN(n632) );
  INV_X1 U511 ( .A(G902), .ZN(n476) );
  NAND2_X1 U512 ( .A1(n476), .A2(n418), .ZN(n419) );
  NAND2_X1 U513 ( .A1(n419), .A2(G214), .ZN(n726) );
  INV_X1 U514 ( .A(n726), .ZN(n573) );
  NAND2_X1 U515 ( .A1(G237), .A2(G234), .ZN(n420) );
  XNOR2_X1 U516 ( .A(n356), .B(n420), .ZN(n425) );
  NAND2_X1 U517 ( .A1(n425), .A2(G902), .ZN(n422) );
  INV_X1 U518 ( .A(n564), .ZN(n424) );
  XOR2_X1 U519 ( .A(G898), .B(KEYINPUT92), .Z(n556) );
  NAND2_X1 U520 ( .A1(G953), .A2(n556), .ZN(n559) );
  INV_X1 U521 ( .A(n559), .ZN(n423) );
  NAND2_X1 U522 ( .A1(n424), .A2(n423), .ZN(n428) );
  NAND2_X1 U523 ( .A1(n425), .A2(G952), .ZN(n426) );
  XNOR2_X1 U524 ( .A(n426), .B(KEYINPUT90), .ZN(n739) );
  NOR2_X1 U525 ( .A1(n739), .A2(G953), .ZN(n427) );
  XNOR2_X1 U526 ( .A(n427), .B(KEYINPUT91), .ZN(n567) );
  NAND2_X1 U527 ( .A1(n428), .A2(n567), .ZN(n429) );
  XOR2_X1 U528 ( .A(KEYINPUT12), .B(G131), .Z(n434) );
  XNOR2_X1 U529 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U530 ( .A(n753), .B(n435), .Z(n437) );
  NAND2_X1 U531 ( .A1(n495), .A2(G214), .ZN(n436) );
  XNOR2_X1 U532 ( .A(n437), .B(n436), .ZN(n441) );
  INV_X1 U533 ( .A(KEYINPUT11), .ZN(n438) );
  XNOR2_X1 U534 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U535 ( .A(n441), .B(n440), .ZN(n658) );
  NAND2_X1 U536 ( .A1(n658), .A2(n476), .ZN(n443) );
  XNOR2_X1 U537 ( .A(KEYINPUT13), .B(G475), .ZN(n442) );
  XNOR2_X1 U538 ( .A(n443), .B(n442), .ZN(n537) );
  XOR2_X1 U539 ( .A(G134), .B(G116), .Z(n445) );
  XNOR2_X1 U540 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U541 ( .A(n447), .B(n446), .ZN(n453) );
  NAND2_X1 U542 ( .A1(G234), .A2(n760), .ZN(n448) );
  XOR2_X1 U543 ( .A(KEYINPUT8), .B(n448), .Z(n484) );
  NAND2_X1 U544 ( .A1(G217), .A2(n484), .ZN(n451) );
  INV_X1 U545 ( .A(KEYINPUT7), .ZN(n449) );
  XNOR2_X1 U546 ( .A(n449), .B(KEYINPUT9), .ZN(n450) );
  XNOR2_X1 U547 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U548 ( .A(n453), .B(n452), .ZN(n645) );
  NOR2_X1 U549 ( .A1(n645), .A2(G902), .ZN(n454) );
  XOR2_X1 U550 ( .A(KEYINPUT99), .B(n454), .Z(n456) );
  INV_X1 U551 ( .A(G478), .ZN(n455) );
  XNOR2_X1 U552 ( .A(n456), .B(n455), .ZN(n536) );
  INV_X1 U553 ( .A(n536), .ZN(n514) );
  NAND2_X1 U554 ( .A1(n632), .A2(G234), .ZN(n458) );
  NAND2_X1 U555 ( .A1(G221), .A2(n489), .ZN(n462) );
  XOR2_X1 U556 ( .A(KEYINPUT96), .B(KEYINPUT97), .Z(n460) );
  INV_X1 U557 ( .A(KEYINPUT21), .ZN(n459) );
  XNOR2_X1 U558 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U559 ( .A(n462), .B(n461), .ZN(n710) );
  INV_X1 U560 ( .A(n710), .ZN(n463) );
  INV_X1 U561 ( .A(KEYINPUT66), .ZN(n465) );
  INV_X1 U562 ( .A(KEYINPUT70), .ZN(n467) );
  XNOR2_X1 U563 ( .A(n467), .B(G137), .ZN(n483) );
  INV_X1 U564 ( .A(n483), .ZN(n468) );
  XNOR2_X1 U565 ( .A(n470), .B(n469), .ZN(n474) );
  NAND2_X1 U566 ( .A1(n760), .A2(G227), .ZN(n471) );
  XNOR2_X1 U567 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U568 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X1 U569 ( .A(n754), .B(n475), .ZN(n665) );
  INV_X1 U570 ( .A(G469), .ZN(n477) );
  XNOR2_X1 U571 ( .A(KEYINPUT67), .B(KEYINPUT1), .ZN(n478) );
  INV_X1 U572 ( .A(n542), .ZN(n605) );
  XOR2_X1 U573 ( .A(KEYINPUT24), .B(G119), .Z(n480) );
  XNOR2_X1 U574 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U575 ( .A(n753), .B(n481), .ZN(n482) );
  XOR2_X1 U576 ( .A(n483), .B(KEYINPUT71), .Z(n486) );
  NAND2_X1 U577 ( .A1(G221), .A2(n484), .ZN(n485) );
  XNOR2_X1 U578 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U579 ( .A(n488), .B(n487), .ZN(n748) );
  NOR2_X1 U580 ( .A1(n748), .A2(G902), .ZN(n494) );
  NAND2_X1 U581 ( .A1(G217), .A2(n489), .ZN(n492) );
  XOR2_X1 U582 ( .A(KEYINPUT25), .B(KEYINPUT76), .Z(n490) );
  XNOR2_X2 U583 ( .A(n494), .B(n493), .ZN(n711) );
  NAND2_X1 U584 ( .A1(n495), .A2(G210), .ZN(n496) );
  XNOR2_X1 U585 ( .A(n496), .B(G137), .ZN(n498) );
  XNOR2_X1 U586 ( .A(G146), .B(KEYINPUT5), .ZN(n497) );
  XNOR2_X1 U587 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U588 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U589 ( .A(n502), .B(n501), .ZN(n652) );
  OR2_X1 U590 ( .A1(n652), .A2(G902), .ZN(n503) );
  XNOR2_X1 U591 ( .A(n503), .B(G472), .ZN(n593) );
  NOR2_X1 U592 ( .A1(n711), .A2(n593), .ZN(n504) );
  NAND2_X1 U593 ( .A1(n605), .A2(n504), .ZN(n505) );
  OR2_X1 U594 ( .A1(n506), .A2(n505), .ZN(n539) );
  XNOR2_X1 U595 ( .A(n539), .B(G110), .ZN(G12) );
  NAND2_X1 U596 ( .A1(n711), .A2(n710), .ZN(n508) );
  INV_X1 U597 ( .A(KEYINPUT68), .ZN(n507) );
  XNOR2_X2 U598 ( .A(n508), .B(n507), .ZN(n708) );
  INV_X1 U599 ( .A(KEYINPUT100), .ZN(n509) );
  XNOR2_X1 U600 ( .A(n509), .B(KEYINPUT6), .ZN(n510) );
  XNOR2_X1 U601 ( .A(n593), .B(n510), .ZN(n571) );
  INV_X1 U602 ( .A(KEYINPUT72), .ZN(n511) );
  INV_X1 U603 ( .A(n512), .ZN(n534) );
  NOR2_X1 U604 ( .A1(n537), .A2(n514), .ZN(n515) );
  XNOR2_X1 U605 ( .A(n515), .B(KEYINPUT102), .ZN(n614) );
  INV_X1 U606 ( .A(KEYINPUT78), .ZN(n516) );
  XNOR2_X1 U607 ( .A(KEYINPUT83), .B(KEYINPUT35), .ZN(n517) );
  INV_X1 U608 ( .A(n677), .ZN(n522) );
  OR2_X1 U609 ( .A1(n605), .A2(n711), .ZN(n518) );
  XNOR2_X1 U610 ( .A(n518), .B(KEYINPUT101), .ZN(n519) );
  INV_X1 U611 ( .A(KEYINPUT32), .ZN(n520) );
  XNOR2_X2 U612 ( .A(n521), .B(n520), .ZN(n563) );
  NAND2_X1 U613 ( .A1(n522), .A2(n526), .ZN(n525) );
  NOR2_X1 U614 ( .A1(KEYINPUT65), .A2(KEYINPUT44), .ZN(n523) );
  AND2_X1 U615 ( .A1(n523), .A2(KEYINPUT86), .ZN(n524) );
  NAND2_X1 U616 ( .A1(n525), .A2(n524), .ZN(n529) );
  NAND2_X1 U617 ( .A1(n677), .A2(KEYINPUT86), .ZN(n527) );
  NAND2_X1 U618 ( .A1(n527), .A2(n358), .ZN(n528) );
  NAND2_X1 U619 ( .A1(n529), .A2(n528), .ZN(n551) );
  NOR2_X1 U620 ( .A1(n677), .A2(KEYINPUT86), .ZN(n549) );
  NAND2_X1 U621 ( .A1(n530), .A2(n593), .ZN(n531) );
  XNOR2_X1 U622 ( .A(n531), .B(KEYINPUT98), .ZN(n719) );
  NOR2_X1 U623 ( .A1(n719), .A2(n512), .ZN(n532) );
  XNOR2_X1 U624 ( .A(n532), .B(KEYINPUT31), .ZN(n695) );
  NAND2_X1 U625 ( .A1(n708), .A2(n714), .ZN(n533) );
  NOR2_X1 U626 ( .A1(n533), .A2(n591), .ZN(n535) );
  NAND2_X1 U627 ( .A1(n535), .A2(n534), .ZN(n679) );
  NAND2_X1 U628 ( .A1(n695), .A2(n679), .ZN(n538) );
  OR2_X1 U629 ( .A1(n536), .A2(n537), .ZN(n692) );
  NAND2_X1 U630 ( .A1(n537), .A2(n536), .ZN(n696) );
  NAND2_X1 U631 ( .A1(n692), .A2(n696), .ZN(n725) );
  NAND2_X1 U632 ( .A1(n538), .A2(n725), .ZN(n547) );
  NAND2_X1 U633 ( .A1(n539), .A2(KEYINPUT65), .ZN(n540) );
  NOR2_X1 U634 ( .A1(n563), .A2(n540), .ZN(n545) );
  INV_X1 U635 ( .A(n711), .ZN(n544) );
  NAND2_X1 U636 ( .A1(n547), .A2(n546), .ZN(n548) );
  NOR2_X1 U637 ( .A1(n549), .A2(n548), .ZN(n550) );
  NAND2_X1 U638 ( .A1(n551), .A2(n550), .ZN(n552) );
  BUF_X1 U639 ( .A(n580), .Z(n553) );
  NOR2_X1 U640 ( .A1(n703), .A2(G953), .ZN(n558) );
  NAND2_X1 U641 ( .A1(G953), .A2(G224), .ZN(n554) );
  XOR2_X1 U642 ( .A(KEYINPUT61), .B(n554), .Z(n555) );
  NOR2_X1 U643 ( .A1(n556), .A2(n555), .ZN(n557) );
  NOR2_X1 U644 ( .A1(n558), .A2(n557), .ZN(n562) );
  NAND2_X1 U645 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U646 ( .A(n562), .B(n561), .ZN(G69) );
  XOR2_X1 U647 ( .A(n563), .B(G119), .Z(G21) );
  OR2_X2 U648 ( .A1(n760), .A2(n564), .ZN(n565) );
  NOR2_X2 U649 ( .A1(G900), .A2(n565), .ZN(n566) );
  INV_X1 U650 ( .A(n567), .ZN(n568) );
  NOR2_X1 U651 ( .A1(n357), .A2(n568), .ZN(n590) );
  INV_X1 U652 ( .A(n590), .ZN(n569) );
  NAND2_X1 U653 ( .A1(n710), .A2(n569), .ZN(n570) );
  OR2_X1 U654 ( .A1(n711), .A2(n570), .ZN(n584) );
  NOR2_X1 U655 ( .A1(n584), .A2(n692), .ZN(n572) );
  NAND2_X1 U656 ( .A1(n572), .A2(n571), .ZN(n599) );
  NOR2_X1 U657 ( .A1(n599), .A2(n573), .ZN(n574) );
  NAND2_X1 U658 ( .A1(n574), .A2(n605), .ZN(n576) );
  XNOR2_X1 U659 ( .A(KEYINPUT43), .B(KEYINPUT104), .ZN(n575) );
  XNOR2_X1 U660 ( .A(n576), .B(n575), .ZN(n577) );
  XOR2_X1 U661 ( .A(G140), .B(KEYINPUT117), .Z(n578) );
  XNOR2_X1 U662 ( .A(n627), .B(n578), .ZN(G42) );
  XOR2_X1 U663 ( .A(G101), .B(n579), .Z(G3) );
  NAND2_X1 U664 ( .A1(n580), .A2(n384), .ZN(n581) );
  XNOR2_X1 U665 ( .A(n581), .B(KEYINPUT82), .ZN(n630) );
  XOR2_X1 U666 ( .A(KEYINPUT108), .B(KEYINPUT42), .Z(n589) );
  NOR2_X2 U667 ( .A1(n584), .A2(n714), .ZN(n585) );
  XNOR2_X1 U668 ( .A(n585), .B(KEYINPUT28), .ZN(n588) );
  INV_X1 U669 ( .A(KEYINPUT106), .ZN(n586) );
  XNOR2_X1 U670 ( .A(n591), .B(n586), .ZN(n587) );
  AND2_X2 U671 ( .A1(n588), .A2(n587), .ZN(n608) );
  INV_X1 U672 ( .A(n692), .ZN(n689) );
  XNOR2_X1 U673 ( .A(n404), .B(KEYINPUT75), .ZN(n596) );
  NAND2_X1 U674 ( .A1(n593), .A2(n726), .ZN(n594) );
  XNOR2_X1 U675 ( .A(n594), .B(KEYINPUT30), .ZN(n595) );
  NAND2_X1 U676 ( .A1(n612), .A2(n727), .ZN(n597) );
  XNOR2_X1 U677 ( .A(n598), .B(KEYINPUT46), .ZN(n625) );
  XNOR2_X1 U678 ( .A(n599), .B(KEYINPUT109), .ZN(n602) );
  INV_X1 U679 ( .A(n600), .ZN(n601) );
  NAND2_X1 U680 ( .A1(n602), .A2(n601), .ZN(n604) );
  XNOR2_X1 U681 ( .A(KEYINPUT110), .B(KEYINPUT36), .ZN(n603) );
  XNOR2_X1 U682 ( .A(n604), .B(n603), .ZN(n606) );
  OR2_X1 U683 ( .A1(n606), .A2(n605), .ZN(n699) );
  INV_X1 U684 ( .A(n699), .ZN(n619) );
  NAND2_X1 U685 ( .A1(n608), .A2(n607), .ZN(n684) );
  INV_X1 U686 ( .A(n725), .ZN(n609) );
  NOR2_X2 U687 ( .A1(n684), .A2(n609), .ZN(n620) );
  INV_X1 U688 ( .A(KEYINPUT47), .ZN(n610) );
  OR2_X1 U689 ( .A1(n620), .A2(n610), .ZN(n616) );
  NAND2_X1 U690 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U691 ( .A(n613), .B(KEYINPUT105), .ZN(n615) );
  NAND2_X1 U692 ( .A1(n616), .A2(n688), .ZN(n617) );
  XNOR2_X1 U693 ( .A(n617), .B(KEYINPUT80), .ZN(n618) );
  OR2_X2 U694 ( .A1(n619), .A2(n618), .ZN(n623) );
  XNOR2_X1 U695 ( .A(KEYINPUT47), .B(KEYINPUT69), .ZN(n621) );
  NAND2_X1 U696 ( .A1(n621), .A2(n620), .ZN(n622) );
  NAND2_X1 U697 ( .A1(n625), .A2(n624), .ZN(n626) );
  XNOR2_X1 U698 ( .A(n626), .B(n401), .ZN(n628) );
  INV_X1 U699 ( .A(n696), .ZN(n685) );
  NAND2_X1 U700 ( .A1(n629), .A2(n685), .ZN(n701) );
  NOR2_X1 U701 ( .A1(n630), .A2(n759), .ZN(n634) );
  INV_X1 U702 ( .A(KEYINPUT2), .ZN(n631) );
  NOR2_X1 U703 ( .A1(n632), .A2(n631), .ZN(n633) );
  NOR2_X1 U704 ( .A1(n634), .A2(n633), .ZN(n644) );
  INV_X1 U705 ( .A(KEYINPUT79), .ZN(n635) );
  NAND2_X1 U706 ( .A1(n635), .A2(KEYINPUT2), .ZN(n636) );
  NOR2_X1 U707 ( .A1(n637), .A2(n636), .ZN(n642) );
  NAND2_X1 U708 ( .A1(n701), .A2(KEYINPUT2), .ZN(n638) );
  NAND2_X1 U709 ( .A1(n638), .A2(KEYINPUT79), .ZN(n639) );
  NOR2_X1 U710 ( .A1(n640), .A2(n639), .ZN(n641) );
  OR2_X2 U711 ( .A1(n642), .A2(n641), .ZN(n643) );
  AND2_X2 U712 ( .A1(n643), .A2(n553), .ZN(n706) );
  NOR2_X4 U713 ( .A1(n644), .A2(n706), .ZN(n747) );
  NAND2_X1 U714 ( .A1(n747), .A2(G478), .ZN(n646) );
  XNOR2_X1 U715 ( .A(n646), .B(n645), .ZN(n648) );
  INV_X1 U716 ( .A(G952), .ZN(n647) );
  NOR2_X2 U717 ( .A1(n648), .A2(n752), .ZN(n649) );
  XNOR2_X1 U718 ( .A(n649), .B(KEYINPUT124), .ZN(G63) );
  NAND2_X1 U719 ( .A1(n747), .A2(G472), .ZN(n654) );
  XOR2_X1 U720 ( .A(KEYINPUT111), .B(KEYINPUT112), .Z(n650) );
  XNOR2_X1 U721 ( .A(n650), .B(KEYINPUT62), .ZN(n651) );
  XNOR2_X1 U722 ( .A(n652), .B(n651), .ZN(n653) );
  XNOR2_X1 U723 ( .A(n654), .B(n653), .ZN(n655) );
  NOR2_X2 U724 ( .A1(n655), .A2(n752), .ZN(n657) );
  XNOR2_X1 U725 ( .A(KEYINPUT87), .B(KEYINPUT63), .ZN(n656) );
  XNOR2_X1 U726 ( .A(n657), .B(n656), .ZN(G57) );
  NAND2_X1 U727 ( .A1(n747), .A2(G475), .ZN(n660) );
  XNOR2_X1 U728 ( .A(n658), .B(KEYINPUT59), .ZN(n659) );
  XNOR2_X1 U729 ( .A(n660), .B(n659), .ZN(n661) );
  NOR2_X2 U730 ( .A1(n661), .A2(n752), .ZN(n663) );
  XOR2_X1 U731 ( .A(KEYINPUT123), .B(KEYINPUT60), .Z(n662) );
  XNOR2_X1 U732 ( .A(n663), .B(n662), .ZN(G60) );
  NAND2_X1 U733 ( .A1(n747), .A2(G469), .ZN(n667) );
  XOR2_X1 U734 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n664) );
  XNOR2_X1 U735 ( .A(n665), .B(n664), .ZN(n666) );
  XNOR2_X1 U736 ( .A(n667), .B(n666), .ZN(n668) );
  NOR2_X2 U737 ( .A1(n668), .A2(n752), .ZN(n669) );
  XNOR2_X1 U738 ( .A(n669), .B(KEYINPUT122), .ZN(G54) );
  NAND2_X1 U739 ( .A1(n747), .A2(G210), .ZN(n673) );
  XOR2_X1 U740 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n670) );
  XNOR2_X1 U741 ( .A(n671), .B(n670), .ZN(n672) );
  XNOR2_X1 U742 ( .A(n673), .B(n672), .ZN(n674) );
  NOR2_X2 U743 ( .A1(n674), .A2(n752), .ZN(n675) );
  XNOR2_X1 U744 ( .A(n675), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U745 ( .A(G122), .B(KEYINPUT127), .ZN(n676) );
  XNOR2_X1 U746 ( .A(n351), .B(n676), .ZN(G24) );
  NOR2_X1 U747 ( .A1(n679), .A2(n692), .ZN(n678) );
  XOR2_X1 U748 ( .A(G104), .B(n678), .Z(G6) );
  NOR2_X1 U749 ( .A1(n679), .A2(n696), .ZN(n683) );
  XOR2_X1 U750 ( .A(KEYINPUT26), .B(KEYINPUT27), .Z(n681) );
  XNOR2_X1 U751 ( .A(G107), .B(KEYINPUT113), .ZN(n680) );
  XNOR2_X1 U752 ( .A(n681), .B(n680), .ZN(n682) );
  XNOR2_X1 U753 ( .A(n683), .B(n682), .ZN(G9) );
  XOR2_X1 U754 ( .A(G128), .B(KEYINPUT29), .Z(n687) );
  INV_X1 U755 ( .A(n684), .ZN(n690) );
  NAND2_X1 U756 ( .A1(n690), .A2(n685), .ZN(n686) );
  XNOR2_X1 U757 ( .A(n687), .B(n686), .ZN(G30) );
  XNOR2_X1 U758 ( .A(G143), .B(n688), .ZN(G45) );
  NAND2_X1 U759 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U760 ( .A(G146), .B(n691), .ZN(G48) );
  NOR2_X1 U761 ( .A1(n692), .A2(n695), .ZN(n693) );
  XOR2_X1 U762 ( .A(KEYINPUT114), .B(n693), .Z(n694) );
  XNOR2_X1 U763 ( .A(G113), .B(n694), .ZN(G15) );
  NOR2_X1 U764 ( .A1(n696), .A2(n695), .ZN(n697) );
  XOR2_X1 U765 ( .A(G116), .B(n697), .Z(G18) );
  XNOR2_X1 U766 ( .A(KEYINPUT115), .B(KEYINPUT37), .ZN(n698) );
  XNOR2_X1 U767 ( .A(n699), .B(n698), .ZN(n700) );
  XNOR2_X1 U768 ( .A(G125), .B(n700), .ZN(G27) );
  XNOR2_X1 U769 ( .A(G134), .B(KEYINPUT116), .ZN(n702) );
  XNOR2_X1 U770 ( .A(n702), .B(n701), .ZN(G36) );
  NOR2_X1 U771 ( .A1(n759), .A2(n703), .ZN(n704) );
  NOR2_X1 U772 ( .A1(n704), .A2(KEYINPUT2), .ZN(n705) );
  NOR2_X1 U773 ( .A1(n706), .A2(n705), .ZN(n744) );
  XOR2_X1 U774 ( .A(KEYINPUT121), .B(KEYINPUT52), .Z(n737) );
  NOR2_X1 U775 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U776 ( .A(n709), .B(KEYINPUT50), .ZN(n717) );
  XNOR2_X1 U777 ( .A(KEYINPUT49), .B(KEYINPUT118), .ZN(n713) );
  NOR2_X1 U778 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U779 ( .A(n713), .B(n712), .ZN(n715) );
  NAND2_X1 U780 ( .A1(n715), .A2(n714), .ZN(n716) );
  NOR2_X1 U781 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U782 ( .A(n718), .B(KEYINPUT119), .ZN(n720) );
  NAND2_X1 U783 ( .A1(n720), .A2(n719), .ZN(n721) );
  XOR2_X1 U784 ( .A(KEYINPUT51), .B(n721), .Z(n722) );
  NAND2_X1 U785 ( .A1(n740), .A2(n722), .ZN(n735) );
  NAND2_X1 U786 ( .A1(n725), .A2(n724), .ZN(n732) );
  NOR2_X1 U787 ( .A1(n727), .A2(n726), .ZN(n728) );
  NOR2_X1 U788 ( .A1(n729), .A2(n728), .ZN(n730) );
  XOR2_X1 U789 ( .A(KEYINPUT120), .B(n730), .Z(n731) );
  NAND2_X1 U790 ( .A1(n732), .A2(n731), .ZN(n733) );
  NAND2_X1 U791 ( .A1(n723), .A2(n733), .ZN(n734) );
  NAND2_X1 U792 ( .A1(n735), .A2(n734), .ZN(n736) );
  XOR2_X1 U793 ( .A(n737), .B(n736), .Z(n738) );
  NOR2_X1 U794 ( .A1(n739), .A2(n738), .ZN(n742) );
  AND2_X1 U795 ( .A1(n740), .A2(n723), .ZN(n741) );
  OR2_X1 U796 ( .A1(n742), .A2(n741), .ZN(n743) );
  OR2_X1 U797 ( .A1(n744), .A2(n743), .ZN(n745) );
  NOR2_X1 U798 ( .A1(n745), .A2(G953), .ZN(n746) );
  XNOR2_X1 U799 ( .A(n746), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U800 ( .A1(n747), .A2(G217), .ZN(n750) );
  XOR2_X1 U801 ( .A(n748), .B(KEYINPUT125), .Z(n749) );
  XNOR2_X1 U802 ( .A(n750), .B(n749), .ZN(n751) );
  NOR2_X1 U803 ( .A1(n752), .A2(n751), .ZN(G66) );
  XNOR2_X1 U804 ( .A(n754), .B(n753), .ZN(n758) );
  XNOR2_X1 U805 ( .A(n758), .B(G227), .ZN(n755) );
  NAND2_X1 U806 ( .A1(n755), .A2(G900), .ZN(n756) );
  NAND2_X1 U807 ( .A1(n756), .A2(G953), .ZN(n757) );
  XNOR2_X1 U808 ( .A(n757), .B(KEYINPUT126), .ZN(n763) );
  XNOR2_X1 U809 ( .A(n759), .B(n758), .ZN(n761) );
  NAND2_X1 U810 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U811 ( .A1(n763), .A2(n762), .ZN(G72) );
  XOR2_X1 U812 ( .A(G137), .B(n764), .Z(G39) );
  XOR2_X1 U813 ( .A(G131), .B(n765), .Z(G33) );
endmodule

