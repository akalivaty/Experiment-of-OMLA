

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722;

  XNOR2_X2 U369 ( .A(n420), .B(n368), .ZN(n709) );
  INV_X2 U370 ( .A(G953), .ZN(n701) );
  AND2_X1 U371 ( .A1(n692), .A2(n576), .ZN(n577) );
  XNOR2_X1 U372 ( .A(n712), .B(n533), .ZN(n578) );
  AND2_X1 U373 ( .A1(n527), .A2(n526), .ZN(n528) );
  NOR2_X1 U374 ( .A1(n536), .A2(n535), .ZN(n538) );
  BUF_X1 U375 ( .A(n466), .Z(n517) );
  XNOR2_X1 U376 ( .A(n442), .B(n441), .ZN(n494) );
  XOR2_X1 U377 ( .A(n700), .B(n456), .Z(n457) );
  XNOR2_X1 U378 ( .A(n371), .B(n458), .ZN(n605) );
  XNOR2_X1 U379 ( .A(n450), .B(n449), .ZN(n700) );
  XNOR2_X1 U380 ( .A(n381), .B(n380), .ZN(n450) );
  INV_X1 U381 ( .A(KEYINPUT63), .ZN(n347) );
  XNOR2_X1 U382 ( .A(G131), .B(KEYINPUT69), .ZN(n362) );
  XNOR2_X1 U383 ( .A(n347), .B(n623), .ZN(G57) );
  AND2_X2 U384 ( .A1(n568), .A2(KEYINPUT85), .ZN(n552) );
  NOR2_X1 U385 ( .A1(n673), .A2(n647), .ZN(n509) );
  NOR2_X1 U386 ( .A1(n721), .A2(n722), .ZN(n505) );
  XNOR2_X1 U387 ( .A(n385), .B(G472), .ZN(n496) );
  XNOR2_X1 U388 ( .A(n379), .B(KEYINPUT3), .ZN(n381) );
  XNOR2_X1 U389 ( .A(G119), .B(G116), .ZN(n379) );
  XNOR2_X1 U390 ( .A(n358), .B(n357), .ZN(n356) );
  INV_X1 U391 ( .A(KEYINPUT34), .ZN(n357) );
  XNOR2_X1 U392 ( .A(n472), .B(n361), .ZN(n476) );
  NOR2_X1 U393 ( .A1(n564), .A2(n471), .ZN(n472) );
  NOR2_X1 U394 ( .A1(n701), .A2(G952), .ZN(n621) );
  XNOR2_X1 U395 ( .A(n525), .B(n524), .ZN(n526) );
  XOR2_X1 U396 ( .A(G137), .B(KEYINPUT70), .Z(n427) );
  INV_X1 U397 ( .A(KEYINPUT76), .ZN(n533) );
  XNOR2_X1 U398 ( .A(n543), .B(n542), .ZN(n558) );
  INV_X1 U399 ( .A(KEYINPUT75), .ZN(n542) );
  OR2_X1 U400 ( .A1(n485), .A2(n484), .ZN(n486) );
  XNOR2_X1 U401 ( .A(G128), .B(G119), .ZN(n425) );
  XNOR2_X1 U402 ( .A(n378), .B(n363), .ZN(n710) );
  INV_X1 U403 ( .A(n427), .ZN(n363) );
  XNOR2_X1 U404 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U405 ( .A(n467), .B(KEYINPUT19), .ZN(n359) );
  OR2_X1 U406 ( .A1(n466), .A2(n465), .ZN(n467) );
  NAND2_X1 U407 ( .A1(G953), .A2(G900), .ZN(n716) );
  XNOR2_X1 U408 ( .A(n491), .B(KEYINPUT107), .ZN(n492) );
  INV_X1 U409 ( .A(KEYINPUT35), .ZN(n353) );
  INV_X1 U410 ( .A(n548), .ZN(n355) );
  XNOR2_X1 U411 ( .A(n538), .B(n537), .ZN(n614) );
  INV_X1 U412 ( .A(KEYINPUT32), .ZN(n537) );
  NOR2_X1 U413 ( .A1(n594), .A2(n621), .ZN(n596) );
  NOR2_X1 U414 ( .A1(n612), .A2(n621), .ZN(n613) );
  NOR2_X1 U415 ( .A1(n602), .A2(n621), .ZN(n604) );
  AND2_X1 U416 ( .A1(n617), .A2(n615), .ZN(n348) );
  AND2_X1 U417 ( .A1(n469), .A2(n468), .ZN(n349) );
  AND2_X1 U418 ( .A1(n615), .A2(G469), .ZN(n350) );
  AND2_X1 U419 ( .A1(n615), .A2(G475), .ZN(n351) );
  AND2_X1 U420 ( .A1(n615), .A2(G210), .ZN(n352) );
  NAND2_X1 U421 ( .A1(n617), .A2(n352), .ZN(n601) );
  NAND2_X1 U422 ( .A1(n617), .A2(n350), .ZN(n611) );
  NAND2_X1 U423 ( .A1(n617), .A2(n351), .ZN(n593) );
  XNOR2_X2 U424 ( .A(n354), .B(n353), .ZN(n568) );
  NAND2_X1 U425 ( .A1(n356), .A2(n355), .ZN(n354) );
  OR2_X2 U426 ( .A1(n650), .A2(n564), .ZN(n358) );
  NAND2_X1 U427 ( .A1(n359), .A2(n349), .ZN(n470) );
  NAND2_X1 U428 ( .A1(n360), .A2(n359), .ZN(n673) );
  INV_X1 U429 ( .A(n506), .ZN(n360) );
  NAND2_X2 U430 ( .A1(n581), .A2(n580), .ZN(n617) );
  XOR2_X1 U431 ( .A(KEYINPUT73), .B(KEYINPUT22), .Z(n361) );
  INV_X1 U432 ( .A(KEYINPUT71), .ZN(n524) );
  INV_X1 U433 ( .A(KEYINPUT2), .ZN(n576) );
  INV_X1 U434 ( .A(n698), .ZN(n370) );
  XNOR2_X1 U435 ( .A(KEYINPUT102), .B(KEYINPUT30), .ZN(n497) );
  XNOR2_X1 U436 ( .A(n710), .B(n366), .ZN(n371) );
  XNOR2_X1 U437 ( .A(n708), .B(n433), .ZN(n434) );
  BUF_X1 U438 ( .A(n496), .Z(n637) );
  XNOR2_X1 U439 ( .A(n483), .B(n482), .ZN(n626) );
  XNOR2_X1 U440 ( .A(n440), .B(n439), .ZN(n441) );
  BUF_X1 U441 ( .A(n541), .Z(n627) );
  XNOR2_X1 U442 ( .A(n493), .B(n492), .ZN(n721) );
  INV_X1 U443 ( .A(n362), .ZN(n393) );
  XOR2_X1 U444 ( .A(G134), .B(n393), .Z(n378) );
  XOR2_X1 U445 ( .A(G146), .B(G140), .Z(n365) );
  NAND2_X1 U446 ( .A1(G227), .A2(n701), .ZN(n364) );
  XNOR2_X1 U447 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X2 U448 ( .A(KEYINPUT65), .B(G143), .ZN(n367) );
  XNOR2_X2 U449 ( .A(n367), .B(G128), .ZN(n420) );
  XNOR2_X1 U450 ( .A(KEYINPUT64), .B(KEYINPUT4), .ZN(n368) );
  XNOR2_X2 U451 ( .A(n709), .B(G101), .ZN(n383) );
  XNOR2_X1 U452 ( .A(G110), .B(G107), .ZN(n369) );
  XNOR2_X1 U453 ( .A(n369), .B(G104), .ZN(n698) );
  XNOR2_X2 U454 ( .A(n383), .B(n370), .ZN(n458) );
  INV_X1 U455 ( .A(G902), .ZN(n422) );
  NAND2_X1 U456 ( .A1(n605), .A2(n422), .ZN(n372) );
  XNOR2_X2 U457 ( .A(n372), .B(G469), .ZN(n488) );
  XNOR2_X1 U458 ( .A(n488), .B(KEYINPUT1), .ZN(n541) );
  XOR2_X1 U459 ( .A(KEYINPUT92), .B(KEYINPUT5), .Z(n374) );
  XNOR2_X1 U460 ( .A(G146), .B(G137), .ZN(n373) );
  XNOR2_X1 U461 ( .A(n374), .B(n373), .ZN(n376) );
  NOR2_X1 U462 ( .A1(G953), .A2(G237), .ZN(n394) );
  NAND2_X1 U463 ( .A1(n394), .A2(G210), .ZN(n375) );
  XNOR2_X1 U464 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U465 ( .A(n378), .B(n377), .ZN(n382) );
  XNOR2_X1 U466 ( .A(G113), .B(KEYINPUT72), .ZN(n380) );
  XNOR2_X1 U467 ( .A(n382), .B(n450), .ZN(n384) );
  XNOR2_X1 U468 ( .A(n384), .B(n383), .ZN(n618) );
  NAND2_X1 U469 ( .A1(n618), .A2(n422), .ZN(n385) );
  XNOR2_X1 U470 ( .A(n637), .B(KEYINPUT6), .ZN(n544) );
  NAND2_X1 U471 ( .A1(G234), .A2(G237), .ZN(n386) );
  XNOR2_X1 U472 ( .A(n386), .B(KEYINPUT14), .ZN(n656) );
  NOR2_X1 U473 ( .A1(G953), .A2(G952), .ZN(n388) );
  NOR2_X1 U474 ( .A1(G902), .A2(n701), .ZN(n387) );
  NOR2_X1 U475 ( .A1(n388), .A2(n387), .ZN(n389) );
  AND2_X1 U476 ( .A1(n656), .A2(n389), .ZN(n469) );
  NAND2_X1 U477 ( .A1(n469), .A2(n716), .ZN(n390) );
  XNOR2_X1 U478 ( .A(KEYINPUT79), .B(n390), .ZN(n501) );
  INV_X1 U479 ( .A(G237), .ZN(n391) );
  NAND2_X1 U480 ( .A1(n422), .A2(n391), .ZN(n460) );
  NAND2_X1 U481 ( .A1(n460), .A2(G214), .ZN(n642) );
  NAND2_X1 U482 ( .A1(n501), .A2(n642), .ZN(n392) );
  NOR2_X1 U483 ( .A1(n544), .A2(n392), .ZN(n447) );
  XNOR2_X1 U484 ( .A(n362), .B(KEYINPUT95), .ZN(n396) );
  NAND2_X1 U485 ( .A1(G214), .A2(n394), .ZN(n395) );
  XNOR2_X1 U486 ( .A(n396), .B(n395), .ZN(n400) );
  XOR2_X1 U487 ( .A(KEYINPUT11), .B(KEYINPUT96), .Z(n398) );
  XNOR2_X1 U488 ( .A(KEYINPUT94), .B(KEYINPUT12), .ZN(n397) );
  XNOR2_X1 U489 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U490 ( .A(n400), .B(n399), .Z(n408) );
  XOR2_X1 U491 ( .A(KEYINPUT68), .B(KEYINPUT10), .Z(n403) );
  INV_X1 U492 ( .A(G146), .ZN(n401) );
  XNOR2_X1 U493 ( .A(n401), .B(G125), .ZN(n454) );
  XNOR2_X1 U494 ( .A(n454), .B(G140), .ZN(n402) );
  XNOR2_X1 U495 ( .A(n403), .B(n402), .ZN(n708) );
  XOR2_X1 U496 ( .A(G122), .B(G104), .Z(n405) );
  XNOR2_X1 U497 ( .A(G143), .B(G113), .ZN(n404) );
  XNOR2_X1 U498 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U499 ( .A(n708), .B(n406), .ZN(n407) );
  XNOR2_X1 U500 ( .A(n408), .B(n407), .ZN(n591) );
  NOR2_X1 U501 ( .A1(n591), .A2(G902), .ZN(n410) );
  XNOR2_X1 U502 ( .A(KEYINPUT13), .B(G475), .ZN(n409) );
  XNOR2_X1 U503 ( .A(n410), .B(n409), .ZN(n514) );
  XOR2_X1 U504 ( .A(KEYINPUT97), .B(n514), .Z(n507) );
  XOR2_X1 U505 ( .A(G122), .B(G107), .Z(n412) );
  XNOR2_X1 U506 ( .A(G116), .B(G134), .ZN(n411) );
  XNOR2_X1 U507 ( .A(n412), .B(n411), .ZN(n416) );
  XOR2_X1 U508 ( .A(KEYINPUT98), .B(KEYINPUT99), .Z(n414) );
  XNOR2_X1 U509 ( .A(KEYINPUT9), .B(KEYINPUT7), .ZN(n413) );
  XNOR2_X1 U510 ( .A(n414), .B(n413), .ZN(n415) );
  XOR2_X1 U511 ( .A(n416), .B(n415), .Z(n419) );
  NAND2_X1 U512 ( .A1(n701), .A2(G234), .ZN(n417) );
  XOR2_X1 U513 ( .A(KEYINPUT8), .B(n417), .Z(n432) );
  NAND2_X1 U514 ( .A1(G217), .A2(n432), .ZN(n418) );
  XNOR2_X1 U515 ( .A(n419), .B(n418), .ZN(n421) );
  XNOR2_X1 U516 ( .A(n421), .B(n420), .ZN(n583) );
  NAND2_X1 U517 ( .A1(n583), .A2(n422), .ZN(n423) );
  XNOR2_X1 U518 ( .A(n423), .B(G478), .ZN(n513) );
  INV_X1 U519 ( .A(n513), .ZN(n424) );
  NAND2_X1 U520 ( .A1(n507), .A2(n424), .ZN(n681) );
  XOR2_X1 U521 ( .A(KEYINPUT24), .B(G110), .Z(n426) );
  XNOR2_X1 U522 ( .A(n426), .B(n425), .ZN(n431) );
  XOR2_X1 U523 ( .A(KEYINPUT23), .B(KEYINPUT81), .Z(n429) );
  XNOR2_X1 U524 ( .A(n427), .B(KEYINPUT89), .ZN(n428) );
  XNOR2_X1 U525 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U526 ( .A(n431), .B(n430), .Z(n435) );
  NAND2_X1 U527 ( .A1(G221), .A2(n432), .ZN(n433) );
  XNOR2_X1 U528 ( .A(n435), .B(n434), .ZN(n587) );
  NOR2_X1 U529 ( .A1(G902), .A2(n587), .ZN(n442) );
  XNOR2_X1 U530 ( .A(KEYINPUT15), .B(G902), .ZN(n582) );
  NAND2_X1 U531 ( .A1(n582), .A2(G234), .ZN(n437) );
  XNOR2_X1 U532 ( .A(KEYINPUT20), .B(KEYINPUT90), .ZN(n436) );
  XNOR2_X1 U533 ( .A(n437), .B(n436), .ZN(n443) );
  NAND2_X1 U534 ( .A1(n443), .A2(G217), .ZN(n438) );
  XOR2_X1 U535 ( .A(KEYINPUT25), .B(n438), .Z(n440) );
  XNOR2_X1 U536 ( .A(KEYINPUT91), .B(KEYINPUT77), .ZN(n439) );
  NAND2_X1 U537 ( .A1(n443), .A2(G221), .ZN(n445) );
  INV_X1 U538 ( .A(KEYINPUT21), .ZN(n444) );
  XNOR2_X1 U539 ( .A(n445), .B(n444), .ZN(n630) );
  NAND2_X1 U540 ( .A1(n494), .A2(n630), .ZN(n485) );
  NOR2_X1 U541 ( .A1(n681), .A2(n485), .ZN(n446) );
  NAND2_X1 U542 ( .A1(n447), .A2(n446), .ZN(n510) );
  OR2_X1 U543 ( .A1(n627), .A2(n510), .ZN(n448) );
  XNOR2_X1 U544 ( .A(KEYINPUT43), .B(n448), .ZN(n464) );
  XNOR2_X1 U545 ( .A(KEYINPUT16), .B(G122), .ZN(n449) );
  NAND2_X1 U546 ( .A1(n701), .A2(G224), .ZN(n451) );
  XNOR2_X1 U547 ( .A(n451), .B(KEYINPUT88), .ZN(n453) );
  XNOR2_X1 U548 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n452) );
  XNOR2_X1 U549 ( .A(n453), .B(n452), .ZN(n455) );
  XNOR2_X1 U550 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U551 ( .A(n458), .B(n457), .ZN(n597) );
  INV_X1 U552 ( .A(n597), .ZN(n459) );
  NAND2_X1 U553 ( .A1(n459), .A2(n582), .ZN(n463) );
  NAND2_X1 U554 ( .A1(n460), .A2(G210), .ZN(n461) );
  XNOR2_X1 U555 ( .A(n461), .B(KEYINPUT78), .ZN(n462) );
  XNOR2_X1 U556 ( .A(n463), .B(n462), .ZN(n466) );
  AND2_X1 U557 ( .A1(n464), .A2(n517), .ZN(n530) );
  XOR2_X1 U558 ( .A(n530), .B(G140), .Z(G42) );
  INV_X1 U559 ( .A(n642), .ZN(n465) );
  NAND2_X1 U560 ( .A1(G953), .A2(G898), .ZN(n468) );
  XNOR2_X2 U561 ( .A(n470), .B(KEYINPUT0), .ZN(n564) );
  NOR2_X1 U562 ( .A1(n514), .A2(n513), .ZN(n481) );
  NAND2_X1 U563 ( .A1(n481), .A2(n630), .ZN(n471) );
  NOR2_X1 U564 ( .A1(n627), .A2(n637), .ZN(n473) );
  NAND2_X1 U565 ( .A1(n476), .A2(n473), .ZN(n474) );
  XOR2_X1 U566 ( .A(KEYINPUT66), .B(n474), .Z(n475) );
  NAND2_X1 U567 ( .A1(n475), .A2(n494), .ZN(n539) );
  XNOR2_X1 U568 ( .A(n539), .B(G110), .ZN(G12) );
  NAND2_X1 U569 ( .A1(n476), .A2(n544), .ZN(n536) );
  XNOR2_X1 U570 ( .A(n536), .B(KEYINPUT84), .ZN(n479) );
  XOR2_X1 U571 ( .A(KEYINPUT100), .B(n494), .Z(n631) );
  INV_X1 U572 ( .A(n627), .ZN(n477) );
  NAND2_X1 U573 ( .A1(n631), .A2(n477), .ZN(n478) );
  NOR2_X1 U574 ( .A1(n479), .A2(n478), .ZN(n567) );
  XOR2_X1 U575 ( .A(G101), .B(n567), .Z(G3) );
  XNOR2_X1 U576 ( .A(KEYINPUT74), .B(KEYINPUT38), .ZN(n480) );
  XOR2_X1 U577 ( .A(n480), .B(n517), .Z(n502) );
  INV_X1 U578 ( .A(n502), .ZN(n643) );
  NAND2_X1 U579 ( .A1(n643), .A2(n642), .ZN(n646) );
  INV_X1 U580 ( .A(n481), .ZN(n645) );
  NOR2_X1 U581 ( .A1(n646), .A2(n645), .ZN(n483) );
  XNOR2_X1 U582 ( .A(KEYINPUT106), .B(KEYINPUT41), .ZN(n482) );
  NAND2_X1 U583 ( .A1(n496), .A2(n501), .ZN(n484) );
  XNOR2_X1 U584 ( .A(n486), .B(KEYINPUT105), .ZN(n487) );
  XNOR2_X1 U585 ( .A(n487), .B(KEYINPUT28), .ZN(n490) );
  XNOR2_X1 U586 ( .A(n488), .B(KEYINPUT104), .ZN(n489) );
  NAND2_X1 U587 ( .A1(n490), .A2(n489), .ZN(n506) );
  NOR2_X1 U588 ( .A1(n626), .A2(n506), .ZN(n493) );
  INV_X1 U589 ( .A(KEYINPUT42), .ZN(n491) );
  INV_X1 U590 ( .A(n630), .ZN(n495) );
  NOR2_X1 U591 ( .A1(n495), .A2(n494), .ZN(n540) );
  NAND2_X1 U592 ( .A1(n488), .A2(n540), .ZN(n562) );
  NAND2_X1 U593 ( .A1(n642), .A2(n496), .ZN(n498) );
  NOR2_X1 U594 ( .A1(n562), .A2(n499), .ZN(n500) );
  NAND2_X1 U595 ( .A1(n501), .A2(n500), .ZN(n518) );
  NOR2_X1 U596 ( .A1(n518), .A2(n502), .ZN(n503) );
  XNOR2_X1 U597 ( .A(n503), .B(KEYINPUT39), .ZN(n529) );
  NOR2_X1 U598 ( .A1(n681), .A2(n529), .ZN(n504) );
  XNOR2_X1 U599 ( .A(KEYINPUT40), .B(n504), .ZN(n722) );
  XNOR2_X1 U600 ( .A(n505), .B(KEYINPUT46), .ZN(n527) );
  INV_X1 U601 ( .A(n507), .ZN(n508) );
  NAND2_X1 U602 ( .A1(n508), .A2(n513), .ZN(n674) );
  AND2_X1 U603 ( .A1(n674), .A2(n681), .ZN(n647) );
  XOR2_X1 U604 ( .A(n509), .B(KEYINPUT47), .Z(n523) );
  NOR2_X1 U605 ( .A1(n510), .A2(n517), .ZN(n511) );
  XNOR2_X1 U606 ( .A(n511), .B(KEYINPUT36), .ZN(n512) );
  NAND2_X1 U607 ( .A1(n512), .A2(n627), .ZN(n690) );
  NAND2_X1 U608 ( .A1(n514), .A2(n513), .ZN(n516) );
  INV_X1 U609 ( .A(KEYINPUT101), .ZN(n515) );
  XNOR2_X1 U610 ( .A(n516), .B(n515), .ZN(n548) );
  NOR2_X1 U611 ( .A1(n518), .A2(n517), .ZN(n519) );
  XNOR2_X1 U612 ( .A(n519), .B(KEYINPUT103), .ZN(n520) );
  NOR2_X1 U613 ( .A1(n548), .A2(n520), .ZN(n679) );
  INV_X1 U614 ( .A(n679), .ZN(n521) );
  NAND2_X1 U615 ( .A1(n690), .A2(n521), .ZN(n522) );
  NOR2_X1 U616 ( .A1(n523), .A2(n522), .ZN(n525) );
  XNOR2_X1 U617 ( .A(n528), .B(KEYINPUT48), .ZN(n532) );
  NOR2_X1 U618 ( .A1(n674), .A2(n529), .ZN(n691) );
  NOR2_X1 U619 ( .A1(n691), .A2(n530), .ZN(n531) );
  NAND2_X1 U620 ( .A1(n532), .A2(n531), .ZN(n712) );
  INV_X1 U621 ( .A(n631), .ZN(n534) );
  NAND2_X1 U622 ( .A1(n534), .A2(n627), .ZN(n535) );
  NAND2_X1 U623 ( .A1(n614), .A2(n539), .ZN(n553) );
  INV_X1 U624 ( .A(n553), .ZN(n551) );
  NAND2_X1 U625 ( .A1(n541), .A2(n540), .ZN(n543) );
  NOR2_X1 U626 ( .A1(n558), .A2(n544), .ZN(n547) );
  INV_X1 U627 ( .A(KEYINPUT87), .ZN(n545) );
  XNOR2_X1 U628 ( .A(n545), .B(KEYINPUT33), .ZN(n546) );
  XNOR2_X1 U629 ( .A(n547), .B(n546), .ZN(n650) );
  NOR2_X1 U630 ( .A1(KEYINPUT44), .A2(KEYINPUT85), .ZN(n549) );
  NAND2_X1 U631 ( .A1(n568), .A2(n549), .ZN(n550) );
  NAND2_X1 U632 ( .A1(n551), .A2(n550), .ZN(n556) );
  NOR2_X1 U633 ( .A1(n552), .A2(KEYINPUT44), .ZN(n554) );
  NAND2_X1 U634 ( .A1(n554), .A2(n553), .ZN(n555) );
  NAND2_X1 U635 ( .A1(n556), .A2(n555), .ZN(n573) );
  INV_X1 U636 ( .A(n637), .ZN(n557) );
  NOR2_X1 U637 ( .A1(n558), .A2(n557), .ZN(n639) );
  INV_X1 U638 ( .A(n564), .ZN(n559) );
  NAND2_X1 U639 ( .A1(n639), .A2(n559), .ZN(n561) );
  XOR2_X1 U640 ( .A(KEYINPUT31), .B(KEYINPUT93), .Z(n560) );
  XNOR2_X1 U641 ( .A(n561), .B(n560), .ZN(n687) );
  OR2_X1 U642 ( .A1(n562), .A2(n637), .ZN(n563) );
  NOR2_X1 U643 ( .A1(n564), .A2(n563), .ZN(n670) );
  NOR2_X1 U644 ( .A1(n687), .A2(n670), .ZN(n565) );
  NOR2_X1 U645 ( .A1(n565), .A2(n647), .ZN(n566) );
  NOR2_X1 U646 ( .A1(n567), .A2(n566), .ZN(n571) );
  INV_X1 U647 ( .A(n568), .ZN(n569) );
  NAND2_X1 U648 ( .A1(n569), .A2(KEYINPUT44), .ZN(n570) );
  AND2_X1 U649 ( .A1(n571), .A2(n570), .ZN(n572) );
  NAND2_X1 U650 ( .A1(n573), .A2(n572), .ZN(n575) );
  XNOR2_X1 U651 ( .A(KEYINPUT82), .B(KEYINPUT45), .ZN(n574) );
  XNOR2_X2 U652 ( .A(n575), .B(n574), .ZN(n692) );
  NAND2_X1 U653 ( .A1(n578), .A2(n577), .ZN(n581) );
  INV_X1 U654 ( .A(n712), .ZN(n579) );
  NAND2_X1 U655 ( .A1(n692), .A2(n579), .ZN(n624) );
  NAND2_X1 U656 ( .A1(n624), .A2(KEYINPUT2), .ZN(n580) );
  INV_X1 U657 ( .A(n582), .ZN(n615) );
  NAND2_X1 U658 ( .A1(n348), .A2(G478), .ZN(n585) );
  XNOR2_X1 U659 ( .A(n583), .B(KEYINPUT121), .ZN(n584) );
  XNOR2_X1 U660 ( .A(n585), .B(n584), .ZN(n586) );
  NOR2_X1 U661 ( .A1(n586), .A2(n621), .ZN(G63) );
  NAND2_X1 U662 ( .A1(n348), .A2(G217), .ZN(n589) );
  XNOR2_X1 U663 ( .A(n587), .B(KEYINPUT122), .ZN(n588) );
  XNOR2_X1 U664 ( .A(n589), .B(n588), .ZN(n590) );
  NOR2_X1 U665 ( .A1(n590), .A2(n621), .ZN(G66) );
  XOR2_X1 U666 ( .A(KEYINPUT59), .B(n591), .Z(n592) );
  XNOR2_X1 U667 ( .A(n593), .B(n592), .ZN(n594) );
  XOR2_X1 U668 ( .A(KEYINPUT67), .B(KEYINPUT60), .Z(n595) );
  XNOR2_X1 U669 ( .A(n596), .B(n595), .ZN(G60) );
  XOR2_X1 U670 ( .A(KEYINPUT86), .B(KEYINPUT54), .Z(n598) );
  XNOR2_X1 U671 ( .A(n598), .B(KEYINPUT55), .ZN(n599) );
  XNOR2_X1 U672 ( .A(n597), .B(n599), .ZN(n600) );
  XNOR2_X1 U673 ( .A(n601), .B(n600), .ZN(n602) );
  XOR2_X1 U674 ( .A(KEYINPUT83), .B(KEYINPUT56), .Z(n603) );
  XNOR2_X1 U675 ( .A(n604), .B(n603), .ZN(G51) );
  XOR2_X1 U676 ( .A(KEYINPUT118), .B(KEYINPUT57), .Z(n606) );
  XNOR2_X1 U677 ( .A(n606), .B(KEYINPUT58), .ZN(n608) );
  XOR2_X1 U678 ( .A(KEYINPUT117), .B(KEYINPUT119), .Z(n607) );
  XNOR2_X1 U679 ( .A(n608), .B(n607), .ZN(n609) );
  XNOR2_X1 U680 ( .A(n605), .B(n609), .ZN(n610) );
  XNOR2_X1 U681 ( .A(n611), .B(n610), .ZN(n612) );
  XNOR2_X1 U682 ( .A(n613), .B(KEYINPUT120), .ZN(G54) );
  XNOR2_X1 U683 ( .A(n614), .B(G119), .ZN(G21) );
  AND2_X1 U684 ( .A1(G472), .A2(n615), .ZN(n616) );
  NAND2_X1 U685 ( .A1(n617), .A2(n616), .ZN(n620) );
  XOR2_X1 U686 ( .A(n618), .B(KEYINPUT62), .Z(n619) );
  XNOR2_X1 U687 ( .A(n620), .B(n619), .ZN(n622) );
  NOR2_X1 U688 ( .A1(n622), .A2(n621), .ZN(n623) );
  XNOR2_X1 U689 ( .A(n568), .B(G122), .ZN(G24) );
  NAND2_X1 U690 ( .A1(n624), .A2(KEYINPUT80), .ZN(n625) );
  XOR2_X1 U691 ( .A(KEYINPUT2), .B(n625), .Z(n664) );
  NOR2_X1 U692 ( .A1(n540), .A2(n627), .ZN(n629) );
  XNOR2_X1 U693 ( .A(KEYINPUT115), .B(KEYINPUT50), .ZN(n628) );
  XNOR2_X1 U694 ( .A(n629), .B(n628), .ZN(n635) );
  NOR2_X1 U695 ( .A1(n631), .A2(n630), .ZN(n633) );
  XNOR2_X1 U696 ( .A(KEYINPUT49), .B(KEYINPUT114), .ZN(n632) );
  XNOR2_X1 U697 ( .A(n633), .B(n632), .ZN(n634) );
  NAND2_X1 U698 ( .A1(n635), .A2(n634), .ZN(n636) );
  NOR2_X1 U699 ( .A1(n637), .A2(n636), .ZN(n638) );
  NOR2_X1 U700 ( .A1(n639), .A2(n638), .ZN(n640) );
  XOR2_X1 U701 ( .A(KEYINPUT51), .B(n640), .Z(n641) );
  NOR2_X1 U702 ( .A1(n626), .A2(n641), .ZN(n654) );
  NOR2_X1 U703 ( .A1(n643), .A2(n642), .ZN(n644) );
  NOR2_X1 U704 ( .A1(n645), .A2(n644), .ZN(n649) );
  NOR2_X1 U705 ( .A1(n647), .A2(n646), .ZN(n648) );
  NOR2_X1 U706 ( .A1(n649), .A2(n648), .ZN(n652) );
  BUF_X1 U707 ( .A(n650), .Z(n651) );
  NOR2_X1 U708 ( .A1(n652), .A2(n651), .ZN(n653) );
  NOR2_X1 U709 ( .A1(n654), .A2(n653), .ZN(n655) );
  XNOR2_X1 U710 ( .A(KEYINPUT52), .B(n655), .ZN(n658) );
  NAND2_X1 U711 ( .A1(G952), .A2(n656), .ZN(n657) );
  NOR2_X1 U712 ( .A1(n658), .A2(n657), .ZN(n659) );
  NOR2_X1 U713 ( .A1(n659), .A2(G953), .ZN(n662) );
  NOR2_X1 U714 ( .A1(n651), .A2(n626), .ZN(n660) );
  XOR2_X1 U715 ( .A(KEYINPUT116), .B(n660), .Z(n661) );
  NAND2_X1 U716 ( .A1(n662), .A2(n661), .ZN(n663) );
  NOR2_X1 U717 ( .A1(n664), .A2(n663), .ZN(n665) );
  XNOR2_X1 U718 ( .A(n665), .B(KEYINPUT53), .ZN(G75) );
  INV_X1 U719 ( .A(n681), .ZN(n684) );
  NAND2_X1 U720 ( .A1(n670), .A2(n684), .ZN(n666) );
  XNOR2_X1 U721 ( .A(n666), .B(G104), .ZN(G6) );
  XOR2_X1 U722 ( .A(KEYINPUT27), .B(KEYINPUT109), .Z(n668) );
  XNOR2_X1 U723 ( .A(G107), .B(KEYINPUT108), .ZN(n667) );
  XNOR2_X1 U724 ( .A(n668), .B(n667), .ZN(n669) );
  XOR2_X1 U725 ( .A(KEYINPUT26), .B(n669), .Z(n672) );
  INV_X1 U726 ( .A(n674), .ZN(n686) );
  NAND2_X1 U727 ( .A1(n670), .A2(n686), .ZN(n671) );
  XNOR2_X1 U728 ( .A(n672), .B(n671), .ZN(G9) );
  NOR2_X1 U729 ( .A1(n673), .A2(n674), .ZN(n678) );
  XOR2_X1 U730 ( .A(KEYINPUT110), .B(KEYINPUT29), .Z(n676) );
  XNOR2_X1 U731 ( .A(G128), .B(KEYINPUT111), .ZN(n675) );
  XNOR2_X1 U732 ( .A(n676), .B(n675), .ZN(n677) );
  XNOR2_X1 U733 ( .A(n678), .B(n677), .ZN(G30) );
  XOR2_X1 U734 ( .A(G143), .B(n679), .Z(n680) );
  XNOR2_X1 U735 ( .A(KEYINPUT112), .B(n680), .ZN(G45) );
  NOR2_X1 U736 ( .A1(n673), .A2(n681), .ZN(n683) );
  XNOR2_X1 U737 ( .A(G146), .B(KEYINPUT113), .ZN(n682) );
  XNOR2_X1 U738 ( .A(n683), .B(n682), .ZN(G48) );
  NAND2_X1 U739 ( .A1(n687), .A2(n684), .ZN(n685) );
  XNOR2_X1 U740 ( .A(n685), .B(G113), .ZN(G15) );
  NAND2_X1 U741 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U742 ( .A(n688), .B(G116), .ZN(G18) );
  XOR2_X1 U743 ( .A(G125), .B(KEYINPUT37), .Z(n689) );
  XNOR2_X1 U744 ( .A(n690), .B(n689), .ZN(G27) );
  XOR2_X1 U745 ( .A(G134), .B(n691), .Z(G36) );
  NAND2_X1 U746 ( .A1(n692), .A2(n701), .ZN(n697) );
  XOR2_X1 U747 ( .A(KEYINPUT123), .B(KEYINPUT61), .Z(n694) );
  NAND2_X1 U748 ( .A1(G224), .A2(G953), .ZN(n693) );
  XNOR2_X1 U749 ( .A(n694), .B(n693), .ZN(n695) );
  NAND2_X1 U750 ( .A1(n695), .A2(G898), .ZN(n696) );
  NAND2_X1 U751 ( .A1(n697), .A2(n696), .ZN(n706) );
  XNOR2_X1 U752 ( .A(n698), .B(G101), .ZN(n699) );
  XNOR2_X1 U753 ( .A(n700), .B(n699), .ZN(n703) );
  NOR2_X1 U754 ( .A1(G898), .A2(n701), .ZN(n702) );
  NOR2_X1 U755 ( .A1(n703), .A2(n702), .ZN(n704) );
  XOR2_X1 U756 ( .A(KEYINPUT124), .B(n704), .Z(n705) );
  XNOR2_X1 U757 ( .A(n706), .B(n705), .ZN(n707) );
  XNOR2_X1 U758 ( .A(KEYINPUT125), .B(n707), .ZN(G69) );
  XNOR2_X1 U759 ( .A(n709), .B(n708), .ZN(n711) );
  XNOR2_X1 U760 ( .A(n711), .B(n710), .ZN(n714) );
  XOR2_X1 U761 ( .A(n714), .B(n712), .Z(n713) );
  NOR2_X1 U762 ( .A1(G953), .A2(n713), .ZN(n719) );
  XNOR2_X1 U763 ( .A(n714), .B(KEYINPUT126), .ZN(n715) );
  XNOR2_X1 U764 ( .A(G227), .B(n715), .ZN(n717) );
  NOR2_X1 U765 ( .A1(n717), .A2(n716), .ZN(n718) );
  NOR2_X1 U766 ( .A1(n719), .A2(n718), .ZN(n720) );
  XOR2_X1 U767 ( .A(KEYINPUT127), .B(n720), .Z(G72) );
  XOR2_X1 U768 ( .A(n721), .B(G137), .Z(G39) );
  XOR2_X1 U769 ( .A(G131), .B(n722), .Z(G33) );
endmodule

