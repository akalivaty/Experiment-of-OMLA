//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 0 1 1 0 0 0 0 1 0 0 1 0 0 0 1 0 0 1 0 0 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 1 0 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:16 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n559, new_n560, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n588,
    new_n589, new_n590, new_n591, new_n594, new_n595, new_n596, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n629, new_n631, new_n632, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1188, new_n1189;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT65), .B(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g018(.A(KEYINPUT66), .B(G452), .ZN(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n446));
  AND2_X1   g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND2_X1  g023(.A1(new_n447), .A2(G567), .ZN(G234));
  NAND2_X1  g024(.A1(new_n447), .A2(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OAI22_X1  g032(.A1(new_n452), .A2(new_n456), .B1(new_n457), .B2(new_n453), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  AND2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  OAI21_X1  g037(.A(G125), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n460), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  OAI211_X1 g040(.A(G137), .B(new_n460), .C1(new_n461), .C2(new_n462), .ZN(new_n466));
  AND2_X1   g041(.A1(new_n460), .A2(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G101), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n465), .A2(new_n469), .ZN(G160));
  XNOR2_X1  g045(.A(KEYINPUT3), .B(G2104), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT68), .ZN(new_n472));
  XNOR2_X1  g047(.A(new_n471), .B(new_n472), .ZN(new_n473));
  AND2_X1   g048(.A1(new_n473), .A2(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G124), .ZN(new_n475));
  XNOR2_X1  g050(.A(new_n475), .B(KEYINPUT69), .ZN(new_n476));
  OAI21_X1  g051(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n477));
  INV_X1    g052(.A(G112), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n477), .B1(new_n478), .B2(G2105), .ZN(new_n479));
  AND2_X1   g054(.A1(new_n473), .A2(new_n460), .ZN(new_n480));
  AND2_X1   g055(.A1(new_n480), .A2(G136), .ZN(new_n481));
  NOR3_X1   g056(.A1(new_n476), .A2(new_n479), .A3(new_n481), .ZN(G162));
  NAND3_X1  g057(.A1(new_n471), .A2(G126), .A3(G2105), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT71), .ZN(new_n484));
  OAI21_X1  g059(.A(KEYINPUT70), .B1(new_n460), .B2(G114), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT70), .ZN(new_n486));
  INV_X1    g061(.A(G114), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n486), .A2(new_n487), .A3(G2105), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n485), .A2(new_n488), .ZN(new_n489));
  OAI21_X1  g064(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n484), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  AOI211_X1 g067(.A(KEYINPUT71), .B(new_n490), .C1(new_n485), .C2(new_n488), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n483), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT72), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  OAI211_X1 g071(.A(G138), .B(new_n460), .C1(new_n461), .C2(new_n462), .ZN(new_n497));
  XNOR2_X1  g072(.A(new_n497), .B(KEYINPUT4), .ZN(new_n498));
  OAI211_X1 g073(.A(KEYINPUT72), .B(new_n483), .C1(new_n492), .C2(new_n493), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n496), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(G164));
  INV_X1    g076(.A(KEYINPUT73), .ZN(new_n502));
  INV_X1    g077(.A(G651), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n502), .B1(new_n503), .B2(KEYINPUT6), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT6), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n505), .A2(KEYINPUT73), .A3(G651), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n503), .A2(KEYINPUT6), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT5), .ZN(new_n510));
  INV_X1    g085(.A(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(KEYINPUT5), .A2(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(new_n514), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n509), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G88), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n507), .A2(G543), .A3(new_n508), .ZN(new_n518));
  INV_X1    g093(.A(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G50), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n514), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n521));
  OR2_X1    g096(.A1(new_n521), .A2(new_n503), .ZN(new_n522));
  AND3_X1   g097(.A1(new_n517), .A2(new_n520), .A3(new_n522), .ZN(G166));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  XOR2_X1   g099(.A(new_n524), .B(KEYINPUT7), .Z(new_n525));
  NAND2_X1  g100(.A1(G63), .A2(G651), .ZN(new_n526));
  INV_X1    g101(.A(G89), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n526), .B1(new_n509), .B2(new_n527), .ZN(new_n528));
  AOI21_X1  g103(.A(new_n525), .B1(new_n528), .B2(new_n514), .ZN(new_n529));
  INV_X1    g104(.A(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(G51), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n518), .A2(KEYINPUT74), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT74), .ZN(new_n533));
  NAND4_X1  g108(.A1(new_n507), .A2(new_n533), .A3(G543), .A4(new_n508), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n531), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n530), .A2(new_n535), .ZN(G168));
  NAND2_X1  g111(.A1(new_n532), .A2(new_n534), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G52), .ZN(new_n538));
  NAND2_X1  g113(.A1(G77), .A2(G543), .ZN(new_n539));
  INV_X1    g114(.A(G64), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n539), .B1(new_n515), .B2(new_n540), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n516), .A2(G90), .B1(new_n541), .B2(G651), .ZN(new_n542));
  AND2_X1   g117(.A1(new_n538), .A2(new_n542), .ZN(G171));
  NAND2_X1  g118(.A1(new_n537), .A2(G43), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT75), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n516), .A2(G81), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(new_n546), .ZN(new_n548));
  INV_X1    g123(.A(G43), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n549), .B1(new_n532), .B2(new_n534), .ZN(new_n550));
  OAI21_X1  g125(.A(KEYINPUT75), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n547), .A2(new_n551), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n514), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n553));
  OR2_X1    g128(.A1(new_n553), .A2(new_n503), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(G153));
  NAND4_X1  g132(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND4_X1  g135(.A1(G319), .A2(G483), .A3(G661), .A4(new_n560), .ZN(G188));
  INV_X1    g136(.A(KEYINPUT80), .ZN(new_n562));
  INV_X1    g137(.A(G65), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT78), .ZN(new_n564));
  INV_X1    g139(.A(new_n513), .ZN(new_n565));
  NOR2_X1   g140(.A1(KEYINPUT5), .A2(G543), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n564), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n512), .A2(KEYINPUT78), .A3(new_n513), .ZN(new_n568));
  AOI21_X1  g143(.A(new_n563), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(G78), .A2(G543), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT77), .ZN(new_n571));
  OAI21_X1  g146(.A(G651), .B1(new_n569), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(KEYINPUT79), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT79), .ZN(new_n574));
  OAI211_X1 g149(.A(new_n574), .B(G651), .C1(new_n569), .C2(new_n571), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(KEYINPUT76), .A2(KEYINPUT9), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n519), .A2(G53), .A3(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(G53), .ZN(new_n579));
  OAI211_X1 g154(.A(KEYINPUT76), .B(KEYINPUT9), .C1(new_n518), .C2(new_n579), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n578), .A2(new_n580), .B1(G91), .B2(new_n516), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n562), .B1(new_n576), .B2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(new_n582), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n576), .A2(new_n581), .A3(new_n562), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(G299));
  INV_X1    g161(.A(G171), .ZN(G301));
  NOR3_X1   g162(.A1(new_n530), .A2(new_n535), .A3(KEYINPUT81), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT81), .ZN(new_n589));
  INV_X1    g164(.A(new_n535), .ZN(new_n590));
  AOI21_X1  g165(.A(new_n589), .B1(new_n590), .B2(new_n529), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n588), .A2(new_n591), .ZN(G286));
  NAND3_X1  g167(.A1(new_n517), .A2(new_n520), .A3(new_n522), .ZN(G303));
  NAND4_X1  g168(.A1(new_n507), .A2(G87), .A3(new_n508), .A4(new_n514), .ZN(new_n594));
  OAI21_X1  g169(.A(G651), .B1(new_n514), .B2(G74), .ZN(new_n595));
  INV_X1    g170(.A(G49), .ZN(new_n596));
  OAI211_X1 g171(.A(new_n594), .B(new_n595), .C1(new_n518), .C2(new_n596), .ZN(G288));
  INV_X1    g172(.A(G61), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n598), .B1(new_n512), .B2(new_n513), .ZN(new_n599));
  AND2_X1   g174(.A1(G73), .A2(G543), .ZN(new_n600));
  OAI21_X1  g175(.A(G651), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND4_X1  g176(.A1(new_n507), .A2(G48), .A3(G543), .A4(new_n508), .ZN(new_n602));
  NAND4_X1  g177(.A1(new_n507), .A2(G86), .A3(new_n508), .A4(new_n514), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(G305));
  XOR2_X1   g179(.A(KEYINPUT82), .B(G47), .Z(new_n605));
  NAND2_X1  g180(.A1(new_n537), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(G72), .A2(G543), .ZN(new_n607));
  INV_X1    g182(.A(G60), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n515), .B2(new_n608), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n516), .A2(G85), .B1(new_n609), .B2(G651), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n606), .A2(new_n610), .ZN(G290));
  NAND2_X1  g186(.A1(G301), .A2(G868), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n516), .A2(G92), .ZN(new_n613));
  INV_X1    g188(.A(KEYINPUT10), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n613), .B(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n537), .A2(G54), .ZN(new_n616));
  NAND2_X1  g191(.A1(G79), .A2(G543), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT83), .ZN(new_n618));
  AND2_X1   g193(.A1(new_n567), .A2(new_n568), .ZN(new_n619));
  INV_X1    g194(.A(G66), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n618), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n621), .A2(G651), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n615), .A2(new_n616), .A3(new_n622), .ZN(new_n623));
  INV_X1    g198(.A(new_n623), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n612), .B1(new_n624), .B2(G868), .ZN(G321));
  XOR2_X1   g200(.A(G321), .B(KEYINPUT84), .Z(G284));
  MUX2_X1   g201(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g202(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g203(.A(G559), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n624), .B1(new_n629), .B2(G860), .ZN(G148));
  NAND2_X1  g205(.A1(new_n624), .A2(new_n629), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n631), .A2(G868), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n632), .B1(G868), .B2(new_n556), .ZN(G323));
  XNOR2_X1  g208(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OAI21_X1  g209(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n635));
  INV_X1    g210(.A(G111), .ZN(new_n636));
  AOI21_X1  g211(.A(new_n635), .B1(new_n636), .B2(G2105), .ZN(new_n637));
  AOI21_X1  g212(.A(new_n637), .B1(new_n480), .B2(G135), .ZN(new_n638));
  AND3_X1   g213(.A1(new_n474), .A2(KEYINPUT85), .A3(G123), .ZN(new_n639));
  AOI21_X1  g214(.A(KEYINPUT85), .B1(new_n474), .B2(G123), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n638), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n641), .A2(G2096), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n641), .A2(G2096), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n471), .A2(new_n467), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT12), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT13), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(G2100), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n642), .A2(new_n643), .A3(new_n647), .ZN(G156));
  INV_X1    g223(.A(KEYINPUT14), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2427), .B(G2438), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(G2430), .ZN(new_n651));
  XNOR2_X1  g226(.A(KEYINPUT15), .B(G2435), .ZN(new_n652));
  AOI21_X1  g227(.A(new_n649), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n653), .B1(new_n652), .B2(new_n651), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2451), .B(G2454), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT16), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1341), .B(G1348), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n654), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2443), .B(G2446), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n659), .A2(new_n660), .ZN(new_n662));
  AND3_X1   g237(.A1(new_n661), .A2(G14), .A3(new_n662), .ZN(G401));
  INV_X1    g238(.A(KEYINPUT18), .ZN(new_n664));
  XOR2_X1   g239(.A(G2084), .B(G2090), .Z(new_n665));
  XNOR2_X1  g240(.A(G2067), .B(G2678), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n667), .A2(KEYINPUT17), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n665), .A2(new_n666), .ZN(new_n669));
  OAI21_X1  g244(.A(new_n664), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(KEYINPUT86), .B(G2100), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(G2072), .B(G2078), .Z(new_n673));
  AOI21_X1  g248(.A(new_n673), .B1(new_n667), .B2(KEYINPUT18), .ZN(new_n674));
  XOR2_X1   g249(.A(new_n674), .B(G2096), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n672), .B(new_n675), .ZN(G227));
  XNOR2_X1  g251(.A(G1971), .B(G1976), .ZN(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT87), .B(KEYINPUT19), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1956), .B(G2474), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1961), .B(G1966), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT20), .ZN(new_n684));
  INV_X1    g259(.A(new_n679), .ZN(new_n685));
  INV_X1    g260(.A(new_n682), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n680), .A2(new_n681), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n685), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  OAI211_X1 g263(.A(new_n684), .B(new_n688), .C1(new_n685), .C2(new_n687), .ZN(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1991), .B(G1996), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1981), .B(G1986), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(G229));
  NAND2_X1  g270(.A1(G162), .A2(G29), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n696), .B1(G29), .B2(G35), .ZN(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT98), .B(KEYINPUT29), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  XOR2_X1   g275(.A(KEYINPUT27), .B(G1996), .Z(new_n701));
  NOR2_X1   g276(.A1(G29), .A2(G32), .ZN(new_n702));
  NAND3_X1  g277(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(KEYINPUT26), .Z(new_n704));
  AND3_X1   g279(.A1(new_n467), .A2(KEYINPUT95), .A3(G105), .ZN(new_n705));
  AOI21_X1  g280(.A(KEYINPUT95), .B1(new_n467), .B2(G105), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n704), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n707), .B1(new_n480), .B2(G141), .ZN(new_n708));
  AND3_X1   g283(.A1(new_n474), .A2(KEYINPUT94), .A3(G129), .ZN(new_n709));
  AOI21_X1  g284(.A(KEYINPUT94), .B1(new_n474), .B2(G129), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n708), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT96), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n702), .B1(new_n712), .B2(G29), .ZN(new_n713));
  AOI22_X1  g288(.A1(new_n700), .A2(G2090), .B1(new_n701), .B2(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(G16), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n715), .A2(G20), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT99), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT23), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(new_n585), .B2(new_n715), .ZN(new_n719));
  INV_X1    g294(.A(G1956), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n713), .A2(new_n701), .ZN(new_n722));
  INV_X1    g297(.A(G2090), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n722), .B1(new_n699), .B2(new_n723), .ZN(new_n724));
  NAND3_X1  g299(.A1(new_n714), .A2(new_n721), .A3(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(G29), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n726), .A2(G26), .ZN(new_n727));
  XOR2_X1   g302(.A(new_n727), .B(KEYINPUT28), .Z(new_n728));
  NAND2_X1  g303(.A1(new_n480), .A2(G140), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n729), .B(KEYINPUT92), .Z(new_n730));
  OAI21_X1  g305(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n731));
  INV_X1    g306(.A(G116), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n731), .B1(new_n732), .B2(G2105), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(new_n474), .B2(G128), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n730), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n728), .B1(new_n735), .B2(G29), .ZN(new_n736));
  INV_X1    g311(.A(G2067), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n715), .A2(G21), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(G168), .B2(new_n715), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n715), .A2(G5), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(G171), .B2(new_n715), .ZN(new_n742));
  AOI22_X1  g317(.A1(G1966), .A2(new_n740), .B1(new_n742), .B2(G1961), .ZN(new_n743));
  OR2_X1    g318(.A1(new_n740), .A2(G1966), .ZN(new_n744));
  OAI211_X1 g319(.A(new_n743), .B(new_n744), .C1(G1961), .C2(new_n742), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n726), .A2(G33), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n460), .A2(G103), .A3(G2104), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(KEYINPUT25), .Z(new_n748));
  AOI22_X1  g323(.A1(new_n471), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n748), .B1(new_n749), .B2(new_n460), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(new_n480), .B2(G139), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n746), .B1(new_n751), .B2(new_n726), .ZN(new_n752));
  XOR2_X1   g327(.A(KEYINPUT93), .B(G2072), .Z(new_n753));
  XNOR2_X1  g328(.A(new_n752), .B(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(G28), .ZN(new_n755));
  OR2_X1    g330(.A1(new_n755), .A2(KEYINPUT30), .ZN(new_n756));
  AOI21_X1  g331(.A(G29), .B1(new_n755), .B2(KEYINPUT30), .ZN(new_n757));
  OR2_X1    g332(.A1(KEYINPUT31), .A2(G11), .ZN(new_n758));
  NAND2_X1  g333(.A1(KEYINPUT31), .A2(G11), .ZN(new_n759));
  AOI22_X1  g334(.A1(new_n756), .A2(new_n757), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(G34), .ZN(new_n761));
  AOI21_X1  g336(.A(G29), .B1(new_n761), .B2(KEYINPUT24), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(KEYINPUT24), .B2(new_n761), .ZN(new_n763));
  INV_X1    g338(.A(G160), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n763), .B1(new_n764), .B2(new_n726), .ZN(new_n765));
  INV_X1    g340(.A(G2084), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n760), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(new_n766), .B2(new_n765), .ZN(new_n768));
  OAI211_X1 g343(.A(new_n754), .B(new_n768), .C1(new_n726), .C2(new_n641), .ZN(new_n769));
  NOR3_X1   g344(.A1(new_n738), .A2(new_n745), .A3(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n726), .A2(G27), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT97), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(G164), .B2(new_n726), .ZN(new_n773));
  INV_X1    g348(.A(G2078), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NOR2_X1   g350(.A1(G4), .A2(G16), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(new_n624), .B2(G16), .ZN(new_n777));
  INV_X1    g352(.A(G1348), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NAND3_X1  g354(.A1(new_n770), .A2(new_n775), .A3(new_n779), .ZN(new_n780));
  NOR2_X1   g355(.A1(G16), .A2(G19), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(new_n556), .B2(G16), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(G1341), .ZN(new_n783));
  NOR3_X1   g358(.A1(new_n725), .A2(new_n780), .A3(new_n783), .ZN(new_n784));
  NOR2_X1   g359(.A1(G6), .A2(G16), .ZN(new_n785));
  AND3_X1   g360(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n785), .B1(new_n786), .B2(G16), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT32), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(G1981), .ZN(new_n789));
  NOR2_X1   g364(.A1(G16), .A2(G23), .ZN(new_n790));
  XOR2_X1   g365(.A(new_n790), .B(KEYINPUT89), .Z(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(G288), .B2(new_n715), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT33), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(G1976), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n715), .A2(G22), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT90), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(G303), .B2(G16), .ZN(new_n797));
  INV_X1    g372(.A(G1971), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  NOR3_X1   g374(.A1(new_n789), .A2(new_n794), .A3(new_n799), .ZN(new_n800));
  XNOR2_X1  g375(.A(KEYINPUT88), .B(KEYINPUT34), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n480), .A2(G131), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n474), .A2(G119), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n460), .A2(G107), .ZN(new_n805));
  OAI21_X1  g380(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n806));
  OAI211_X1 g381(.A(new_n803), .B(new_n804), .C1(new_n805), .C2(new_n806), .ZN(new_n807));
  MUX2_X1   g382(.A(G25), .B(new_n807), .S(G29), .Z(new_n808));
  XOR2_X1   g383(.A(KEYINPUT35), .B(G1991), .Z(new_n809));
  INV_X1    g384(.A(new_n809), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n808), .B(new_n810), .ZN(new_n811));
  MUX2_X1   g386(.A(G24), .B(G290), .S(G16), .Z(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(G1986), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  AND3_X1   g389(.A1(new_n802), .A2(KEYINPUT91), .A3(new_n814), .ZN(new_n815));
  AOI21_X1  g390(.A(KEYINPUT91), .B1(new_n802), .B2(new_n814), .ZN(new_n816));
  OAI22_X1  g391(.A1(new_n815), .A2(new_n816), .B1(new_n801), .B2(new_n800), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT36), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n784), .A2(new_n818), .ZN(G150));
  INV_X1    g394(.A(G150), .ZN(G311));
  NOR2_X1   g395(.A1(new_n623), .A2(new_n629), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT38), .ZN(new_n822));
  AND2_X1   g397(.A1(new_n537), .A2(G55), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n516), .A2(G93), .ZN(new_n824));
  AOI22_X1  g399(.A1(new_n514), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n824), .B1(new_n503), .B2(new_n825), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n823), .A2(new_n826), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n827), .B1(new_n552), .B2(new_n554), .ZN(new_n828));
  INV_X1    g403(.A(new_n828), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n552), .A2(new_n554), .A3(new_n827), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n822), .B(new_n831), .ZN(new_n832));
  OR2_X1    g407(.A1(new_n832), .A2(KEYINPUT39), .ZN(new_n833));
  INV_X1    g408(.A(G860), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n832), .A2(KEYINPUT39), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n833), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n827), .A2(new_n834), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT37), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n836), .A2(new_n838), .ZN(G145));
  XNOR2_X1  g414(.A(new_n641), .B(new_n764), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(G162), .ZN(new_n841));
  INV_X1    g416(.A(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT100), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT4), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n497), .B(new_n844), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n843), .B1(new_n494), .B2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(new_n483), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n486), .B1(new_n487), .B2(G2105), .ZN(new_n848));
  NOR3_X1   g423(.A1(new_n460), .A2(KEYINPUT70), .A3(G114), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n491), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n850), .A2(KEYINPUT71), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n489), .A2(new_n484), .A3(new_n491), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n847), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n853), .A2(KEYINPUT100), .A3(new_n498), .ZN(new_n854));
  AND2_X1   g429(.A1(new_n846), .A2(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n735), .B(new_n855), .ZN(new_n856));
  OR2_X1    g431(.A1(new_n711), .A2(new_n751), .ZN(new_n857));
  INV_X1    g432(.A(new_n751), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n857), .B1(new_n712), .B2(new_n858), .ZN(new_n859));
  OR2_X1    g434(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n480), .A2(G142), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n474), .A2(G130), .ZN(new_n862));
  OAI21_X1  g437(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT101), .ZN(new_n864));
  INV_X1    g439(.A(G118), .ZN(new_n865));
  AOI22_X1  g440(.A1(new_n863), .A2(new_n864), .B1(new_n865), .B2(G2105), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n866), .B1(new_n864), .B2(new_n863), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n861), .A2(new_n862), .A3(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(new_n645), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(new_n807), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n856), .A2(new_n859), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n860), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT102), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n860), .A2(new_n871), .ZN(new_n875));
  INV_X1    g450(.A(new_n870), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n872), .A2(new_n873), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n842), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n841), .B(KEYINPUT103), .ZN(new_n881));
  AND2_X1   g456(.A1(new_n881), .A2(new_n872), .ZN(new_n882));
  AOI21_X1  g457(.A(G37), .B1(new_n882), .B2(new_n877), .ZN(new_n883));
  AND3_X1   g458(.A1(new_n880), .A2(new_n883), .A3(KEYINPUT40), .ZN(new_n884));
  AOI21_X1  g459(.A(KEYINPUT40), .B1(new_n880), .B2(new_n883), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n884), .A2(new_n885), .ZN(G395));
  NAND2_X1  g461(.A1(G166), .A2(KEYINPUT104), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT104), .ZN(new_n888));
  NAND2_X1  g463(.A1(G303), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n890), .A2(new_n786), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n887), .A2(new_n889), .A3(G305), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(G290), .A2(G288), .ZN(new_n894));
  INV_X1    g469(.A(G288), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n606), .A2(new_n895), .A3(new_n610), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n897), .A2(KEYINPUT105), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT105), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n894), .A2(new_n899), .A3(new_n896), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n893), .A2(new_n898), .A3(new_n900), .ZN(new_n901));
  NAND4_X1  g476(.A1(new_n891), .A2(KEYINPUT105), .A3(new_n897), .A4(new_n892), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n903), .B(KEYINPUT106), .ZN(new_n904));
  MUX2_X1   g479(.A(new_n903), .B(new_n904), .S(KEYINPUT42), .Z(new_n905));
  XNOR2_X1  g480(.A(new_n831), .B(new_n631), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n624), .A2(new_n583), .A3(new_n584), .ZN(new_n907));
  INV_X1    g482(.A(new_n584), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n623), .B1(new_n908), .B2(new_n582), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n907), .A2(KEYINPUT41), .A3(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  AOI21_X1  g486(.A(KEYINPUT41), .B1(new_n907), .B2(new_n909), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n906), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n907), .A2(new_n909), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n914), .B1(new_n906), .B2(new_n915), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n905), .B(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(G868), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n918), .B1(G868), .B2(new_n827), .ZN(G295));
  OAI21_X1  g494(.A(new_n918), .B1(G868), .B2(new_n827), .ZN(G331));
  OAI21_X1  g495(.A(G171), .B1(new_n588), .B2(new_n591), .ZN(new_n921));
  INV_X1    g496(.A(G168), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(G301), .ZN(new_n923));
  INV_X1    g498(.A(new_n830), .ZN(new_n924));
  OAI211_X1 g499(.A(new_n921), .B(new_n923), .C1(new_n924), .C2(new_n828), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n921), .A2(new_n923), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n926), .A2(new_n829), .A3(new_n830), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g503(.A(KEYINPUT107), .B1(new_n913), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n915), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT41), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n915), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(new_n910), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT107), .ZN(new_n934));
  NAND4_X1  g509(.A1(new_n933), .A2(new_n934), .A3(new_n927), .A4(new_n925), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n904), .A2(new_n929), .A3(new_n930), .A4(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(G37), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n928), .B1(new_n910), .B2(new_n932), .ZN(new_n939));
  AOI22_X1  g514(.A1(new_n939), .A2(new_n934), .B1(new_n915), .B2(new_n928), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n904), .B1(new_n940), .B2(new_n929), .ZN(new_n941));
  OAI21_X1  g516(.A(KEYINPUT43), .B1(new_n938), .B2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT106), .ZN(new_n943));
  XNOR2_X1  g518(.A(new_n903), .B(new_n943), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n930), .B1(new_n913), .B2(new_n928), .ZN(new_n945));
  AOI21_X1  g520(.A(G37), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT43), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n936), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(KEYINPUT108), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT108), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n936), .A2(new_n946), .A3(new_n950), .A4(new_n947), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n942), .A2(new_n949), .A3(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT44), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(new_n938), .ZN(new_n955));
  INV_X1    g530(.A(new_n941), .ZN(new_n956));
  AOI21_X1  g531(.A(KEYINPUT43), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  AND3_X1   g532(.A1(new_n936), .A2(new_n946), .A3(KEYINPUT43), .ZN(new_n958));
  OAI21_X1  g533(.A(KEYINPUT44), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n954), .A2(new_n959), .ZN(G397));
  INV_X1    g535(.A(G1384), .ZN(new_n961));
  AOI21_X1  g536(.A(KEYINPUT45), .B1(new_n855), .B2(new_n961), .ZN(new_n962));
  XNOR2_X1  g537(.A(KEYINPUT109), .B(G40), .ZN(new_n963));
  NOR3_X1   g538(.A1(new_n465), .A2(new_n469), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n965), .A2(G1996), .ZN(new_n966));
  XOR2_X1   g541(.A(new_n966), .B(KEYINPUT46), .Z(new_n967));
  XNOR2_X1  g542(.A(new_n965), .B(KEYINPUT110), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n735), .A2(G2067), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n730), .A2(new_n737), .A3(new_n734), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n968), .B1(new_n711), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n967), .A2(new_n972), .ZN(new_n973));
  XNOR2_X1  g548(.A(new_n973), .B(KEYINPUT47), .ZN(new_n974));
  AOI22_X1  g549(.A1(new_n968), .A2(new_n971), .B1(new_n712), .B2(new_n966), .ZN(new_n975));
  XNOR2_X1  g550(.A(new_n807), .B(new_n809), .ZN(new_n976));
  INV_X1    g551(.A(new_n968), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n968), .A2(G1996), .A3(new_n711), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT111), .ZN(new_n979));
  AND2_X1   g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n978), .A2(new_n979), .ZN(new_n981));
  OAI221_X1 g556(.A(new_n975), .B1(new_n976), .B2(new_n977), .C1(new_n980), .C2(new_n981), .ZN(new_n982));
  NOR3_X1   g557(.A1(new_n965), .A2(G1986), .A3(G290), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n983), .B(KEYINPUT48), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n974), .B1(new_n982), .B2(new_n984), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n807), .A2(new_n810), .ZN(new_n986));
  OAI211_X1 g561(.A(new_n986), .B(new_n975), .C1(new_n980), .C2(new_n981), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n977), .B1(new_n987), .B2(new_n970), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n985), .A2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(new_n964), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n961), .B1(new_n494), .B2(new_n845), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT45), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n990), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n992), .A2(G1384), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n499), .A2(new_n498), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n851), .A2(new_n852), .ZN(new_n996));
  AOI21_X1  g571(.A(KEYINPUT72), .B1(new_n996), .B2(new_n483), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n994), .B1(new_n995), .B2(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n993), .A2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(G1966), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g576(.A(G1384), .B1(new_n853), .B2(new_n498), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT50), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n990), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n845), .B1(new_n853), .B2(KEYINPUT72), .ZN(new_n1005));
  AOI21_X1  g580(.A(G1384), .B1(new_n1005), .B2(new_n496), .ZN(new_n1006));
  OAI211_X1 g581(.A(new_n766), .B(new_n1004), .C1(new_n1006), .C2(new_n1003), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1001), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(G8), .ZN(new_n1009));
  OR3_X1    g584(.A1(new_n1009), .A2(KEYINPUT116), .A3(G286), .ZN(new_n1010));
  OAI21_X1  g585(.A(KEYINPUT116), .B1(new_n1009), .B2(G286), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(G303), .A2(G8), .ZN(new_n1013));
  XNOR2_X1  g588(.A(new_n1013), .B(KEYINPUT55), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n846), .A2(new_n854), .A3(new_n994), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(new_n964), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1017), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n961), .B1(new_n995), .B2(new_n997), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(new_n992), .ZN(new_n1020));
  AOI21_X1  g595(.A(G1971), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1004), .B1(new_n1006), .B2(new_n1003), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1022), .A2(G2090), .ZN(new_n1023));
  OAI211_X1 g598(.A(G8), .B(new_n1015), .C1(new_n1021), .C2(new_n1023), .ZN(new_n1024));
  OAI211_X1 g599(.A(new_n961), .B(new_n964), .C1(new_n494), .C2(new_n845), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n895), .A2(G1976), .ZN(new_n1026));
  INV_X1    g601(.A(G1976), .ZN(new_n1027));
  AOI21_X1  g602(.A(KEYINPUT52), .B1(G288), .B2(new_n1027), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n1025), .A2(new_n1026), .A3(G8), .A4(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT113), .ZN(new_n1030));
  XNOR2_X1  g605(.A(new_n1029), .B(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(G8), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1032), .B1(new_n1002), .B2(new_n964), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT112), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1033), .A2(new_n1034), .A3(new_n1026), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1025), .A2(new_n1026), .A3(G8), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(KEYINPUT112), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1035), .A2(KEYINPUT52), .A3(new_n1037), .ZN(new_n1038));
  XNOR2_X1  g613(.A(KEYINPUT114), .B(G1981), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n786), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(G305), .A2(G1981), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT49), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1040), .A2(new_n1041), .A3(KEYINPUT49), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1044), .A2(new_n1033), .A3(new_n1045), .ZN(new_n1046));
  AND3_X1   g621(.A1(new_n1031), .A2(new_n1038), .A3(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1024), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT63), .ZN(new_n1050));
  OAI21_X1  g625(.A(G8), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1050), .B1(new_n1051), .B2(new_n1014), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1012), .A2(new_n1049), .A3(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1046), .A2(new_n1027), .A3(new_n895), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(new_n1040), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(new_n1033), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1031), .A2(new_n1038), .A3(new_n1046), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1056), .B1(new_n1024), .B2(new_n1057), .ZN(new_n1058));
  OR2_X1    g633(.A1(new_n1058), .A2(KEYINPUT115), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1058), .A2(KEYINPUT115), .ZN(new_n1060));
  AOI22_X1  g635(.A1(new_n1053), .A2(KEYINPUT63), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  AOI22_X1  g636(.A1(new_n1049), .A2(new_n1052), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT51), .ZN(new_n1063));
  NOR2_X1   g638(.A1(G168), .A2(new_n1032), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT123), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1063), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1064), .ZN(new_n1068));
  OAI211_X1 g643(.A(new_n1003), .B(new_n961), .C1(new_n494), .C2(new_n845), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(new_n964), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1070), .B1(new_n1019), .B2(KEYINPUT50), .ZN(new_n1071));
  AOI22_X1  g646(.A1(new_n1071), .A2(new_n766), .B1(new_n999), .B2(new_n1000), .ZN(new_n1072));
  OAI211_X1 g647(.A(new_n1067), .B(new_n1068), .C1(new_n1072), .C2(new_n1032), .ZN(new_n1073));
  OAI211_X1 g648(.A(G8), .B(new_n1066), .C1(new_n1008), .C2(new_n922), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  OAI21_X1  g650(.A(KEYINPUT122), .B1(new_n1072), .B2(new_n1068), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT122), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1008), .A2(new_n1077), .A3(new_n1064), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1076), .A2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1075), .A2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n993), .A2(new_n998), .A3(new_n774), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT124), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n993), .A2(new_n998), .A3(KEYINPUT124), .A4(new_n774), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1083), .A2(KEYINPUT53), .A3(new_n1084), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1020), .A2(new_n774), .A3(new_n964), .A4(new_n1016), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT53), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  XNOR2_X1  g663(.A(KEYINPUT125), .B(G1961), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1022), .A2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1085), .A2(new_n1088), .A3(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(G171), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(KEYINPUT126), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT126), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1091), .A2(new_n1094), .A3(G171), .ZN(new_n1095));
  AOI22_X1  g670(.A1(KEYINPUT62), .A2(new_n1080), .B1(new_n1093), .B2(new_n1095), .ZN(new_n1096));
  OR2_X1    g671(.A1(new_n1080), .A2(KEYINPUT62), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1062), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1006), .A2(KEYINPUT45), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n798), .B1(new_n1099), .B2(new_n1017), .ZN(new_n1100));
  OAI211_X1 g675(.A(new_n1003), .B(new_n961), .C1(new_n995), .C2(new_n997), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n990), .B1(new_n991), .B2(KEYINPUT50), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1101), .A2(new_n1102), .A3(new_n723), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1100), .A2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1015), .B1(new_n1104), .B2(G8), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1048), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1106), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1061), .B1(new_n1098), .B2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT57), .ZN(new_n1109));
  AND3_X1   g684(.A1(new_n576), .A2(new_n1109), .A3(new_n581), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1109), .B1(new_n576), .B2(new_n581), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  XNOR2_X1  g687(.A(KEYINPUT56), .B(G2072), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1020), .A2(new_n964), .A3(new_n1016), .A4(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(new_n720), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT118), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1112), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1114), .A2(KEYINPUT118), .A3(new_n1116), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1025), .A2(KEYINPUT117), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n853), .A2(new_n498), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT117), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1122), .A2(new_n1123), .A3(new_n961), .A4(new_n964), .ZN(new_n1124));
  AOI21_X1  g699(.A(G2067), .B1(new_n1121), .B2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1125), .B1(new_n1022), .B2(new_n778), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1126), .A2(new_n623), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1114), .A2(new_n1112), .A3(new_n1116), .ZN(new_n1128));
  AOI22_X1  g703(.A1(new_n1119), .A2(new_n1120), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT61), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1130), .A2(KEYINPUT119), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1128), .A2(new_n1132), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1114), .A2(new_n1116), .A3(new_n1112), .A4(new_n1131), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  OAI211_X1 g710(.A(new_n1117), .B(new_n1130), .C1(new_n1111), .C2(new_n1110), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT59), .ZN(new_n1137));
  INV_X1    g712(.A(G1996), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1018), .A2(new_n1138), .A3(new_n1020), .ZN(new_n1139));
  XOR2_X1   g714(.A(KEYINPUT58), .B(G1341), .Z(new_n1140));
  NAND3_X1  g715(.A1(new_n1121), .A2(new_n1124), .A3(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1137), .B1(new_n1142), .B2(new_n556), .ZN(new_n1143));
  AOI211_X1 g718(.A(KEYINPUT59), .B(new_n555), .C1(new_n1139), .C2(new_n1141), .ZN(new_n1144));
  OAI211_X1 g719(.A(new_n1135), .B(new_n1136), .C1(new_n1143), .C2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n624), .B1(new_n1126), .B2(KEYINPUT60), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT120), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1147), .B1(new_n1126), .B2(KEYINPUT60), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1003), .B1(new_n500), .B2(new_n961), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n778), .B1(new_n1149), .B2(new_n1070), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1125), .ZN(new_n1151));
  AND4_X1   g726(.A1(new_n1147), .A2(new_n1150), .A3(KEYINPUT60), .A4(new_n1151), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1146), .B1(new_n1148), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT60), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n623), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1150), .A2(new_n1151), .A3(KEYINPUT60), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1157), .A2(KEYINPUT120), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1126), .A2(new_n1147), .A3(KEYINPUT60), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1156), .A2(new_n1158), .A3(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1153), .A2(new_n1160), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1129), .B1(new_n1145), .B2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1162), .A2(KEYINPUT121), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT121), .ZN(new_n1164));
  OAI211_X1 g739(.A(new_n1129), .B(new_n1164), .C1(new_n1145), .C2(new_n1161), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1163), .A2(new_n1165), .ZN(new_n1166));
  AND3_X1   g741(.A1(new_n774), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1016), .A2(G160), .A3(new_n1167), .ZN(new_n1168));
  OR2_X1    g743(.A1(new_n962), .A2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1088), .A2(new_n1169), .A3(new_n1090), .ZN(new_n1170));
  OR2_X1    g745(.A1(new_n1170), .A2(G171), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1093), .A2(new_n1095), .A3(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT54), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1170), .A2(G171), .ZN(new_n1175));
  NAND4_X1  g750(.A1(new_n1085), .A2(new_n1088), .A3(G301), .A4(new_n1090), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1175), .A2(KEYINPUT54), .A3(new_n1176), .ZN(new_n1177));
  AND3_X1   g752(.A1(new_n1106), .A2(new_n1177), .A3(new_n1080), .ZN(new_n1178));
  AOI21_X1  g753(.A(KEYINPUT127), .B1(new_n1174), .B2(new_n1178), .ZN(new_n1179));
  NOR2_X1   g754(.A1(new_n1166), .A2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1174), .A2(new_n1178), .A3(KEYINPUT127), .ZN(new_n1181));
  AOI21_X1  g756(.A(new_n1108), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  XOR2_X1   g757(.A(G290), .B(G1986), .Z(new_n1183));
  NOR2_X1   g758(.A1(new_n965), .A2(new_n1183), .ZN(new_n1184));
  OR2_X1    g759(.A1(new_n982), .A2(new_n1184), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n989), .B1(new_n1182), .B2(new_n1185), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g761(.A1(new_n880), .A2(new_n883), .ZN(new_n1188));
  NOR4_X1   g762(.A1(G229), .A2(new_n458), .A3(G401), .A4(G227), .ZN(new_n1189));
  NAND3_X1  g763(.A1(new_n952), .A2(new_n1188), .A3(new_n1189), .ZN(G225));
  INV_X1    g764(.A(G225), .ZN(G308));
endmodule


