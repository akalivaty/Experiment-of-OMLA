//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 0 1 0 1 0 0 0 1 0 1 0 0 1 1 0 0 1 0 0 1 0 0 0 0 0 1 1 0 1 0 0 1 0 1 1 1 1 0 0 0 1 1 1 0 1 1 1 0 1 1 0 1 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:17 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1227,
    new_n1228, new_n1229, new_n1230, new_n1231, new_n1232, new_n1233,
    new_n1234, new_n1235, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1287, new_n1288,
    new_n1289, new_n1290, new_n1291, new_n1292, new_n1293, new_n1294,
    new_n1295, new_n1296, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1308, new_n1309, new_n1310, new_n1311, new_n1312, new_n1313,
    new_n1314, new_n1315, new_n1316, new_n1317, new_n1318, new_n1319,
    new_n1320, new_n1321, new_n1322, new_n1323, new_n1325, new_n1326,
    new_n1327, new_n1329, new_n1330, new_n1331, new_n1332, new_n1333,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1390, new_n1391, new_n1392, new_n1393, new_n1394,
    new_n1395, new_n1396, new_n1397, new_n1398, new_n1399, new_n1400,
    new_n1401, new_n1402, new_n1403, new_n1404, new_n1405, new_n1406,
    new_n1407, new_n1408, new_n1409, new_n1410, new_n1411, new_n1412,
    new_n1413, new_n1414, new_n1415, new_n1416, new_n1417, new_n1418,
    new_n1419, new_n1420, new_n1422, new_n1423, new_n1424, new_n1425,
    new_n1426, new_n1427;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  OAI21_X1  g0015(.A(G50), .B1(G58), .B2(G68), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  AND2_X1   g0017(.A1(G1), .A2(G13), .ZN(new_n218));
  NAND3_X1  g0018(.A1(new_n217), .A2(G20), .A3(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT64), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G116), .B2(G270), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n224));
  NAND3_X1  g0024(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n212), .B1(new_n221), .B2(new_n225), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n215), .B(new_n219), .C1(KEYINPUT1), .C2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XOR2_X1   g0028(.A(G238), .B(G244), .Z(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G226), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n233), .B(new_n236), .Z(G358));
  XNOR2_X1  g0037(.A(G50), .B(G68), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G58), .B(G77), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n238), .B(new_n239), .Z(new_n240));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G351));
  INV_X1    g0044(.A(KEYINPUT66), .ZN(new_n245));
  AND2_X1   g0045(.A1(G33), .A2(G41), .ZN(new_n246));
  NAND2_X1  g0046(.A1(G1), .A2(G13), .ZN(new_n247));
  OAI21_X1  g0047(.A(new_n245), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g0048(.A1(G33), .A2(G41), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n218), .A2(KEYINPUT66), .A3(new_n249), .ZN(new_n250));
  OAI21_X1  g0050(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n251));
  NAND4_X1  g0051(.A1(new_n248), .A2(new_n250), .A3(G226), .A4(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G274), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n254), .A2(new_n248), .A3(new_n250), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n252), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(KEYINPUT3), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT3), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(G33), .ZN(new_n261));
  INV_X1    g0061(.A(G1698), .ZN(new_n262));
  NAND4_X1  g0062(.A1(new_n259), .A2(new_n261), .A3(G222), .A4(new_n262), .ZN(new_n263));
  NAND4_X1  g0063(.A1(new_n259), .A2(new_n261), .A3(G223), .A4(G1698), .ZN(new_n264));
  INV_X1    g0064(.A(G77), .ZN(new_n265));
  XNOR2_X1  g0065(.A(KEYINPUT3), .B(G33), .ZN(new_n266));
  OAI211_X1 g0066(.A(new_n263), .B(new_n264), .C1(new_n265), .C2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n218), .A2(new_n249), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n257), .A2(new_n270), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n271), .A2(G179), .ZN(new_n272));
  NAND3_X1  g0072(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(new_n247), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G58), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(KEYINPUT8), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT8), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G58), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n210), .A2(G33), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NOR2_X1   g0082(.A1(G20), .A2(G33), .ZN(new_n283));
  AOI22_X1  g0083(.A1(new_n280), .A2(new_n282), .B1(G150), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n203), .A2(G20), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n275), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n209), .A2(G13), .A3(G20), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n275), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n209), .A2(G20), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G50), .ZN(new_n290));
  OAI22_X1  g0090(.A1(new_n288), .A2(new_n290), .B1(G50), .B2(new_n287), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n286), .A2(new_n291), .ZN(new_n292));
  AOI21_X1  g0092(.A(G169), .B1(new_n257), .B2(new_n270), .ZN(new_n293));
  NOR3_X1   g0093(.A1(new_n272), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n271), .A2(G200), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n292), .A2(KEYINPUT9), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n257), .A2(new_n270), .A3(G190), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT9), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n298), .B1(new_n286), .B2(new_n291), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n295), .A2(new_n296), .A3(new_n297), .A4(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(KEYINPUT10), .ZN(new_n301));
  NOR3_X1   g0101(.A1(new_n286), .A2(new_n291), .A3(new_n298), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n283), .A2(G150), .ZN(new_n303));
  XNOR2_X1  g0103(.A(KEYINPUT8), .B(G58), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n303), .B1(new_n304), .B2(new_n281), .ZN(new_n305));
  INV_X1    g0105(.A(new_n285), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n274), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n287), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n308), .A2(new_n274), .ZN(new_n309));
  INV_X1    g0109(.A(new_n290), .ZN(new_n310));
  AOI22_X1  g0110(.A1(new_n309), .A2(new_n310), .B1(new_n202), .B2(new_n308), .ZN(new_n311));
  AOI21_X1  g0111(.A(KEYINPUT9), .B1(new_n307), .B2(new_n311), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n302), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT10), .ZN(new_n314));
  NAND4_X1  g0114(.A1(new_n313), .A2(new_n314), .A3(new_n297), .A4(new_n295), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n294), .B1(new_n301), .B2(new_n315), .ZN(new_n316));
  NAND4_X1  g0116(.A1(new_n248), .A2(new_n250), .A3(G244), .A4(new_n251), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(new_n255), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n266), .A2(G232), .A3(new_n262), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n266), .A2(G238), .A3(G1698), .ZN(new_n320));
  OAI211_X1 g0120(.A(new_n319), .B(new_n320), .C1(new_n206), .C2(new_n266), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n318), .B1(new_n269), .B2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(G179), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n321), .A2(new_n269), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n325), .A2(new_n255), .A3(new_n317), .ZN(new_n326));
  INV_X1    g0126(.A(G169), .ZN(new_n327));
  AOI22_X1  g0127(.A1(new_n280), .A2(new_n283), .B1(G20), .B2(G77), .ZN(new_n328));
  XNOR2_X1  g0128(.A(KEYINPUT15), .B(G87), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n328), .B1(new_n281), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(new_n274), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n289), .A2(G77), .ZN(new_n332));
  OAI22_X1  g0132(.A1(new_n288), .A2(new_n332), .B1(G77), .B2(new_n287), .ZN(new_n333));
  INV_X1    g0133(.A(new_n333), .ZN(new_n334));
  AOI22_X1  g0134(.A1(new_n326), .A2(new_n327), .B1(new_n331), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n331), .A2(new_n334), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n336), .B1(G190), .B2(new_n322), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n326), .A2(G200), .ZN(new_n338));
  AOI22_X1  g0138(.A1(new_n324), .A2(new_n335), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND4_X1  g0139(.A1(new_n259), .A2(new_n261), .A3(G232), .A4(G1698), .ZN(new_n340));
  NAND4_X1  g0140(.A1(new_n259), .A2(new_n261), .A3(G226), .A4(new_n262), .ZN(new_n341));
  NAND2_X1  g0141(.A1(G33), .A2(G97), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n340), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(new_n269), .ZN(new_n344));
  NAND4_X1  g0144(.A1(new_n248), .A2(new_n250), .A3(G238), .A4(new_n251), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n344), .A2(new_n255), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(KEYINPUT13), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT13), .ZN(new_n348));
  NAND4_X1  g0148(.A1(new_n344), .A2(new_n348), .A3(new_n255), .A4(new_n345), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n347), .A2(KEYINPUT67), .A3(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT67), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n346), .A2(new_n351), .A3(KEYINPUT13), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n350), .A2(G200), .A3(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(G68), .ZN(new_n354));
  AOI22_X1  g0154(.A1(new_n283), .A2(G50), .B1(G20), .B2(new_n354), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n355), .B1(new_n265), .B2(new_n281), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(new_n274), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT11), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n308), .A2(new_n354), .ZN(new_n360));
  XNOR2_X1  g0160(.A(new_n360), .B(KEYINPUT12), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n356), .A2(KEYINPUT11), .A3(new_n274), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n309), .A2(G68), .A3(new_n289), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n359), .A2(new_n361), .A3(new_n362), .A4(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(G190), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n365), .B1(new_n346), .B2(KEYINPUT13), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n364), .B1(new_n366), .B2(new_n349), .ZN(new_n367));
  AND3_X1   g0167(.A1(new_n353), .A2(KEYINPUT68), .A3(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(KEYINPUT68), .B1(new_n353), .B2(new_n367), .ZN(new_n369));
  OAI211_X1 g0169(.A(new_n316), .B(new_n339), .C1(new_n368), .C2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n280), .A2(new_n289), .ZN(new_n372));
  OAI22_X1  g0172(.A1(new_n288), .A2(new_n372), .B1(new_n287), .B2(new_n280), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT71), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n259), .A2(new_n261), .ZN(new_n375));
  AOI21_X1  g0175(.A(KEYINPUT7), .B1(new_n375), .B2(new_n210), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT7), .ZN(new_n377));
  AOI211_X1 g0177(.A(new_n377), .B(G20), .C1(new_n259), .C2(new_n261), .ZN(new_n378));
  OAI21_X1  g0178(.A(G68), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT69), .ZN(new_n380));
  AND2_X1   g0180(.A1(G58), .A2(G68), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n380), .B(G20), .C1(new_n381), .C2(new_n201), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n283), .A2(G159), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  XNOR2_X1  g0184(.A(G58), .B(G68), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n380), .B1(new_n385), .B2(G20), .ZN(new_n386));
  OAI21_X1  g0186(.A(KEYINPUT70), .B1(new_n384), .B2(new_n386), .ZN(new_n387));
  OAI21_X1  g0187(.A(G20), .B1(new_n381), .B2(new_n201), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(KEYINPUT69), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT70), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n389), .A2(new_n390), .A3(new_n383), .A4(new_n382), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n379), .A2(new_n387), .A3(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT16), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n374), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n379), .A2(new_n387), .A3(KEYINPUT16), .A4(new_n391), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(new_n274), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n392), .A2(new_n374), .A3(new_n393), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n373), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n259), .A2(new_n261), .A3(G226), .A4(G1698), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n259), .A2(new_n261), .A3(G223), .A4(new_n262), .ZN(new_n401));
  NAND2_X1  g0201(.A1(G33), .A2(G87), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n400), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(new_n269), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT72), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n403), .A2(KEYINPUT72), .A3(new_n269), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n248), .A2(new_n250), .A3(G232), .A4(new_n251), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(new_n255), .ZN(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n406), .A2(new_n323), .A3(new_n407), .A4(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(KEYINPUT73), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n410), .A2(new_n404), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(new_n327), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n409), .B1(new_n404), .B2(new_n405), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT73), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n415), .A2(new_n416), .A3(new_n323), .A4(new_n407), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n412), .A2(new_n414), .A3(new_n417), .ZN(new_n418));
  NOR3_X1   g0218(.A1(new_n399), .A2(KEYINPUT18), .A3(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT18), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n392), .A2(new_n393), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(KEYINPUT71), .ZN(new_n422));
  AND2_X1   g0222(.A1(new_n395), .A2(new_n274), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n422), .A2(new_n423), .A3(new_n398), .ZN(new_n424));
  INV_X1    g0224(.A(new_n373), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  AND3_X1   g0226(.A1(new_n412), .A2(new_n414), .A3(new_n417), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n420), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n419), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n350), .A2(G169), .A3(new_n352), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT14), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n350), .A2(new_n352), .A3(KEYINPUT14), .A4(G169), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n347), .A2(G179), .A3(new_n349), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(new_n364), .ZN(new_n437));
  AND2_X1   g0237(.A1(new_n365), .A2(KEYINPUT74), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n365), .A2(KEYINPUT74), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n415), .A2(new_n407), .A3(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(G200), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n413), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(KEYINPUT17), .B1(new_n399), .B2(new_n444), .ZN(new_n445));
  AND4_X1   g0245(.A1(KEYINPUT17), .A2(new_n424), .A3(new_n425), .A4(new_n444), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n371), .A2(new_n429), .A3(new_n437), .A4(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT19), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n210), .B1(new_n342), .B2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(G87), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n451), .A2(new_n205), .A3(new_n206), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n259), .A2(new_n261), .A3(new_n210), .A4(G68), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n449), .B1(new_n281), .B2(new_n205), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n453), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(new_n274), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n209), .A2(G33), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n309), .A2(G87), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n329), .A2(new_n308), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n457), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n259), .A2(new_n261), .A3(G244), .A4(G1698), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n259), .A2(new_n261), .A3(G238), .A4(new_n262), .ZN(new_n463));
  NAND2_X1  g0263(.A1(G33), .A2(G116), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n462), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  NOR3_X1   g0265(.A1(new_n246), .A2(new_n245), .A3(new_n247), .ZN(new_n466));
  AOI21_X1  g0266(.A(KEYINPUT66), .B1(new_n218), .B2(new_n249), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  AOI21_X1  g0268(.A(G250), .B1(new_n209), .B2(G45), .ZN(new_n469));
  INV_X1    g0269(.A(G45), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n470), .A2(G1), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n469), .B1(new_n253), .B2(new_n471), .ZN(new_n472));
  AOI22_X1  g0272(.A1(new_n465), .A2(new_n269), .B1(new_n468), .B2(new_n472), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n461), .B1(G190), .B2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(new_n473), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(G200), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  AOI22_X1  g0277(.A1(new_n456), .A2(new_n274), .B1(new_n308), .B2(new_n329), .ZN(new_n478));
  AND3_X1   g0278(.A1(new_n275), .A2(new_n287), .A3(new_n458), .ZN(new_n479));
  INV_X1    g0279(.A(new_n329), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  AOI22_X1  g0281(.A1(new_n323), .A2(new_n473), .B1(new_n478), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n475), .A2(new_n327), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n477), .A2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(G41), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(KEYINPUT5), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT5), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(G41), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n471), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  AND4_X1   g0290(.A1(G257), .A2(new_n490), .A3(new_n248), .A4(new_n250), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n471), .A2(G274), .A3(new_n489), .ZN(new_n493));
  OAI21_X1  g0293(.A(KEYINPUT78), .B1(new_n488), .B2(G41), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT78), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n495), .A2(new_n486), .A3(KEYINPUT5), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n493), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  AOI21_X1  g0297(.A(KEYINPUT79), .B1(new_n497), .B2(new_n468), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n494), .A2(new_n496), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n486), .A2(KEYINPUT5), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n209), .A2(G45), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n499), .A2(new_n502), .A3(G274), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n248), .A2(new_n250), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT79), .ZN(new_n505));
  NOR3_X1   g0305(.A1(new_n503), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n492), .B1(new_n498), .B2(new_n506), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n259), .A2(new_n261), .A3(G244), .A4(new_n262), .ZN(new_n508));
  AND2_X1   g0308(.A1(KEYINPUT76), .A2(KEYINPUT4), .ZN(new_n509));
  NOR2_X1   g0309(.A1(KEYINPUT76), .A2(KEYINPUT4), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(G33), .A2(G283), .ZN(new_n513));
  INV_X1    g0313(.A(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(G250), .A2(G1698), .ZN(new_n515));
  NAND2_X1  g0315(.A1(KEYINPUT4), .A2(G244), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n515), .B1(new_n516), .B2(G1698), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n514), .B1(new_n266), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n512), .A2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT77), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n512), .A2(new_n518), .A3(KEYINPUT77), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n268), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n327), .B1(new_n507), .B2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(new_n522), .ZN(new_n525));
  AOI21_X1  g0325(.A(KEYINPUT77), .B1(new_n512), .B2(new_n518), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n269), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n505), .B1(new_n503), .B2(new_n504), .ZN(new_n528));
  INV_X1    g0328(.A(new_n493), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n468), .A2(KEYINPUT79), .A3(new_n499), .A4(new_n529), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n491), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n527), .A2(new_n531), .A3(new_n323), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT6), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(KEYINPUT75), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT75), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(KEYINPUT6), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n206), .A2(G97), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(G97), .A2(G107), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n207), .A2(new_n534), .A3(new_n536), .A4(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n539), .A2(G20), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n283), .A2(G77), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n377), .B1(new_n266), .B2(G20), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n375), .A2(KEYINPUT7), .A3(new_n210), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n206), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n274), .B1(new_n544), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n287), .A2(G97), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n549), .B1(new_n479), .B2(G97), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n524), .A2(new_n532), .A3(new_n551), .ZN(new_n552));
  OAI21_X1  g0352(.A(G200), .B1(new_n507), .B2(new_n523), .ZN(new_n553));
  INV_X1    g0353(.A(new_n551), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n527), .A2(new_n531), .A3(G190), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n552), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n479), .A2(G107), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT25), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n559), .B1(new_n287), .B2(G107), .ZN(new_n560));
  INV_X1    g0360(.A(new_n560), .ZN(new_n561));
  NOR3_X1   g0361(.A1(new_n287), .A2(new_n559), .A3(G107), .ZN(new_n562));
  OR2_X1    g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n259), .A2(new_n261), .A3(new_n210), .A4(G87), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT22), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n564), .A2(KEYINPUT81), .A3(new_n565), .ZN(new_n566));
  XNOR2_X1  g0366(.A(KEYINPUT81), .B(KEYINPUT22), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n266), .A2(new_n567), .A3(new_n210), .A4(G87), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT23), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n569), .A2(new_n206), .A3(G20), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(KEYINPUT82), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT82), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n572), .A2(new_n569), .A3(new_n206), .A4(G20), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(KEYINPUT83), .A2(KEYINPUT24), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n575), .B1(new_n464), .B2(G20), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n569), .B1(G20), .B2(new_n206), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n566), .A2(new_n568), .A3(new_n574), .A4(new_n578), .ZN(new_n579));
  NOR2_X1   g0379(.A1(KEYINPUT83), .A2(KEYINPUT24), .ZN(new_n580));
  XNOR2_X1  g0380(.A(new_n579), .B(new_n580), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n558), .B(new_n563), .C1(new_n581), .C2(new_n275), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n528), .A2(new_n530), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT84), .ZN(new_n584));
  OR2_X1    g0384(.A1(G250), .A2(G1698), .ZN(new_n585));
  OR2_X1    g0385(.A1(new_n262), .A2(G257), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n266), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(G33), .A2(G294), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n268), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  AND4_X1   g0389(.A1(G264), .A2(new_n490), .A3(new_n248), .A4(new_n250), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  AND3_X1   g0391(.A1(new_n583), .A2(new_n584), .A3(new_n591), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n584), .B1(new_n583), .B2(new_n591), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n365), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n583), .A2(new_n591), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(new_n442), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n582), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n558), .A2(new_n563), .ZN(new_n598));
  INV_X1    g0398(.A(new_n580), .ZN(new_n599));
  XNOR2_X1  g0399(.A(new_n579), .B(new_n599), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n598), .B1(new_n600), .B2(new_n274), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n595), .A2(KEYINPUT84), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n583), .A2(new_n584), .A3(new_n591), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n602), .A2(G169), .A3(new_n603), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n595), .A2(new_n323), .ZN(new_n605));
  INV_X1    g0405(.A(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n601), .B1(new_n604), .B2(new_n606), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n597), .A2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT21), .ZN(new_n609));
  INV_X1    g0409(.A(G116), .ZN(new_n610));
  AOI22_X1  g0410(.A1(new_n273), .A2(new_n247), .B1(G20), .B2(new_n610), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n513), .B(new_n210), .C1(G33), .C2(new_n205), .ZN(new_n612));
  AND3_X1   g0412(.A1(new_n611), .A2(KEYINPUT20), .A3(new_n612), .ZN(new_n613));
  AOI21_X1  g0413(.A(KEYINPUT20), .B1(new_n611), .B2(new_n612), .ZN(new_n614));
  OR2_X1    g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n287), .A2(G116), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n616), .B1(new_n479), .B2(G116), .ZN(new_n617));
  AOI211_X1 g0417(.A(new_n609), .B(new_n327), .C1(new_n615), .C2(new_n617), .ZN(new_n618));
  AND4_X1   g0418(.A1(G270), .A2(new_n490), .A3(new_n248), .A4(new_n250), .ZN(new_n619));
  INV_X1    g0419(.A(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(G303), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n268), .B1(new_n375), .B2(new_n621), .ZN(new_n622));
  NOR2_X1   g0422(.A1(G257), .A2(G1698), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n262), .A2(G264), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n266), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n622), .A2(new_n625), .ZN(new_n626));
  AND4_X1   g0426(.A1(KEYINPUT80), .A2(new_n583), .A3(new_n620), .A4(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n619), .B1(new_n528), .B2(new_n530), .ZN(new_n628));
  AOI21_X1  g0428(.A(KEYINPUT80), .B1(new_n628), .B2(new_n626), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n618), .B1(new_n627), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n615), .A2(new_n617), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n323), .B1(new_n622), .B2(new_n625), .ZN(new_n633));
  OAI211_X1 g0433(.A(new_n620), .B(new_n633), .C1(new_n498), .C2(new_n506), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n630), .A2(new_n636), .ZN(new_n637));
  OAI211_X1 g0437(.A(new_n620), .B(new_n626), .C1(new_n498), .C2(new_n506), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT80), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n628), .A2(KEYINPUT80), .A3(new_n626), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n631), .A2(G169), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  AOI21_X1  g0444(.A(KEYINPUT21), .B1(new_n642), .B2(new_n644), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n637), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n642), .A2(G200), .ZN(new_n647));
  OAI211_X1 g0447(.A(new_n647), .B(new_n632), .C1(new_n440), .C2(new_n642), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n608), .A2(new_n646), .A3(new_n648), .ZN(new_n649));
  NOR4_X1   g0449(.A1(new_n448), .A2(new_n485), .A3(new_n557), .A4(new_n649), .ZN(G372));
  INV_X1    g0450(.A(new_n294), .ZN(new_n651));
  INV_X1    g0451(.A(new_n429), .ZN(new_n652));
  AND2_X1   g0452(.A1(new_n353), .A2(new_n367), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n335), .A2(new_n324), .ZN(new_n654));
  OR2_X1    g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n437), .A2(new_n655), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n652), .B1(new_n656), .B2(new_n447), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n301), .A2(new_n315), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n651), .B1(new_n657), .B2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n604), .A2(new_n606), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(new_n582), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n644), .B1(new_n627), .B2(new_n629), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(new_n609), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n635), .B1(new_n642), .B2(new_n618), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT86), .ZN(new_n667));
  AND3_X1   g0467(.A1(new_n665), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n667), .B1(new_n665), .B2(new_n666), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n663), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n465), .A2(new_n269), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT85), .ZN(new_n672));
  INV_X1    g0472(.A(new_n469), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n471), .A2(new_n253), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n672), .B1(new_n504), .B2(new_n675), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n468), .A2(KEYINPUT85), .A3(new_n472), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n671), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(G200), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n474), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n678), .A2(new_n327), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n482), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n594), .A2(new_n596), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n683), .B1(new_n684), .B2(new_n601), .ZN(new_n685));
  INV_X1    g0485(.A(new_n557), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  AOI22_X1  g0488(.A1(new_n474), .A2(new_n679), .B1(new_n482), .B2(new_n681), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT26), .ZN(new_n690));
  AOI211_X1 g0490(.A(G179), .B(new_n491), .C1(new_n528), .C2(new_n530), .ZN(new_n691));
  AOI22_X1  g0491(.A1(new_n691), .A2(new_n527), .B1(new_n548), .B2(new_n550), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n689), .A2(new_n690), .A3(new_n692), .A4(new_n524), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(new_n682), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n583), .A2(new_n323), .A3(new_n492), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n551), .B1(new_n695), .B2(new_n523), .ZN(new_n696));
  AOI21_X1  g0496(.A(G169), .B1(new_n527), .B2(new_n531), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  AOI22_X1  g0498(.A1(new_n474), .A2(new_n476), .B1(new_n482), .B2(new_n483), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n690), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  OAI21_X1  g0500(.A(KEYINPUT87), .B1(new_n694), .B2(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(KEYINPUT26), .B1(new_n552), .B2(new_n485), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT87), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n702), .A2(new_n703), .A3(new_n682), .A4(new_n693), .ZN(new_n704));
  AOI22_X1  g0504(.A1(new_n670), .A2(new_n688), .B1(new_n701), .B2(new_n704), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n661), .B1(new_n448), .B2(new_n705), .ZN(G369));
  INV_X1    g0506(.A(G330), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n643), .B1(new_n640), .B2(new_n641), .ZN(new_n708));
  OAI211_X1 g0508(.A(new_n630), .B(new_n636), .C1(new_n708), .C2(KEYINPUT21), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(KEYINPUT86), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n665), .A2(new_n666), .A3(new_n667), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n209), .A2(new_n210), .A3(G13), .ZN(new_n712));
  OR2_X1    g0512(.A1(new_n712), .A2(KEYINPUT27), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(KEYINPUT27), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n713), .A2(G213), .A3(new_n714), .ZN(new_n715));
  XOR2_X1   g0515(.A(new_n715), .B(KEYINPUT88), .Z(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(G343), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(new_n631), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n710), .A2(new_n711), .A3(new_n720), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n646), .A2(new_n648), .A3(new_n719), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n707), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  AOI21_X1  g0523(.A(G190), .B1(new_n602), .B2(new_n603), .ZN(new_n724));
  INV_X1    g0524(.A(new_n596), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n601), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n582), .A2(new_n718), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n663), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n607), .A2(new_n718), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n723), .A2(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n718), .B1(new_n665), .B2(new_n666), .ZN(new_n732));
  AOI22_X1  g0532(.A1(new_n608), .A2(new_n732), .B1(new_n607), .B2(new_n717), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n731), .A2(new_n733), .ZN(G399));
  INV_X1    g0534(.A(new_n213), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n735), .A2(G41), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n452), .A2(G116), .ZN(new_n738));
  XOR2_X1   g0538(.A(new_n738), .B(KEYINPUT89), .Z(new_n739));
  NAND3_X1  g0539(.A1(new_n737), .A2(G1), .A3(new_n739), .ZN(new_n740));
  OAI22_X1  g0540(.A1(new_n740), .A2(KEYINPUT90), .B1(new_n216), .B2(new_n737), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n741), .B1(KEYINPUT90), .B2(new_n740), .ZN(new_n742));
  XNOR2_X1  g0542(.A(new_n742), .B(KEYINPUT28), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT29), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n744), .B1(new_n705), .B2(new_n718), .ZN(new_n745));
  OAI211_X1 g0545(.A(new_n685), .B(new_n686), .C1(new_n607), .C2(new_n709), .ZN(new_n746));
  OAI21_X1  g0546(.A(KEYINPUT26), .B1(new_n552), .B2(new_n683), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n699), .A2(new_n690), .A3(new_n692), .A4(new_n524), .ZN(new_n748));
  AND3_X1   g0548(.A1(new_n747), .A2(new_n682), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n746), .A2(new_n749), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n750), .A2(KEYINPUT29), .A3(new_n717), .ZN(new_n751));
  AND4_X1   g0551(.A1(new_n699), .A2(new_n552), .A3(new_n556), .A4(new_n717), .ZN(new_n752));
  NAND4_X1  g0552(.A1(new_n608), .A2(new_n646), .A3(new_n752), .A4(new_n648), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n591), .A2(new_n473), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n634), .A2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n507), .A2(new_n523), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n755), .A2(new_n756), .A3(KEYINPUT30), .ZN(new_n757));
  INV_X1    g0557(.A(KEYINPUT30), .ZN(new_n758));
  NAND4_X1  g0558(.A1(new_n628), .A2(new_n473), .A3(new_n591), .A4(new_n633), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n527), .A2(new_n531), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n758), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n627), .A2(new_n629), .ZN(new_n762));
  NAND4_X1  g0562(.A1(new_n760), .A2(new_n323), .A3(new_n595), .A4(new_n678), .ZN(new_n763));
  OAI211_X1 g0563(.A(new_n757), .B(new_n761), .C1(new_n762), .C2(new_n763), .ZN(new_n764));
  AOI21_X1  g0564(.A(KEYINPUT31), .B1(new_n764), .B2(new_n718), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n764), .A2(KEYINPUT31), .A3(new_n718), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n753), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(G330), .ZN(new_n769));
  INV_X1    g0569(.A(KEYINPUT91), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  AND3_X1   g0571(.A1(new_n764), .A2(KEYINPUT31), .A3(new_n718), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(new_n765), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n707), .B1(new_n773), .B2(new_n753), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(KEYINPUT91), .ZN(new_n775));
  AOI22_X1  g0575(.A1(new_n745), .A2(new_n751), .B1(new_n771), .B2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n743), .B1(new_n777), .B2(new_n209), .ZN(new_n778));
  XNOR2_X1  g0578(.A(new_n778), .B(KEYINPUT92), .ZN(G364));
  INV_X1    g0579(.A(G13), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(G20), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n209), .B1(new_n781), .B2(G45), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n736), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n213), .A2(new_n266), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n785), .B1(KEYINPUT93), .B2(G355), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n786), .B1(KEYINPUT93), .B2(G355), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n787), .B1(G116), .B2(new_n213), .ZN(new_n788));
  OR2_X1    g0588(.A1(new_n240), .A2(new_n470), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n735), .A2(new_n266), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n791), .B1(new_n470), .B2(new_n217), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n788), .B1(new_n789), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(G13), .A2(G33), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n795), .A2(G20), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n247), .B1(G20), .B2(new_n327), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n784), .B1(new_n793), .B2(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(G179), .A2(G200), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n210), .B1(new_n801), .B2(G190), .ZN(new_n802));
  XOR2_X1   g0602(.A(new_n802), .B(KEYINPUT95), .Z(new_n803));
  NAND2_X1  g0603(.A1(new_n803), .A2(G97), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n210), .A2(new_n323), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n805), .A2(G200), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n440), .A2(new_n806), .ZN(new_n807));
  NOR3_X1   g0607(.A1(new_n210), .A2(new_n442), .A3(G179), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n808), .A2(new_n365), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  AOI22_X1  g0610(.A1(new_n807), .A2(G50), .B1(new_n810), .B2(G107), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n808), .A2(G190), .ZN(new_n812));
  OAI211_X1 g0612(.A(new_n804), .B(new_n811), .C1(new_n451), .C2(new_n812), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n801), .A2(G20), .A3(new_n365), .ZN(new_n814));
  INV_X1    g0614(.A(G159), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  XNOR2_X1  g0616(.A(KEYINPUT94), .B(KEYINPUT32), .ZN(new_n817));
  XNOR2_X1  g0617(.A(new_n816), .B(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n805), .A2(new_n442), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n440), .A2(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n806), .A2(G190), .ZN(new_n821));
  AOI22_X1  g0621(.A1(new_n820), .A2(G58), .B1(new_n821), .B2(G68), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n819), .A2(G190), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n375), .B1(new_n823), .B2(G77), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n818), .A2(new_n822), .A3(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(G283), .ZN(new_n826));
  INV_X1    g0626(.A(G329), .ZN(new_n827));
  OAI22_X1  g0627(.A1(new_n809), .A2(new_n826), .B1(new_n827), .B2(new_n814), .ZN(new_n828));
  XOR2_X1   g0628(.A(new_n828), .B(KEYINPUT96), .Z(new_n829));
  INV_X1    g0629(.A(new_n812), .ZN(new_n830));
  AOI22_X1  g0630(.A1(new_n807), .A2(G326), .B1(new_n830), .B2(G303), .ZN(new_n831));
  AOI22_X1  g0631(.A1(new_n820), .A2(G322), .B1(new_n823), .B2(G311), .ZN(new_n832));
  INV_X1    g0632(.A(G317), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(KEYINPUT33), .ZN(new_n834));
  OR2_X1    g0634(.A1(new_n833), .A2(KEYINPUT33), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n821), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n802), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n266), .B1(new_n837), .B2(G294), .ZN(new_n838));
  NAND4_X1  g0638(.A1(new_n831), .A2(new_n832), .A3(new_n836), .A4(new_n838), .ZN(new_n839));
  OAI22_X1  g0639(.A1(new_n813), .A2(new_n825), .B1(new_n829), .B2(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n800), .B1(new_n840), .B2(new_n797), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n721), .A2(new_n722), .ZN(new_n842));
  INV_X1    g0642(.A(new_n796), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n841), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  OR2_X1    g0644(.A1(new_n723), .A2(new_n784), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n842), .A2(G330), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n844), .B1(new_n845), .B2(new_n846), .ZN(G396));
  INV_X1    g0647(.A(new_n654), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n337), .A2(new_n338), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n718), .A2(new_n336), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n848), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n654), .A2(new_n718), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n854), .B1(new_n705), .B2(new_n718), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n701), .A2(new_n704), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n710), .A2(new_n711), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n687), .B1(new_n858), .B2(new_n663), .ZN(new_n859));
  OAI211_X1 g0659(.A(new_n717), .B(new_n853), .C1(new_n857), .C2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n855), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n771), .A2(new_n775), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n784), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n863), .B1(new_n862), .B2(new_n861), .ZN(new_n864));
  INV_X1    g0664(.A(G311), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n375), .B1(new_n814), .B2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n823), .ZN(new_n867));
  OAI22_X1  g0667(.A1(new_n867), .A2(new_n610), .B1(new_n812), .B2(new_n206), .ZN(new_n868));
  AOI211_X1 g0668(.A(new_n866), .B(new_n868), .C1(G283), .C2(new_n821), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n809), .A2(new_n451), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  AOI22_X1  g0671(.A1(G294), .A2(new_n820), .B1(new_n807), .B2(G303), .ZN(new_n872));
  NAND4_X1  g0672(.A1(new_n869), .A2(new_n804), .A3(new_n871), .A4(new_n872), .ZN(new_n873));
  AOI22_X1  g0673(.A1(new_n820), .A2(G143), .B1(new_n821), .B2(G150), .ZN(new_n874));
  INV_X1    g0674(.A(G137), .ZN(new_n875));
  INV_X1    g0675(.A(new_n807), .ZN(new_n876));
  OAI221_X1 g0676(.A(new_n874), .B1(new_n875), .B2(new_n876), .C1(new_n815), .C2(new_n867), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT34), .ZN(new_n878));
  AND2_X1   g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(new_n814), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n375), .B1(new_n880), .B2(G132), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n881), .B1(new_n354), .B2(new_n809), .ZN(new_n882));
  OAI22_X1  g0682(.A1(new_n812), .A2(new_n202), .B1(new_n276), .B2(new_n802), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n884), .B1(new_n877), .B2(new_n878), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n873), .B1(new_n879), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(new_n797), .ZN(new_n887));
  INV_X1    g0687(.A(new_n784), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n797), .A2(new_n794), .ZN(new_n889));
  XOR2_X1   g0689(.A(new_n889), .B(KEYINPUT97), .Z(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n888), .B1(new_n891), .B2(new_n265), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n887), .B(new_n892), .C1(new_n853), .C2(new_n795), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n864), .A2(new_n893), .ZN(G384));
  NOR2_X1   g0694(.A1(new_n781), .A2(new_n209), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT38), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n424), .A2(new_n425), .A3(new_n444), .ZN(new_n897));
  AND2_X1   g0697(.A1(new_n417), .A2(new_n414), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n384), .A2(new_n386), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n545), .A2(new_n546), .ZN(new_n900));
  AOI22_X1  g0700(.A1(new_n899), .A2(new_n390), .B1(new_n900), .B2(G68), .ZN(new_n901));
  AOI21_X1  g0701(.A(KEYINPUT16), .B1(new_n901), .B2(new_n387), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n425), .B1(new_n902), .B2(new_n396), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n898), .A2(new_n903), .A3(new_n412), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n897), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(KEYINPUT100), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT100), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n897), .A2(new_n904), .A3(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT99), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n903), .A2(new_n909), .A3(new_n716), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n909), .B1(new_n903), .B2(new_n716), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n906), .A2(new_n908), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n426), .A2(new_n427), .ZN(new_n915));
  AOI21_X1  g0715(.A(KEYINPUT37), .B1(new_n915), .B2(KEYINPUT101), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT101), .ZN(new_n917));
  AND3_X1   g0717(.A1(new_n392), .A2(new_n374), .A3(new_n393), .ZN(new_n918));
  NOR3_X1   g0718(.A1(new_n918), .A2(new_n394), .A3(new_n396), .ZN(new_n919));
  OAI211_X1 g0719(.A(new_n427), .B(new_n917), .C1(new_n919), .C2(new_n373), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n716), .B1(new_n919), .B2(new_n373), .ZN(new_n921));
  AND3_X1   g0721(.A1(new_n920), .A2(new_n897), .A3(new_n921), .ZN(new_n922));
  AOI22_X1  g0722(.A1(new_n914), .A2(KEYINPUT37), .B1(new_n916), .B2(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n913), .B1(new_n429), .B2(new_n447), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n896), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n418), .B1(new_n424), .B2(new_n425), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(new_n420), .ZN(new_n927));
  OAI21_X1  g0727(.A(KEYINPUT18), .B1(new_n399), .B2(new_n418), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT17), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n897), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n399), .A2(KEYINPUT17), .A3(new_n444), .ZN(new_n931));
  NAND4_X1  g0731(.A1(new_n927), .A2(new_n928), .A3(new_n930), .A4(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n373), .B1(new_n423), .B2(new_n421), .ZN(new_n933));
  INV_X1    g0733(.A(new_n716), .ZN(new_n934));
  OAI21_X1  g0734(.A(KEYINPUT99), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(new_n910), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n932), .A2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT37), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n907), .B1(new_n897), .B2(new_n904), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n939), .A2(new_n936), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n938), .B1(new_n940), .B2(new_n908), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n920), .A2(new_n897), .A3(new_n921), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n938), .B1(new_n926), .B2(new_n917), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  OAI211_X1 g0744(.A(KEYINPUT38), .B(new_n937), .C1(new_n941), .C2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n925), .A2(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(new_n364), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n717), .A2(new_n947), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n653), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n437), .A2(new_n949), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n368), .A2(new_n369), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n948), .B1(new_n951), .B2(new_n436), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n953), .A2(new_n768), .A3(new_n853), .ZN(new_n954));
  INV_X1    g0754(.A(new_n954), .ZN(new_n955));
  AOI21_X1  g0755(.A(KEYINPUT40), .B1(new_n946), .B2(new_n955), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n915), .A2(new_n897), .A3(new_n921), .ZN(new_n957));
  AOI22_X1  g0757(.A1(new_n922), .A2(new_n916), .B1(KEYINPUT37), .B2(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n921), .B1(new_n429), .B2(new_n447), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n896), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n945), .A2(new_n960), .ZN(new_n961));
  NAND4_X1  g0761(.A1(new_n953), .A2(KEYINPUT40), .A3(new_n768), .A4(new_n853), .ZN(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n956), .B1(new_n961), .B2(new_n963), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n964), .B(KEYINPUT103), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n947), .B1(new_n434), .B2(new_n435), .ZN(new_n966));
  NOR3_X1   g0766(.A1(new_n932), .A2(new_n370), .A3(new_n966), .ZN(new_n967));
  AND2_X1   g0767(.A1(new_n967), .A2(new_n768), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n707), .B1(new_n965), .B2(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n969), .B1(new_n965), .B2(new_n968), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT39), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n961), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n966), .A2(new_n717), .ZN(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n925), .A2(KEYINPUT39), .A3(new_n945), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n972), .A2(new_n974), .A3(new_n975), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n429), .A2(new_n716), .ZN(new_n977));
  INV_X1    g0777(.A(new_n953), .ZN(new_n978));
  INV_X1    g0778(.A(new_n852), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n978), .B1(new_n860), .B2(new_n979), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n977), .B1(new_n980), .B2(new_n946), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n976), .A2(new_n981), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n607), .B1(new_n710), .B2(new_n711), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n856), .B1(new_n983), .B2(new_n687), .ZN(new_n984));
  AOI21_X1  g0784(.A(KEYINPUT29), .B1(new_n984), .B2(new_n717), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n751), .A2(new_n967), .ZN(new_n986));
  NOR3_X1   g0786(.A1(new_n985), .A2(KEYINPUT102), .A3(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT102), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n718), .B1(new_n746), .B2(new_n749), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n448), .B1(KEYINPUT29), .B2(new_n989), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n988), .B1(new_n745), .B2(new_n990), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n661), .B1(new_n987), .B2(new_n991), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n982), .B(new_n992), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n895), .B1(new_n970), .B2(new_n993), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n994), .B1(new_n993), .B2(new_n970), .ZN(new_n995));
  NOR3_X1   g0795(.A1(new_n247), .A2(new_n210), .A3(new_n610), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n539), .A2(new_n541), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT35), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n996), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n999), .B1(new_n998), .B2(new_n997), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(KEYINPUT98), .B(KEYINPUT36), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1000), .B(new_n1001), .ZN(new_n1002));
  NOR3_X1   g0802(.A1(new_n216), .A2(new_n381), .A3(new_n265), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n354), .A2(G50), .ZN(new_n1004));
  OAI211_X1 g0804(.A(G1), .B(new_n780), .C1(new_n1003), .C2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n995), .A2(new_n1002), .A3(new_n1005), .ZN(G367));
  INV_X1    g0806(.A(KEYINPUT105), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n745), .A2(new_n751), .ZN(new_n1008));
  NAND4_X1  g0808(.A1(new_n709), .A2(new_n663), .A3(new_n726), .A4(new_n717), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1009), .B1(new_n730), .B2(new_n732), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n723), .B(new_n1010), .ZN(new_n1011));
  AND3_X1   g0811(.A1(new_n1008), .A2(new_n862), .A3(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n607), .A2(new_n717), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1009), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n698), .A2(new_n718), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n554), .A2(new_n717), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1015), .B1(new_n557), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(KEYINPUT44), .B1(new_n1014), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT44), .ZN(new_n1020));
  AOI211_X1 g0820(.A(new_n1020), .B(new_n1017), .C1(new_n1009), .C2(new_n1013), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1022));
  AOI221_X4 g0822(.A(new_n707), .B1(new_n728), .B2(new_n729), .C1(new_n721), .C2(new_n722), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1009), .A2(new_n1013), .A3(new_n1017), .ZN(new_n1024));
  XOR2_X1   g0824(.A(KEYINPUT104), .B(KEYINPUT45), .Z(new_n1025));
  INV_X1    g0825(.A(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1027));
  NAND4_X1  g0827(.A1(new_n1009), .A2(new_n1013), .A3(new_n1017), .A4(new_n1025), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NOR3_X1   g0829(.A1(new_n1022), .A2(new_n1023), .A3(new_n1029), .ZN(new_n1030));
  AND2_X1   g0830(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1020), .B1(new_n733), .B2(new_n1017), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1014), .A2(new_n1018), .A3(KEYINPUT44), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n731), .B1(new_n1031), .B2(new_n1034), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n1030), .A2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1007), .B1(new_n1012), .B2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n1008), .A2(new_n862), .A3(new_n1011), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1023), .B1(new_n1022), .B2(new_n1029), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1031), .A2(new_n1034), .A3(new_n731), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NOR3_X1   g0841(.A1(new_n1038), .A2(new_n1041), .A3(KEYINPUT105), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n776), .B1(new_n1037), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT106), .ZN(new_n1044));
  XOR2_X1   g0844(.A(new_n736), .B(KEYINPUT41), .Z(new_n1045));
  INV_X1    g0845(.A(new_n1045), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1043), .A2(new_n1044), .A3(new_n1046), .ZN(new_n1047));
  NAND4_X1  g0847(.A1(new_n1036), .A2(new_n1007), .A3(new_n776), .A4(new_n1011), .ZN(new_n1048));
  OAI21_X1  g0848(.A(KEYINPUT105), .B1(new_n1038), .B2(new_n1041), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n777), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g0850(.A(KEYINPUT106), .B1(new_n1050), .B2(new_n1045), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1047), .A2(new_n1051), .A3(new_n782), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1017), .A2(new_n608), .A3(new_n732), .ZN(new_n1053));
  OR2_X1    g0853(.A1(new_n1053), .A2(KEYINPUT42), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n607), .A2(new_n556), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n718), .B1(new_n1055), .B2(new_n552), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1056), .B1(new_n1053), .B2(KEYINPUT42), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n718), .A2(new_n461), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1058), .A2(new_n689), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1059), .B1(new_n682), .B2(new_n1058), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n1054), .A2(new_n1057), .B1(KEYINPUT43), .B2(new_n1060), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n1060), .A2(KEYINPUT43), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1061), .B(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1023), .A2(new_n1017), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1063), .B(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1052), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n790), .A2(new_n236), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n1067), .B(new_n798), .C1(new_n213), .C2(new_n329), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n784), .B1(new_n1068), .B2(KEYINPUT107), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1069), .B1(KEYINPUT107), .B2(new_n1068), .ZN(new_n1070));
  XOR2_X1   g0870(.A(new_n1070), .B(KEYINPUT108), .Z(new_n1071));
  NOR2_X1   g0871(.A1(new_n812), .A2(new_n610), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(new_n1072), .B(KEYINPUT46), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n375), .B1(new_n814), .B2(new_n833), .C1(new_n206), .C2(new_n802), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n821), .ZN(new_n1075));
  INV_X1    g0875(.A(G294), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n1075), .A2(new_n1076), .B1(new_n809), .B2(new_n205), .ZN(new_n1077));
  NOR3_X1   g0877(.A1(new_n1073), .A2(new_n1074), .A3(new_n1077), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(G303), .A2(new_n820), .B1(new_n807), .B2(G311), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n1078), .B(new_n1079), .C1(new_n826), .C2(new_n867), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n803), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n1081), .A2(new_n354), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(G77), .A2(new_n810), .B1(new_n823), .B2(G50), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n830), .A2(G58), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n820), .A2(G150), .B1(new_n821), .B2(G159), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n266), .B1(new_n814), .B2(new_n875), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1086), .B1(new_n807), .B2(G143), .ZN(new_n1087));
  NAND4_X1  g0887(.A1(new_n1083), .A2(new_n1084), .A3(new_n1085), .A4(new_n1087), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1080), .B1(new_n1082), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(KEYINPUT47), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1092), .A2(new_n797), .ZN(new_n1093));
  OAI221_X1 g0893(.A(new_n1071), .B1(new_n843), .B2(new_n1060), .C1(new_n1091), .C2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1066), .A2(new_n1094), .ZN(G387));
  NAND2_X1  g0895(.A1(new_n1011), .A2(new_n783), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n790), .B1(new_n233), .B2(new_n470), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1097), .B1(new_n739), .B2(new_n785), .ZN(new_n1098));
  OR3_X1    g0898(.A1(new_n304), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1099));
  OAI21_X1  g0899(.A(KEYINPUT50), .B1(new_n304), .B2(G50), .ZN(new_n1100));
  AOI21_X1  g0900(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1101));
  NAND4_X1  g0901(.A1(new_n739), .A2(new_n1099), .A3(new_n1100), .A4(new_n1101), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n1098), .A2(new_n1102), .B1(new_n206), .B2(new_n735), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n784), .B1(new_n1103), .B2(new_n799), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(KEYINPUT109), .B(G322), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(G317), .A2(new_n820), .B1(new_n807), .B2(new_n1105), .ZN(new_n1106));
  OAI221_X1 g0906(.A(new_n1106), .B1(new_n621), .B2(new_n867), .C1(new_n865), .C2(new_n1075), .ZN(new_n1107));
  INV_X1    g0907(.A(KEYINPUT48), .ZN(new_n1108));
  OR2_X1    g0908(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n830), .A2(G294), .B1(new_n837), .B2(G283), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1109), .A2(new_n1110), .A3(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(KEYINPUT49), .ZN(new_n1113));
  OR2_X1    g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n809), .A2(new_n610), .ZN(new_n1116));
  AOI211_X1 g0916(.A(new_n266), .B(new_n1116), .C1(G326), .C2(new_n880), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1114), .A2(new_n1115), .A3(new_n1117), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n1075), .A2(new_n304), .B1(new_n265), .B2(new_n812), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1119), .B1(G159), .B2(new_n807), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n803), .A2(new_n480), .ZN(new_n1121));
  INV_X1    g0921(.A(G150), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n266), .B1(new_n814), .B2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1123), .B1(new_n810), .B2(G97), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n820), .A2(G50), .B1(new_n823), .B2(G68), .ZN(new_n1125));
  NAND4_X1  g0925(.A1(new_n1120), .A2(new_n1121), .A3(new_n1124), .A4(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1118), .A2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1104), .B1(new_n1127), .B2(new_n797), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1128), .B1(new_n730), .B2(new_n843), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1038), .A2(new_n736), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n776), .A2(new_n1011), .ZN(new_n1131));
  OAI211_X1 g0931(.A(new_n1096), .B(new_n1129), .C1(new_n1130), .C2(new_n1131), .ZN(G393));
  NAND2_X1  g0932(.A1(new_n1036), .A2(new_n783), .ZN(new_n1133));
  OAI221_X1 g0933(.A(new_n798), .B1(new_n205), .B2(new_n213), .C1(new_n791), .C2(new_n243), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1134), .A2(new_n784), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(G311), .A2(new_n820), .B1(new_n807), .B2(G317), .ZN(new_n1136));
  AND2_X1   g0936(.A1(new_n1136), .A2(KEYINPUT52), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n1136), .A2(KEYINPUT52), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n266), .B1(new_n880), .B2(new_n1105), .ZN(new_n1139));
  OAI221_X1 g0939(.A(new_n1139), .B1(new_n206), .B2(new_n809), .C1(new_n826), .C2(new_n812), .ZN(new_n1140));
  OR3_X1    g0940(.A1(new_n1137), .A2(new_n1138), .A3(new_n1140), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n823), .A2(G294), .B1(G116), .B2(new_n837), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1142), .B1(new_n621), .B2(new_n1075), .ZN(new_n1143));
  XNOR2_X1  g0943(.A(new_n1143), .B(KEYINPUT110), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(G150), .A2(new_n807), .B1(new_n820), .B2(G159), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(new_n1145), .B(KEYINPUT51), .ZN(new_n1146));
  AOI211_X1 g0946(.A(new_n375), .B(new_n870), .C1(G143), .C2(new_n880), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n803), .A2(G77), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n821), .A2(G50), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(G68), .A2(new_n830), .B1(new_n823), .B2(new_n280), .ZN(new_n1150));
  NAND4_X1  g0950(.A1(new_n1147), .A2(new_n1148), .A3(new_n1149), .A4(new_n1150), .ZN(new_n1151));
  OAI22_X1  g0951(.A1(new_n1141), .A2(new_n1144), .B1(new_n1146), .B2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1135), .B1(new_n1152), .B2(new_n797), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1153), .B1(new_n1017), .B2(new_n843), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT111), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n737), .B1(new_n1038), .B2(new_n1041), .ZN(new_n1157));
  AND3_X1   g0957(.A1(new_n1155), .A2(new_n1156), .A3(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1156), .B1(new_n1155), .B2(new_n1157), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n1133), .B(new_n1154), .C1(new_n1158), .C2(new_n1159), .ZN(G390));
  AND3_X1   g0960(.A1(new_n925), .A2(KEYINPUT39), .A3(new_n945), .ZN(new_n1161));
  AOI21_X1  g0961(.A(KEYINPUT39), .B1(new_n945), .B2(new_n960), .ZN(new_n1162));
  OAI22_X1  g0962(.A1(new_n1161), .A2(new_n1162), .B1(new_n974), .B2(new_n980), .ZN(new_n1163));
  AOI211_X1 g0963(.A(new_n770), .B(new_n707), .C1(new_n773), .C2(new_n753), .ZN(new_n1164));
  AOI21_X1  g0964(.A(KEYINPUT91), .B1(new_n768), .B2(G330), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n978), .A2(new_n854), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  AND2_X1   g0968(.A1(new_n945), .A2(new_n960), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n851), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n852), .B1(new_n989), .B2(new_n1170), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n973), .B1(new_n1171), .B2(new_n978), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1169), .A2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1163), .A2(new_n1168), .A3(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n980), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1176), .A2(new_n973), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n972), .A2(new_n975), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1173), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n768), .A2(G330), .A3(new_n853), .ZN(new_n1180));
  OAI21_X1  g0980(.A(KEYINPUT112), .B1(new_n1180), .B2(new_n978), .ZN(new_n1181));
  INV_X1    g0981(.A(KEYINPUT112), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n774), .A2(new_n1182), .A3(new_n953), .A4(new_n853), .ZN(new_n1183));
  AND2_X1   g0983(.A1(new_n1181), .A2(new_n1183), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n1175), .B(new_n783), .C1(new_n1179), .C2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1185), .A2(KEYINPUT113), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1181), .A2(new_n1183), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(new_n1176), .A2(new_n973), .B1(new_n972), .B2(new_n975), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1187), .B1(new_n1188), .B2(new_n1173), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT113), .ZN(new_n1190));
  NAND4_X1  g0990(.A1(new_n1189), .A2(new_n1190), .A3(new_n783), .A4(new_n1175), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1186), .A2(new_n1191), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n769), .A2(new_n448), .ZN(new_n1193));
  OAI21_X1  g0993(.A(KEYINPUT102), .B1(new_n985), .B2(new_n986), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n745), .A2(new_n990), .A3(new_n988), .ZN(new_n1195));
  AOI211_X1 g0995(.A(new_n660), .B(new_n1193), .C1(new_n1194), .C2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n771), .A2(new_n775), .A3(new_n853), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1197), .A2(new_n978), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(new_n1184), .A2(new_n1198), .B1(new_n979), .B2(new_n860), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1180), .A2(new_n978), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1200), .A2(new_n1171), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1201), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1196), .B1(new_n1199), .B2(new_n1202), .ZN(new_n1203));
  AND3_X1   g1003(.A1(new_n1163), .A2(new_n1168), .A3(new_n1174), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1184), .B1(new_n1163), .B2(new_n1174), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1203), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n860), .A2(new_n979), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n953), .B1(new_n1166), .B2(new_n853), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1207), .B1(new_n1208), .B2(new_n1187), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1168), .A2(new_n1171), .A3(new_n1200), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n1189), .A2(new_n1175), .A3(new_n1211), .A4(new_n1196), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1206), .A2(new_n1212), .A3(new_n736), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n795), .B1(new_n972), .B2(new_n975), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n812), .A2(new_n1122), .ZN(new_n1215));
  XNOR2_X1  g1015(.A(new_n1215), .B(KEYINPUT53), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1216), .B1(new_n815), .B2(new_n1081), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(new_n820), .A2(G132), .B1(new_n810), .B2(G50), .ZN(new_n1218));
  XOR2_X1   g1018(.A(KEYINPUT54), .B(G143), .Z(new_n1219));
  AOI22_X1  g1019(.A1(new_n807), .A2(G128), .B1(new_n823), .B2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n821), .A2(G137), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n375), .B1(new_n880), .B2(G125), .ZN(new_n1222));
  NAND4_X1  g1022(.A1(new_n1218), .A2(new_n1220), .A3(new_n1221), .A4(new_n1222), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n820), .A2(G116), .B1(new_n821), .B2(G107), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n807), .A2(G283), .B1(new_n823), .B2(G97), .ZN(new_n1225));
  OAI22_X1  g1025(.A1(new_n809), .A2(new_n354), .B1(new_n1076), .B2(new_n814), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1226), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1148), .A2(new_n1224), .A3(new_n1225), .A4(new_n1227), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n375), .B1(new_n812), .B2(new_n451), .ZN(new_n1229));
  XNOR2_X1  g1029(.A(new_n1229), .B(KEYINPUT114), .ZN(new_n1230));
  OAI22_X1  g1030(.A1(new_n1217), .A2(new_n1223), .B1(new_n1228), .B2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1231), .A2(new_n797), .ZN(new_n1232));
  OAI211_X1 g1032(.A(new_n1232), .B(new_n784), .C1(new_n280), .C2(new_n890), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n1214), .A2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1192), .A2(new_n1213), .A3(new_n1235), .ZN(G378));
  INV_X1    g1036(.A(new_n889), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n784), .B1(G50), .B2(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n316), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n934), .A2(new_n292), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1241), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1243));
  XNOR2_X1  g1043(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1244), .ZN(new_n1245));
  OR3_X1    g1045(.A1(new_n1242), .A2(new_n1243), .A3(new_n1245), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1245), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1248), .A2(new_n795), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n266), .A2(G41), .ZN(new_n1250));
  AOI211_X1 g1050(.A(G50), .B(new_n1250), .C1(new_n258), .C2(new_n486), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n820), .A2(G107), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1252), .B1(new_n876), .B2(new_n610), .ZN(new_n1253));
  OAI22_X1  g1053(.A1(new_n205), .A2(new_n1075), .B1(new_n867), .B2(new_n329), .ZN(new_n1254));
  OAI221_X1 g1054(.A(new_n1250), .B1(new_n826), .B2(new_n814), .C1(new_n812), .C2(new_n265), .ZN(new_n1255));
  NOR3_X1   g1055(.A1(new_n1253), .A2(new_n1254), .A3(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n810), .A2(G58), .ZN(new_n1257));
  XNOR2_X1  g1057(.A(new_n1257), .B(KEYINPUT115), .ZN(new_n1258));
  OAI211_X1 g1058(.A(new_n1256), .B(new_n1258), .C1(new_n354), .C2(new_n1081), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT58), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1251), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n803), .A2(G150), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(new_n807), .A2(G125), .B1(new_n821), .B2(G132), .ZN(new_n1263));
  AOI22_X1  g1063(.A1(new_n830), .A2(new_n1219), .B1(new_n823), .B2(G137), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n820), .A2(G128), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1262), .A2(new_n1263), .A3(new_n1264), .A4(new_n1265), .ZN(new_n1266));
  XNOR2_X1  g1066(.A(new_n1266), .B(KEYINPUT59), .ZN(new_n1267));
  AOI211_X1 g1067(.A(G33), .B(G41), .C1(new_n880), .C2(G124), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1268), .B1(new_n815), .B2(new_n809), .ZN(new_n1269));
  OAI221_X1 g1069(.A(new_n1261), .B1(new_n1260), .B2(new_n1259), .C1(new_n1267), .C2(new_n1269), .ZN(new_n1270));
  AOI211_X1 g1070(.A(new_n1238), .B(new_n1249), .C1(new_n797), .C2(new_n1270), .ZN(new_n1271));
  OAI21_X1  g1071(.A(G330), .B1(new_n1169), .B2(new_n962), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1248), .ZN(new_n1273));
  NOR3_X1   g1073(.A1(new_n1272), .A2(new_n956), .A3(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n946), .A2(new_n955), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT40), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n707), .B1(new_n961), .B2(new_n963), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1248), .B1(new_n1277), .B2(new_n1278), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n982), .B1(new_n1274), .B2(new_n1279), .ZN(new_n1280));
  AND2_X1   g1080(.A1(new_n976), .A2(new_n981), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1277), .A2(new_n1278), .A3(new_n1248), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1273), .B1(new_n1272), .B2(new_n956), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1281), .A2(new_n1282), .A3(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1280), .A2(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1271), .B1(new_n1285), .B2(new_n783), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1193), .ZN(new_n1287));
  OAI211_X1 g1087(.A(new_n661), .B(new_n1287), .C1(new_n987), .C2(new_n991), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1288), .B1(new_n1289), .B2(new_n1211), .ZN(new_n1290));
  AND3_X1   g1090(.A1(new_n1281), .A2(new_n1282), .A3(new_n1283), .ZN(new_n1291));
  AOI22_X1  g1091(.A1(new_n1282), .A2(new_n1283), .B1(new_n976), .B2(new_n981), .ZN(new_n1292));
  OAI21_X1  g1092(.A(KEYINPUT57), .B1(new_n1291), .B2(new_n1292), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n736), .B1(new_n1290), .B2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1212), .A2(new_n1196), .ZN(new_n1295));
  AOI21_X1  g1095(.A(KEYINPUT57), .B1(new_n1295), .B2(new_n1285), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1286), .B1(new_n1294), .B2(new_n1296), .ZN(G375));
  XNOR2_X1  g1097(.A(new_n782), .B(KEYINPUT116), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1211), .A2(new_n1298), .ZN(new_n1299));
  OAI22_X1  g1099(.A1(new_n1075), .A2(new_n610), .B1(new_n205), .B2(new_n812), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1300), .B1(G283), .B2(new_n820), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n375), .B1(new_n814), .B2(new_n621), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1302), .B1(new_n810), .B2(G77), .ZN(new_n1303));
  AOI22_X1  g1103(.A1(new_n807), .A2(G294), .B1(new_n823), .B2(G107), .ZN(new_n1304));
  NAND4_X1  g1104(.A1(new_n1301), .A2(new_n1121), .A3(new_n1303), .A4(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n807), .A2(G132), .ZN(new_n1306));
  XNOR2_X1  g1106(.A(new_n1306), .B(KEYINPUT117), .ZN(new_n1307));
  OAI211_X1 g1107(.A(new_n1307), .B(new_n1258), .C1(new_n202), .C2(new_n1081), .ZN(new_n1308));
  AOI22_X1  g1108(.A1(G159), .A2(new_n830), .B1(new_n821), .B2(new_n1219), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n820), .A2(G137), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n375), .B1(new_n880), .B2(G128), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n823), .A2(G150), .ZN(new_n1312));
  NAND4_X1  g1112(.A1(new_n1309), .A2(new_n1310), .A3(new_n1311), .A4(new_n1312), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1305), .B1(new_n1308), .B2(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1314), .A2(new_n797), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n888), .B1(new_n891), .B2(new_n354), .ZN(new_n1316));
  OAI211_X1 g1116(.A(new_n1315), .B(new_n1316), .C1(new_n953), .C2(new_n795), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1299), .A2(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1184), .A2(new_n1198), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1202), .B1(new_n1320), .B2(new_n1207), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1321), .A2(new_n1288), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1322), .A2(new_n1046), .A3(new_n1203), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1319), .A2(new_n1323), .ZN(G381));
  INV_X1    g1124(.A(G390), .ZN(new_n1325));
  NOR3_X1   g1125(.A1(G393), .A2(G384), .A3(G396), .ZN(new_n1326));
  NAND4_X1  g1126(.A1(new_n1325), .A2(new_n1319), .A3(new_n1323), .A4(new_n1326), .ZN(new_n1327));
  OR4_X1    g1127(.A1(G387), .A2(G375), .A3(new_n1327), .A4(G378), .ZN(G407));
  INV_X1    g1128(.A(G378), .ZN(new_n1329));
  INV_X1    g1129(.A(G213), .ZN(new_n1330));
  NOR2_X1   g1130(.A1(new_n1330), .A2(G343), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1329), .A2(new_n1331), .ZN(new_n1332));
  OAI211_X1 g1132(.A(G407), .B(G213), .C1(G375), .C2(new_n1332), .ZN(new_n1333));
  XNOR2_X1  g1133(.A(new_n1333), .B(KEYINPUT118), .ZN(G409));
  XOR2_X1   g1134(.A(G393), .B(G396), .Z(new_n1335));
  INV_X1    g1135(.A(new_n1335), .ZN(new_n1336));
  INV_X1    g1136(.A(KEYINPUT123), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(G387), .A2(new_n1325), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1066), .A2(new_n1094), .A3(G390), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1338), .A2(new_n1339), .ZN(new_n1340));
  INV_X1    g1140(.A(KEYINPUT124), .ZN(new_n1341));
  AOI21_X1  g1141(.A(new_n1337), .B1(new_n1340), .B2(new_n1341), .ZN(new_n1342));
  AND3_X1   g1142(.A1(new_n1066), .A2(new_n1094), .A3(G390), .ZN(new_n1343));
  AOI21_X1  g1143(.A(G390), .B1(new_n1066), .B2(new_n1094), .ZN(new_n1344));
  OAI211_X1 g1144(.A(new_n1337), .B(new_n1341), .C1(new_n1343), .C2(new_n1344), .ZN(new_n1345));
  INV_X1    g1145(.A(new_n1345), .ZN(new_n1346));
  OAI21_X1  g1146(.A(new_n1336), .B1(new_n1342), .B2(new_n1346), .ZN(new_n1347));
  OAI21_X1  g1147(.A(new_n1341), .B1(new_n1343), .B2(new_n1344), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1348), .A2(KEYINPUT123), .ZN(new_n1349));
  NAND3_X1  g1149(.A1(new_n1349), .A2(new_n1335), .A3(new_n1345), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1347), .A2(new_n1350), .ZN(new_n1351));
  OAI211_X1 g1151(.A(G378), .B(new_n1286), .C1(new_n1294), .C2(new_n1296), .ZN(new_n1352));
  NAND3_X1  g1152(.A1(new_n1295), .A2(new_n1046), .A3(new_n1285), .ZN(new_n1353));
  AOI21_X1  g1153(.A(new_n1271), .B1(new_n1285), .B2(new_n1298), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1353), .A2(new_n1354), .ZN(new_n1355));
  AND2_X1   g1155(.A1(new_n1213), .A2(new_n1235), .ZN(new_n1356));
  NAND3_X1  g1156(.A1(new_n1355), .A2(new_n1192), .A3(new_n1356), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1352), .A2(new_n1357), .ZN(new_n1358));
  INV_X1    g1158(.A(new_n1331), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1358), .A2(new_n1359), .ZN(new_n1360));
  INV_X1    g1160(.A(G2897), .ZN(new_n1361));
  NOR2_X1   g1161(.A1(new_n1359), .A2(new_n1361), .ZN(new_n1362));
  INV_X1    g1162(.A(new_n1362), .ZN(new_n1363));
  INV_X1    g1163(.A(G384), .ZN(new_n1364));
  OR2_X1    g1164(.A1(new_n1364), .A2(KEYINPUT120), .ZN(new_n1365));
  NAND2_X1  g1165(.A1(new_n1364), .A2(KEYINPUT120), .ZN(new_n1366));
  NAND4_X1  g1166(.A1(new_n1209), .A2(KEYINPUT60), .A3(new_n1288), .A4(new_n1210), .ZN(new_n1367));
  NAND2_X1  g1167(.A1(new_n1367), .A2(new_n736), .ZN(new_n1368));
  XOR2_X1   g1168(.A(KEYINPUT119), .B(KEYINPUT60), .Z(new_n1369));
  OAI21_X1  g1169(.A(new_n1369), .B1(new_n1321), .B2(new_n1288), .ZN(new_n1370));
  AOI21_X1  g1170(.A(new_n1368), .B1(new_n1322), .B2(new_n1370), .ZN(new_n1371));
  OAI211_X1 g1171(.A(new_n1365), .B(new_n1366), .C1(new_n1371), .C2(new_n1318), .ZN(new_n1372));
  INV_X1    g1172(.A(new_n1369), .ZN(new_n1373));
  AOI21_X1  g1173(.A(new_n1373), .B1(new_n1211), .B2(new_n1196), .ZN(new_n1374));
  NOR2_X1   g1174(.A1(new_n1211), .A2(new_n1196), .ZN(new_n1375));
  OAI211_X1 g1175(.A(new_n736), .B(new_n1367), .C1(new_n1374), .C2(new_n1375), .ZN(new_n1376));
  NAND4_X1  g1176(.A1(new_n1376), .A2(KEYINPUT120), .A3(new_n1364), .A4(new_n1319), .ZN(new_n1377));
  AND3_X1   g1177(.A1(new_n1372), .A2(KEYINPUT121), .A3(new_n1377), .ZN(new_n1378));
  AOI21_X1  g1178(.A(KEYINPUT121), .B1(new_n1372), .B2(new_n1377), .ZN(new_n1379));
  OAI21_X1  g1179(.A(new_n1363), .B1(new_n1378), .B2(new_n1379), .ZN(new_n1380));
  NAND2_X1  g1180(.A1(new_n1372), .A2(new_n1377), .ZN(new_n1381));
  NOR2_X1   g1181(.A1(new_n1381), .A2(new_n1363), .ZN(new_n1382));
  INV_X1    g1182(.A(new_n1382), .ZN(new_n1383));
  NAND3_X1  g1183(.A1(new_n1360), .A2(new_n1380), .A3(new_n1383), .ZN(new_n1384));
  INV_X1    g1184(.A(KEYINPUT61), .ZN(new_n1385));
  AOI21_X1  g1185(.A(KEYINPUT125), .B1(new_n1384), .B2(new_n1385), .ZN(new_n1386));
  NOR2_X1   g1186(.A1(new_n1378), .A2(new_n1379), .ZN(new_n1387));
  OAI21_X1  g1187(.A(KEYINPUT62), .B1(new_n1360), .B2(new_n1387), .ZN(new_n1388));
  INV_X1    g1188(.A(KEYINPUT121), .ZN(new_n1389));
  NAND2_X1  g1189(.A1(new_n1381), .A2(new_n1389), .ZN(new_n1390));
  NAND3_X1  g1190(.A1(new_n1372), .A2(KEYINPUT121), .A3(new_n1377), .ZN(new_n1391));
  NAND2_X1  g1191(.A1(new_n1390), .A2(new_n1391), .ZN(new_n1392));
  AOI21_X1  g1192(.A(new_n1331), .B1(new_n1352), .B2(new_n1357), .ZN(new_n1393));
  INV_X1    g1193(.A(KEYINPUT62), .ZN(new_n1394));
  NAND3_X1  g1194(.A1(new_n1392), .A2(new_n1393), .A3(new_n1394), .ZN(new_n1395));
  NAND2_X1  g1195(.A1(new_n1388), .A2(new_n1395), .ZN(new_n1396));
  NOR2_X1   g1196(.A1(new_n1386), .A2(new_n1396), .ZN(new_n1397));
  NAND3_X1  g1197(.A1(new_n1384), .A2(KEYINPUT125), .A3(new_n1385), .ZN(new_n1398));
  AOI21_X1  g1198(.A(new_n1351), .B1(new_n1397), .B2(new_n1398), .ZN(new_n1399));
  INV_X1    g1199(.A(KEYINPUT63), .ZN(new_n1400));
  OAI21_X1  g1200(.A(new_n1400), .B1(new_n1360), .B2(new_n1387), .ZN(new_n1401));
  NAND3_X1  g1201(.A1(new_n1392), .A2(new_n1393), .A3(KEYINPUT63), .ZN(new_n1402));
  AND3_X1   g1202(.A1(new_n1349), .A2(new_n1335), .A3(new_n1345), .ZN(new_n1403));
  AOI21_X1  g1203(.A(new_n1335), .B1(new_n1349), .B2(new_n1345), .ZN(new_n1404));
  OAI211_X1 g1204(.A(new_n1401), .B(new_n1402), .C1(new_n1403), .C2(new_n1404), .ZN(new_n1405));
  AOI21_X1  g1205(.A(new_n1362), .B1(new_n1390), .B2(new_n1391), .ZN(new_n1406));
  OAI21_X1  g1206(.A(KEYINPUT122), .B1(new_n1406), .B2(new_n1382), .ZN(new_n1407));
  INV_X1    g1207(.A(KEYINPUT122), .ZN(new_n1408));
  NAND3_X1  g1208(.A1(new_n1380), .A2(new_n1383), .A3(new_n1408), .ZN(new_n1409));
  NAND3_X1  g1209(.A1(new_n1407), .A2(new_n1409), .A3(new_n1360), .ZN(new_n1410));
  NAND2_X1  g1210(.A1(new_n1410), .A2(new_n1385), .ZN(new_n1411));
  NOR2_X1   g1211(.A1(new_n1405), .A2(new_n1411), .ZN(new_n1412));
  OAI21_X1  g1212(.A(KEYINPUT126), .B1(new_n1399), .B2(new_n1412), .ZN(new_n1413));
  INV_X1    g1213(.A(new_n1402), .ZN(new_n1414));
  AOI21_X1  g1214(.A(new_n1414), .B1(new_n1347), .B2(new_n1350), .ZN(new_n1415));
  NAND4_X1  g1215(.A1(new_n1415), .A2(new_n1385), .A3(new_n1410), .A4(new_n1401), .ZN(new_n1416));
  INV_X1    g1216(.A(KEYINPUT126), .ZN(new_n1417));
  AND3_X1   g1217(.A1(new_n1384), .A2(KEYINPUT125), .A3(new_n1385), .ZN(new_n1418));
  NOR3_X1   g1218(.A1(new_n1418), .A2(new_n1386), .A3(new_n1396), .ZN(new_n1419));
  OAI211_X1 g1219(.A(new_n1416), .B(new_n1417), .C1(new_n1351), .C2(new_n1419), .ZN(new_n1420));
  NAND2_X1  g1220(.A1(new_n1413), .A2(new_n1420), .ZN(G405));
  NAND2_X1  g1221(.A1(G375), .A2(new_n1329), .ZN(new_n1422));
  NAND4_X1  g1222(.A1(new_n1422), .A2(new_n1377), .A3(new_n1372), .A4(new_n1352), .ZN(new_n1423));
  OR2_X1    g1223(.A1(new_n1423), .A2(KEYINPUT127), .ZN(new_n1424));
  AOI21_X1  g1224(.A(new_n1387), .B1(new_n1422), .B2(new_n1352), .ZN(new_n1425));
  NAND2_X1  g1225(.A1(new_n1423), .A2(KEYINPUT127), .ZN(new_n1426));
  OAI21_X1  g1226(.A(new_n1424), .B1(new_n1425), .B2(new_n1426), .ZN(new_n1427));
  XNOR2_X1  g1227(.A(new_n1427), .B(new_n1351), .ZN(G402));
endmodule


