//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 0 0 0 0 0 0 1 0 1 1 0 1 0 0 1 1 0 0 0 0 0 1 0 0 1 1 0 0 0 0 0 0 0 1 0 1 0 0 1 0 0 0 1 1 1 1 1 1 1 1 0 0 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:10 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n555, new_n557, new_n558,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n576, new_n577, new_n578, new_n580, new_n581, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n622, new_n625,
    new_n626, new_n628, new_n629, new_n630, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n836,
    new_n837, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n962, new_n963, new_n964, new_n965, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1224, new_n1225, new_n1226;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT64), .B(G96), .Z(G221));
  XOR2_X1   g012(.A(KEYINPUT65), .B(G69), .Z(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  AOI22_X1  g030(.A1(new_n451), .A2(G2106), .B1(G567), .B2(new_n453), .ZN(new_n456));
  XOR2_X1   g031(.A(new_n456), .B(KEYINPUT66), .Z(G319));
  INV_X1    g032(.A(G2104), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n458), .A2(KEYINPUT3), .ZN(new_n459));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G2104), .ZN(new_n461));
  NAND3_X1  g036(.A1(new_n459), .A2(new_n461), .A3(G137), .ZN(new_n462));
  NAND2_X1  g037(.A1(G101), .A2(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(G2105), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n459), .A2(new_n461), .A3(G125), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(KEYINPUT67), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT67), .ZN(new_n467));
  NAND4_X1  g042(.A1(new_n459), .A2(new_n461), .A3(new_n467), .A4(G125), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT68), .ZN(new_n470));
  XNOR2_X1  g045(.A(new_n469), .B(new_n470), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n466), .A2(new_n468), .A3(new_n471), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n464), .B1(new_n472), .B2(G2105), .ZN(G160));
  NAND2_X1  g048(.A1(new_n459), .A2(new_n461), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT69), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  XNOR2_X1  g051(.A(KEYINPUT3), .B(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(KEYINPUT69), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n476), .A2(new_n478), .A3(G2105), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  INV_X1    g056(.A(G2105), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n476), .A2(new_n478), .A3(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G136), .ZN(new_n485));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n482), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n481), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  INV_X1    g064(.A(G138), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n490), .A2(G2105), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n491), .A2(new_n459), .A3(new_n461), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(KEYINPUT4), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n477), .A2(new_n494), .A3(new_n491), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n459), .A2(new_n461), .A3(G126), .ZN(new_n497));
  NAND2_X1  g072(.A1(G114), .A2(G2104), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(G2105), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n482), .A2(G102), .A3(G2104), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n496), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(G164));
  INV_X1    g078(.A(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(KEYINPUT5), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT5), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(G543), .ZN(new_n507));
  AND2_X1   g082(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  XNOR2_X1  g083(.A(KEYINPUT6), .B(G651), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G88), .ZN(new_n511));
  INV_X1    g086(.A(G50), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n509), .A2(G543), .ZN(new_n513));
  OAI22_X1  g088(.A1(new_n510), .A2(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT70), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n508), .A2(new_n515), .A3(G62), .ZN(new_n516));
  NAND2_X1  g091(.A1(G75), .A2(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n505), .A2(new_n507), .ZN(new_n518));
  INV_X1    g093(.A(G62), .ZN(new_n519));
  OAI21_X1  g094(.A(KEYINPUT70), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n516), .A2(new_n517), .A3(new_n520), .ZN(new_n521));
  AOI21_X1  g096(.A(new_n514), .B1(G651), .B2(new_n521), .ZN(G166));
  NAND2_X1  g097(.A1(new_n513), .A2(KEYINPUT71), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT71), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n509), .A2(new_n524), .A3(G543), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G51), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n508), .A2(G63), .A3(G651), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n508), .A2(G89), .A3(new_n509), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT72), .ZN(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n531), .B(KEYINPUT7), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n529), .A2(new_n530), .A3(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(new_n533), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n530), .B1(new_n529), .B2(new_n532), .ZN(new_n535));
  OAI211_X1 g110(.A(new_n527), .B(new_n528), .C1(new_n534), .C2(new_n535), .ZN(G286));
  INV_X1    g111(.A(G286), .ZN(G168));
  NAND2_X1  g112(.A1(new_n526), .A2(G52), .ZN(new_n538));
  INV_X1    g113(.A(new_n510), .ZN(new_n539));
  NAND2_X1  g114(.A1(G77), .A2(G543), .ZN(new_n540));
  INV_X1    g115(.A(G64), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n540), .B1(new_n518), .B2(new_n541), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n539), .A2(G90), .B1(G651), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n538), .A2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(new_n544), .ZN(G171));
  AND2_X1   g120(.A1(new_n526), .A2(G43), .ZN(new_n546));
  NAND2_X1  g121(.A1(G68), .A2(G543), .ZN(new_n547));
  INV_X1    g122(.A(G56), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n547), .B1(new_n518), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G651), .ZN(new_n550));
  INV_X1    g125(.A(G81), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n550), .B1(new_n551), .B2(new_n510), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n546), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G860), .ZN(G153));
  AND3_X1   g129(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G36), .ZN(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n555), .A2(new_n558), .ZN(G188));
  XNOR2_X1  g134(.A(KEYINPUT73), .B(KEYINPUT9), .ZN(new_n560));
  INV_X1    g135(.A(G53), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n560), .B1(new_n513), .B2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT9), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n563), .A2(KEYINPUT73), .ZN(new_n564));
  NAND4_X1  g139(.A1(new_n509), .A2(G53), .A3(G543), .A4(new_n564), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n508), .A2(G91), .A3(new_n509), .ZN(new_n566));
  AND3_X1   g141(.A1(new_n562), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT74), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n505), .A2(new_n507), .A3(G65), .ZN(new_n569));
  NAND2_X1  g144(.A1(G78), .A2(G543), .ZN(new_n570));
  AOI21_X1  g145(.A(new_n568), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(new_n571), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n569), .A2(new_n568), .A3(new_n570), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n572), .A2(G651), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n567), .A2(new_n574), .ZN(G299));
  NAND2_X1  g150(.A1(new_n544), .A2(KEYINPUT75), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT75), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n538), .A2(new_n543), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n576), .A2(new_n578), .ZN(G301));
  NAND2_X1  g154(.A1(new_n521), .A2(G651), .ZN(new_n580));
  INV_X1    g155(.A(new_n514), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(new_n581), .ZN(G303));
  OAI21_X1  g157(.A(G651), .B1(new_n508), .B2(G74), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n509), .A2(G49), .A3(G543), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n508), .A2(G87), .A3(new_n509), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(G288));
  INV_X1    g161(.A(KEYINPUT76), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n508), .A2(new_n587), .A3(G61), .ZN(new_n588));
  NAND2_X1  g163(.A1(G73), .A2(G543), .ZN(new_n589));
  INV_X1    g164(.A(G61), .ZN(new_n590));
  OAI21_X1  g165(.A(KEYINPUT76), .B1(new_n518), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n588), .A2(new_n589), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n592), .A2(G651), .ZN(new_n593));
  INV_X1    g168(.A(G86), .ZN(new_n594));
  INV_X1    g169(.A(G48), .ZN(new_n595));
  OAI22_X1  g170(.A1(new_n510), .A2(new_n594), .B1(new_n595), .B2(new_n513), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n593), .A2(new_n597), .ZN(G305));
  XNOR2_X1  g173(.A(KEYINPUT77), .B(G47), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n526), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(G72), .A2(G543), .ZN(new_n601));
  INV_X1    g176(.A(G60), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n518), .B2(new_n602), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n539), .A2(G85), .B1(G651), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n600), .A2(new_n604), .ZN(G290));
  XOR2_X1   g180(.A(KEYINPUT78), .B(KEYINPUT10), .Z(new_n606));
  INV_X1    g181(.A(new_n606), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n539), .A2(G92), .A3(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(G92), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n606), .B1(new_n510), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n526), .A2(G54), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n508), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n613));
  INV_X1    g188(.A(G651), .ZN(new_n614));
  OR2_X1    g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n611), .A2(new_n612), .A3(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(G868), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(G301), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n619), .B2(new_n617), .ZN(G284));
  OAI21_X1  g195(.A(new_n618), .B1(new_n619), .B2(new_n617), .ZN(G321));
  NAND2_X1  g196(.A1(G299), .A2(new_n617), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(G168), .B2(new_n617), .ZN(G297));
  OAI21_X1  g198(.A(new_n622), .B1(G168), .B2(new_n617), .ZN(G280));
  INV_X1    g199(.A(new_n616), .ZN(new_n625));
  INV_X1    g200(.A(G559), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n625), .B1(new_n626), .B2(G860), .ZN(G148));
  INV_X1    g202(.A(new_n553), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(new_n617), .ZN(new_n629));
  NOR2_X1   g204(.A1(new_n616), .A2(G559), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n629), .B1(new_n630), .B2(new_n617), .ZN(G323));
  XNOR2_X1  g206(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g207(.A1(new_n480), .A2(G123), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n484), .A2(G135), .ZN(new_n634));
  NOR2_X1   g209(.A1(G99), .A2(G2105), .ZN(new_n635));
  OAI21_X1  g210(.A(G2104), .B1(new_n482), .B2(G111), .ZN(new_n636));
  OAI211_X1 g211(.A(new_n633), .B(new_n634), .C1(new_n635), .C2(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(G2096), .Z(new_n638));
  NAND3_X1  g213(.A1(new_n482), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT12), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT13), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2100), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n638), .A2(new_n642), .ZN(G156));
  XNOR2_X1  g218(.A(G2451), .B(G2454), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT16), .ZN(new_n645));
  XOR2_X1   g220(.A(G2443), .B(G2446), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G1341), .B(G1348), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(KEYINPUT15), .B(G2435), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(G2438), .ZN(new_n651));
  XOR2_X1   g226(.A(G2427), .B(G2430), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT79), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n651), .B(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n654), .A2(KEYINPUT14), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n649), .B(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n656), .A2(G14), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(G401));
  XNOR2_X1  g233(.A(G2067), .B(G2678), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT80), .ZN(new_n660));
  XOR2_X1   g235(.A(G2084), .B(G2090), .Z(new_n661));
  XNOR2_X1  g236(.A(G2072), .B(G2078), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n660), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n663), .B(KEYINPUT81), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT18), .ZN(new_n665));
  INV_X1    g240(.A(KEYINPUT17), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n660), .B(KEYINPUT82), .ZN(new_n667));
  INV_X1    g242(.A(new_n661), .ZN(new_n668));
  AOI21_X1  g243(.A(new_n666), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n669), .B(new_n662), .Z(new_n670));
  OR2_X1    g245(.A1(new_n667), .A2(new_n668), .ZN(new_n671));
  AOI21_X1  g246(.A(new_n665), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G2096), .B(G2100), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(G227));
  INV_X1    g249(.A(KEYINPUT20), .ZN(new_n675));
  XOR2_X1   g250(.A(G1961), .B(G1966), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT83), .ZN(new_n677));
  XOR2_X1   g252(.A(G1956), .B(G2474), .Z(new_n678));
  NAND2_X1  g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1971), .B(G1976), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT19), .ZN(new_n681));
  OAI21_X1  g256(.A(new_n675), .B1(new_n679), .B2(new_n681), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n677), .A2(new_n678), .ZN(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n684), .A2(new_n681), .A3(new_n679), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n679), .A2(new_n675), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n686), .A2(new_n683), .ZN(new_n687));
  OAI211_X1 g262(.A(new_n682), .B(new_n685), .C1(new_n687), .C2(new_n681), .ZN(new_n688));
  XOR2_X1   g263(.A(G1991), .B(G1996), .Z(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n688), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT84), .B(G1986), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(G1981), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n692), .B(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(G229));
  MUX2_X1   g271(.A(G24), .B(G290), .S(G16), .Z(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(G1986), .ZN(new_n698));
  INV_X1    g273(.A(G16), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G23), .ZN(new_n700));
  AND3_X1   g275(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n700), .B1(new_n701), .B2(new_n699), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT33), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(G1976), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n699), .A2(G22), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(G166), .B2(new_n699), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT85), .B(G1971), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n699), .A2(G6), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n596), .B1(G651), .B2(new_n592), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n709), .B1(new_n710), .B2(new_n699), .ZN(new_n711));
  XOR2_X1   g286(.A(KEYINPUT32), .B(G1981), .Z(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n704), .A2(new_n708), .A3(new_n713), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n698), .B1(new_n714), .B2(KEYINPUT34), .ZN(new_n715));
  INV_X1    g290(.A(G29), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(G25), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n480), .A2(G119), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n484), .A2(G131), .ZN(new_n719));
  OR2_X1    g294(.A1(G95), .A2(G2105), .ZN(new_n720));
  OAI211_X1 g295(.A(new_n720), .B(G2104), .C1(G107), .C2(new_n482), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n718), .A2(new_n719), .A3(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n717), .B1(new_n723), .B2(new_n716), .ZN(new_n724));
  XNOR2_X1  g299(.A(KEYINPUT35), .B(G1991), .ZN(new_n725));
  INV_X1    g300(.A(new_n725), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n724), .B(new_n726), .ZN(new_n727));
  OAI211_X1 g302(.A(new_n715), .B(new_n727), .C1(KEYINPUT34), .C2(new_n714), .ZN(new_n728));
  INV_X1    g303(.A(KEYINPUT86), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n729), .A2(KEYINPUT36), .ZN(new_n730));
  OR2_X1    g305(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(KEYINPUT92), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(G16), .B2(G21), .ZN(new_n733));
  NOR2_X1   g308(.A1(G286), .A2(new_n699), .ZN(new_n734));
  MUX2_X1   g309(.A(new_n733), .B(new_n732), .S(new_n734), .Z(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(G1966), .ZN(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT31), .B(G11), .ZN(new_n737));
  INV_X1    g312(.A(KEYINPUT30), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n716), .B1(new_n738), .B2(G28), .ZN(new_n739));
  OR2_X1    g314(.A1(new_n739), .A2(KEYINPUT93), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n738), .A2(G28), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n739), .A2(KEYINPUT93), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n740), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(new_n637), .B2(new_n716), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n699), .A2(G5), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(G171), .B2(new_n699), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT94), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n744), .B1(new_n747), .B2(G1961), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n736), .A2(new_n737), .A3(new_n748), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT95), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n716), .A2(G27), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(G164), .B2(new_n716), .ZN(new_n752));
  XNOR2_X1  g327(.A(KEYINPUT96), .B(G2078), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n752), .B(new_n753), .ZN(new_n754));
  OR2_X1    g329(.A1(new_n747), .A2(G1961), .ZN(new_n755));
  NAND2_X1  g330(.A1(G115), .A2(G2104), .ZN(new_n756));
  INV_X1    g331(.A(G127), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n756), .B1(new_n474), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n758), .A2(G2105), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n482), .A2(G103), .A3(G2104), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT25), .Z(new_n761));
  INV_X1    g336(.A(G139), .ZN(new_n762));
  OAI211_X1 g337(.A(new_n759), .B(new_n761), .C1(new_n483), .C2(new_n762), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT88), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n764), .A2(new_n716), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(new_n716), .B2(G33), .ZN(new_n766));
  INV_X1    g341(.A(G2072), .ZN(new_n767));
  OR2_X1    g342(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(G2084), .ZN(new_n769));
  XOR2_X1   g344(.A(KEYINPUT89), .B(KEYINPUT24), .Z(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(G34), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n771), .A2(new_n716), .ZN(new_n772));
  INV_X1    g347(.A(G160), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n772), .B1(new_n773), .B2(new_n716), .ZN(new_n774));
  AOI22_X1  g349(.A1(new_n766), .A2(new_n767), .B1(new_n769), .B2(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n716), .A2(G35), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(G162), .B2(new_n716), .ZN(new_n777));
  XOR2_X1   g352(.A(KEYINPUT29), .B(G2090), .Z(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NAND4_X1  g354(.A1(new_n755), .A2(new_n768), .A3(new_n775), .A4(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(KEYINPUT28), .ZN(new_n781));
  INV_X1    g356(.A(G26), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n781), .B1(new_n782), .B2(G29), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n782), .A2(G29), .ZN(new_n784));
  OR2_X1    g359(.A1(G104), .A2(G2105), .ZN(new_n785));
  OAI211_X1 g360(.A(new_n785), .B(G2104), .C1(G116), .C2(new_n482), .ZN(new_n786));
  INV_X1    g361(.A(G128), .ZN(new_n787));
  INV_X1    g362(.A(G140), .ZN(new_n788));
  OAI221_X1 g363(.A(new_n786), .B1(new_n479), .B2(new_n787), .C1(new_n788), .C2(new_n483), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n784), .B1(new_n789), .B2(G29), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n783), .B1(new_n790), .B2(new_n781), .ZN(new_n791));
  OR2_X1    g366(.A1(new_n791), .A2(G2067), .ZN(new_n792));
  INV_X1    g367(.A(new_n792), .ZN(new_n793));
  INV_X1    g368(.A(G19), .ZN(new_n794));
  OAI21_X1  g369(.A(KEYINPUT87), .B1(new_n794), .B2(G16), .ZN(new_n795));
  OR3_X1    g370(.A1(new_n794), .A2(KEYINPUT87), .A3(G16), .ZN(new_n796));
  OAI211_X1 g371(.A(new_n795), .B(new_n796), .C1(new_n553), .C2(new_n699), .ZN(new_n797));
  XOR2_X1   g372(.A(new_n797), .B(G1341), .Z(new_n798));
  NAND2_X1  g373(.A1(new_n699), .A2(G4), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(new_n625), .B2(new_n699), .ZN(new_n800));
  INV_X1    g375(.A(G1348), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n800), .B(new_n801), .ZN(new_n802));
  OR2_X1    g377(.A1(new_n774), .A2(new_n769), .ZN(new_n803));
  AND3_X1   g378(.A1(new_n699), .A2(KEYINPUT23), .A3(G20), .ZN(new_n804));
  INV_X1    g379(.A(new_n573), .ZN(new_n805));
  NOR3_X1   g380(.A1(new_n805), .A2(new_n571), .A3(new_n614), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n562), .A2(new_n565), .A3(new_n566), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  OAI21_X1  g383(.A(KEYINPUT23), .B1(new_n808), .B2(new_n699), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n699), .A2(G20), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n804), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(G1956), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND4_X1  g388(.A1(new_n798), .A2(new_n802), .A3(new_n803), .A4(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n791), .A2(G2067), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(new_n811), .B2(new_n812), .ZN(new_n816));
  NOR4_X1   g391(.A1(new_n780), .A2(new_n793), .A3(new_n814), .A4(new_n816), .ZN(new_n817));
  NAND4_X1  g392(.A1(new_n731), .A2(new_n750), .A3(new_n754), .A4(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n484), .A2(G141), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n480), .A2(G129), .ZN(new_n820));
  NAND3_X1  g395(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n821));
  XOR2_X1   g396(.A(new_n821), .B(KEYINPUT26), .Z(new_n822));
  NAND3_X1  g397(.A1(new_n482), .A2(G105), .A3(G2104), .ZN(new_n823));
  NAND4_X1  g398(.A1(new_n819), .A2(new_n820), .A3(new_n822), .A4(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n825), .A2(G29), .ZN(new_n826));
  OAI211_X1 g401(.A(new_n826), .B(KEYINPUT90), .C1(G29), .C2(G32), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n827), .B1(KEYINPUT90), .B2(new_n826), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n828), .B(KEYINPUT91), .Z(new_n829));
  XOR2_X1   g404(.A(KEYINPUT27), .B(G1996), .Z(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(KEYINPUT86), .B(KEYINPUT36), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n728), .A2(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(new_n833), .ZN(new_n834));
  NOR3_X1   g409(.A1(new_n818), .A2(new_n831), .A3(new_n834), .ZN(G311));
  AND3_X1   g410(.A1(new_n750), .A2(new_n754), .A3(new_n817), .ZN(new_n836));
  INV_X1    g411(.A(new_n831), .ZN(new_n837));
  NAND4_X1  g412(.A1(new_n836), .A2(new_n837), .A3(new_n833), .A4(new_n731), .ZN(G150));
  NAND2_X1  g413(.A1(new_n526), .A2(G55), .ZN(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(new_n840));
  AOI22_X1  g415(.A1(new_n508), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n841));
  INV_X1    g416(.A(G93), .ZN(new_n842));
  OAI22_X1  g417(.A1(new_n841), .A2(new_n614), .B1(new_n842), .B2(new_n510), .ZN(new_n843));
  NOR3_X1   g418(.A1(new_n840), .A2(KEYINPUT97), .A3(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT97), .ZN(new_n845));
  INV_X1    g420(.A(new_n843), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n845), .B1(new_n846), .B2(new_n839), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n844), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(G860), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(KEYINPUT99), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT37), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n625), .A2(G559), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT38), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n628), .B1(new_n844), .B2(new_n847), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n553), .B1(new_n840), .B2(new_n843), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n853), .B(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n857), .A2(KEYINPUT39), .ZN(new_n858));
  AOI21_X1  g433(.A(G860), .B1(new_n858), .B2(KEYINPUT98), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n859), .B1(KEYINPUT98), .B2(new_n858), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n857), .A2(KEYINPUT39), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n851), .B1(new_n860), .B2(new_n861), .ZN(G145));
  XNOR2_X1  g437(.A(new_n789), .B(G164), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT88), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n763), .B(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n865), .A2(KEYINPUT100), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT100), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n764), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n863), .A2(new_n866), .A3(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n863), .B1(new_n866), .B2(new_n868), .ZN(new_n871));
  NOR3_X1   g446(.A1(new_n870), .A2(new_n871), .A3(new_n824), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n866), .A2(new_n868), .ZN(new_n873));
  INV_X1    g448(.A(new_n863), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n825), .B1(new_n875), .B2(new_n869), .ZN(new_n876));
  OAI21_X1  g451(.A(KEYINPUT102), .B1(new_n872), .B2(new_n876), .ZN(new_n877));
  OR2_X1    g452(.A1(G106), .A2(G2105), .ZN(new_n878));
  OAI211_X1 g453(.A(new_n878), .B(G2104), .C1(G118), .C2(new_n482), .ZN(new_n879));
  INV_X1    g454(.A(G130), .ZN(new_n880));
  INV_X1    g455(.A(G142), .ZN(new_n881));
  OAI221_X1 g456(.A(new_n879), .B1(new_n479), .B2(new_n880), .C1(new_n881), .C2(new_n483), .ZN(new_n882));
  INV_X1    g457(.A(new_n640), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n480), .A2(G130), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n484), .A2(G142), .ZN(new_n886));
  NAND4_X1  g461(.A1(new_n885), .A2(new_n886), .A3(new_n640), .A4(new_n879), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n723), .A2(new_n884), .A3(new_n887), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n824), .B1(new_n870), .B2(new_n871), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT102), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n875), .A2(new_n825), .A3(new_n869), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n723), .B1(new_n884), .B2(new_n887), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  NAND4_X1  g469(.A1(new_n877), .A2(new_n888), .A3(new_n892), .A4(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n894), .A2(KEYINPUT101), .A3(new_n888), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT101), .ZN(new_n897));
  INV_X1    g472(.A(new_n888), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n897), .B1(new_n898), .B2(new_n893), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n896), .A2(new_n899), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n900), .B1(new_n872), .B2(new_n876), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n637), .B(new_n773), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n902), .B(new_n488), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n895), .A2(new_n901), .A3(new_n904), .ZN(new_n905));
  NAND4_X1  g480(.A1(new_n889), .A2(new_n896), .A3(new_n891), .A4(new_n899), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n901), .A2(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(G37), .B1(new_n907), .B2(new_n903), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n905), .A2(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n909), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g485(.A(G303), .B(KEYINPUT104), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n911), .A2(new_n710), .ZN(new_n912));
  XNOR2_X1  g487(.A(G166), .B(KEYINPUT104), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n913), .A2(G305), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(G290), .A2(new_n701), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n600), .A2(new_n604), .A3(G288), .ZN(new_n917));
  AND3_X1   g492(.A1(new_n916), .A2(KEYINPUT105), .A3(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(KEYINPUT105), .B1(new_n916), .B2(new_n917), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n915), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n912), .A2(new_n914), .A3(new_n919), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  OAI211_X1 g498(.A(new_n854), .B(new_n855), .C1(G559), .C2(new_n616), .ZN(new_n924));
  INV_X1    g499(.A(new_n855), .ZN(new_n925));
  OAI21_X1  g500(.A(KEYINPUT97), .B1(new_n840), .B2(new_n843), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n846), .A2(new_n845), .A3(new_n839), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n553), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n630), .B1(new_n925), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n924), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT41), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n616), .A2(G299), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n808), .A2(new_n611), .A3(new_n612), .A4(new_n615), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n931), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(KEYINPUT103), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n932), .A2(new_n933), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(KEYINPUT41), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT103), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n932), .A2(new_n933), .A3(new_n931), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n937), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n930), .B1(new_n935), .B2(new_n940), .ZN(new_n941));
  XNOR2_X1  g516(.A(KEYINPUT106), .B(KEYINPUT42), .ZN(new_n942));
  INV_X1    g517(.A(new_n936), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n943), .B1(new_n924), .B2(new_n929), .ZN(new_n944));
  NOR3_X1   g519(.A1(new_n941), .A2(new_n942), .A3(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(new_n942), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n940), .A2(new_n935), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n947), .A2(new_n929), .A3(new_n924), .ZN(new_n948));
  INV_X1    g523(.A(new_n944), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n946), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n923), .B1(new_n945), .B2(new_n950), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n942), .B1(new_n941), .B2(new_n944), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n948), .A2(new_n946), .A3(new_n949), .ZN(new_n953));
  INV_X1    g528(.A(new_n923), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n952), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n951), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(G868), .ZN(new_n957));
  INV_X1    g532(.A(new_n848), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n958), .A2(G868), .ZN(new_n959));
  INV_X1    g534(.A(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n957), .A2(new_n960), .ZN(G295));
  INV_X1    g536(.A(KEYINPUT107), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n957), .A2(new_n962), .A3(new_n960), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n617), .B1(new_n951), .B2(new_n955), .ZN(new_n964));
  OAI21_X1  g539(.A(KEYINPUT107), .B1(new_n964), .B2(new_n959), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n963), .A2(new_n965), .ZN(G331));
  INV_X1    g541(.A(KEYINPUT44), .ZN(new_n967));
  NOR2_X1   g542(.A1(G168), .A2(new_n544), .ZN(new_n968));
  AOI21_X1  g543(.A(G286), .B1(new_n576), .B2(new_n578), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(new_n856), .ZN(new_n971));
  OAI211_X1 g546(.A(new_n854), .B(new_n855), .C1(new_n968), .C2(new_n969), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n936), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(new_n947), .ZN(new_n974));
  AND2_X1   g549(.A1(new_n971), .A2(new_n972), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n973), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  AOI21_X1  g551(.A(G37), .B1(new_n976), .B2(new_n954), .ZN(new_n977));
  AOI21_X1  g552(.A(KEYINPUT109), .B1(new_n921), .B2(new_n922), .ZN(new_n978));
  INV_X1    g553(.A(new_n978), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n921), .A2(KEYINPUT109), .A3(new_n922), .ZN(new_n980));
  AND2_X1   g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT110), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n973), .A2(new_n982), .ZN(new_n983));
  AOI211_X1 g558(.A(KEYINPUT110), .B(new_n936), .C1(new_n971), .C2(new_n972), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n937), .A2(new_n939), .ZN(new_n985));
  AND3_X1   g560(.A1(new_n971), .A2(new_n985), .A3(new_n972), .ZN(new_n986));
  NOR3_X1   g561(.A1(new_n983), .A2(new_n984), .A3(new_n986), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n977), .B1(new_n981), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n988), .A2(KEYINPUT43), .ZN(new_n989));
  XOR2_X1   g564(.A(KEYINPUT108), .B(KEYINPUT43), .Z(new_n990));
  INV_X1    g565(.A(new_n990), .ZN(new_n991));
  OAI211_X1 g566(.A(new_n977), .B(new_n991), .C1(new_n976), .C2(new_n981), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n967), .B1(new_n989), .B2(new_n992), .ZN(new_n993));
  OAI211_X1 g568(.A(new_n977), .B(new_n991), .C1(new_n987), .C2(new_n981), .ZN(new_n994));
  INV_X1    g569(.A(G37), .ZN(new_n995));
  INV_X1    g570(.A(new_n973), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n940), .A2(new_n971), .A3(new_n935), .A4(new_n972), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n995), .B1(new_n998), .B2(new_n923), .ZN(new_n999));
  AOI22_X1  g574(.A1(new_n979), .A2(new_n980), .B1(new_n996), .B2(new_n997), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n990), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  AND3_X1   g576(.A1(new_n994), .A2(new_n1001), .A3(new_n967), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n993), .A2(new_n1002), .ZN(G397));
  XNOR2_X1  g578(.A(KEYINPUT112), .B(KEYINPUT45), .ZN(new_n1004));
  XOR2_X1   g579(.A(KEYINPUT111), .B(G1384), .Z(new_n1005));
  AOI21_X1  g580(.A(new_n1004), .B1(new_n502), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(G40), .ZN(new_n1007));
  AOI211_X1 g582(.A(new_n1007), .B(new_n464), .C1(new_n472), .C2(G2105), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  NOR3_X1   g584(.A1(new_n1009), .A2(G1986), .A3(G290), .ZN(new_n1010));
  XOR2_X1   g585(.A(new_n1010), .B(KEYINPUT48), .Z(new_n1011));
  INV_X1    g586(.A(G1996), .ZN(new_n1012));
  XNOR2_X1  g587(.A(new_n824), .B(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(G2067), .ZN(new_n1014));
  XNOR2_X1  g589(.A(new_n789), .B(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1016), .B1(new_n725), .B2(new_n722), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n723), .A2(new_n726), .ZN(new_n1018));
  AND2_X1   g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1011), .B1(new_n1019), .B2(new_n1009), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1009), .B1(new_n1015), .B2(new_n825), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1009), .ZN(new_n1022));
  AND3_X1   g597(.A1(new_n1022), .A2(KEYINPUT46), .A3(new_n1012), .ZN(new_n1023));
  AOI21_X1  g598(.A(KEYINPUT46), .B1(new_n1022), .B2(new_n1012), .ZN(new_n1024));
  NOR3_X1   g599(.A1(new_n1021), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1025));
  XOR2_X1   g600(.A(new_n1025), .B(KEYINPUT47), .Z(new_n1026));
  OAI22_X1  g601(.A1(new_n1016), .A2(new_n1018), .B1(G2067), .B2(new_n789), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(new_n1022), .ZN(new_n1028));
  AND3_X1   g603(.A1(new_n1020), .A2(new_n1026), .A3(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(G1966), .ZN(new_n1030));
  INV_X1    g605(.A(G1384), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n502), .A2(new_n1031), .A3(new_n1004), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(new_n1008), .ZN(new_n1033));
  AOI21_X1  g608(.A(KEYINPUT45), .B1(new_n502), .B2(new_n1031), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1030), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n502), .A2(new_n1031), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(KEYINPUT50), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT50), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n502), .A2(new_n1038), .A3(new_n1031), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n1037), .A2(new_n769), .A3(new_n1008), .A4(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1035), .A2(new_n1040), .ZN(new_n1041));
  XNOR2_X1  g616(.A(KEYINPUT113), .B(G8), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT124), .ZN(new_n1044));
  AOI21_X1  g619(.A(KEYINPUT51), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1042), .ZN(new_n1046));
  NOR2_X1   g621(.A1(G168), .A2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1046), .B1(new_n1035), .B2(new_n1040), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1047), .B1(new_n1048), .B2(KEYINPUT124), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1047), .ZN(new_n1050));
  AND3_X1   g625(.A1(new_n502), .A2(new_n1038), .A3(new_n1031), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1038), .B1(new_n502), .B2(new_n1031), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n472), .A2(G2105), .ZN(new_n1053));
  INV_X1    g628(.A(new_n464), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1053), .A2(G40), .A3(new_n1054), .ZN(new_n1055));
  NOR3_X1   g630(.A1(new_n1051), .A2(new_n1052), .A3(new_n1055), .ZN(new_n1056));
  AOI22_X1  g631(.A1(new_n493), .A2(new_n495), .B1(new_n499), .B2(G2105), .ZN(new_n1057));
  AOI21_X1  g632(.A(G1384), .B1(new_n1057), .B2(new_n501), .ZN(new_n1058));
  OAI211_X1 g633(.A(new_n1032), .B(new_n1008), .C1(new_n1058), .C2(KEYINPUT45), .ZN(new_n1059));
  AOI22_X1  g634(.A1(new_n1056), .A2(new_n769), .B1(new_n1030), .B2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(G8), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1050), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  AOI22_X1  g637(.A1(new_n1045), .A2(new_n1049), .B1(KEYINPUT51), .B2(new_n1062), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1060), .A2(new_n1050), .ZN(new_n1064));
  OAI21_X1  g639(.A(KEYINPUT62), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g640(.A(KEYINPUT125), .B1(new_n1059), .B2(G2078), .ZN(new_n1066));
  AND2_X1   g641(.A1(new_n1032), .A2(new_n1008), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT125), .ZN(new_n1068));
  INV_X1    g643(.A(G2078), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1034), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1067), .A2(new_n1068), .A3(new_n1069), .A4(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1066), .A2(new_n1071), .A3(KEYINPUT53), .ZN(new_n1072));
  OR2_X1    g647(.A1(new_n1056), .A2(G1961), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(KEYINPUT126), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT126), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1072), .A2(new_n1076), .A3(new_n1073), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1075), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT53), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1004), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1036), .A2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n502), .A2(KEYINPUT45), .A3(new_n1005), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1081), .A2(new_n1008), .A3(new_n1082), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1079), .B1(new_n1083), .B2(G2078), .ZN(new_n1084));
  AOI21_X1  g659(.A(G301), .B1(new_n1078), .B2(new_n1084), .ZN(new_n1085));
  OAI21_X1  g660(.A(KEYINPUT55), .B1(G166), .B2(new_n1061), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT55), .ZN(new_n1087));
  NAND3_X1  g662(.A1(G303), .A2(new_n1087), .A3(G8), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(G2090), .ZN(new_n1090));
  INV_X1    g665(.A(G1971), .ZN(new_n1091));
  AOI22_X1  g666(.A1(new_n1056), .A2(new_n1090), .B1(new_n1083), .B2(new_n1091), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1089), .B1(new_n1092), .B2(new_n1046), .ZN(new_n1093));
  NAND2_X1  g668(.A1(G305), .A2(G1981), .ZN(new_n1094));
  INV_X1    g669(.A(G1981), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n710), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(KEYINPUT49), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT49), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1094), .A2(new_n1096), .A3(new_n1099), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1042), .B1(new_n1055), .B2(new_n1036), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT114), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NAND4_X1  g678(.A1(G160), .A2(G40), .A3(new_n502), .A4(new_n1031), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1104), .A2(KEYINPUT114), .A3(new_n1042), .ZN(new_n1105));
  AOI22_X1  g680(.A1(new_n1098), .A2(new_n1100), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n701), .A2(G1976), .ZN(new_n1107));
  XNOR2_X1  g682(.A(new_n1107), .B(KEYINPUT115), .ZN(new_n1108));
  INV_X1    g683(.A(G1976), .ZN(new_n1109));
  AOI21_X1  g684(.A(KEYINPUT52), .B1(G288), .B2(new_n1109), .ZN(new_n1110));
  XNOR2_X1  g685(.A(new_n1110), .B(KEYINPUT116), .ZN(new_n1111));
  AND3_X1   g686(.A1(new_n1104), .A2(KEYINPUT114), .A3(new_n1042), .ZN(new_n1112));
  AOI21_X1  g687(.A(KEYINPUT114), .B1(new_n1104), .B2(new_n1042), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n1108), .B(new_n1111), .C1(new_n1112), .C2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(KEYINPUT117), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT117), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1116), .A2(new_n1117), .A3(new_n1108), .A4(new_n1111), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1106), .B1(new_n1115), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1083), .A2(new_n1091), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1037), .A2(new_n1090), .A3(new_n1008), .A4(new_n1039), .ZN(new_n1121));
  AOI211_X1 g696(.A(new_n1061), .B(new_n1089), .C1(new_n1120), .C2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1116), .A2(new_n1108), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(KEYINPUT52), .ZN(new_n1125));
  AND4_X1   g700(.A1(new_n1093), .A2(new_n1119), .A3(new_n1123), .A4(new_n1125), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1061), .B1(new_n1035), .B2(new_n1040), .ZN(new_n1127));
  OAI21_X1  g702(.A(KEYINPUT51), .B1(new_n1127), .B2(new_n1047), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1050), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT51), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1130), .B1(new_n1048), .B2(KEYINPUT124), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1128), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT62), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1064), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1132), .A2(new_n1133), .A3(new_n1134), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1065), .A2(new_n1085), .A3(new_n1126), .A4(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1106), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1137), .A2(new_n1109), .A3(new_n701), .ZN(new_n1138));
  AOI22_X1  g713(.A1(new_n1138), .A2(new_n1096), .B1(new_n1105), .B2(new_n1103), .ZN(new_n1139));
  XOR2_X1   g714(.A(KEYINPUT118), .B(KEYINPUT63), .Z(new_n1140));
  NAND2_X1  g715(.A1(new_n1115), .A2(new_n1118), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1141), .A2(new_n1125), .A3(new_n1137), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1043), .A2(G286), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1122), .B1(new_n1143), .B2(new_n1093), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1140), .B1(new_n1142), .B2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1048), .A2(KEYINPUT63), .A3(G168), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1147), .A2(G8), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1146), .B1(new_n1089), .B2(new_n1148), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n1149), .A2(new_n1123), .A3(new_n1125), .A4(new_n1119), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1139), .B1(new_n1145), .B2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1136), .A2(new_n1151), .ZN(new_n1152));
  AND2_X1   g727(.A1(new_n1084), .A2(G301), .ZN(new_n1153));
  AOI21_X1  g728(.A(KEYINPUT127), .B1(new_n1078), .B2(new_n1153), .ZN(new_n1154));
  AND3_X1   g729(.A1(new_n1072), .A2(new_n1076), .A3(new_n1073), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1076), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1156));
  OAI211_X1 g731(.A(KEYINPUT127), .B(new_n1153), .C1(new_n1155), .C2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1157), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n1154), .A2(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT54), .ZN(new_n1160));
  NOR3_X1   g735(.A1(new_n1006), .A2(new_n1079), .A3(G2078), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1161), .A2(new_n1008), .A3(new_n1082), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1073), .A2(new_n1084), .A3(new_n1162), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1160), .B1(new_n1163), .B2(G171), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT122), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT119), .ZN(new_n1166));
  OAI211_X1 g741(.A(new_n1166), .B(KEYINPUT57), .C1(new_n806), .C2(new_n807), .ZN(new_n1167));
  OR2_X1    g742(.A1(new_n1166), .A2(KEYINPUT57), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1166), .A2(KEYINPUT57), .ZN(new_n1169));
  NAND4_X1  g744(.A1(new_n567), .A2(new_n574), .A3(new_n1168), .A4(new_n1169), .ZN(new_n1170));
  AND2_X1   g745(.A1(new_n1167), .A2(new_n1170), .ZN(new_n1171));
  XNOR2_X1  g746(.A(KEYINPUT56), .B(G2072), .ZN(new_n1172));
  NAND4_X1  g747(.A1(new_n1081), .A2(new_n1008), .A3(new_n1082), .A4(new_n1172), .ZN(new_n1173));
  OAI211_X1 g748(.A(new_n1171), .B(new_n1173), .C1(new_n1056), .C2(G1956), .ZN(new_n1174));
  INV_X1    g749(.A(new_n1174), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1037), .A2(new_n1008), .A3(new_n1039), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1176), .A2(new_n812), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1171), .B1(new_n1177), .B2(new_n1173), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1165), .B1(new_n1175), .B2(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT61), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  OAI211_X1 g756(.A(new_n1165), .B(KEYINPUT61), .C1(new_n1175), .C2(new_n1178), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1176), .A2(new_n801), .ZN(new_n1184));
  INV_X1    g759(.A(KEYINPUT120), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1104), .A2(new_n1185), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n1008), .A2(new_n1058), .A3(KEYINPUT120), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1186), .A2(new_n1187), .A3(new_n1014), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1184), .A2(new_n1188), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT60), .ZN(new_n1190));
  NOR2_X1   g765(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  INV_X1    g766(.A(new_n1191), .ZN(new_n1192));
  AOI21_X1  g767(.A(new_n616), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1193));
  INV_X1    g768(.A(KEYINPUT123), .ZN(new_n1194));
  NOR2_X1   g769(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  AOI21_X1  g770(.A(KEYINPUT60), .B1(new_n1184), .B2(new_n1188), .ZN(new_n1196));
  NOR3_X1   g771(.A1(new_n1196), .A2(KEYINPUT123), .A3(new_n616), .ZN(new_n1197));
  OAI21_X1  g772(.A(new_n1192), .B1(new_n1195), .B2(new_n1197), .ZN(new_n1198));
  NOR2_X1   g773(.A1(new_n1083), .A2(G1996), .ZN(new_n1199));
  XNOR2_X1  g774(.A(KEYINPUT58), .B(G1341), .ZN(new_n1200));
  AOI21_X1  g775(.A(new_n1200), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1201));
  OAI21_X1  g776(.A(new_n553), .B1(new_n1199), .B2(new_n1201), .ZN(new_n1202));
  XNOR2_X1  g777(.A(new_n1202), .B(KEYINPUT59), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1204));
  OAI21_X1  g779(.A(KEYINPUT123), .B1(new_n1196), .B2(new_n616), .ZN(new_n1205));
  NAND3_X1  g780(.A1(new_n1204), .A2(new_n1191), .A3(new_n1205), .ZN(new_n1206));
  NAND4_X1  g781(.A1(new_n1183), .A2(new_n1198), .A3(new_n1203), .A4(new_n1206), .ZN(new_n1207));
  INV_X1    g782(.A(new_n1178), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1189), .A2(new_n625), .ZN(new_n1209));
  AOI21_X1  g784(.A(new_n1175), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  XNOR2_X1  g785(.A(new_n1210), .B(KEYINPUT121), .ZN(new_n1211));
  AOI22_X1  g786(.A1(new_n1159), .A2(new_n1164), .B1(new_n1207), .B2(new_n1211), .ZN(new_n1212));
  OAI21_X1  g787(.A(new_n1084), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1213), .A2(new_n619), .ZN(new_n1214));
  OR2_X1    g789(.A1(new_n1163), .A2(new_n619), .ZN(new_n1215));
  AOI21_X1  g790(.A(KEYINPUT54), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1216));
  OAI21_X1  g791(.A(new_n1126), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1217));
  NOR2_X1   g792(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  AOI21_X1  g793(.A(new_n1152), .B1(new_n1212), .B2(new_n1218), .ZN(new_n1219));
  XOR2_X1   g794(.A(G290), .B(G1986), .Z(new_n1220));
  AOI21_X1  g795(.A(new_n1009), .B1(new_n1019), .B2(new_n1220), .ZN(new_n1221));
  OAI21_X1  g796(.A(new_n1029), .B1(new_n1219), .B2(new_n1221), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g797(.A1(new_n657), .A2(G319), .ZN(new_n1224));
  AOI211_X1 g798(.A(G227), .B(new_n1224), .C1(new_n905), .C2(new_n908), .ZN(new_n1225));
  AOI21_X1  g799(.A(G229), .B1(new_n994), .B2(new_n1001), .ZN(new_n1226));
  AND2_X1   g800(.A1(new_n1225), .A2(new_n1226), .ZN(G308));
  NAND2_X1  g801(.A1(new_n1225), .A2(new_n1226), .ZN(G225));
endmodule


