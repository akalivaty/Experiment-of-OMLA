

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U552 ( .A1(n634), .A2(n564), .ZN(n655) );
  NOR2_X2 U553 ( .A1(n808), .A2(n809), .ZN(n726) );
  AND2_X1 U554 ( .A1(n1007), .A2(G138), .ZN(n555) );
  XNOR2_X1 U555 ( .A(n535), .B(KEYINPUT32), .ZN(n534) );
  NAND2_X1 U556 ( .A1(n539), .A2(n538), .ZN(n808) );
  INV_X1 U557 ( .A(G1384), .ZN(n538) );
  XNOR2_X1 U558 ( .A(n787), .B(n786), .ZN(n533) );
  NAND2_X1 U559 ( .A1(n547), .A2(n551), .ZN(n540) );
  INV_X1 U560 ( .A(n520), .ZN(n530) );
  NAND2_X1 U561 ( .A1(n528), .A2(n526), .ZN(n525) );
  NAND2_X1 U562 ( .A1(n527), .A2(n530), .ZN(n526) );
  NAND2_X1 U563 ( .A1(n529), .A2(n842), .ZN(n528) );
  INV_X1 U564 ( .A(n842), .ZN(n527) );
  OR2_X1 U565 ( .A1(n762), .A2(n740), .ZN(n741) );
  AND2_X1 U566 ( .A1(n730), .A2(n542), .ZN(n541) );
  XNOR2_X1 U567 ( .A(n764), .B(n763), .ZN(n769) );
  NAND2_X1 U568 ( .A1(n534), .A2(n546), .ZN(n764) );
  NAND2_X1 U569 ( .A1(n531), .A2(n530), .ZN(n529) );
  INV_X1 U570 ( .A(n834), .ZN(n531) );
  NOR2_X1 U571 ( .A1(G651), .A2(n634), .ZN(n661) );
  OR2_X1 U572 ( .A1(n556), .A2(n557), .ZN(n539) );
  NAND2_X1 U573 ( .A1(n523), .A2(n519), .ZN(n522) );
  NOR2_X2 U574 ( .A1(n547), .A2(n551), .ZN(n625) );
  OR2_X1 U575 ( .A1(n769), .A2(n766), .ZN(n518) );
  NOR2_X2 U576 ( .A1(G2104), .A2(n547), .ZN(n695) );
  AND2_X1 U577 ( .A1(n842), .A2(n530), .ZN(n519) );
  XOR2_X1 U578 ( .A(KEYINPUT40), .B(n843), .Z(n520) );
  AND2_X1 U579 ( .A1(n521), .A2(n525), .ZN(n524) );
  NAND2_X1 U580 ( .A1(n533), .A2(n532), .ZN(n521) );
  NAND2_X1 U581 ( .A1(n524), .A2(n522), .ZN(G329) );
  INV_X1 U582 ( .A(n533), .ZN(n523) );
  AND2_X1 U583 ( .A1(n834), .A2(n520), .ZN(n532) );
  NAND2_X1 U584 ( .A1(n536), .A2(G8), .ZN(n535) );
  XNOR2_X1 U585 ( .A(n756), .B(n537), .ZN(n536) );
  INV_X1 U586 ( .A(KEYINPUT97), .ZN(n537) );
  INV_X1 U587 ( .A(n539), .ZN(G164) );
  NAND2_X1 U588 ( .A1(n726), .A2(G1996), .ZN(n711) );
  XNOR2_X2 U589 ( .A(n540), .B(KEYINPUT17), .ZN(n1007) );
  NAND2_X1 U590 ( .A1(n543), .A2(n541), .ZN(n544) );
  NAND2_X1 U591 ( .A1(n721), .A2(n724), .ZN(n542) );
  NAND2_X1 U592 ( .A1(n722), .A2(n724), .ZN(n543) );
  NAND2_X1 U593 ( .A1(n733), .A2(n544), .ZN(n736) );
  NAND2_X1 U594 ( .A1(n749), .A2(n748), .ZN(n757) );
  NOR2_X1 U595 ( .A1(n704), .A2(n703), .ZN(n545) );
  OR2_X1 U596 ( .A1(n762), .A2(n761), .ZN(n546) );
  INV_X1 U597 ( .A(n758), .ZN(n739) );
  XNOR2_X1 U598 ( .A(n734), .B(KEYINPUT29), .ZN(n735) );
  INV_X1 U599 ( .A(KEYINPUT31), .ZN(n746) );
  INV_X1 U600 ( .A(KEYINPUT98), .ZN(n763) );
  INV_X1 U601 ( .A(n705), .ZN(n706) );
  NAND2_X1 U602 ( .A1(n545), .A2(n706), .ZN(n809) );
  INV_X1 U603 ( .A(KEYINPUT83), .ZN(n554) );
  INV_X1 U604 ( .A(G2105), .ZN(n547) );
  NAND2_X1 U605 ( .A1(G126), .A2(n695), .ZN(n549) );
  INV_X1 U606 ( .A(G2104), .ZN(n551) );
  NAND2_X1 U607 ( .A1(G114), .A2(n625), .ZN(n548) );
  NAND2_X1 U608 ( .A1(n549), .A2(n548), .ZN(n550) );
  XOR2_X1 U609 ( .A(KEYINPUT82), .B(n550), .Z(n553) );
  NOR2_X1 U610 ( .A1(G2105), .A2(n551), .ZN(n697) );
  NAND2_X1 U611 ( .A1(n697), .A2(G102), .ZN(n552) );
  NAND2_X1 U612 ( .A1(n553), .A2(n552), .ZN(n557) );
  XNOR2_X1 U613 ( .A(n555), .B(n554), .ZN(n556) );
  XOR2_X1 U614 ( .A(G543), .B(KEYINPUT0), .Z(n634) );
  NAND2_X1 U615 ( .A1(G51), .A2(n661), .ZN(n561) );
  INV_X1 U616 ( .A(G651), .ZN(n564) );
  NOR2_X1 U617 ( .A1(G543), .A2(n564), .ZN(n558) );
  XOR2_X1 U618 ( .A(KEYINPUT1), .B(n558), .Z(n559) );
  NAND2_X1 U619 ( .A1(G63), .A2(n559), .ZN(n560) );
  NAND2_X1 U620 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U621 ( .A(KEYINPUT6), .B(n562), .ZN(n570) );
  NOR2_X1 U622 ( .A1(G651), .A2(G543), .ZN(n654) );
  NAND2_X1 U623 ( .A1(n654), .A2(G89), .ZN(n563) );
  XNOR2_X1 U624 ( .A(KEYINPUT4), .B(n563), .ZN(n567) );
  NAND2_X1 U625 ( .A1(n655), .A2(G76), .ZN(n565) );
  XOR2_X1 U626 ( .A(KEYINPUT67), .B(n565), .Z(n566) );
  NAND2_X1 U627 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U628 ( .A(n568), .B(KEYINPUT5), .Z(n569) );
  NOR2_X1 U629 ( .A1(n570), .A2(n569), .ZN(n571) );
  XOR2_X1 U630 ( .A(KEYINPUT68), .B(n571), .Z(n572) );
  XNOR2_X1 U631 ( .A(KEYINPUT7), .B(n572), .ZN(G168) );
  XOR2_X1 U632 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U633 ( .A1(G85), .A2(n654), .ZN(n574) );
  NAND2_X1 U634 ( .A1(G72), .A2(n655), .ZN(n573) );
  NAND2_X1 U635 ( .A1(n574), .A2(n573), .ZN(n578) );
  NAND2_X1 U636 ( .A1(G47), .A2(n661), .ZN(n576) );
  NAND2_X1 U637 ( .A1(G60), .A2(n559), .ZN(n575) );
  NAND2_X1 U638 ( .A1(n576), .A2(n575), .ZN(n577) );
  OR2_X1 U639 ( .A1(n578), .A2(n577), .ZN(G290) );
  NAND2_X1 U640 ( .A1(G52), .A2(n661), .ZN(n580) );
  NAND2_X1 U641 ( .A1(G64), .A2(n559), .ZN(n579) );
  NAND2_X1 U642 ( .A1(n580), .A2(n579), .ZN(n585) );
  NAND2_X1 U643 ( .A1(G90), .A2(n654), .ZN(n582) );
  NAND2_X1 U644 ( .A1(G77), .A2(n655), .ZN(n581) );
  NAND2_X1 U645 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U646 ( .A(KEYINPUT9), .B(n583), .Z(n584) );
  NOR2_X1 U647 ( .A1(n585), .A2(n584), .ZN(G171) );
  AND2_X1 U648 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U649 ( .A(G120), .ZN(G236) );
  INV_X1 U650 ( .A(G132), .ZN(G219) );
  INV_X1 U651 ( .A(G82), .ZN(G220) );
  NAND2_X1 U652 ( .A1(G7), .A2(G661), .ZN(n586) );
  XNOR2_X1 U653 ( .A(n586), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U654 ( .A(G223), .ZN(n844) );
  NAND2_X1 U655 ( .A1(n844), .A2(G567), .ZN(n587) );
  XOR2_X1 U656 ( .A(KEYINPUT11), .B(n587), .Z(G234) );
  NAND2_X1 U657 ( .A1(G56), .A2(n559), .ZN(n588) );
  XOR2_X1 U658 ( .A(KEYINPUT14), .B(n588), .Z(n594) );
  NAND2_X1 U659 ( .A1(n654), .A2(G81), .ZN(n589) );
  XNOR2_X1 U660 ( .A(n589), .B(KEYINPUT12), .ZN(n591) );
  NAND2_X1 U661 ( .A1(G68), .A2(n655), .ZN(n590) );
  NAND2_X1 U662 ( .A1(n591), .A2(n590), .ZN(n592) );
  XOR2_X1 U663 ( .A(KEYINPUT13), .B(n592), .Z(n593) );
  NOR2_X1 U664 ( .A1(n594), .A2(n593), .ZN(n596) );
  NAND2_X1 U665 ( .A1(n661), .A2(G43), .ZN(n595) );
  NAND2_X1 U666 ( .A1(n596), .A2(n595), .ZN(n977) );
  INV_X1 U667 ( .A(G860), .ZN(n618) );
  OR2_X1 U668 ( .A1(n977), .A2(n618), .ZN(G153) );
  INV_X1 U669 ( .A(G171), .ZN(G301) );
  NAND2_X1 U670 ( .A1(G92), .A2(n654), .ZN(n598) );
  NAND2_X1 U671 ( .A1(G79), .A2(n655), .ZN(n597) );
  NAND2_X1 U672 ( .A1(n598), .A2(n597), .ZN(n602) );
  NAND2_X1 U673 ( .A1(G54), .A2(n661), .ZN(n600) );
  NAND2_X1 U674 ( .A1(G66), .A2(n559), .ZN(n599) );
  NAND2_X1 U675 ( .A1(n600), .A2(n599), .ZN(n601) );
  NOR2_X1 U676 ( .A1(n602), .A2(n601), .ZN(n603) );
  XOR2_X1 U677 ( .A(KEYINPUT15), .B(n603), .Z(n604) );
  XNOR2_X2 U678 ( .A(KEYINPUT65), .B(n604), .ZN(n1026) );
  INV_X1 U679 ( .A(G868), .ZN(n614) );
  NAND2_X1 U680 ( .A1(n1026), .A2(n614), .ZN(n605) );
  XNOR2_X1 U681 ( .A(n605), .B(KEYINPUT66), .ZN(n607) );
  NAND2_X1 U682 ( .A1(G868), .A2(G301), .ZN(n606) );
  NAND2_X1 U683 ( .A1(n607), .A2(n606), .ZN(G284) );
  NAND2_X1 U684 ( .A1(G53), .A2(n661), .ZN(n609) );
  NAND2_X1 U685 ( .A1(G65), .A2(n559), .ZN(n608) );
  NAND2_X1 U686 ( .A1(n609), .A2(n608), .ZN(n613) );
  NAND2_X1 U687 ( .A1(G91), .A2(n654), .ZN(n611) );
  NAND2_X1 U688 ( .A1(G78), .A2(n655), .ZN(n610) );
  NAND2_X1 U689 ( .A1(n611), .A2(n610), .ZN(n612) );
  NOR2_X1 U690 ( .A1(n613), .A2(n612), .ZN(n920) );
  INV_X1 U691 ( .A(n920), .ZN(G299) );
  NAND2_X1 U692 ( .A1(G299), .A2(n614), .ZN(n616) );
  NAND2_X1 U693 ( .A1(G868), .A2(G286), .ZN(n615) );
  NAND2_X1 U694 ( .A1(n616), .A2(n615), .ZN(n617) );
  XOR2_X1 U695 ( .A(KEYINPUT69), .B(n617), .Z(G297) );
  NAND2_X1 U696 ( .A1(n618), .A2(G559), .ZN(n619) );
  INV_X1 U697 ( .A(n1026), .ZN(n675) );
  NAND2_X1 U698 ( .A1(n619), .A2(n675), .ZN(n620) );
  XNOR2_X1 U699 ( .A(n620), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U700 ( .A1(G868), .A2(n977), .ZN(n623) );
  NAND2_X1 U701 ( .A1(n675), .A2(G868), .ZN(n621) );
  NOR2_X1 U702 ( .A1(G559), .A2(n621), .ZN(n622) );
  NOR2_X1 U703 ( .A1(n623), .A2(n622), .ZN(G282) );
  NAND2_X1 U704 ( .A1(n695), .A2(G123), .ZN(n624) );
  XNOR2_X1 U705 ( .A(n624), .B(KEYINPUT18), .ZN(n627) );
  NAND2_X1 U706 ( .A1(G111), .A2(n625), .ZN(n626) );
  NAND2_X1 U707 ( .A1(n627), .A2(n626), .ZN(n631) );
  NAND2_X1 U708 ( .A1(G135), .A2(n1007), .ZN(n629) );
  NAND2_X1 U709 ( .A1(G99), .A2(n697), .ZN(n628) );
  NAND2_X1 U710 ( .A1(n629), .A2(n628), .ZN(n630) );
  NOR2_X1 U711 ( .A1(n631), .A2(n630), .ZN(n1015) );
  XOR2_X1 U712 ( .A(G2096), .B(n1015), .Z(n632) );
  NOR2_X1 U713 ( .A1(G2100), .A2(n632), .ZN(n633) );
  XOR2_X1 U714 ( .A(KEYINPUT70), .B(n633), .Z(G156) );
  NAND2_X1 U715 ( .A1(G49), .A2(n661), .ZN(n636) );
  NAND2_X1 U716 ( .A1(G87), .A2(n634), .ZN(n635) );
  NAND2_X1 U717 ( .A1(n636), .A2(n635), .ZN(n637) );
  NOR2_X1 U718 ( .A1(n559), .A2(n637), .ZN(n639) );
  NAND2_X1 U719 ( .A1(G651), .A2(G74), .ZN(n638) );
  NAND2_X1 U720 ( .A1(n639), .A2(n638), .ZN(G288) );
  NAND2_X1 U721 ( .A1(G86), .A2(n654), .ZN(n641) );
  NAND2_X1 U722 ( .A1(G48), .A2(n661), .ZN(n640) );
  NAND2_X1 U723 ( .A1(n641), .A2(n640), .ZN(n644) );
  NAND2_X1 U724 ( .A1(n655), .A2(G73), .ZN(n642) );
  XOR2_X1 U725 ( .A(KEYINPUT2), .B(n642), .Z(n643) );
  NOR2_X1 U726 ( .A1(n644), .A2(n643), .ZN(n646) );
  NAND2_X1 U727 ( .A1(n559), .A2(G61), .ZN(n645) );
  NAND2_X1 U728 ( .A1(n646), .A2(n645), .ZN(G305) );
  NAND2_X1 U729 ( .A1(G50), .A2(n661), .ZN(n648) );
  NAND2_X1 U730 ( .A1(G62), .A2(n559), .ZN(n647) );
  NAND2_X1 U731 ( .A1(n648), .A2(n647), .ZN(n652) );
  NAND2_X1 U732 ( .A1(G88), .A2(n654), .ZN(n650) );
  NAND2_X1 U733 ( .A1(G75), .A2(n655), .ZN(n649) );
  NAND2_X1 U734 ( .A1(n650), .A2(n649), .ZN(n651) );
  NOR2_X1 U735 ( .A1(n652), .A2(n651), .ZN(n653) );
  XNOR2_X1 U736 ( .A(n653), .B(KEYINPUT74), .ZN(G166) );
  INV_X1 U737 ( .A(G166), .ZN(G303) );
  NAND2_X1 U738 ( .A1(G93), .A2(n654), .ZN(n657) );
  NAND2_X1 U739 ( .A1(G80), .A2(n655), .ZN(n656) );
  NAND2_X1 U740 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U741 ( .A(n658), .B(KEYINPUT71), .ZN(n660) );
  NAND2_X1 U742 ( .A1(G67), .A2(n559), .ZN(n659) );
  NAND2_X1 U743 ( .A1(n660), .A2(n659), .ZN(n664) );
  NAND2_X1 U744 ( .A1(n661), .A2(G55), .ZN(n662) );
  XOR2_X1 U745 ( .A(KEYINPUT72), .B(n662), .Z(n663) );
  NOR2_X1 U746 ( .A1(n664), .A2(n663), .ZN(n665) );
  XOR2_X1 U747 ( .A(KEYINPUT73), .B(n665), .Z(n979) );
  NOR2_X1 U748 ( .A1(G868), .A2(n979), .ZN(n666) );
  XNOR2_X1 U749 ( .A(n666), .B(KEYINPUT77), .ZN(n678) );
  XNOR2_X1 U750 ( .A(n920), .B(G290), .ZN(n667) );
  XNOR2_X1 U751 ( .A(n667), .B(G288), .ZN(n668) );
  XOR2_X1 U752 ( .A(n668), .B(KEYINPUT76), .Z(n670) );
  XNOR2_X1 U753 ( .A(KEYINPUT19), .B(KEYINPUT75), .ZN(n669) );
  XNOR2_X1 U754 ( .A(n670), .B(n669), .ZN(n671) );
  XNOR2_X1 U755 ( .A(n979), .B(n671), .ZN(n673) );
  XNOR2_X1 U756 ( .A(G305), .B(G303), .ZN(n672) );
  XNOR2_X1 U757 ( .A(n673), .B(n672), .ZN(n674) );
  XOR2_X1 U758 ( .A(n674), .B(n977), .Z(n1027) );
  NAND2_X1 U759 ( .A1(n675), .A2(G559), .ZN(n976) );
  XNOR2_X1 U760 ( .A(n1027), .B(n976), .ZN(n676) );
  NAND2_X1 U761 ( .A1(G868), .A2(n676), .ZN(n677) );
  NAND2_X1 U762 ( .A1(n678), .A2(n677), .ZN(G295) );
  NAND2_X1 U763 ( .A1(G2078), .A2(G2084), .ZN(n681) );
  XNOR2_X1 U764 ( .A(KEYINPUT78), .B(KEYINPUT20), .ZN(n679) );
  XNOR2_X1 U765 ( .A(n679), .B(KEYINPUT79), .ZN(n680) );
  XNOR2_X1 U766 ( .A(n681), .B(n680), .ZN(n682) );
  NAND2_X1 U767 ( .A1(n682), .A2(G2090), .ZN(n683) );
  XNOR2_X1 U768 ( .A(KEYINPUT21), .B(n683), .ZN(n684) );
  NAND2_X1 U769 ( .A1(n684), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U770 ( .A(KEYINPUT80), .B(G44), .ZN(n685) );
  XNOR2_X1 U771 ( .A(n685), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U772 ( .A1(G220), .A2(G219), .ZN(n686) );
  XOR2_X1 U773 ( .A(KEYINPUT22), .B(n686), .Z(n687) );
  NOR2_X1 U774 ( .A1(G218), .A2(n687), .ZN(n688) );
  XOR2_X1 U775 ( .A(KEYINPUT81), .B(n688), .Z(n689) );
  NAND2_X1 U776 ( .A1(G96), .A2(n689), .ZN(n974) );
  NAND2_X1 U777 ( .A1(n974), .A2(G2106), .ZN(n693) );
  NAND2_X1 U778 ( .A1(G69), .A2(G108), .ZN(n690) );
  NOR2_X1 U779 ( .A1(G236), .A2(n690), .ZN(n691) );
  NAND2_X1 U780 ( .A1(G57), .A2(n691), .ZN(n975) );
  NAND2_X1 U781 ( .A1(n975), .A2(G567), .ZN(n692) );
  NAND2_X1 U782 ( .A1(n693), .A2(n692), .ZN(n981) );
  NAND2_X1 U783 ( .A1(G661), .A2(G483), .ZN(n694) );
  NOR2_X1 U784 ( .A1(n981), .A2(n694), .ZN(n847) );
  NAND2_X1 U785 ( .A1(n847), .A2(G36), .ZN(G176) );
  NAND2_X1 U786 ( .A1(G125), .A2(n695), .ZN(n696) );
  XNOR2_X1 U787 ( .A(n696), .B(KEYINPUT64), .ZN(n700) );
  NAND2_X1 U788 ( .A1(G101), .A2(n697), .ZN(n698) );
  XOR2_X1 U789 ( .A(KEYINPUT23), .B(n698), .Z(n699) );
  NAND2_X1 U790 ( .A1(n700), .A2(n699), .ZN(n705) );
  NAND2_X1 U791 ( .A1(G113), .A2(n625), .ZN(n702) );
  NAND2_X1 U792 ( .A1(G137), .A2(n1007), .ZN(n701) );
  NAND2_X1 U793 ( .A1(n702), .A2(n701), .ZN(n704) );
  NOR2_X1 U794 ( .A1(n705), .A2(n704), .ZN(G160) );
  INV_X1 U795 ( .A(G40), .ZN(n703) );
  INV_X1 U796 ( .A(n726), .ZN(n750) );
  NAND2_X2 U797 ( .A1(n750), .A2(G8), .ZN(n790) );
  NOR2_X1 U798 ( .A1(n726), .A2(G1961), .ZN(n707) );
  XOR2_X1 U799 ( .A(KEYINPUT90), .B(n707), .Z(n709) );
  XNOR2_X1 U800 ( .A(G2078), .B(KEYINPUT25), .ZN(n900) );
  NAND2_X1 U801 ( .A1(n726), .A2(n900), .ZN(n708) );
  NAND2_X1 U802 ( .A1(n709), .A2(n708), .ZN(n743) );
  NAND2_X1 U803 ( .A1(n743), .A2(G171), .ZN(n738) );
  NAND2_X1 U804 ( .A1(KEYINPUT26), .A2(G1341), .ZN(n710) );
  OR2_X1 U805 ( .A1(n726), .A2(n710), .ZN(n715) );
  XNOR2_X1 U806 ( .A(KEYINPUT26), .B(n711), .ZN(n712) );
  NAND2_X1 U807 ( .A1(n715), .A2(n712), .ZN(n714) );
  INV_X1 U808 ( .A(KEYINPUT93), .ZN(n713) );
  NAND2_X1 U809 ( .A1(n714), .A2(n713), .ZN(n717) );
  NAND2_X1 U810 ( .A1(KEYINPUT93), .A2(n715), .ZN(n716) );
  NAND2_X1 U811 ( .A1(n717), .A2(n716), .ZN(n718) );
  NOR2_X1 U812 ( .A1(n718), .A2(n977), .ZN(n722) );
  NAND2_X1 U813 ( .A1(G1348), .A2(n750), .ZN(n720) );
  NAND2_X1 U814 ( .A1(G2067), .A2(n726), .ZN(n719) );
  NAND2_X1 U815 ( .A1(n720), .A2(n719), .ZN(n723) );
  NOR2_X1 U816 ( .A1(n1026), .A2(n723), .ZN(n721) );
  NAND2_X1 U817 ( .A1(n1026), .A2(n723), .ZN(n724) );
  NAND2_X1 U818 ( .A1(n726), .A2(G2072), .ZN(n725) );
  XNOR2_X1 U819 ( .A(KEYINPUT27), .B(n725), .ZN(n729) );
  XNOR2_X1 U820 ( .A(G1956), .B(KEYINPUT91), .ZN(n945) );
  NOR2_X1 U821 ( .A1(n726), .A2(n945), .ZN(n727) );
  XNOR2_X1 U822 ( .A(n727), .B(KEYINPUT92), .ZN(n728) );
  NOR2_X1 U823 ( .A1(n729), .A2(n728), .ZN(n731) );
  NAND2_X1 U824 ( .A1(n920), .A2(n731), .ZN(n730) );
  NOR2_X1 U825 ( .A1(n731), .A2(n920), .ZN(n732) );
  XOR2_X1 U826 ( .A(n732), .B(KEYINPUT28), .Z(n733) );
  XNOR2_X1 U827 ( .A(KEYINPUT94), .B(KEYINPUT95), .ZN(n734) );
  XNOR2_X1 U828 ( .A(n736), .B(n735), .ZN(n737) );
  NAND2_X1 U829 ( .A1(n738), .A2(n737), .ZN(n749) );
  NOR2_X1 U830 ( .A1(G1966), .A2(n790), .ZN(n762) );
  NOR2_X1 U831 ( .A1(G2084), .A2(n750), .ZN(n758) );
  NAND2_X1 U832 ( .A1(n739), .A2(G8), .ZN(n740) );
  XNOR2_X1 U833 ( .A(KEYINPUT30), .B(n741), .ZN(n742) );
  NOR2_X1 U834 ( .A1(n742), .A2(G168), .ZN(n745) );
  NOR2_X1 U835 ( .A1(G171), .A2(n743), .ZN(n744) );
  NOR2_X1 U836 ( .A1(n745), .A2(n744), .ZN(n747) );
  XNOR2_X1 U837 ( .A(n747), .B(n746), .ZN(n748) );
  NAND2_X1 U838 ( .A1(n757), .A2(G286), .ZN(n755) );
  NOR2_X1 U839 ( .A1(G1971), .A2(n790), .ZN(n752) );
  NOR2_X1 U840 ( .A1(G2090), .A2(n750), .ZN(n751) );
  NOR2_X1 U841 ( .A1(n752), .A2(n751), .ZN(n753) );
  NAND2_X1 U842 ( .A1(G303), .A2(n753), .ZN(n754) );
  NAND2_X1 U843 ( .A1(n755), .A2(n754), .ZN(n756) );
  XNOR2_X1 U844 ( .A(n757), .B(KEYINPUT96), .ZN(n760) );
  NAND2_X1 U845 ( .A1(n758), .A2(G8), .ZN(n759) );
  NAND2_X1 U846 ( .A1(n760), .A2(n759), .ZN(n761) );
  NAND2_X1 U847 ( .A1(G8), .A2(G166), .ZN(n765) );
  NOR2_X1 U848 ( .A1(n765), .A2(G2090), .ZN(n766) );
  NAND2_X1 U849 ( .A1(n790), .A2(n518), .ZN(n768) );
  INV_X1 U850 ( .A(KEYINPUT99), .ZN(n767) );
  XNOR2_X1 U851 ( .A(n768), .B(n767), .ZN(n785) );
  INV_X1 U852 ( .A(n769), .ZN(n772) );
  NOR2_X1 U853 ( .A1(G1976), .A2(G288), .ZN(n776) );
  NOR2_X1 U854 ( .A1(G1971), .A2(G303), .ZN(n770) );
  NOR2_X1 U855 ( .A1(n776), .A2(n770), .ZN(n919) );
  INV_X1 U856 ( .A(KEYINPUT33), .ZN(n775) );
  AND2_X1 U857 ( .A1(n919), .A2(n775), .ZN(n771) );
  NAND2_X1 U858 ( .A1(n772), .A2(n771), .ZN(n783) );
  NAND2_X1 U859 ( .A1(G1976), .A2(G288), .ZN(n918) );
  INV_X1 U860 ( .A(n790), .ZN(n773) );
  NAND2_X1 U861 ( .A1(n918), .A2(n773), .ZN(n774) );
  AND2_X1 U862 ( .A1(n775), .A2(n774), .ZN(n781) );
  NAND2_X1 U863 ( .A1(n776), .A2(KEYINPUT33), .ZN(n777) );
  NOR2_X1 U864 ( .A1(n777), .A2(n790), .ZN(n779) );
  XOR2_X1 U865 ( .A(G1981), .B(G305), .Z(n928) );
  INV_X1 U866 ( .A(n928), .ZN(n778) );
  OR2_X1 U867 ( .A1(n779), .A2(n778), .ZN(n780) );
  NOR2_X1 U868 ( .A1(n781), .A2(n780), .ZN(n782) );
  NAND2_X1 U869 ( .A1(n783), .A2(n782), .ZN(n784) );
  NAND2_X1 U870 ( .A1(n785), .A2(n784), .ZN(n787) );
  INV_X1 U871 ( .A(KEYINPUT100), .ZN(n786) );
  NOR2_X1 U872 ( .A1(G1981), .A2(G305), .ZN(n788) );
  XOR2_X1 U873 ( .A(n788), .B(KEYINPUT24), .Z(n789) );
  NOR2_X1 U874 ( .A1(n790), .A2(n789), .ZN(n833) );
  NAND2_X1 U875 ( .A1(G105), .A2(n697), .ZN(n791) );
  XNOR2_X1 U876 ( .A(n791), .B(KEYINPUT38), .ZN(n799) );
  NAND2_X1 U877 ( .A1(G129), .A2(n695), .ZN(n793) );
  NAND2_X1 U878 ( .A1(G117), .A2(n625), .ZN(n792) );
  NAND2_X1 U879 ( .A1(n793), .A2(n792), .ZN(n794) );
  XNOR2_X1 U880 ( .A(KEYINPUT88), .B(n794), .ZN(n797) );
  NAND2_X1 U881 ( .A1(G141), .A2(n1007), .ZN(n795) );
  XNOR2_X1 U882 ( .A(KEYINPUT89), .B(n795), .ZN(n796) );
  NOR2_X1 U883 ( .A1(n797), .A2(n796), .ZN(n798) );
  NAND2_X1 U884 ( .A1(n799), .A2(n798), .ZN(n1020) );
  NOR2_X1 U885 ( .A1(G1996), .A2(n1020), .ZN(n800) );
  XOR2_X1 U886 ( .A(KEYINPUT101), .B(n800), .Z(n868) );
  AND2_X1 U887 ( .A1(n1020), .A2(G1996), .ZN(n863) );
  NAND2_X1 U888 ( .A1(G119), .A2(n695), .ZN(n802) );
  NAND2_X1 U889 ( .A1(G107), .A2(n625), .ZN(n801) );
  NAND2_X1 U890 ( .A1(n802), .A2(n801), .ZN(n803) );
  XNOR2_X1 U891 ( .A(KEYINPUT87), .B(n803), .ZN(n807) );
  NAND2_X1 U892 ( .A1(G131), .A2(n1007), .ZN(n805) );
  NAND2_X1 U893 ( .A1(G95), .A2(n697), .ZN(n804) );
  AND2_X1 U894 ( .A1(n805), .A2(n804), .ZN(n806) );
  NAND2_X1 U895 ( .A1(n807), .A2(n806), .ZN(n1002) );
  AND2_X1 U896 ( .A1(n1002), .A2(G1991), .ZN(n856) );
  OR2_X1 U897 ( .A1(n863), .A2(n856), .ZN(n811) );
  INV_X1 U898 ( .A(n808), .ZN(n810) );
  NOR2_X1 U899 ( .A1(n810), .A2(n809), .ZN(n837) );
  NAND2_X1 U900 ( .A1(n811), .A2(n837), .ZN(n835) );
  INV_X1 U901 ( .A(n835), .ZN(n814) );
  NOR2_X1 U902 ( .A1(G1986), .A2(G290), .ZN(n812) );
  NOR2_X1 U903 ( .A1(G1991), .A2(n1002), .ZN(n859) );
  NOR2_X1 U904 ( .A1(n812), .A2(n859), .ZN(n813) );
  NOR2_X1 U905 ( .A1(n814), .A2(n813), .ZN(n815) );
  NOR2_X1 U906 ( .A1(n868), .A2(n815), .ZN(n816) );
  XNOR2_X1 U907 ( .A(n816), .B(KEYINPUT39), .ZN(n829) );
  NAND2_X1 U908 ( .A1(n697), .A2(G104), .ZN(n817) );
  XOR2_X1 U909 ( .A(KEYINPUT85), .B(n817), .Z(n819) );
  NAND2_X1 U910 ( .A1(n1007), .A2(G140), .ZN(n818) );
  NAND2_X1 U911 ( .A1(n819), .A2(n818), .ZN(n820) );
  XNOR2_X1 U912 ( .A(KEYINPUT34), .B(n820), .ZN(n825) );
  NAND2_X1 U913 ( .A1(G128), .A2(n695), .ZN(n822) );
  NAND2_X1 U914 ( .A1(G116), .A2(n625), .ZN(n821) );
  NAND2_X1 U915 ( .A1(n822), .A2(n821), .ZN(n823) );
  XOR2_X1 U916 ( .A(n823), .B(KEYINPUT35), .Z(n824) );
  NOR2_X1 U917 ( .A1(n825), .A2(n824), .ZN(n826) );
  XOR2_X1 U918 ( .A(KEYINPUT36), .B(n826), .Z(n827) );
  XOR2_X1 U919 ( .A(KEYINPUT86), .B(n827), .Z(n1024) );
  XNOR2_X1 U920 ( .A(G2067), .B(KEYINPUT37), .ZN(n828) );
  XNOR2_X1 U921 ( .A(n828), .B(KEYINPUT84), .ZN(n830) );
  NOR2_X1 U922 ( .A1(n1024), .A2(n830), .ZN(n865) );
  NAND2_X1 U923 ( .A1(n837), .A2(n865), .ZN(n836) );
  NAND2_X1 U924 ( .A1(n829), .A2(n836), .ZN(n831) );
  NAND2_X1 U925 ( .A1(n1024), .A2(n830), .ZN(n874) );
  NAND2_X1 U926 ( .A1(n831), .A2(n874), .ZN(n832) );
  AND2_X1 U927 ( .A1(n832), .A2(n837), .ZN(n841) );
  NOR2_X1 U928 ( .A1(n833), .A2(n841), .ZN(n834) );
  NAND2_X1 U929 ( .A1(n836), .A2(n835), .ZN(n839) );
  XNOR2_X1 U930 ( .A(G1986), .B(G290), .ZN(n915) );
  AND2_X1 U931 ( .A1(n915), .A2(n837), .ZN(n838) );
  NOR2_X1 U932 ( .A1(n839), .A2(n838), .ZN(n840) );
  OR2_X1 U933 ( .A1(n841), .A2(n840), .ZN(n842) );
  XOR2_X1 U934 ( .A(KEYINPUT102), .B(KEYINPUT103), .Z(n843) );
  NAND2_X1 U935 ( .A1(G2106), .A2(n844), .ZN(G217) );
  AND2_X1 U936 ( .A1(G15), .A2(G2), .ZN(n845) );
  NAND2_X1 U937 ( .A1(G661), .A2(n845), .ZN(G259) );
  NAND2_X1 U938 ( .A1(G3), .A2(G1), .ZN(n846) );
  NAND2_X1 U939 ( .A1(n847), .A2(n846), .ZN(G188) );
  XOR2_X1 U940 ( .A(G69), .B(KEYINPUT106), .Z(G235) );
  XNOR2_X1 U941 ( .A(G108), .B(KEYINPUT113), .ZN(G238) );
  NAND2_X1 U943 ( .A1(G112), .A2(n625), .ZN(n849) );
  NAND2_X1 U944 ( .A1(G100), .A2(n697), .ZN(n848) );
  NAND2_X1 U945 ( .A1(n849), .A2(n848), .ZN(n850) );
  XNOR2_X1 U946 ( .A(n850), .B(KEYINPUT109), .ZN(n852) );
  NAND2_X1 U947 ( .A1(G136), .A2(n1007), .ZN(n851) );
  NAND2_X1 U948 ( .A1(n852), .A2(n851), .ZN(n855) );
  NAND2_X1 U949 ( .A1(n695), .A2(G124), .ZN(n853) );
  XOR2_X1 U950 ( .A(KEYINPUT44), .B(n853), .Z(n854) );
  NOR2_X1 U951 ( .A1(n855), .A2(n854), .ZN(G162) );
  NOR2_X1 U952 ( .A1(n856), .A2(n1015), .ZN(n861) );
  XOR2_X1 U953 ( .A(G160), .B(G2084), .Z(n857) );
  XNOR2_X1 U954 ( .A(KEYINPUT114), .B(n857), .ZN(n858) );
  NOR2_X1 U955 ( .A1(n859), .A2(n858), .ZN(n860) );
  NAND2_X1 U956 ( .A1(n861), .A2(n860), .ZN(n862) );
  OR2_X1 U957 ( .A1(n863), .A2(n862), .ZN(n864) );
  NOR2_X1 U958 ( .A1(n865), .A2(n864), .ZN(n866) );
  XOR2_X1 U959 ( .A(KEYINPUT115), .B(n866), .Z(n872) );
  XOR2_X1 U960 ( .A(G2090), .B(G162), .Z(n867) );
  NOR2_X1 U961 ( .A1(n868), .A2(n867), .ZN(n869) );
  XOR2_X1 U962 ( .A(KEYINPUT116), .B(n869), .Z(n870) );
  XNOR2_X1 U963 ( .A(KEYINPUT51), .B(n870), .ZN(n871) );
  NAND2_X1 U964 ( .A1(n872), .A2(n871), .ZN(n873) );
  XNOR2_X1 U965 ( .A(n873), .B(KEYINPUT117), .ZN(n875) );
  NAND2_X1 U966 ( .A1(n875), .A2(n874), .ZN(n888) );
  NAND2_X1 U967 ( .A1(G139), .A2(n1007), .ZN(n877) );
  NAND2_X1 U968 ( .A1(G103), .A2(n697), .ZN(n876) );
  NAND2_X1 U969 ( .A1(n877), .A2(n876), .ZN(n883) );
  NAND2_X1 U970 ( .A1(G127), .A2(n695), .ZN(n879) );
  NAND2_X1 U971 ( .A1(G115), .A2(n625), .ZN(n878) );
  NAND2_X1 U972 ( .A1(n879), .A2(n878), .ZN(n880) );
  XNOR2_X1 U973 ( .A(KEYINPUT47), .B(n880), .ZN(n881) );
  XNOR2_X1 U974 ( .A(KEYINPUT111), .B(n881), .ZN(n882) );
  NOR2_X1 U975 ( .A1(n883), .A2(n882), .ZN(n1001) );
  XOR2_X1 U976 ( .A(G2072), .B(n1001), .Z(n885) );
  XOR2_X1 U977 ( .A(G164), .B(G2078), .Z(n884) );
  NOR2_X1 U978 ( .A1(n885), .A2(n884), .ZN(n886) );
  XOR2_X1 U979 ( .A(KEYINPUT50), .B(n886), .Z(n887) );
  NOR2_X1 U980 ( .A1(n888), .A2(n887), .ZN(n889) );
  XNOR2_X1 U981 ( .A(KEYINPUT52), .B(n889), .ZN(n890) );
  INV_X1 U982 ( .A(KEYINPUT55), .ZN(n910) );
  NAND2_X1 U983 ( .A1(n890), .A2(n910), .ZN(n891) );
  NAND2_X1 U984 ( .A1(n891), .A2(G29), .ZN(n972) );
  XNOR2_X1 U985 ( .A(G2090), .B(G35), .ZN(n905) );
  XNOR2_X1 U986 ( .A(G2067), .B(G26), .ZN(n893) );
  XNOR2_X1 U987 ( .A(G33), .B(G2072), .ZN(n892) );
  NOR2_X1 U988 ( .A1(n893), .A2(n892), .ZN(n899) );
  XOR2_X1 U989 ( .A(G32), .B(G1996), .Z(n894) );
  NAND2_X1 U990 ( .A1(n894), .A2(G28), .ZN(n897) );
  XNOR2_X1 U991 ( .A(KEYINPUT118), .B(G1991), .ZN(n895) );
  XNOR2_X1 U992 ( .A(G25), .B(n895), .ZN(n896) );
  NOR2_X1 U993 ( .A1(n897), .A2(n896), .ZN(n898) );
  NAND2_X1 U994 ( .A1(n899), .A2(n898), .ZN(n902) );
  XOR2_X1 U995 ( .A(G27), .B(n900), .Z(n901) );
  NOR2_X1 U996 ( .A1(n902), .A2(n901), .ZN(n903) );
  XNOR2_X1 U997 ( .A(KEYINPUT53), .B(n903), .ZN(n904) );
  NOR2_X1 U998 ( .A1(n905), .A2(n904), .ZN(n908) );
  XOR2_X1 U999 ( .A(G2084), .B(G34), .Z(n906) );
  XNOR2_X1 U1000 ( .A(KEYINPUT54), .B(n906), .ZN(n907) );
  NAND2_X1 U1001 ( .A1(n908), .A2(n907), .ZN(n909) );
  XNOR2_X1 U1002 ( .A(n910), .B(n909), .ZN(n912) );
  INV_X1 U1003 ( .A(G29), .ZN(n911) );
  NAND2_X1 U1004 ( .A1(n912), .A2(n911), .ZN(n913) );
  NAND2_X1 U1005 ( .A1(G11), .A2(n913), .ZN(n970) );
  XNOR2_X1 U1006 ( .A(G16), .B(KEYINPUT56), .ZN(n936) );
  XNOR2_X1 U1007 ( .A(G1348), .B(n1026), .ZN(n914) );
  NOR2_X1 U1008 ( .A1(n915), .A2(n914), .ZN(n934) );
  XNOR2_X1 U1009 ( .A(G301), .B(G1961), .ZN(n917) );
  XNOR2_X1 U1010 ( .A(n977), .B(G1341), .ZN(n916) );
  NOR2_X1 U1011 ( .A1(n917), .A2(n916), .ZN(n927) );
  NAND2_X1 U1012 ( .A1(n919), .A2(n918), .ZN(n924) );
  XNOR2_X1 U1013 ( .A(G1956), .B(n920), .ZN(n922) );
  NAND2_X1 U1014 ( .A1(G303), .A2(G1971), .ZN(n921) );
  NAND2_X1 U1015 ( .A1(n922), .A2(n921), .ZN(n923) );
  NOR2_X1 U1016 ( .A1(n924), .A2(n923), .ZN(n925) );
  XOR2_X1 U1017 ( .A(KEYINPUT119), .B(n925), .Z(n926) );
  NAND2_X1 U1018 ( .A1(n927), .A2(n926), .ZN(n932) );
  XNOR2_X1 U1019 ( .A(G1966), .B(G168), .ZN(n929) );
  NAND2_X1 U1020 ( .A1(n929), .A2(n928), .ZN(n930) );
  XOR2_X1 U1021 ( .A(KEYINPUT57), .B(n930), .Z(n931) );
  NOR2_X1 U1022 ( .A1(n932), .A2(n931), .ZN(n933) );
  NAND2_X1 U1023 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1024 ( .A1(n936), .A2(n935), .ZN(n968) );
  INV_X1 U1025 ( .A(G16), .ZN(n966) );
  XOR2_X1 U1026 ( .A(G1981), .B(G6), .Z(n937) );
  XNOR2_X1 U1027 ( .A(KEYINPUT121), .B(n937), .ZN(n939) );
  XNOR2_X1 U1028 ( .A(G19), .B(G1341), .ZN(n938) );
  NOR2_X1 U1029 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1030 ( .A(KEYINPUT122), .B(n940), .ZN(n944) );
  XOR2_X1 U1031 ( .A(KEYINPUT123), .B(G4), .Z(n942) );
  XNOR2_X1 U1032 ( .A(G1348), .B(KEYINPUT59), .ZN(n941) );
  XNOR2_X1 U1033 ( .A(n942), .B(n941), .ZN(n943) );
  NAND2_X1 U1034 ( .A1(n944), .A2(n943), .ZN(n948) );
  XOR2_X1 U1035 ( .A(G20), .B(n945), .Z(n946) );
  XNOR2_X1 U1036 ( .A(KEYINPUT120), .B(n946), .ZN(n947) );
  NOR2_X1 U1037 ( .A1(n948), .A2(n947), .ZN(n949) );
  XNOR2_X1 U1038 ( .A(KEYINPUT60), .B(n949), .ZN(n950) );
  XNOR2_X1 U1039 ( .A(n950), .B(KEYINPUT124), .ZN(n954) );
  XNOR2_X1 U1040 ( .A(G1966), .B(G21), .ZN(n952) );
  XNOR2_X1 U1041 ( .A(G5), .B(G1961), .ZN(n951) );
  NOR2_X1 U1042 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1043 ( .A1(n954), .A2(n953), .ZN(n962) );
  XNOR2_X1 U1044 ( .A(G1986), .B(G24), .ZN(n959) );
  XNOR2_X1 U1045 ( .A(G1976), .B(G23), .ZN(n956) );
  XNOR2_X1 U1046 ( .A(G22), .B(G1971), .ZN(n955) );
  NOR2_X1 U1047 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1048 ( .A(KEYINPUT125), .B(n957), .ZN(n958) );
  NOR2_X1 U1049 ( .A1(n959), .A2(n958), .ZN(n960) );
  XOR2_X1 U1050 ( .A(n960), .B(KEYINPUT58), .Z(n961) );
  NOR2_X1 U1051 ( .A1(n962), .A2(n961), .ZN(n963) );
  XOR2_X1 U1052 ( .A(KEYINPUT126), .B(n963), .Z(n964) );
  XOR2_X1 U1053 ( .A(KEYINPUT61), .B(n964), .Z(n965) );
  NAND2_X1 U1054 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1055 ( .A1(n968), .A2(n967), .ZN(n969) );
  NOR2_X1 U1056 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1057 ( .A1(n972), .A2(n971), .ZN(n973) );
  XOR2_X1 U1058 ( .A(KEYINPUT62), .B(n973), .Z(G311) );
  XNOR2_X1 U1059 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1060 ( .A(G96), .ZN(G221) );
  NOR2_X1 U1061 ( .A1(n975), .A2(n974), .ZN(G325) );
  INV_X1 U1062 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U1063 ( .A(n977), .B(n976), .ZN(n978) );
  NOR2_X1 U1064 ( .A1(n978), .A2(G860), .ZN(n980) );
  XNOR2_X1 U1065 ( .A(n980), .B(n979), .ZN(G145) );
  INV_X1 U1066 ( .A(n981), .ZN(G319) );
  XNOR2_X1 U1067 ( .A(G1986), .B(G1976), .ZN(n991) );
  XOR2_X1 U1068 ( .A(G1966), .B(G1971), .Z(n983) );
  XNOR2_X1 U1069 ( .A(G1996), .B(G1981), .ZN(n982) );
  XNOR2_X1 U1070 ( .A(n983), .B(n982), .ZN(n987) );
  XOR2_X1 U1071 ( .A(KEYINPUT108), .B(G2474), .Z(n985) );
  XNOR2_X1 U1072 ( .A(G1991), .B(G1961), .ZN(n984) );
  XNOR2_X1 U1073 ( .A(n985), .B(n984), .ZN(n986) );
  XOR2_X1 U1074 ( .A(n987), .B(n986), .Z(n989) );
  XNOR2_X1 U1075 ( .A(G1956), .B(KEYINPUT41), .ZN(n988) );
  XNOR2_X1 U1076 ( .A(n989), .B(n988), .ZN(n990) );
  XNOR2_X1 U1077 ( .A(n991), .B(n990), .ZN(G229) );
  XOR2_X1 U1078 ( .A(KEYINPUT107), .B(G2078), .Z(n993) );
  XNOR2_X1 U1079 ( .A(G2067), .B(G2084), .ZN(n992) );
  XNOR2_X1 U1080 ( .A(n993), .B(n992), .ZN(n994) );
  XOR2_X1 U1081 ( .A(n994), .B(G2678), .Z(n996) );
  XNOR2_X1 U1082 ( .A(G2072), .B(KEYINPUT42), .ZN(n995) );
  XNOR2_X1 U1083 ( .A(n996), .B(n995), .ZN(n1000) );
  XOR2_X1 U1084 ( .A(G2100), .B(G2096), .Z(n998) );
  XNOR2_X1 U1085 ( .A(G2090), .B(KEYINPUT43), .ZN(n997) );
  XNOR2_X1 U1086 ( .A(n998), .B(n997), .ZN(n999) );
  XOR2_X1 U1087 ( .A(n1000), .B(n999), .Z(G227) );
  XOR2_X1 U1088 ( .A(G162), .B(n1001), .Z(n1004) );
  XOR2_X1 U1089 ( .A(G160), .B(n1002), .Z(n1003) );
  XNOR2_X1 U1090 ( .A(n1004), .B(n1003), .ZN(n1019) );
  XOR2_X1 U1091 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n1017) );
  NAND2_X1 U1092 ( .A1(G130), .A2(n695), .ZN(n1006) );
  NAND2_X1 U1093 ( .A1(G118), .A2(n625), .ZN(n1005) );
  NAND2_X1 U1094 ( .A1(n1006), .A2(n1005), .ZN(n1013) );
  NAND2_X1 U1095 ( .A1(G142), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1096 ( .A1(G106), .A2(n697), .ZN(n1008) );
  NAND2_X1 U1097 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XOR2_X1 U1098 ( .A(KEYINPUT45), .B(n1010), .Z(n1011) );
  XNOR2_X1 U1099 ( .A(KEYINPUT110), .B(n1011), .ZN(n1012) );
  NOR2_X1 U1100 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1101 ( .A(n1015), .B(n1014), .ZN(n1016) );
  XNOR2_X1 U1102 ( .A(n1017), .B(n1016), .ZN(n1018) );
  XOR2_X1 U1103 ( .A(n1019), .B(n1018), .Z(n1022) );
  XOR2_X1 U1104 ( .A(G164), .B(n1020), .Z(n1021) );
  XNOR2_X1 U1105 ( .A(n1022), .B(n1021), .ZN(n1023) );
  XOR2_X1 U1106 ( .A(n1024), .B(n1023), .Z(n1025) );
  NOR2_X1 U1107 ( .A1(G37), .A2(n1025), .ZN(G395) );
  XNOR2_X1 U1108 ( .A(KEYINPUT112), .B(n1026), .ZN(n1028) );
  XNOR2_X1 U1109 ( .A(n1028), .B(n1027), .ZN(n1030) );
  XNOR2_X1 U1110 ( .A(G286), .B(G171), .ZN(n1029) );
  XNOR2_X1 U1111 ( .A(n1030), .B(n1029), .ZN(n1031) );
  NOR2_X1 U1112 ( .A1(G37), .A2(n1031), .ZN(G397) );
  XNOR2_X1 U1113 ( .A(G1341), .B(G2446), .ZN(n1041) );
  XOR2_X1 U1114 ( .A(G2451), .B(G2430), .Z(n1033) );
  XNOR2_X1 U1115 ( .A(G1348), .B(KEYINPUT105), .ZN(n1032) );
  XNOR2_X1 U1116 ( .A(n1033), .B(n1032), .ZN(n1037) );
  XOR2_X1 U1117 ( .A(G2435), .B(G2454), .Z(n1035) );
  XNOR2_X1 U1118 ( .A(KEYINPUT104), .B(G2438), .ZN(n1034) );
  XNOR2_X1 U1119 ( .A(n1035), .B(n1034), .ZN(n1036) );
  XOR2_X1 U1120 ( .A(n1037), .B(n1036), .Z(n1039) );
  XNOR2_X1 U1121 ( .A(G2443), .B(G2427), .ZN(n1038) );
  XNOR2_X1 U1122 ( .A(n1039), .B(n1038), .ZN(n1040) );
  XNOR2_X1 U1123 ( .A(n1041), .B(n1040), .ZN(n1042) );
  NAND2_X1 U1124 ( .A1(n1042), .A2(G14), .ZN(n1048) );
  NAND2_X1 U1125 ( .A1(G319), .A2(n1048), .ZN(n1045) );
  NOR2_X1 U1126 ( .A1(G229), .A2(G227), .ZN(n1043) );
  XNOR2_X1 U1127 ( .A(KEYINPUT49), .B(n1043), .ZN(n1044) );
  NOR2_X1 U1128 ( .A1(n1045), .A2(n1044), .ZN(n1047) );
  NOR2_X1 U1129 ( .A1(G395), .A2(G397), .ZN(n1046) );
  NAND2_X1 U1130 ( .A1(n1047), .A2(n1046), .ZN(G225) );
  INV_X1 U1131 ( .A(G225), .ZN(G308) );
  INV_X1 U1132 ( .A(G57), .ZN(G237) );
  INV_X1 U1133 ( .A(n1048), .ZN(G401) );
endmodule

