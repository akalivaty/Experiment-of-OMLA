//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 1 1 0 0 1 1 0 1 0 0 1 1 1 1 1 0 1 0 1 1 1 1 0 1 0 1 0 1 1 1 0 1 0 0 1 0 0 1 1 0 0 0 1 0 1 0 0 0 1 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:38 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n614, new_n615, new_n616, new_n617,
    new_n618, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n661, new_n662, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n709, new_n710,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n863,
    new_n864, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938;
  INV_X1    g000(.A(KEYINPUT96), .ZN(new_n187));
  INV_X1    g001(.A(G140), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G125), .ZN(new_n189));
  INV_X1    g003(.A(G125), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G140), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n189), .A2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT16), .ZN(new_n193));
  OAI21_X1  g007(.A(KEYINPUT81), .B1(new_n192), .B2(new_n193), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n193), .A2(new_n188), .A3(G125), .ZN(new_n195));
  XNOR2_X1  g009(.A(G125), .B(G140), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT81), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n196), .A2(new_n197), .A3(KEYINPUT16), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n194), .A2(new_n195), .A3(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G146), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n194), .A2(G146), .A3(new_n198), .A4(new_n195), .ZN(new_n202));
  INV_X1    g016(.A(G237), .ZN(new_n203));
  INV_X1    g017(.A(G953), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n203), .A2(new_n204), .A3(G214), .ZN(new_n205));
  INV_X1    g019(.A(G143), .ZN(new_n206));
  XNOR2_X1  g020(.A(new_n205), .B(new_n206), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n207), .A2(KEYINPUT17), .A3(G131), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n201), .A2(new_n202), .A3(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(KEYINPUT90), .ZN(new_n210));
  INV_X1    g024(.A(new_n207), .ZN(new_n211));
  INV_X1    g025(.A(G131), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n211), .A2(KEYINPUT88), .A3(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT17), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n207), .A2(G131), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT88), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n216), .B1(new_n207), .B2(G131), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n213), .A2(new_n214), .A3(new_n215), .A4(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT90), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n201), .A2(new_n219), .A3(new_n202), .A4(new_n208), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n210), .A2(new_n218), .A3(new_n220), .ZN(new_n221));
  XNOR2_X1  g035(.A(G113), .B(G122), .ZN(new_n222));
  INV_X1    g036(.A(G104), .ZN(new_n223));
  XNOR2_X1  g037(.A(new_n222), .B(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT18), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n211), .B1(new_n225), .B2(new_n212), .ZN(new_n226));
  XNOR2_X1  g040(.A(new_n196), .B(new_n200), .ZN(new_n227));
  OAI211_X1 g041(.A(new_n226), .B(new_n227), .C1(new_n225), .C2(new_n215), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n221), .A2(new_n224), .A3(new_n228), .ZN(new_n229));
  AND3_X1   g043(.A1(new_n213), .A2(new_n215), .A3(new_n217), .ZN(new_n230));
  NOR2_X1   g044(.A1(KEYINPUT89), .A2(KEYINPUT19), .ZN(new_n231));
  AND2_X1   g045(.A1(KEYINPUT89), .A2(KEYINPUT19), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n196), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n233), .B1(new_n196), .B2(new_n231), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n202), .B1(new_n234), .B2(G146), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n228), .B1(new_n230), .B2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n224), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n229), .A2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(G475), .ZN(new_n240));
  INV_X1    g054(.A(G902), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n239), .A2(new_n240), .A3(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT20), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(new_n229), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n224), .B1(new_n221), .B2(new_n228), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n241), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(G475), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n239), .A2(KEYINPUT20), .A3(new_n240), .A4(new_n241), .ZN(new_n249));
  AND3_X1   g063(.A1(new_n244), .A2(new_n248), .A3(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(G234), .A2(G237), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n251), .A2(G952), .A3(new_n204), .ZN(new_n252));
  XOR2_X1   g066(.A(KEYINPUT21), .B(G898), .Z(new_n253));
  NAND3_X1  g067(.A1(new_n251), .A2(G902), .A3(G953), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n252), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT92), .ZN(new_n256));
  INV_X1    g070(.A(G116), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G122), .ZN(new_n258));
  INV_X1    g072(.A(G122), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G116), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT91), .ZN(new_n261));
  AND3_X1   g075(.A1(new_n258), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n261), .B1(new_n258), .B2(new_n260), .ZN(new_n263));
  NOR3_X1   g077(.A1(new_n262), .A2(new_n263), .A3(G107), .ZN(new_n264));
  INV_X1    g078(.A(G107), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n259), .A2(G116), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n257), .A2(G122), .ZN(new_n267));
  OAI21_X1  g081(.A(KEYINPUT91), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n258), .A2(new_n260), .A3(new_n261), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n265), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n256), .B1(new_n264), .B2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT94), .ZN(new_n272));
  OAI21_X1  g086(.A(KEYINPUT93), .B1(new_n206), .B2(G128), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT93), .ZN(new_n274));
  INV_X1    g088(.A(G128), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n274), .A2(new_n275), .A3(G143), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n273), .A2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(G134), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n275), .A2(G143), .ZN(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  AND4_X1   g094(.A1(new_n272), .A2(new_n277), .A3(new_n278), .A4(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n279), .B1(new_n273), .B2(new_n276), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n272), .B1(new_n282), .B2(new_n278), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  OAI21_X1  g098(.A(G107), .B1(new_n262), .B2(new_n263), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n268), .A2(new_n265), .A3(new_n269), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n285), .A2(new_n286), .A3(KEYINPUT92), .ZN(new_n287));
  XNOR2_X1  g101(.A(new_n279), .B(KEYINPUT13), .ZN(new_n288));
  INV_X1    g102(.A(new_n277), .ZN(new_n289));
  OAI21_X1  g103(.A(G134), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND4_X1  g104(.A1(new_n271), .A2(new_n284), .A3(new_n287), .A4(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n266), .A2(KEYINPUT14), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n258), .A2(new_n260), .ZN(new_n293));
  OAI211_X1 g107(.A(new_n292), .B(G107), .C1(new_n293), .C2(KEYINPUT14), .ZN(new_n294));
  AND2_X1   g108(.A1(new_n282), .A2(new_n278), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n282), .A2(new_n278), .ZN(new_n296));
  OAI211_X1 g110(.A(new_n294), .B(new_n286), .C1(new_n295), .C2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n291), .A2(new_n297), .ZN(new_n298));
  XOR2_X1   g112(.A(KEYINPUT9), .B(G234), .Z(new_n299));
  NAND3_X1  g113(.A1(new_n299), .A2(G217), .A3(new_n204), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(new_n300), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n291), .A2(new_n297), .A3(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(G478), .ZN(new_n305));
  OR2_X1    g119(.A1(new_n305), .A2(KEYINPUT15), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n304), .A2(new_n241), .A3(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n306), .B1(new_n304), .B2(new_n241), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND4_X1  g124(.A1(new_n250), .A2(KEYINPUT95), .A3(new_n255), .A4(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT95), .ZN(new_n312));
  NAND4_X1  g126(.A1(new_n310), .A2(new_n244), .A3(new_n248), .A4(new_n249), .ZN(new_n313));
  INV_X1    g127(.A(new_n255), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n312), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  AND2_X1   g129(.A1(new_n311), .A2(new_n315), .ZN(new_n316));
  OAI21_X1  g130(.A(G214), .B1(G237), .B2(G902), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(KEYINPUT3), .B1(new_n223), .B2(G107), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT3), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n320), .A2(new_n265), .A3(G104), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n223), .A2(G107), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n319), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G101), .ZN(new_n324));
  INV_X1    g138(.A(G101), .ZN(new_n325));
  NAND4_X1  g139(.A1(new_n319), .A2(new_n321), .A3(new_n325), .A4(new_n322), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n324), .A2(KEYINPUT4), .A3(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT83), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  XOR2_X1   g143(.A(G116), .B(G119), .Z(new_n330));
  XNOR2_X1  g144(.A(KEYINPUT2), .B(G113), .ZN(new_n331));
  XNOR2_X1  g145(.A(new_n330), .B(new_n331), .ZN(new_n332));
  OR2_X1    g146(.A1(new_n324), .A2(KEYINPUT4), .ZN(new_n333));
  NAND4_X1  g147(.A1(new_n324), .A2(KEYINPUT83), .A3(KEYINPUT4), .A4(new_n326), .ZN(new_n334));
  NAND4_X1  g148(.A1(new_n329), .A2(new_n332), .A3(new_n333), .A4(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(new_n322), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n223), .A2(G107), .ZN(new_n337));
  OAI21_X1  g151(.A(G101), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  AND2_X1   g152(.A1(new_n338), .A2(new_n326), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT5), .ZN(new_n340));
  INV_X1    g154(.A(G119), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n340), .A2(new_n341), .A3(G116), .ZN(new_n342));
  OAI211_X1 g156(.A(G113), .B(new_n342), .C1(new_n330), .C2(new_n340), .ZN(new_n343));
  OAI211_X1 g157(.A(new_n339), .B(new_n343), .C1(new_n331), .C2(new_n330), .ZN(new_n344));
  XOR2_X1   g158(.A(G110), .B(G122), .Z(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  AND3_X1   g160(.A1(new_n335), .A2(new_n344), .A3(new_n346), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n346), .B1(new_n335), .B2(new_n344), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT6), .ZN(new_n349));
  NOR3_X1   g163(.A1(new_n347), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n335), .A2(new_n344), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(new_n345), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n352), .A2(KEYINPUT6), .ZN(new_n353));
  OAI21_X1  g167(.A(KEYINPUT84), .B1(new_n350), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n200), .A2(G143), .ZN(new_n355));
  AND3_X1   g169(.A1(new_n206), .A2(KEYINPUT65), .A3(G146), .ZN(new_n356));
  AOI21_X1  g170(.A(KEYINPUT65), .B1(new_n206), .B2(G146), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n355), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n275), .B1(new_n355), .B2(KEYINPUT1), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n206), .A2(G146), .ZN(new_n361));
  AND3_X1   g175(.A1(new_n355), .A2(new_n361), .A3(G128), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT1), .ZN(new_n363));
  AOI22_X1  g177(.A1(new_n358), .A2(new_n360), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(new_n190), .ZN(new_n365));
  NOR2_X1   g179(.A1(KEYINPUT0), .A2(G128), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(KEYINPUT0), .A2(G128), .ZN(new_n368));
  XNOR2_X1  g182(.A(new_n368), .B(KEYINPUT64), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n358), .A2(new_n367), .A3(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT66), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND4_X1  g186(.A1(new_n358), .A2(KEYINPUT66), .A3(new_n367), .A4(new_n369), .ZN(new_n373));
  INV_X1    g187(.A(new_n368), .ZN(new_n374));
  AND2_X1   g188(.A1(new_n355), .A2(new_n361), .ZN(new_n375));
  AOI22_X1  g189(.A1(new_n372), .A2(new_n373), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n365), .B1(new_n376), .B2(new_n190), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n204), .A2(G224), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  XNOR2_X1  g193(.A(new_n377), .B(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n335), .A2(new_n344), .A3(new_n346), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n352), .A2(KEYINPUT6), .A3(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT84), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n354), .A2(new_n380), .A3(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT7), .ZN(new_n386));
  OR3_X1    g200(.A1(new_n377), .A2(new_n386), .A3(new_n379), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(KEYINPUT87), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n339), .A2(KEYINPUT85), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n343), .B1(new_n331), .B2(new_n330), .ZN(new_n390));
  XNOR2_X1  g204(.A(new_n389), .B(new_n390), .ZN(new_n391));
  XOR2_X1   g205(.A(new_n345), .B(KEYINPUT8), .Z(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(KEYINPUT86), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT86), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n391), .A2(new_n395), .A3(new_n392), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n347), .B1(new_n394), .B2(new_n396), .ZN(new_n397));
  OR4_X1    g211(.A1(KEYINPUT87), .A2(new_n377), .A3(new_n386), .A4(new_n379), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n377), .B1(new_n386), .B2(new_n379), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n388), .A2(new_n397), .A3(new_n398), .A4(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n385), .A2(new_n241), .A3(new_n400), .ZN(new_n401));
  OAI21_X1  g215(.A(G210), .B1(G237), .B2(G902), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n385), .A2(new_n400), .A3(new_n241), .A4(new_n402), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n318), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(G221), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n407), .B1(new_n299), .B2(new_n241), .ZN(new_n408));
  INV_X1    g222(.A(G469), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n409), .A2(new_n241), .ZN(new_n410));
  OAI21_X1  g224(.A(KEYINPUT67), .B1(new_n278), .B2(G137), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(KEYINPUT11), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n278), .A2(G137), .ZN(new_n413));
  INV_X1    g227(.A(G137), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(G134), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT11), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n415), .A2(KEYINPUT67), .A3(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n412), .A2(new_n413), .A3(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT69), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n412), .A2(new_n417), .A3(KEYINPUT69), .A4(new_n413), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n420), .A2(G131), .A3(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT70), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n412), .A2(new_n417), .A3(new_n212), .A4(new_n413), .ZN(new_n425));
  OR2_X1    g239(.A1(new_n425), .A2(KEYINPUT68), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(KEYINPUT68), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND4_X1  g242(.A1(new_n420), .A2(KEYINPUT70), .A3(G131), .A4(new_n421), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n424), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n362), .A2(new_n363), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n432), .B1(new_n375), .B2(new_n359), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(new_n339), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT10), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n376), .A2(new_n333), .A3(new_n329), .A4(new_n334), .ZN(new_n437));
  INV_X1    g251(.A(new_n364), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n438), .A2(KEYINPUT10), .A3(new_n339), .ZN(new_n439));
  NAND4_X1  g253(.A1(new_n431), .A2(new_n436), .A3(new_n437), .A4(new_n439), .ZN(new_n440));
  XNOR2_X1  g254(.A(G110), .B(G140), .ZN(new_n441));
  AND2_X1   g255(.A1(new_n204), .A2(G227), .ZN(new_n442));
  XOR2_X1   g256(.A(new_n441), .B(new_n442), .Z(new_n443));
  NAND2_X1  g257(.A1(new_n440), .A2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n376), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n329), .A2(new_n333), .A3(new_n334), .ZN(new_n447));
  OAI211_X1 g261(.A(new_n436), .B(new_n439), .C1(new_n446), .C2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(new_n430), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n434), .B1(new_n438), .B2(new_n339), .ZN(new_n450));
  AND3_X1   g264(.A1(new_n430), .A2(KEYINPUT12), .A3(new_n450), .ZN(new_n451));
  AOI21_X1  g265(.A(KEYINPUT12), .B1(new_n430), .B2(new_n450), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n440), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(new_n443), .ZN(new_n454));
  AOI22_X1  g268(.A1(new_n445), .A2(new_n449), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n410), .B1(new_n455), .B2(G469), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n451), .A2(new_n452), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n444), .A2(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n443), .B1(new_n449), .B2(new_n440), .ZN(new_n459));
  OAI211_X1 g273(.A(new_n409), .B(new_n241), .C1(new_n458), .C2(new_n459), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n408), .B1(new_n456), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n406), .A2(new_n461), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n187), .B1(new_n316), .B2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT32), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT30), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT72), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n413), .A2(new_n415), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n466), .B1(new_n467), .B2(G131), .ZN(new_n468));
  AOI211_X1 g282(.A(KEYINPUT72), .B(new_n212), .C1(new_n413), .C2(new_n415), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  AOI211_X1 g284(.A(new_n470), .B(new_n364), .C1(new_n426), .C2(new_n427), .ZN(new_n471));
  AOI211_X1 g285(.A(new_n465), .B(new_n471), .C1(new_n376), .C2(new_n430), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT71), .ZN(new_n474));
  AND3_X1   g288(.A1(new_n430), .A2(new_n474), .A3(new_n376), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n474), .B1(new_n430), .B2(new_n376), .ZN(new_n476));
  NOR3_X1   g290(.A1(new_n475), .A2(new_n476), .A3(new_n471), .ZN(new_n477));
  OAI211_X1 g291(.A(new_n332), .B(new_n473), .C1(new_n477), .C2(KEYINPUT30), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n471), .B1(new_n430), .B2(new_n376), .ZN(new_n479));
  INV_X1    g293(.A(new_n332), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n203), .A2(new_n204), .A3(G210), .ZN(new_n482));
  XNOR2_X1  g296(.A(new_n482), .B(new_n325), .ZN(new_n483));
  XNOR2_X1  g297(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n484));
  XOR2_X1   g298(.A(new_n483), .B(new_n484), .Z(new_n485));
  NAND3_X1  g299(.A1(new_n478), .A2(new_n481), .A3(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT31), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(new_n481), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n430), .A2(new_n376), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(KEYINPUT71), .ZN(new_n491));
  INV_X1    g305(.A(new_n471), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n430), .A2(new_n474), .A3(new_n376), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n491), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n472), .B1(new_n494), .B2(new_n465), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n489), .B1(new_n495), .B2(new_n332), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n496), .A2(KEYINPUT31), .A3(new_n485), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT28), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n481), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n479), .A2(KEYINPUT28), .A3(new_n480), .ZN(new_n500));
  OAI211_X1 g314(.A(new_n499), .B(new_n500), .C1(new_n477), .C2(new_n480), .ZN(new_n501));
  INV_X1    g315(.A(new_n485), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(KEYINPUT73), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT73), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n501), .A2(new_n505), .A3(new_n502), .ZN(new_n506));
  AOI22_X1  g320(.A1(new_n488), .A2(new_n497), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  NOR2_X1   g321(.A1(G472), .A2(G902), .ZN(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n464), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(KEYINPUT31), .B1(new_n496), .B2(new_n485), .ZN(new_n511));
  AND4_X1   g325(.A1(KEYINPUT31), .A2(new_n478), .A3(new_n481), .A4(new_n485), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n505), .B1(new_n501), .B2(new_n502), .ZN(new_n513));
  AND3_X1   g327(.A1(new_n501), .A2(new_n505), .A3(new_n502), .ZN(new_n514));
  OAI22_X1  g328(.A1(new_n511), .A2(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n515), .A2(KEYINPUT32), .A3(new_n508), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n481), .A2(KEYINPUT76), .A3(new_n498), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT76), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n499), .A2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT74), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n481), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n479), .A2(KEYINPUT74), .A3(new_n480), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n490), .A2(new_n492), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n523), .A2(KEYINPUT75), .A3(new_n332), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT75), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n525), .B1(new_n479), .B2(new_n480), .ZN(new_n526));
  AOI22_X1  g340(.A1(new_n521), .A2(new_n522), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n517), .B(new_n519), .C1(new_n527), .C2(new_n498), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n485), .B1(new_n501), .B2(KEYINPUT29), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n241), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n478), .A2(new_n481), .A3(new_n502), .ZN(new_n531));
  AOI21_X1  g345(.A(KEYINPUT29), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  OAI21_X1  g346(.A(G472), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n510), .A2(new_n516), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n201), .A2(new_n202), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT80), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n536), .B1(new_n341), .B2(G128), .ZN(new_n537));
  OR2_X1    g351(.A1(new_n537), .A2(KEYINPUT23), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(KEYINPUT23), .ZN(new_n539));
  OAI211_X1 g353(.A(new_n538), .B(new_n539), .C1(G119), .C2(new_n275), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT79), .ZN(new_n541));
  XOR2_X1   g355(.A(KEYINPUT24), .B(G110), .Z(new_n542));
  XNOR2_X1  g356(.A(G119), .B(G128), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AOI22_X1  g358(.A1(new_n540), .A2(G110), .B1(new_n541), .B2(new_n544), .ZN(new_n545));
  OAI211_X1 g359(.A(new_n535), .B(new_n545), .C1(new_n541), .C2(new_n544), .ZN(new_n546));
  OAI22_X1  g360(.A1(new_n540), .A2(G110), .B1(new_n543), .B2(new_n542), .ZN(new_n547));
  OAI211_X1 g361(.A(new_n547), .B(new_n202), .C1(G146), .C2(new_n192), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  XNOR2_X1  g363(.A(KEYINPUT22), .B(G137), .ZN(new_n550));
  INV_X1    g364(.A(G234), .ZN(new_n551));
  NOR3_X1   g365(.A1(new_n407), .A2(new_n551), .A3(G953), .ZN(new_n552));
  XOR2_X1   g366(.A(new_n550), .B(new_n552), .Z(new_n553));
  XNOR2_X1  g367(.A(new_n549), .B(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  OAI21_X1  g369(.A(G217), .B1(new_n551), .B2(G902), .ZN(new_n556));
  XNOR2_X1  g370(.A(new_n556), .B(KEYINPUT77), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(new_n241), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n555), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n554), .A2(new_n241), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(KEYINPUT82), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n561), .B(KEYINPUT25), .ZN(new_n562));
  XNOR2_X1  g376(.A(new_n557), .B(KEYINPUT78), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n559), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n311), .A2(new_n315), .ZN(new_n565));
  NAND4_X1  g379(.A1(new_n565), .A2(KEYINPUT96), .A3(new_n406), .A4(new_n461), .ZN(new_n566));
  NAND4_X1  g380(.A1(new_n463), .A2(new_n534), .A3(new_n564), .A4(new_n566), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n567), .B(G101), .ZN(G3));
  INV_X1    g382(.A(G472), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n569), .B1(new_n515), .B2(new_n241), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n507), .A2(new_n509), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n462), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n572), .A2(new_n564), .A3(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n244), .A2(new_n248), .A3(new_n249), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT98), .ZN(new_n576));
  AND3_X1   g390(.A1(new_n291), .A2(KEYINPUT97), .A3(new_n297), .ZN(new_n577));
  AOI21_X1  g391(.A(KEYINPUT97), .B1(new_n291), .B2(new_n297), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n576), .B1(new_n579), .B2(new_n300), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT97), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n298), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n291), .A2(new_n297), .A3(KEYINPUT97), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n582), .A2(new_n576), .A3(new_n300), .A4(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(new_n303), .ZN(new_n585));
  OAI21_X1  g399(.A(KEYINPUT33), .B1(new_n580), .B2(new_n585), .ZN(new_n586));
  OR2_X1    g400(.A1(new_n304), .A2(KEYINPUT33), .ZN(new_n587));
  AOI211_X1 g401(.A(new_n305), .B(G902), .C1(new_n586), .C2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n304), .A2(new_n241), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(new_n305), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  OAI211_X1 g405(.A(new_n255), .B(new_n575), .C1(new_n588), .C2(new_n591), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n574), .A2(new_n592), .ZN(new_n593));
  XNOR2_X1  g407(.A(KEYINPUT34), .B(G104), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n593), .B(new_n594), .ZN(G6));
  INV_X1    g409(.A(new_n310), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n250), .A2(new_n596), .ZN(new_n597));
  OR3_X1    g411(.A1(new_n597), .A2(KEYINPUT99), .A3(new_n314), .ZN(new_n598));
  OAI21_X1  g412(.A(KEYINPUT99), .B1(new_n597), .B2(new_n314), .ZN(new_n599));
  AND2_X1   g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n574), .A2(new_n601), .ZN(new_n602));
  XNOR2_X1  g416(.A(KEYINPUT35), .B(G107), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n602), .B(new_n603), .ZN(G9));
  NAND2_X1  g418(.A1(new_n562), .A2(new_n563), .ZN(new_n605));
  INV_X1    g419(.A(new_n553), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n606), .A2(KEYINPUT36), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n549), .B(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n608), .A2(new_n241), .A3(new_n557), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n605), .A2(new_n609), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n463), .A2(new_n572), .A3(new_n566), .A4(new_n610), .ZN(new_n611));
  XOR2_X1   g425(.A(KEYINPUT37), .B(G110), .Z(new_n612));
  XNOR2_X1  g426(.A(new_n611), .B(new_n612), .ZN(G12));
  OR2_X1    g427(.A1(new_n254), .A2(G900), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(new_n252), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n597), .A2(new_n616), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n534), .A2(new_n573), .A3(new_n610), .A4(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(G128), .ZN(G30));
  NAND2_X1  g433(.A1(new_n404), .A2(new_n405), .ZN(new_n620));
  XOR2_X1   g434(.A(KEYINPUT100), .B(KEYINPUT38), .Z(new_n621));
  XNOR2_X1  g435(.A(new_n620), .B(new_n621), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n622), .A2(new_n318), .ZN(new_n623));
  INV_X1    g437(.A(new_n610), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n496), .A2(new_n502), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n527), .A2(new_n502), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(new_n241), .ZN(new_n627));
  OAI21_X1  g441(.A(G472), .B1(new_n625), .B2(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n510), .A2(new_n516), .A3(new_n628), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n250), .A2(new_n310), .ZN(new_n630));
  NAND4_X1  g444(.A1(new_n623), .A2(new_n624), .A3(new_n629), .A4(new_n630), .ZN(new_n631));
  OR2_X1    g445(.A1(new_n631), .A2(KEYINPUT101), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n631), .A2(KEYINPUT101), .ZN(new_n633));
  XNOR2_X1  g447(.A(KEYINPUT102), .B(KEYINPUT39), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n615), .B(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n461), .A2(new_n636), .ZN(new_n637));
  XOR2_X1   g451(.A(new_n637), .B(KEYINPUT40), .Z(new_n638));
  NAND3_X1  g452(.A1(new_n632), .A2(new_n633), .A3(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(KEYINPUT103), .B(G143), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G45));
  NAND2_X1  g455(.A1(new_n586), .A2(new_n587), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n642), .A2(G478), .A3(new_n241), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n250), .B1(new_n643), .B2(new_n590), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(new_n615), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n534), .A2(new_n573), .A3(new_n610), .A4(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(G146), .ZN(G48));
  NOR2_X1   g462(.A1(new_n458), .A2(new_n459), .ZN(new_n649));
  OAI21_X1  g463(.A(G469), .B1(new_n649), .B2(G902), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT104), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n650), .A2(new_n651), .A3(new_n460), .ZN(new_n652));
  OAI211_X1 g466(.A(KEYINPUT104), .B(G469), .C1(new_n649), .C2(G902), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n408), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  AND2_X1   g468(.A1(new_n654), .A2(new_n406), .ZN(new_n655));
  INV_X1    g469(.A(new_n592), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n534), .A2(new_n655), .A3(new_n564), .A4(new_n656), .ZN(new_n657));
  XOR2_X1   g471(.A(KEYINPUT41), .B(G113), .Z(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(KEYINPUT105), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n657), .B(new_n659), .ZN(G15));
  NAND4_X1  g474(.A1(new_n600), .A2(new_n534), .A3(new_n564), .A4(new_n655), .ZN(new_n661));
  XNOR2_X1  g475(.A(KEYINPUT106), .B(G116), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G18));
  NAND4_X1  g477(.A1(new_n534), .A2(new_n655), .A3(new_n565), .A4(new_n610), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(G119), .ZN(G21));
  INV_X1    g479(.A(new_n559), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n605), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n488), .A2(new_n497), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n528), .A2(new_n502), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n509), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NOR3_X1   g484(.A1(new_n570), .A2(new_n667), .A3(new_n670), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n654), .A2(new_n255), .A3(new_n406), .A4(new_n630), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  AOI21_X1  g487(.A(KEYINPUT107), .B1(new_n671), .B2(new_n673), .ZN(new_n674));
  OAI21_X1  g488(.A(G472), .B1(new_n507), .B2(G902), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n669), .B1(new_n511), .B2(new_n512), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(new_n508), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n675), .A2(new_n564), .A3(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT107), .ZN(new_n679));
  NOR3_X1   g493(.A1(new_n678), .A2(new_n679), .A3(new_n672), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n674), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(new_n259), .ZN(G24));
  NOR2_X1   g496(.A1(new_n570), .A2(new_n670), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n683), .A2(new_n655), .A3(new_n610), .A4(new_n646), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G125), .ZN(G27));
  AND2_X1   g499(.A1(new_n534), .A2(new_n564), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n461), .A2(new_n317), .A3(new_n404), .A4(new_n405), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n686), .A2(new_n646), .A3(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT42), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT109), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n510), .A2(new_n516), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT108), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  OR2_X1    g509(.A1(new_n530), .A2(new_n532), .ZN(new_n696));
  AOI22_X1  g510(.A1(new_n516), .A2(KEYINPUT108), .B1(new_n696), .B2(G472), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n667), .B1(new_n695), .B2(new_n697), .ZN(new_n698));
  NOR3_X1   g512(.A1(new_n645), .A2(new_n687), .A3(new_n690), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n692), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NOR3_X1   g514(.A1(new_n507), .A2(new_n464), .A3(new_n509), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n533), .B1(new_n701), .B2(new_n694), .ZN(new_n702));
  AOI21_X1  g516(.A(KEYINPUT108), .B1(new_n510), .B2(new_n516), .ZN(new_n703));
  OAI211_X1 g517(.A(new_n564), .B(new_n699), .C1(new_n702), .C2(new_n703), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n704), .A2(KEYINPUT109), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n691), .B1(new_n700), .B2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(KEYINPUT110), .B(G131), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n706), .B(new_n707), .ZN(G33));
  NAND2_X1  g522(.A1(new_n686), .A2(new_n688), .ZN(new_n709));
  NOR3_X1   g523(.A1(new_n709), .A2(new_n597), .A3(new_n616), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(new_n278), .ZN(G36));
  INV_X1    g525(.A(KEYINPUT46), .ZN(new_n712));
  OR2_X1    g526(.A1(new_n455), .A2(KEYINPUT45), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n455), .A2(KEYINPUT45), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n713), .A2(G469), .A3(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(new_n715), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n712), .B1(new_n716), .B2(new_n410), .ZN(new_n717));
  INV_X1    g531(.A(new_n410), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n715), .A2(KEYINPUT46), .A3(new_n718), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n717), .A2(new_n460), .A3(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(new_n408), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n720), .A2(new_n721), .A3(new_n636), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n588), .A2(new_n591), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n723), .A2(new_n575), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(KEYINPUT43), .ZN(new_n725));
  OAI211_X1 g539(.A(new_n725), .B(new_n610), .C1(new_n571), .C2(new_n570), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT44), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n722), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n404), .A2(new_n317), .A3(new_n405), .ZN(new_n729));
  INV_X1    g543(.A(new_n729), .ZN(new_n730));
  OAI211_X1 g544(.A(new_n728), .B(new_n730), .C1(new_n727), .C2(new_n726), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G137), .ZN(G39));
  NAND2_X1  g546(.A1(new_n720), .A2(new_n721), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT47), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n720), .A2(KEYINPUT47), .A3(new_n721), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n534), .A2(new_n564), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n737), .A2(new_n646), .A3(new_n730), .A4(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G140), .ZN(G42));
  NAND2_X1  g554(.A1(new_n204), .A2(G952), .ZN(new_n741));
  INV_X1    g555(.A(new_n252), .ZN(new_n742));
  AND3_X1   g556(.A1(new_n725), .A2(new_n742), .A3(new_n671), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n741), .B1(new_n743), .B2(new_n655), .ZN(new_n744));
  AND2_X1   g558(.A1(new_n725), .A2(new_n742), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n654), .A2(new_n730), .ZN(new_n746));
  INV_X1    g560(.A(new_n746), .ZN(new_n747));
  AND3_X1   g561(.A1(new_n745), .A2(new_n698), .A3(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT48), .ZN(new_n749));
  AND2_X1   g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n748), .A2(new_n749), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n744), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  AND2_X1   g566(.A1(new_n652), .A2(new_n653), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n753), .A2(new_n721), .ZN(new_n754));
  OAI211_X1 g568(.A(new_n730), .B(new_n743), .C1(new_n737), .C2(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n622), .A2(new_n318), .A3(new_n654), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(KEYINPUT115), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT116), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT50), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n758), .A2(new_n759), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n757), .A2(new_n743), .A3(new_n761), .A4(new_n762), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n629), .A2(new_n746), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n667), .A2(new_n252), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n764), .A2(new_n250), .A3(new_n723), .A4(new_n765), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n745), .A2(new_n610), .A3(new_n683), .A4(new_n747), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n755), .A2(new_n763), .A3(new_n766), .A4(new_n767), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n761), .B1(new_n757), .B2(new_n743), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n755), .A2(KEYINPUT117), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(KEYINPUT51), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  OAI211_X1 g587(.A(KEYINPUT51), .B(new_n771), .C1(new_n768), .C2(new_n769), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n752), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n764), .A2(new_n644), .A3(new_n765), .ZN(new_n776));
  AND3_X1   g590(.A1(new_n775), .A2(KEYINPUT118), .A3(new_n776), .ZN(new_n777));
  AOI21_X1  g591(.A(KEYINPUT118), .B1(new_n775), .B2(new_n776), .ZN(new_n778));
  OR2_X1    g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT114), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT53), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n597), .A2(new_n314), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n572), .A2(new_n564), .A3(new_n573), .A4(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n611), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n620), .A2(new_n317), .ZN(new_n785));
  OAI21_X1  g599(.A(KEYINPUT111), .B1(new_n785), .B2(new_n592), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT111), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n644), .A2(new_n406), .A3(new_n787), .A4(new_n255), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n789), .A2(new_n564), .A3(new_n461), .A4(new_n572), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n790), .A2(new_n567), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(KEYINPUT112), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT112), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n790), .A2(new_n567), .A3(new_n793), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n784), .B1(new_n792), .B2(new_n794), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n657), .B1(new_n674), .B2(new_n680), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT113), .ZN(new_n797));
  INV_X1    g611(.A(new_n313), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n730), .A2(new_n797), .A3(new_n798), .A4(new_n615), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n404), .A2(new_n317), .A3(new_n405), .A4(new_n615), .ZN(new_n800));
  OAI21_X1  g614(.A(KEYINPUT113), .B1(new_n800), .B2(new_n313), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n802), .A2(new_n534), .A3(new_n461), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n683), .A2(new_n646), .A3(new_n688), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n624), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n661), .A2(new_n664), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n796), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n710), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n795), .A2(new_n706), .A3(new_n807), .A4(new_n808), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n462), .A2(new_n616), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n629), .A2(new_n624), .A3(new_n630), .A4(new_n810), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n618), .A2(new_n647), .A3(new_n811), .A4(new_n684), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(KEYINPUT52), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n781), .B1(new_n809), .B2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(new_n681), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n803), .A2(new_n804), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(new_n610), .ZN(new_n817));
  INV_X1    g631(.A(new_n806), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n815), .A2(new_n657), .A3(new_n817), .A4(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(new_n784), .ZN(new_n820));
  AND3_X1   g634(.A1(new_n790), .A2(new_n793), .A3(new_n567), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n793), .B1(new_n790), .B2(new_n567), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n820), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n819), .A2(new_n823), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n704), .B(KEYINPUT109), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n710), .B1(new_n825), .B2(new_n691), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT52), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n812), .B(new_n827), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n824), .A2(KEYINPUT53), .A3(new_n826), .A4(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n814), .A2(KEYINPUT54), .A3(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(new_n830), .ZN(new_n831));
  AOI21_X1  g645(.A(KEYINPUT54), .B1(new_n814), .B2(new_n829), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n780), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(new_n832), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n834), .A2(KEYINPUT114), .A3(new_n830), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  OAI22_X1  g650(.A1(new_n779), .A2(new_n836), .B1(G952), .B2(G953), .ZN(new_n837));
  OR2_X1    g651(.A1(new_n753), .A2(KEYINPUT49), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n753), .A2(KEYINPUT49), .ZN(new_n839));
  AND4_X1   g653(.A1(new_n564), .A2(new_n838), .A3(new_n317), .A4(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(new_n629), .ZN(new_n841));
  NOR3_X1   g655(.A1(new_n723), .A2(new_n575), .A3(new_n408), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n840), .A2(new_n841), .A3(new_n622), .A4(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n837), .A2(new_n843), .ZN(G75));
  AOI21_X1  g658(.A(new_n241), .B1(new_n814), .B2(new_n829), .ZN(new_n845));
  AOI21_X1  g659(.A(KEYINPUT56), .B1(new_n845), .B2(G210), .ZN(new_n846));
  AND2_X1   g660(.A1(new_n354), .A2(new_n384), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n847), .B(new_n380), .ZN(new_n848));
  XNOR2_X1  g662(.A(new_n848), .B(KEYINPUT55), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT56), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n849), .B1(KEYINPUT119), .B2(new_n850), .ZN(new_n851));
  XNOR2_X1  g665(.A(new_n846), .B(new_n851), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n204), .A2(G952), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n852), .A2(new_n853), .ZN(G51));
  NOR2_X1   g668(.A1(new_n831), .A2(new_n832), .ZN(new_n855));
  XOR2_X1   g669(.A(KEYINPUT120), .B(KEYINPUT57), .Z(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(new_n410), .ZN(new_n857));
  OR2_X1    g671(.A1(new_n856), .A2(new_n410), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n855), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n859), .B1(new_n459), .B2(new_n458), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n845), .A2(new_n716), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n853), .B1(new_n860), .B2(new_n861), .ZN(G54));
  NAND3_X1  g676(.A1(new_n845), .A2(KEYINPUT58), .A3(G475), .ZN(new_n863));
  XOR2_X1   g677(.A(new_n863), .B(new_n239), .Z(new_n864));
  NOR2_X1   g678(.A1(new_n864), .A2(new_n853), .ZN(G60));
  INV_X1    g679(.A(new_n853), .ZN(new_n866));
  NAND2_X1  g680(.A1(G478), .A2(G902), .ZN(new_n867));
  XOR2_X1   g681(.A(new_n867), .B(KEYINPUT59), .Z(new_n868));
  INV_X1    g682(.A(new_n868), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n855), .A2(new_n642), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n868), .B1(new_n833), .B2(new_n835), .ZN(new_n871));
  OAI211_X1 g685(.A(new_n866), .B(new_n870), .C1(new_n871), .C2(new_n642), .ZN(new_n872));
  INV_X1    g686(.A(new_n872), .ZN(G63));
  NAND2_X1  g687(.A1(new_n814), .A2(new_n829), .ZN(new_n874));
  NAND2_X1  g688(.A1(G217), .A2(G902), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n875), .B(KEYINPUT122), .ZN(new_n876));
  XNOR2_X1  g690(.A(KEYINPUT121), .B(KEYINPUT60), .ZN(new_n877));
  XOR2_X1   g691(.A(new_n876), .B(new_n877), .Z(new_n878));
  NAND2_X1  g692(.A1(new_n874), .A2(new_n878), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n853), .B1(new_n879), .B2(new_n555), .ZN(new_n880));
  INV_X1    g694(.A(new_n878), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n881), .B1(new_n814), .B2(new_n829), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(new_n608), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  OAI211_X1 g698(.A(KEYINPUT123), .B(new_n866), .C1(new_n882), .C2(new_n554), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT124), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT61), .ZN(new_n887));
  AND3_X1   g701(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n886), .B1(new_n885), .B2(new_n887), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n884), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n885), .A2(new_n887), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n891), .A2(KEYINPUT124), .ZN(new_n892));
  AND2_X1   g706(.A1(new_n880), .A2(new_n883), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  AND2_X1   g709(.A1(new_n890), .A2(new_n895), .ZN(G66));
  AOI21_X1  g710(.A(new_n204), .B1(new_n253), .B2(G224), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n795), .A2(new_n657), .A3(new_n815), .A4(new_n818), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n897), .B1(new_n898), .B2(new_n204), .ZN(new_n899));
  INV_X1    g713(.A(G898), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n847), .B1(new_n900), .B2(G953), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n899), .B(new_n901), .ZN(G69));
  INV_X1    g716(.A(new_n644), .ZN(new_n903));
  AOI211_X1 g717(.A(new_n635), .B(new_n709), .C1(new_n903), .C2(new_n597), .ZN(new_n904));
  AND3_X1   g718(.A1(new_n618), .A2(new_n647), .A3(new_n684), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n639), .A2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT62), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n639), .A2(KEYINPUT62), .A3(new_n905), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n904), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  AND2_X1   g724(.A1(new_n731), .A2(new_n739), .ZN(new_n911));
  AOI21_X1  g725(.A(G953), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  XOR2_X1   g726(.A(new_n495), .B(new_n234), .Z(new_n913));
  OR3_X1    g727(.A1(new_n912), .A2(KEYINPUT125), .A3(new_n913), .ZN(new_n914));
  OAI21_X1  g728(.A(KEYINPUT125), .B1(new_n912), .B2(new_n913), .ZN(new_n915));
  NAND2_X1  g729(.A1(G900), .A2(G953), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n826), .B(KEYINPUT126), .ZN(new_n917));
  INV_X1    g731(.A(new_n905), .ZN(new_n918));
  NOR4_X1   g732(.A1(new_n722), .A2(new_n310), .A3(new_n250), .A4(new_n785), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n918), .B1(new_n698), .B2(new_n919), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n917), .A2(new_n920), .A3(new_n911), .ZN(new_n921));
  OAI211_X1 g735(.A(new_n916), .B(new_n913), .C1(new_n921), .C2(G953), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n914), .A2(new_n915), .A3(new_n922), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n204), .B1(G227), .B2(G900), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n923), .B(new_n924), .ZN(G72));
  NAND2_X1  g739(.A1(G472), .A2(G902), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n926), .B(KEYINPUT63), .Z(new_n927));
  NAND2_X1  g741(.A1(new_n910), .A2(new_n911), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n927), .B1(new_n928), .B2(new_n898), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n929), .A2(new_n625), .ZN(new_n930));
  INV_X1    g744(.A(new_n531), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n625), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n874), .A2(new_n927), .A3(new_n932), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n930), .A2(new_n866), .A3(new_n933), .ZN(new_n934));
  OR2_X1    g748(.A1(new_n921), .A2(new_n898), .ZN(new_n935));
  AND3_X1   g749(.A1(new_n935), .A2(KEYINPUT127), .A3(new_n927), .ZN(new_n936));
  AOI21_X1  g750(.A(KEYINPUT127), .B1(new_n935), .B2(new_n927), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n934), .B1(new_n938), .B2(new_n931), .ZN(G57));
endmodule


