//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 1 0 1 0 1 0 0 0 1 0 0 1 0 1 1 0 0 0 1 0 1 1 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 0 0 0 1 1 0 0 0 0 1 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:35 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n456, new_n457, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n566, new_n568, new_n569, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n581, new_n582,
    new_n583, new_n584, new_n586, new_n587, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n621, new_n623, new_n624, new_n625, new_n626,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1184,
    new_n1185, new_n1187, new_n1188, new_n1189;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT65), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XOR2_X1   g013(.A(KEYINPUT66), .B(G120), .Z(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g018(.A(KEYINPUT67), .B(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  OR4_X1    g026(.A1(G237), .A2(G236), .A3(G235), .A4(G238), .ZN(new_n452));
  NOR2_X1   g027(.A1(new_n451), .A2(new_n452), .ZN(G325));
  INV_X1    g028(.A(G325), .ZN(G261));
  AOI22_X1  g029(.A1(new_n451), .A2(G2106), .B1(G567), .B2(new_n452), .ZN(G319));
  NAND2_X1  g030(.A1(G113), .A2(G2104), .ZN(new_n456));
  XOR2_X1   g031(.A(KEYINPUT3), .B(G2104), .Z(new_n457));
  INV_X1    g032(.A(G125), .ZN(new_n458));
  OAI21_X1  g033(.A(new_n456), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G2105), .ZN(new_n460));
  AND2_X1   g035(.A1(KEYINPUT68), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT68), .A2(G2104), .ZN(new_n462));
  OR2_X1    g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n463), .A2(G2105), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G101), .ZN(new_n465));
  OR2_X1    g040(.A1(KEYINPUT69), .A2(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(KEYINPUT69), .A2(KEYINPUT3), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n466), .A2(G2104), .A3(new_n467), .ZN(new_n468));
  OAI21_X1  g043(.A(KEYINPUT3), .B1(new_n461), .B2(new_n462), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  NAND4_X1  g045(.A1(new_n468), .A2(new_n469), .A3(G137), .A4(new_n470), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n460), .A2(new_n465), .A3(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(new_n472), .ZN(G160));
  NAND3_X1  g048(.A1(new_n468), .A2(new_n469), .A3(G2105), .ZN(new_n474));
  XNOR2_X1  g049(.A(new_n474), .B(KEYINPUT70), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n468), .A2(new_n469), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n476), .A2(G2105), .ZN(new_n477));
  AOI22_X1  g052(.A1(new_n475), .A2(G124), .B1(G136), .B2(new_n477), .ZN(new_n478));
  OAI21_X1  g053(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n479));
  INV_X1    g054(.A(G112), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n479), .B1(new_n480), .B2(G2105), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  AND2_X1   g057(.A1(new_n478), .A2(new_n482), .ZN(G162));
  NAND4_X1  g058(.A1(new_n468), .A2(new_n469), .A3(G138), .A4(new_n470), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(KEYINPUT4), .ZN(new_n485));
  INV_X1    g060(.A(G138), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT4), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(KEYINPUT71), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT71), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(KEYINPUT4), .ZN(new_n490));
  AOI211_X1 g065(.A(new_n486), .B(G2105), .C1(new_n488), .C2(new_n490), .ZN(new_n491));
  XNOR2_X1  g066(.A(KEYINPUT3), .B(G2104), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n485), .A2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT72), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n468), .A2(new_n469), .A3(G126), .A4(G2105), .ZN(new_n496));
  OR2_X1    g071(.A1(G102), .A2(G2105), .ZN(new_n497));
  OAI211_X1 g072(.A(new_n497), .B(G2104), .C1(G114), .C2(new_n470), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n494), .A2(new_n495), .A3(new_n500), .ZN(new_n501));
  AOI22_X1  g076(.A1(new_n484), .A2(KEYINPUT4), .B1(new_n491), .B2(new_n492), .ZN(new_n502));
  OAI21_X1  g077(.A(KEYINPUT72), .B1(new_n502), .B2(new_n499), .ZN(new_n503));
  AND2_X1   g078(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(G164));
  XNOR2_X1  g080(.A(KEYINPUT6), .B(G651), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(G543), .ZN(new_n507));
  INV_X1    g082(.A(G50), .ZN(new_n508));
  INV_X1    g083(.A(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(KEYINPUT5), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT5), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G543), .ZN(new_n512));
  INV_X1    g087(.A(G651), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(KEYINPUT6), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT6), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G651), .ZN(new_n516));
  NAND4_X1  g091(.A1(new_n510), .A2(new_n512), .A3(new_n514), .A4(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(G88), .ZN(new_n518));
  OAI22_X1  g093(.A1(new_n507), .A2(new_n508), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT73), .ZN(new_n520));
  XNOR2_X1  g095(.A(new_n519), .B(new_n520), .ZN(new_n521));
  XNOR2_X1  g096(.A(KEYINPUT5), .B(G543), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n522), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n523));
  OR2_X1    g098(.A1(new_n523), .A2(new_n513), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n521), .A2(new_n524), .ZN(G303));
  INV_X1    g100(.A(G303), .ZN(G166));
  INV_X1    g101(.A(new_n507), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G51), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n522), .A2(G63), .A3(G651), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n522), .A2(new_n506), .A3(G89), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT74), .ZN(new_n531));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(KEYINPUT7), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT7), .ZN(new_n534));
  NAND4_X1  g109(.A1(new_n534), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  AND3_X1   g111(.A1(new_n530), .A2(new_n531), .A3(new_n536), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n531), .B1(new_n530), .B2(new_n536), .ZN(new_n538));
  OAI211_X1 g113(.A(new_n528), .B(new_n529), .C1(new_n537), .C2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT75), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(G89), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n536), .B1(new_n517), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(KEYINPUT74), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n530), .A2(new_n531), .A3(new_n536), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND4_X1  g121(.A1(new_n546), .A2(KEYINPUT75), .A3(new_n528), .A4(new_n529), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n541), .A2(new_n547), .ZN(G168));
  AOI22_X1  g123(.A1(new_n522), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n549), .A2(new_n513), .ZN(new_n550));
  INV_X1    g125(.A(G52), .ZN(new_n551));
  INV_X1    g126(.A(G90), .ZN(new_n552));
  OAI22_X1  g127(.A1(new_n507), .A2(new_n551), .B1(new_n517), .B2(new_n552), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n550), .A2(new_n553), .ZN(G171));
  AOI22_X1  g129(.A1(new_n522), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n555), .A2(new_n513), .ZN(new_n556));
  INV_X1    g131(.A(G43), .ZN(new_n557));
  INV_X1    g132(.A(G81), .ZN(new_n558));
  OAI22_X1  g133(.A1(new_n507), .A2(new_n557), .B1(new_n517), .B2(new_n558), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT76), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  OAI21_X1  g137(.A(KEYINPUT76), .B1(new_n556), .B2(new_n559), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G860), .ZN(G153));
  AND3_X1   g140(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G36), .ZN(G176));
  NAND2_X1  g142(.A1(G1), .A2(G3), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT8), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n566), .A2(new_n569), .ZN(G188));
  AND3_X1   g145(.A1(new_n506), .A2(G53), .A3(G543), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT9), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n571), .B(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT77), .ZN(new_n574));
  XNOR2_X1  g149(.A(new_n517), .B(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(G91), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n522), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n577));
  OR2_X1    g152(.A1(new_n577), .A2(new_n513), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n573), .A2(new_n576), .A3(new_n578), .ZN(G299));
  INV_X1    g154(.A(G171), .ZN(G301));
  INV_X1    g155(.A(KEYINPUT78), .ZN(new_n581));
  AND3_X1   g156(.A1(new_n541), .A2(new_n581), .A3(new_n547), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n581), .B1(new_n541), .B2(new_n547), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(new_n584), .ZN(G286));
  AOI22_X1  g160(.A1(new_n575), .A2(G87), .B1(G49), .B2(new_n527), .ZN(new_n586));
  OAI21_X1  g161(.A(G651), .B1(new_n522), .B2(G74), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(G288));
  NAND2_X1  g163(.A1(new_n522), .A2(G61), .ZN(new_n589));
  NAND2_X1  g164(.A1(G73), .A2(G543), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT79), .ZN(new_n591));
  XNOR2_X1  g166(.A(new_n590), .B(new_n591), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n513), .B1(new_n589), .B2(new_n592), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n506), .A2(G48), .A3(G543), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(new_n595));
  AOI211_X1 g170(.A(new_n593), .B(new_n595), .C1(new_n575), .C2(G86), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(G305));
  AOI22_X1  g172(.A1(new_n522), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n598), .A2(new_n513), .ZN(new_n599));
  XNOR2_X1  g174(.A(new_n599), .B(KEYINPUT80), .ZN(new_n600));
  INV_X1    g175(.A(new_n517), .ZN(new_n601));
  AOI22_X1  g176(.A1(G47), .A2(new_n527), .B1(new_n601), .B2(G85), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n600), .A2(new_n602), .ZN(G290));
  NAND2_X1  g178(.A1(G301), .A2(G868), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n575), .A2(G92), .ZN(new_n605));
  XOR2_X1   g180(.A(KEYINPUT81), .B(KEYINPUT10), .Z(new_n606));
  INV_X1    g181(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(G79), .A2(G543), .ZN(new_n609));
  INV_X1    g184(.A(new_n522), .ZN(new_n610));
  INV_X1    g185(.A(G66), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n609), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n612), .A2(G651), .B1(new_n527), .B2(G54), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n575), .A2(G92), .A3(new_n606), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n608), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n604), .B1(new_n616), .B2(G868), .ZN(G284));
  OAI21_X1  g192(.A(new_n604), .B1(new_n616), .B2(G868), .ZN(G321));
  MUX2_X1   g193(.A(G299), .B(G286), .S(G868), .Z(G297));
  XOR2_X1   g194(.A(G297), .B(KEYINPUT82), .Z(G280));
  INV_X1    g195(.A(G559), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n616), .B1(new_n621), .B2(G860), .ZN(G148));
  NAND2_X1  g197(.A1(new_n616), .A2(new_n621), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n623), .A2(G868), .ZN(new_n624));
  OR2_X1    g199(.A1(new_n624), .A2(KEYINPUT83), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n624), .A2(KEYINPUT83), .ZN(new_n626));
  OAI211_X1 g201(.A(new_n625), .B(new_n626), .C1(G868), .C2(new_n564), .ZN(G323));
  XNOR2_X1  g202(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g203(.A1(new_n475), .A2(G123), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n477), .A2(G135), .ZN(new_n630));
  OR2_X1    g205(.A1(G99), .A2(G2105), .ZN(new_n631));
  OAI211_X1 g206(.A(new_n631), .B(G2104), .C1(G111), .C2(new_n470), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n629), .A2(new_n630), .A3(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(KEYINPUT85), .B(G2096), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  NOR3_X1   g210(.A1(new_n463), .A2(new_n457), .A3(G2105), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT84), .B(KEYINPUT12), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n636), .B(new_n637), .Z(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT13), .B(G2100), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n635), .A2(new_n640), .ZN(G156));
  XNOR2_X1  g216(.A(G2427), .B(G2438), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G2430), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT15), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n644), .B(G2435), .Z(new_n645));
  NAND2_X1  g220(.A1(new_n645), .A2(KEYINPUT14), .ZN(new_n646));
  XOR2_X1   g221(.A(G2443), .B(G2446), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G1341), .B(G1348), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT16), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n648), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2451), .B(G2454), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  INV_X1    g228(.A(G14), .ZN(new_n654));
  OR2_X1    g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(G401));
  XOR2_X1   g231(.A(G2084), .B(G2090), .Z(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(G2067), .B(G2678), .Z(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2072), .B(G2078), .ZN(new_n661));
  OAI21_X1  g236(.A(new_n658), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n662), .B(KEYINPUT86), .Z(new_n663));
  XOR2_X1   g238(.A(new_n661), .B(KEYINPUT17), .Z(new_n664));
  OAI21_X1  g239(.A(new_n663), .B1(new_n659), .B2(new_n664), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n660), .A2(new_n661), .A3(new_n657), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n666), .B(KEYINPUT18), .Z(new_n667));
  NAND3_X1  g242(.A1(new_n664), .A2(new_n659), .A3(new_n657), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n665), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G2096), .B(G2100), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(G227));
  XOR2_X1   g247(.A(G1956), .B(G2474), .Z(new_n673));
  XOR2_X1   g248(.A(G1961), .B(G1966), .Z(new_n674));
  NOR2_X1   g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1971), .B(G1976), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT19), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n679), .B(KEYINPUT87), .Z(new_n680));
  NAND2_X1  g255(.A1(new_n673), .A2(new_n674), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(new_n682), .B(KEYINPUT20), .Z(new_n683));
  NAND3_X1  g258(.A1(new_n676), .A2(new_n678), .A3(new_n681), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n680), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(G1986), .ZN(new_n686));
  XOR2_X1   g261(.A(G1991), .B(G1996), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XOR2_X1   g263(.A(KEYINPUT88), .B(G1981), .Z(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n688), .B(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(G229));
  INV_X1    g268(.A(G16), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n694), .B1(new_n586), .B2(new_n587), .ZN(new_n695));
  AND2_X1   g270(.A1(new_n694), .A2(G23), .ZN(new_n696));
  OAI21_X1  g271(.A(KEYINPUT33), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(new_n698));
  NOR3_X1   g273(.A1(new_n695), .A2(KEYINPUT33), .A3(new_n696), .ZN(new_n699));
  INV_X1    g274(.A(G1976), .ZN(new_n700));
  NOR3_X1   g275(.A1(new_n698), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  OR3_X1    g276(.A1(new_n695), .A2(KEYINPUT33), .A3(new_n696), .ZN(new_n702));
  AOI21_X1  g277(.A(G1976), .B1(new_n702), .B2(new_n697), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(KEYINPUT34), .ZN(new_n705));
  OR2_X1    g280(.A1(G16), .A2(G22), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(G303), .B2(new_n694), .ZN(new_n707));
  XNOR2_X1  g282(.A(KEYINPUT90), .B(G1971), .ZN(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  OAI211_X1 g285(.A(new_n706), .B(new_n708), .C1(G303), .C2(new_n694), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n694), .A2(G6), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(new_n596), .B2(new_n694), .ZN(new_n714));
  XOR2_X1   g289(.A(KEYINPUT32), .B(G1981), .Z(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  NAND4_X1  g291(.A1(new_n704), .A2(new_n705), .A3(new_n712), .A4(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n694), .A2(G24), .ZN(new_n718));
  INV_X1    g293(.A(G290), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n718), .B1(new_n719), .B2(new_n694), .ZN(new_n720));
  INV_X1    g295(.A(G1986), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n700), .B1(new_n698), .B2(new_n699), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n702), .A2(G1976), .A3(new_n697), .ZN(new_n724));
  NAND4_X1  g299(.A1(new_n723), .A2(new_n712), .A3(new_n724), .A4(new_n716), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n725), .A2(KEYINPUT34), .ZN(new_n726));
  INV_X1    g301(.A(G29), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n727), .A2(G25), .ZN(new_n728));
  AOI22_X1  g303(.A1(new_n475), .A2(G119), .B1(G131), .B2(new_n477), .ZN(new_n729));
  OR2_X1    g304(.A1(G95), .A2(G2105), .ZN(new_n730));
  OAI211_X1 g305(.A(new_n730), .B(G2104), .C1(G107), .C2(new_n470), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(KEYINPUT89), .ZN(new_n732));
  INV_X1    g307(.A(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n729), .A2(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(new_n734), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n728), .B1(new_n735), .B2(new_n727), .ZN(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT35), .B(G1991), .ZN(new_n737));
  INV_X1    g312(.A(new_n737), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n736), .B(new_n738), .ZN(new_n739));
  NAND4_X1  g314(.A1(new_n717), .A2(new_n722), .A3(new_n726), .A4(new_n739), .ZN(new_n740));
  XOR2_X1   g315(.A(KEYINPUT91), .B(KEYINPUT36), .Z(new_n741));
  AND2_X1   g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n727), .B1(new_n478), .B2(new_n482), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n727), .A2(G35), .ZN(new_n744));
  INV_X1    g319(.A(new_n744), .ZN(new_n745));
  OR3_X1    g320(.A1(new_n743), .A2(KEYINPUT29), .A3(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(G2090), .ZN(new_n747));
  OAI21_X1  g322(.A(KEYINPUT29), .B1(new_n743), .B2(new_n745), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n746), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n749), .A2(KEYINPUT96), .ZN(new_n750));
  INV_X1    g325(.A(KEYINPUT96), .ZN(new_n751));
  NAND4_X1  g326(.A1(new_n746), .A2(new_n751), .A3(new_n747), .A4(new_n748), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g328(.A1(G16), .A2(G21), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(G168), .B2(G16), .ZN(new_n755));
  INV_X1    g330(.A(G1966), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  NOR2_X1   g332(.A1(G27), .A2(G29), .ZN(new_n758));
  INV_X1    g333(.A(new_n758), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(new_n504), .B2(new_n727), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(G2078), .ZN(new_n761));
  INV_X1    g336(.A(G33), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n762), .A2(G29), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n470), .A2(G103), .A3(G2104), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(KEYINPUT25), .Z(new_n765));
  NAND4_X1  g340(.A1(new_n468), .A2(new_n469), .A3(G139), .A4(new_n470), .ZN(new_n766));
  AOI22_X1  g341(.A1(new_n492), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n767));
  OAI211_X1 g342(.A(new_n765), .B(new_n766), .C1(new_n470), .C2(new_n767), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n763), .B1(new_n768), .B2(G29), .ZN(new_n769));
  INV_X1    g344(.A(G2072), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(KEYINPUT93), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n694), .A2(G19), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(new_n564), .B2(new_n694), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n775), .A2(G1341), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n472), .A2(G29), .ZN(new_n777));
  OR2_X1    g352(.A1(KEYINPUT24), .A2(G34), .ZN(new_n778));
  NAND2_X1  g353(.A1(KEYINPUT24), .A2(G34), .ZN(new_n779));
  NAND3_X1  g354(.A1(new_n778), .A2(new_n727), .A3(new_n779), .ZN(new_n780));
  AND2_X1   g355(.A1(new_n777), .A2(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(G2084), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NOR3_X1   g358(.A1(new_n773), .A2(new_n776), .A3(new_n783), .ZN(new_n784));
  AND2_X1   g359(.A1(new_n781), .A2(new_n782), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n633), .A2(new_n727), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n769), .A2(new_n770), .ZN(new_n787));
  INV_X1    g362(.A(KEYINPUT30), .ZN(new_n788));
  OR2_X1    g363(.A1(new_n788), .A2(G28), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n788), .A2(G28), .ZN(new_n790));
  AND3_X1   g365(.A1(new_n789), .A2(new_n790), .A3(new_n727), .ZN(new_n791));
  NOR4_X1   g366(.A1(new_n785), .A2(new_n786), .A3(new_n787), .A4(new_n791), .ZN(new_n792));
  NAND4_X1  g367(.A1(new_n757), .A2(new_n761), .A3(new_n784), .A4(new_n792), .ZN(new_n793));
  XOR2_X1   g368(.A(KEYINPUT31), .B(G11), .Z(new_n794));
  NOR3_X1   g369(.A1(new_n753), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  XNOR2_X1  g370(.A(KEYINPUT98), .B(KEYINPUT23), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n694), .A2(G20), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(G299), .B2(G16), .ZN(new_n799));
  INV_X1    g374(.A(G1956), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n747), .B1(new_n746), .B2(new_n748), .ZN(new_n802));
  OR2_X1    g377(.A1(new_n802), .A2(KEYINPUT97), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n802), .A2(KEYINPUT97), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n801), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n775), .A2(G1341), .ZN(new_n806));
  INV_X1    g381(.A(KEYINPUT95), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(G5), .B2(G16), .ZN(new_n808));
  OR3_X1    g383(.A1(new_n807), .A2(G5), .A3(G16), .ZN(new_n809));
  OAI211_X1 g384(.A(new_n808), .B(new_n809), .C1(G301), .C2(new_n694), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(G1961), .ZN(new_n811));
  NAND4_X1  g386(.A1(new_n795), .A2(new_n805), .A3(new_n806), .A4(new_n811), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n740), .A2(new_n741), .ZN(new_n813));
  NOR3_X1   g388(.A1(new_n742), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n727), .A2(G32), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n477), .A2(G141), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT94), .ZN(new_n817));
  NAND3_X1  g392(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT26), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n819), .B1(new_n475), .B2(G129), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n464), .A2(G105), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n817), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(new_n822), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n815), .B1(new_n823), .B2(new_n727), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT27), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(G1996), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n727), .A2(G26), .ZN(new_n827));
  AOI22_X1  g402(.A1(new_n475), .A2(G128), .B1(G140), .B2(new_n477), .ZN(new_n828));
  OR2_X1    g403(.A1(G104), .A2(G2105), .ZN(new_n829));
  OAI211_X1 g404(.A(new_n829), .B(G2104), .C1(G116), .C2(new_n470), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(new_n831), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n827), .B1(new_n832), .B2(new_n727), .ZN(new_n833));
  MUX2_X1   g408(.A(new_n827), .B(new_n833), .S(KEYINPUT28), .Z(new_n834));
  XNOR2_X1  g409(.A(KEYINPUT92), .B(G2067), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n834), .B(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n694), .A2(G4), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n837), .B1(new_n616), .B2(new_n694), .ZN(new_n838));
  INV_X1    g413(.A(G1348), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n838), .B(new_n839), .ZN(new_n840));
  NAND4_X1  g415(.A1(new_n814), .A2(new_n826), .A3(new_n836), .A4(new_n840), .ZN(G150));
  NAND2_X1  g416(.A1(G150), .A2(KEYINPUT99), .ZN(new_n842));
  INV_X1    g417(.A(new_n840), .ZN(new_n843));
  NOR4_X1   g418(.A1(new_n742), .A2(new_n812), .A3(new_n813), .A4(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT99), .ZN(new_n845));
  NAND4_X1  g420(.A1(new_n844), .A2(new_n845), .A3(new_n826), .A4(new_n836), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n842), .A2(new_n846), .ZN(G311));
  NAND2_X1  g422(.A1(G80), .A2(G543), .ZN(new_n848));
  INV_X1    g423(.A(G67), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n848), .B1(new_n610), .B2(new_n849), .ZN(new_n850));
  AND2_X1   g425(.A1(new_n850), .A2(G651), .ZN(new_n851));
  INV_X1    g426(.A(G55), .ZN(new_n852));
  INV_X1    g427(.A(G93), .ZN(new_n853));
  OAI22_X1  g428(.A1(new_n507), .A2(new_n852), .B1(new_n517), .B2(new_n853), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n851), .A2(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(KEYINPUT100), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n857), .A2(G860), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n858), .B(KEYINPUT37), .Z(new_n859));
  NOR2_X1   g434(.A1(new_n615), .A2(new_n621), .ZN(new_n860));
  XOR2_X1   g435(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n861));
  XNOR2_X1  g436(.A(new_n860), .B(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n560), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n856), .A2(new_n863), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n564), .B1(new_n851), .B2(new_n854), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n862), .B(new_n866), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n859), .B1(new_n867), .B2(G860), .ZN(G145));
  INV_X1    g443(.A(G37), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n832), .A2(new_n822), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT101), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n768), .A2(new_n872), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n502), .A2(new_n499), .ZN(new_n874));
  XOR2_X1   g449(.A(new_n873), .B(new_n874), .Z(new_n875));
  NAND2_X1  g450(.A1(new_n832), .A2(new_n822), .ZN(new_n876));
  AND3_X1   g451(.A1(new_n871), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n875), .B1(new_n871), .B2(new_n876), .ZN(new_n878));
  OR2_X1    g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  AOI22_X1  g454(.A1(new_n475), .A2(G130), .B1(G142), .B2(new_n477), .ZN(new_n880));
  OR2_X1    g455(.A1(G106), .A2(G2105), .ZN(new_n881));
  OAI211_X1 g456(.A(new_n881), .B(G2104), .C1(G118), .C2(new_n470), .ZN(new_n882));
  AND2_X1   g457(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT102), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n883), .A2(new_n884), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n735), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n887), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n889), .A2(new_n734), .A3(new_n885), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n638), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n888), .A2(new_n890), .A3(new_n638), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n879), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n877), .A2(new_n878), .ZN(new_n895));
  INV_X1    g470(.A(new_n893), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n895), .B1(new_n896), .B2(new_n891), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n633), .B(G160), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n898), .B(G162), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n894), .A2(new_n897), .A3(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT103), .ZN(new_n902));
  AND3_X1   g477(.A1(new_n894), .A2(new_n897), .A3(new_n902), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n899), .B1(new_n897), .B2(new_n902), .ZN(new_n904));
  OAI211_X1 g479(.A(new_n869), .B(new_n901), .C1(new_n903), .C2(new_n904), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n905), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g481(.A(new_n866), .B(new_n623), .ZN(new_n907));
  NAND2_X1  g482(.A1(G299), .A2(KEYINPUT104), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT104), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n573), .A2(new_n576), .A3(new_n909), .A4(new_n578), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n908), .A2(new_n615), .A3(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n910), .B1(new_n908), .B2(new_n615), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n907), .A2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n913), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n916), .A2(KEYINPUT41), .A3(new_n911), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT41), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n918), .B1(new_n912), .B2(new_n913), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n915), .B1(new_n907), .B2(new_n920), .ZN(new_n921));
  OR2_X1    g496(.A1(KEYINPUT105), .A2(KEYINPUT42), .ZN(new_n922));
  OR2_X1    g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(KEYINPUT105), .A2(KEYINPUT42), .ZN(new_n924));
  XNOR2_X1  g499(.A(G303), .B(G288), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(new_n596), .ZN(new_n926));
  INV_X1    g501(.A(G288), .ZN(new_n927));
  NAND2_X1  g502(.A1(G166), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(G303), .A2(G288), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n928), .A2(G305), .A3(new_n929), .ZN(new_n930));
  AND3_X1   g505(.A1(new_n926), .A2(new_n719), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n719), .B1(new_n926), .B2(new_n930), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n924), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n921), .A2(new_n922), .ZN(new_n934));
  AND3_X1   g509(.A1(new_n923), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n933), .B1(new_n923), .B2(new_n934), .ZN(new_n936));
  OAI21_X1  g511(.A(G868), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n937), .B1(G868), .B2(new_n856), .ZN(G295));
  OAI21_X1  g513(.A(new_n937), .B1(G868), .B2(new_n856), .ZN(G331));
  INV_X1    g514(.A(KEYINPUT44), .ZN(new_n940));
  INV_X1    g515(.A(new_n932), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n926), .A2(new_n719), .A3(new_n930), .ZN(new_n942));
  AOI21_X1  g517(.A(KEYINPUT107), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT106), .ZN(new_n944));
  OAI211_X1 g519(.A(new_n944), .B(G171), .C1(new_n582), .C2(new_n583), .ZN(new_n945));
  AOI22_X1  g520(.A1(new_n544), .A2(new_n545), .B1(G51), .B2(new_n527), .ZN(new_n946));
  AOI21_X1  g521(.A(KEYINPUT75), .B1(new_n946), .B2(new_n529), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n539), .A2(new_n540), .ZN(new_n948));
  OAI21_X1  g523(.A(KEYINPUT78), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n541), .A2(new_n547), .A3(new_n581), .ZN(new_n950));
  AOI21_X1  g525(.A(G301), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n947), .A2(new_n948), .ZN(new_n952));
  OAI21_X1  g527(.A(KEYINPUT106), .B1(new_n952), .B2(G171), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n945), .B1(new_n951), .B2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(new_n866), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  OAI211_X1 g531(.A(new_n866), .B(new_n945), .C1(new_n951), .C2(new_n953), .ZN(new_n957));
  AND3_X1   g532(.A1(new_n956), .A2(new_n914), .A3(new_n957), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n920), .B1(new_n956), .B2(new_n957), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n943), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(new_n920), .ZN(new_n961));
  INV_X1    g536(.A(new_n957), .ZN(new_n962));
  OAI21_X1  g537(.A(G171), .B1(new_n582), .B2(new_n583), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n944), .B1(G168), .B2(G301), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n866), .B1(new_n965), .B2(new_n945), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n961), .B1(new_n962), .B2(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n956), .A2(new_n914), .A3(new_n957), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT107), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n969), .B1(new_n931), .B2(new_n932), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n967), .A2(new_n968), .A3(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n960), .A2(new_n869), .A3(new_n971), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n972), .A2(KEYINPUT108), .A3(KEYINPUT43), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n931), .A2(new_n932), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n974), .B1(new_n968), .B2(KEYINPUT109), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n967), .A2(new_n968), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT43), .ZN(new_n978));
  OAI211_X1 g553(.A(new_n967), .B(new_n968), .C1(KEYINPUT109), .C2(new_n974), .ZN(new_n979));
  NAND4_X1  g554(.A1(new_n977), .A2(new_n978), .A3(new_n869), .A4(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n973), .A2(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(KEYINPUT108), .B1(new_n972), .B2(KEYINPUT43), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n940), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT110), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n977), .A2(new_n869), .A3(new_n979), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(KEYINPUT43), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n960), .A2(new_n978), .A3(new_n971), .A4(new_n869), .ZN(new_n987));
  AND4_X1   g562(.A1(new_n984), .A2(new_n986), .A3(KEYINPUT44), .A4(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n940), .B1(new_n985), .B2(KEYINPUT43), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n984), .B1(new_n989), .B2(new_n987), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n983), .B1(new_n988), .B2(new_n990), .ZN(G397));
  NAND2_X1  g566(.A1(G303), .A2(G8), .ZN(new_n992));
  NAND2_X1  g567(.A1(KEYINPUT115), .A2(KEYINPUT55), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  XOR2_X1   g569(.A(KEYINPUT115), .B(KEYINPUT55), .Z(new_n995));
  OAI21_X1  g570(.A(new_n994), .B1(new_n992), .B2(new_n995), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n460), .A2(new_n465), .A3(G40), .A4(new_n471), .ZN(new_n997));
  INV_X1    g572(.A(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(G1384), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n999), .B1(new_n502), .B2(new_n499), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT45), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n998), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n501), .A2(new_n503), .A3(new_n999), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n1002), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n997), .B1(new_n1000), .B2(KEYINPUT50), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1005), .B1(new_n1003), .B2(KEYINPUT50), .ZN(new_n1006));
  OAI22_X1  g581(.A1(new_n1004), .A2(G1971), .B1(new_n1006), .B2(G2090), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n996), .B1(new_n1007), .B2(G8), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT119), .ZN(new_n1009));
  OR2_X1    g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(G8), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1003), .A2(new_n1001), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1002), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(G1971), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n997), .B1(new_n1003), .B2(KEYINPUT50), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT50), .ZN(new_n1018));
  OAI211_X1 g593(.A(new_n1018), .B(new_n999), .C1(new_n502), .C2(new_n499), .ZN(new_n1019));
  XNOR2_X1  g594(.A(new_n1019), .B(KEYINPUT114), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1017), .A2(new_n1020), .A3(new_n747), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1011), .B1(new_n1016), .B2(new_n1021), .ZN(new_n1022));
  AOI22_X1  g597(.A1(new_n1008), .A2(new_n1009), .B1(new_n1022), .B2(new_n996), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n522), .A2(new_n506), .A3(G86), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1024), .A2(new_n594), .A3(KEYINPUT116), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1025), .ZN(new_n1026));
  AOI21_X1  g601(.A(KEYINPUT116), .B1(new_n1024), .B2(new_n594), .ZN(new_n1027));
  OR3_X1    g602(.A1(new_n1026), .A2(new_n593), .A3(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT117), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1028), .A2(new_n1029), .A3(G1981), .ZN(new_n1030));
  INV_X1    g605(.A(G1981), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n596), .A2(new_n1031), .ZN(new_n1032));
  NOR3_X1   g607(.A1(new_n1026), .A2(new_n1027), .A3(new_n593), .ZN(new_n1033));
  OAI21_X1  g608(.A(KEYINPUT117), .B1(new_n1033), .B2(new_n1031), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1030), .A2(new_n1032), .A3(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT49), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1000), .A2(new_n997), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1038), .A2(new_n1011), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n1030), .A2(new_n1032), .A3(new_n1034), .A4(KEYINPUT49), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1037), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT118), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n1037), .A2(KEYINPUT118), .A3(new_n1039), .A4(new_n1040), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1039), .B1(new_n700), .B2(G288), .ZN(new_n1045));
  AOI22_X1  g620(.A1(new_n1043), .A2(new_n1044), .B1(KEYINPUT52), .B2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(KEYINPUT52), .B1(G288), .B2(new_n700), .ZN(new_n1047));
  OAI211_X1 g622(.A(new_n1039), .B(new_n1047), .C1(new_n700), .C2(G288), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1010), .A2(new_n1023), .A3(new_n1046), .A4(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT53), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1050), .B1(new_n1014), .B2(G2078), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n997), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1052), .B1(new_n1003), .B2(new_n1001), .ZN(new_n1053));
  OR2_X1    g628(.A1(new_n1050), .A2(G2078), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1017), .A2(new_n1020), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(KEYINPUT123), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT123), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1017), .A2(new_n1020), .A3(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1059));
  OAI221_X1 g634(.A(new_n1051), .B1(new_n1053), .B2(new_n1054), .C1(new_n1059), .C2(G1961), .ZN(new_n1060));
  XOR2_X1   g635(.A(G171), .B(KEYINPUT54), .Z(new_n1061));
  AOI21_X1  g636(.A(new_n1049), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1053), .A2(new_n756), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT120), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1017), .A2(new_n1020), .A3(new_n782), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1053), .A2(KEYINPUT120), .A3(new_n756), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1065), .A2(new_n1066), .A3(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(G8), .ZN(new_n1069));
  NOR2_X1   g644(.A1(G168), .A2(new_n1011), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(KEYINPUT125), .ZN(new_n1071));
  NAND2_X1  g646(.A1(KEYINPUT125), .A2(KEYINPUT51), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1072), .B1(G168), .B2(new_n1011), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1069), .A2(new_n1071), .A3(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT51), .ZN(new_n1075));
  OAI211_X1 g650(.A(new_n1075), .B(G8), .C1(new_n1068), .C2(new_n952), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1068), .A2(new_n1070), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1074), .A2(new_n1076), .A3(new_n1077), .ZN(new_n1078));
  XNOR2_X1  g653(.A(new_n1000), .B(new_n1001), .ZN(new_n1079));
  XNOR2_X1  g654(.A(new_n459), .B(KEYINPUT127), .ZN(new_n1080));
  OAI21_X1  g655(.A(G40), .B1(new_n1080), .B2(new_n470), .ZN(new_n1081));
  NOR3_X1   g656(.A1(new_n1079), .A2(new_n1054), .A3(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n465), .A2(new_n471), .ZN(new_n1083));
  XOR2_X1   g658(.A(new_n1083), .B(KEYINPUT126), .Z(new_n1084));
  AOI21_X1  g659(.A(new_n1061), .B1(new_n1082), .B2(new_n1084), .ZN(new_n1085));
  OAI211_X1 g660(.A(new_n1051), .B(new_n1085), .C1(new_n1059), .C2(G1961), .ZN(new_n1086));
  AND2_X1   g661(.A1(new_n1078), .A2(new_n1086), .ZN(new_n1087));
  XOR2_X1   g662(.A(KEYINPUT58), .B(G1341), .Z(new_n1088));
  INV_X1    g663(.A(new_n1088), .ZN(new_n1089));
  OAI22_X1  g664(.A1(new_n1014), .A2(G1996), .B1(new_n1038), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(new_n564), .ZN(new_n1091));
  XNOR2_X1  g666(.A(new_n1091), .B(KEYINPUT59), .ZN(new_n1092));
  XNOR2_X1  g667(.A(G299), .B(KEYINPUT57), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1006), .A2(new_n800), .ZN(new_n1095));
  XNOR2_X1  g670(.A(KEYINPUT56), .B(G2072), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1012), .A2(new_n1013), .A3(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1094), .A2(new_n1095), .A3(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT122), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1095), .A2(new_n1097), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(new_n1093), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1094), .A2(new_n1095), .A3(KEYINPUT122), .A4(new_n1097), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1100), .A2(new_n1102), .A3(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT61), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1102), .A2(KEYINPUT61), .A3(new_n1098), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1092), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1056), .A2(new_n839), .A3(new_n1058), .ZN(new_n1109));
  INV_X1    g684(.A(G2067), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1038), .A2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(KEYINPUT60), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1109), .A2(KEYINPUT60), .A3(new_n1111), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(new_n616), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1109), .A2(KEYINPUT60), .A3(new_n615), .A4(new_n1111), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1112), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1108), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1100), .A2(new_n1103), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n615), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT124), .ZN(new_n1120));
  OR2_X1    g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  AOI22_X1  g696(.A1(new_n1119), .A2(new_n1120), .B1(new_n1093), .B2(new_n1101), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1118), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  OAI211_X1 g698(.A(new_n1062), .B(new_n1087), .C1(new_n1117), .C2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1125));
  NOR2_X1   g700(.A1(G288), .A2(G1976), .ZN(new_n1126));
  AOI22_X1  g701(.A1(new_n1125), .A2(new_n1126), .B1(new_n1031), .B2(new_n596), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1039), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1022), .A2(new_n996), .ZN(new_n1130));
  OAI22_X1  g705(.A1(new_n1127), .A2(new_n1128), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT63), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1068), .A2(G8), .A3(new_n584), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT121), .ZN(new_n1134));
  XNOR2_X1  g709(.A(new_n1133), .B(new_n1134), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1132), .B1(new_n1135), .B2(new_n1049), .ZN(new_n1136));
  XNOR2_X1  g711(.A(new_n1133), .B(KEYINPUT121), .ZN(new_n1137));
  OR2_X1    g712(.A1(new_n1022), .A2(new_n996), .ZN(new_n1138));
  AND4_X1   g713(.A1(new_n1046), .A2(new_n1138), .A3(new_n1048), .A4(new_n1130), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1137), .A2(new_n1139), .A3(KEYINPUT63), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1131), .B1(new_n1136), .B2(new_n1140), .ZN(new_n1141));
  OR2_X1    g716(.A1(new_n1078), .A2(KEYINPUT62), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1060), .A2(G171), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1049), .A2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1078), .A2(KEYINPUT62), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1142), .A2(new_n1144), .A3(new_n1145), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1124), .A2(new_n1141), .A3(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1000), .ZN(new_n1148));
  NOR3_X1   g723(.A1(new_n1148), .A2(KEYINPUT45), .A3(new_n997), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1149), .ZN(new_n1150));
  XNOR2_X1  g725(.A(new_n831), .B(new_n1110), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n822), .A2(G1996), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1150), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  OR2_X1    g728(.A1(new_n1150), .A2(G1996), .ZN(new_n1154));
  OR2_X1    g729(.A1(new_n1154), .A2(KEYINPUT112), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1154), .A2(KEYINPUT112), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1153), .B1(new_n1157), .B2(new_n823), .ZN(new_n1158));
  OR2_X1    g733(.A1(new_n1158), .A2(KEYINPUT113), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1158), .A2(KEYINPUT113), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n735), .A2(new_n738), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n734), .A2(new_n737), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1149), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  NOR3_X1   g738(.A1(new_n1150), .A2(G1986), .A3(G290), .ZN(new_n1164));
  NOR3_X1   g739(.A1(new_n1150), .A2(new_n721), .A3(new_n719), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  XOR2_X1   g741(.A(new_n1166), .B(KEYINPUT111), .Z(new_n1167));
  AND4_X1   g742(.A1(new_n1159), .A2(new_n1160), .A3(new_n1163), .A4(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1147), .A2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1159), .A2(new_n1160), .A3(new_n1162), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n832), .A2(new_n1110), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1150), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1150), .B1(new_n1151), .B2(new_n823), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT46), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1157), .A2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1155), .A2(KEYINPUT46), .A3(new_n1156), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1173), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  XNOR2_X1  g752(.A(new_n1177), .B(KEYINPUT47), .ZN(new_n1178));
  XOR2_X1   g753(.A(new_n1164), .B(KEYINPUT48), .Z(new_n1179));
  AND4_X1   g754(.A1(new_n1159), .A2(new_n1160), .A3(new_n1163), .A4(new_n1179), .ZN(new_n1180));
  NOR3_X1   g755(.A1(new_n1172), .A2(new_n1178), .A3(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1169), .A2(new_n1181), .ZN(G329));
  assign    G231 = 1'b0;
  OAI211_X1 g757(.A(new_n655), .B(new_n692), .C1(new_n981), .C2(new_n982), .ZN(new_n1184));
  NAND3_X1  g758(.A1(new_n905), .A2(G319), .A3(new_n671), .ZN(new_n1185));
  NOR2_X1   g759(.A1(new_n1184), .A2(new_n1185), .ZN(G308));
  INV_X1    g760(.A(new_n1185), .ZN(new_n1187));
  INV_X1    g761(.A(new_n982), .ZN(new_n1188));
  NAND3_X1  g762(.A1(new_n1188), .A2(new_n980), .A3(new_n973), .ZN(new_n1189));
  NAND4_X1  g763(.A1(new_n1187), .A2(new_n1189), .A3(new_n655), .A4(new_n692), .ZN(G225));
endmodule


