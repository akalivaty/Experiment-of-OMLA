//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 1 1 0 1 1 0 0 0 1 1 1 1 0 1 1 0 1 1 0 0 1 0 1 1 0 1 0 1 1 1 1 0 0 1 0 0 0 0 1 0 1 0 1 0 1 1 1 0 1 1 1 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:49 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1258, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n216), .A2(new_n210), .ZN(new_n217));
  XNOR2_X1  g0017(.A(new_n217), .B(KEYINPUT65), .ZN(new_n218));
  OAI21_X1  g0018(.A(G50), .B1(G58), .B2(G68), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n221));
  INV_X1    g0021(.A(KEYINPUT66), .ZN(new_n222));
  AND2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n221), .A2(new_n222), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n220), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  OR2_X1    g0025(.A1(new_n225), .A2(KEYINPUT67), .ZN(new_n226));
  INV_X1    g0026(.A(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n225), .A2(KEYINPUT67), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n229));
  AOI22_X1  g0029(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n230));
  NAND3_X1  g0030(.A1(new_n228), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n212), .B1(new_n227), .B2(new_n231), .ZN(new_n232));
  OAI221_X1 g0032(.A(new_n215), .B1(new_n218), .B2(new_n219), .C1(new_n232), .C2(KEYINPUT1), .ZN(new_n233));
  AOI21_X1  g0033(.A(new_n233), .B1(KEYINPUT1), .B2(new_n232), .ZN(G361));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT68), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(KEYINPUT2), .B(G226), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n238), .B(new_n242), .ZN(G358));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT70), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G68), .B(G77), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(KEYINPUT69), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G50), .B(G58), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(new_n247), .B(new_n251), .Z(G351));
  NAND3_X1  g0052(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(new_n216), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  XOR2_X1   g0055(.A(KEYINPUT8), .B(G58), .Z(new_n256));
  NAND2_X1  g0056(.A1(new_n210), .A2(G33), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  NOR2_X1   g0058(.A1(G20), .A2(G33), .ZN(new_n259));
  AOI22_X1  g0059(.A1(new_n256), .A2(new_n258), .B1(G150), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n203), .A2(G20), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n255), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n209), .A2(G13), .A3(G20), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G50), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n255), .B1(G1), .B2(new_n210), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n266), .B1(new_n267), .B2(new_n265), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n262), .A2(new_n268), .ZN(new_n269));
  XOR2_X1   g0069(.A(new_n269), .B(KEYINPUT9), .Z(new_n270));
  XNOR2_X1  g0070(.A(KEYINPUT3), .B(G33), .ZN(new_n271));
  INV_X1    g0071(.A(G1698), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n271), .A2(G222), .A3(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G77), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n271), .A2(G1698), .ZN(new_n275));
  INV_X1    g0075(.A(G223), .ZN(new_n276));
  OAI221_X1 g0076(.A(new_n273), .B1(new_n274), .B2(new_n271), .C1(new_n275), .C2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(G33), .A2(G41), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n278), .A2(G1), .A3(G13), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n277), .A2(new_n280), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n282));
  INV_X1    g0082(.A(G274), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n279), .A2(new_n282), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT72), .ZN(new_n287));
  XNOR2_X1  g0087(.A(new_n286), .B(new_n287), .ZN(new_n288));
  XOR2_X1   g0088(.A(KEYINPUT71), .B(G226), .Z(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n281), .A2(new_n285), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G200), .ZN(new_n292));
  INV_X1    g0092(.A(new_n291), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(G190), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n270), .A2(new_n292), .A3(new_n294), .ZN(new_n295));
  XNOR2_X1  g0095(.A(new_n295), .B(KEYINPUT10), .ZN(new_n296));
  INV_X1    g0096(.A(G179), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n293), .A2(new_n297), .ZN(new_n298));
  XNOR2_X1  g0098(.A(new_n298), .B(KEYINPUT73), .ZN(new_n299));
  INV_X1    g0099(.A(G169), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n269), .B1(new_n291), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n296), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G68), .ZN(new_n304));
  AOI22_X1  g0104(.A1(new_n258), .A2(G77), .B1(G20), .B2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(G33), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n210), .A2(new_n306), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n305), .B1(new_n265), .B2(new_n307), .ZN(new_n308));
  AND3_X1   g0108(.A1(new_n308), .A2(KEYINPUT11), .A3(new_n254), .ZN(new_n309));
  AOI21_X1  g0109(.A(KEYINPUT11), .B1(new_n308), .B2(new_n254), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT12), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n311), .B1(new_n264), .B2(new_n304), .ZN(new_n312));
  NOR3_X1   g0112(.A1(new_n263), .A2(KEYINPUT12), .A3(G68), .ZN(new_n313));
  OAI22_X1  g0113(.A1(new_n267), .A2(new_n304), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NOR3_X1   g0114(.A1(new_n309), .A2(new_n310), .A3(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  AND2_X1   g0116(.A1(KEYINPUT3), .A2(G33), .ZN(new_n317));
  NOR2_X1   g0117(.A1(KEYINPUT3), .A2(G33), .ZN(new_n318));
  OAI211_X1 g0118(.A(G232), .B(G1698), .C1(new_n317), .C2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT75), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND4_X1  g0121(.A1(new_n271), .A2(KEYINPUT75), .A3(G232), .A4(G1698), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  OAI211_X1 g0123(.A(G226), .B(new_n272), .C1(new_n317), .C2(new_n318), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT74), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND4_X1  g0126(.A1(new_n271), .A2(KEYINPUT74), .A3(G226), .A4(new_n272), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(G33), .A2(G97), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(KEYINPUT76), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT76), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n331), .A2(G33), .A3(G97), .ZN(new_n332));
  AND2_X1   g0132(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n323), .A2(new_n328), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(new_n280), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT13), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n284), .B1(new_n288), .B2(G238), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n335), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n330), .A2(new_n332), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n339), .B1(new_n326), .B2(new_n327), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n279), .B1(new_n340), .B2(new_n323), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n286), .A2(new_n287), .ZN(new_n342));
  AOI21_X1  g0142(.A(KEYINPUT72), .B1(new_n279), .B2(new_n282), .ZN(new_n343));
  OAI21_X1  g0143(.A(G238), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(new_n285), .ZN(new_n345));
  OAI21_X1  g0145(.A(KEYINPUT13), .B1(new_n341), .B2(new_n345), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n338), .A2(new_n346), .A3(G179), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n300), .B1(new_n338), .B2(new_n346), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT14), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n347), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  AOI211_X1 g0150(.A(KEYINPUT14), .B(new_n300), .C1(new_n338), .C2(new_n346), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n316), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n338), .A2(new_n346), .A3(G190), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(new_n315), .ZN(new_n355));
  INV_X1    g0155(.A(G200), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n356), .B1(new_n338), .B2(new_n346), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n264), .A2(new_n274), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n359), .B1(new_n267), .B2(new_n274), .ZN(new_n360));
  XNOR2_X1  g0160(.A(KEYINPUT15), .B(G87), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  AOI22_X1  g0162(.A1(new_n362), .A2(new_n258), .B1(G20), .B2(G77), .ZN(new_n363));
  INV_X1    g0163(.A(new_n256), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n363), .B1(new_n364), .B2(new_n307), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n360), .B1(new_n254), .B2(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n284), .B1(new_n288), .B2(G244), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n271), .A2(G232), .A3(new_n272), .ZN(new_n368));
  INV_X1    g0168(.A(G238), .ZN(new_n369));
  OAI221_X1 g0169(.A(new_n368), .B1(new_n206), .B2(new_n271), .C1(new_n275), .C2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(new_n280), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n367), .A2(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n366), .B1(new_n372), .B2(new_n300), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n367), .A2(new_n371), .A3(new_n297), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n356), .B1(new_n367), .B2(new_n371), .ZN(new_n376));
  INV_X1    g0176(.A(G190), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n366), .B1(new_n372), .B2(new_n377), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n375), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  NOR4_X1   g0179(.A1(new_n303), .A2(new_n353), .A3(new_n358), .A4(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(G159), .ZN(new_n381));
  OAI21_X1  g0181(.A(KEYINPUT78), .B1(new_n307), .B2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT78), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n259), .A2(new_n383), .A3(G159), .ZN(new_n384));
  XNOR2_X1  g0184(.A(G58), .B(G68), .ZN(new_n385));
  AOI22_X1  g0185(.A1(new_n382), .A2(new_n384), .B1(new_n385), .B2(G20), .ZN(new_n386));
  NOR3_X1   g0186(.A1(new_n317), .A2(new_n318), .A3(G20), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT7), .ZN(new_n388));
  OAI21_X1  g0188(.A(G68), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  OR2_X1    g0189(.A1(KEYINPUT3), .A2(G33), .ZN(new_n390));
  NAND2_X1  g0190(.A1(KEYINPUT3), .A2(G33), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n390), .A2(new_n210), .A3(new_n391), .ZN(new_n392));
  XNOR2_X1  g0192(.A(KEYINPUT77), .B(KEYINPUT7), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  OAI211_X1 g0194(.A(KEYINPUT16), .B(new_n386), .C1(new_n389), .C2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(new_n254), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n390), .A2(new_n388), .A3(new_n210), .A4(new_n391), .ZN(new_n397));
  XOR2_X1   g0197(.A(KEYINPUT77), .B(KEYINPUT7), .Z(new_n398));
  OAI211_X1 g0198(.A(G68), .B(new_n397), .C1(new_n387), .C2(new_n398), .ZN(new_n399));
  AOI21_X1  g0199(.A(KEYINPUT16), .B1(new_n399), .B2(new_n386), .ZN(new_n400));
  OAI21_X1  g0200(.A(KEYINPUT79), .B1(new_n396), .B2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(new_n400), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT79), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n402), .A2(new_n403), .A3(new_n254), .A4(new_n395), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n401), .A2(new_n404), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n256), .A2(new_n264), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n406), .B1(new_n267), .B2(new_n256), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n276), .A2(new_n272), .ZN(new_n409));
  OAI211_X1 g0209(.A(new_n271), .B(new_n409), .C1(G226), .C2(new_n272), .ZN(new_n410));
  NAND2_X1  g0210(.A1(G33), .A2(G87), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(new_n280), .ZN(new_n413));
  INV_X1    g0213(.A(G232), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n285), .B1(new_n286), .B2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n413), .A2(G190), .A3(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n279), .B1(new_n410), .B2(new_n411), .ZN(new_n418));
  OAI21_X1  g0218(.A(G200), .B1(new_n418), .B2(new_n415), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n405), .A2(new_n408), .A3(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT17), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n407), .B1(new_n401), .B2(new_n404), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n425), .A2(KEYINPUT17), .A3(new_n421), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT81), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT18), .ZN(new_n429));
  NOR3_X1   g0229(.A1(new_n418), .A2(new_n297), .A3(new_n415), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n413), .A2(new_n416), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n430), .B1(G169), .B2(new_n431), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n429), .B1(new_n425), .B2(new_n432), .ZN(new_n433));
  NOR3_X1   g0233(.A1(new_n425), .A2(new_n429), .A3(new_n432), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n433), .B1(new_n434), .B2(KEYINPUT80), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT80), .ZN(new_n436));
  NOR4_X1   g0236(.A1(new_n425), .A2(new_n436), .A3(new_n429), .A4(new_n432), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n428), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  AND2_X1   g0238(.A1(G58), .A2(G68), .ZN(new_n439));
  OAI21_X1  g0239(.A(G20), .B1(new_n439), .B2(new_n202), .ZN(new_n440));
  NOR4_X1   g0240(.A1(new_n381), .A2(KEYINPUT78), .A3(G20), .A4(G33), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n383), .B1(new_n259), .B2(G159), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n440), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n387), .A2(new_n398), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n304), .B1(new_n392), .B2(KEYINPUT7), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n443), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n255), .B1(new_n446), .B2(KEYINPUT16), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n403), .B1(new_n447), .B2(new_n402), .ZN(new_n448));
  NOR3_X1   g0248(.A1(new_n396), .A2(KEYINPUT79), .A3(new_n400), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n408), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(new_n432), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n450), .A2(KEYINPUT18), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(new_n436), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n434), .A2(KEYINPUT80), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n453), .A2(new_n454), .A3(KEYINPUT81), .A4(new_n433), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n427), .B1(new_n438), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n380), .A2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n271), .A2(G250), .A3(new_n272), .ZN(new_n459));
  OAI211_X1 g0259(.A(G257), .B(G1698), .C1(new_n317), .C2(new_n318), .ZN(new_n460));
  NAND2_X1  g0260(.A1(G33), .A2(G294), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n459), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(new_n280), .ZN(new_n463));
  XNOR2_X1  g0263(.A(KEYINPUT5), .B(G41), .ZN(new_n464));
  INV_X1    g0264(.A(G45), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n465), .A2(G1), .ZN(new_n466));
  INV_X1    g0266(.A(new_n216), .ZN(new_n467));
  AOI22_X1  g0267(.A1(new_n464), .A2(new_n466), .B1(new_n467), .B2(new_n278), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(G264), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n209), .A2(G45), .ZN(new_n470));
  NOR2_X1   g0270(.A1(KEYINPUT5), .A2(G41), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(KEYINPUT5), .A2(G41), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n470), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n283), .B1(new_n467), .B2(new_n278), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  AND4_X1   g0276(.A1(G190), .A2(new_n463), .A3(new_n469), .A4(new_n476), .ZN(new_n477));
  AOI22_X1  g0277(.A1(new_n462), .A2(new_n280), .B1(G264), .B2(new_n468), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n356), .B1(new_n478), .B2(new_n476), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n264), .A2(KEYINPUT25), .A3(new_n206), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  AOI21_X1  g0282(.A(KEYINPUT25), .B1(new_n264), .B2(new_n206), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n209), .A2(G33), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n263), .A2(new_n484), .A3(new_n216), .A4(new_n253), .ZN(new_n485));
  OAI22_X1  g0285(.A1(new_n482), .A2(new_n483), .B1(new_n206), .B2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(G20), .B1(new_n390), .B2(new_n391), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n488), .A2(KEYINPUT86), .A3(KEYINPUT22), .A4(G87), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n210), .B(G87), .C1(new_n317), .C2(new_n318), .ZN(new_n490));
  OR2_X1    g0290(.A1(KEYINPUT86), .A2(KEYINPUT22), .ZN(new_n491));
  NAND2_X1  g0291(.A1(KEYINPUT86), .A2(KEYINPUT22), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n490), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(G33), .A2(G116), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n494), .A2(G20), .ZN(new_n495));
  AOI21_X1  g0295(.A(KEYINPUT23), .B1(new_n206), .B2(G20), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n206), .A2(KEYINPUT23), .A3(G20), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n495), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n489), .A2(new_n493), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(KEYINPUT24), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT24), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n489), .A2(new_n493), .A3(new_n502), .A4(new_n499), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  AOI21_X1  g0304(.A(KEYINPUT87), .B1(new_n504), .B2(new_n254), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT87), .ZN(new_n506));
  AOI211_X1 g0306(.A(new_n506), .B(new_n255), .C1(new_n501), .C2(new_n503), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n480), .B(new_n487), .C1(new_n505), .C2(new_n507), .ZN(new_n508));
  AND3_X1   g0308(.A1(new_n206), .A2(KEYINPUT23), .A3(G20), .ZN(new_n509));
  OAI22_X1  g0309(.A1(new_n509), .A2(new_n496), .B1(G20), .B2(new_n494), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n490), .A2(new_n491), .ZN(new_n511));
  INV_X1    g0311(.A(new_n492), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n502), .B1(new_n513), .B2(new_n493), .ZN(new_n514));
  INV_X1    g0314(.A(new_n503), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n254), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(new_n506), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n504), .A2(KEYINPUT87), .A3(new_n254), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n486), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n478), .A2(new_n476), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n300), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n521), .B1(G179), .B2(new_n520), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n508), .B1(new_n519), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(KEYINPUT88), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n487), .B1(new_n505), .B2(new_n507), .ZN(new_n525));
  INV_X1    g0325(.A(new_n522), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT88), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n527), .A2(new_n528), .A3(new_n508), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n524), .A2(new_n529), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n362), .A2(new_n263), .ZN(new_n531));
  INV_X1    g0331(.A(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(new_n485), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(new_n362), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n271), .A2(new_n210), .A3(G68), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT19), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n536), .B1(new_n257), .B2(new_n205), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n210), .B1(new_n333), .B2(new_n536), .ZN(new_n539));
  INV_X1    g0339(.A(G87), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n540), .A2(new_n205), .A3(new_n206), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n538), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n532), .B(new_n534), .C1(new_n542), .C2(new_n255), .ZN(new_n543));
  OAI211_X1 g0343(.A(G238), .B(new_n272), .C1(new_n317), .C2(new_n318), .ZN(new_n544));
  OAI211_X1 g0344(.A(G244), .B(G1698), .C1(new_n317), .C2(new_n318), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n544), .A2(new_n545), .A3(new_n494), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(new_n280), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT83), .ZN(new_n548));
  INV_X1    g0348(.A(G250), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n549), .B1(new_n209), .B2(G45), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n279), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n466), .A2(G274), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n548), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n551), .A2(new_n548), .A3(new_n552), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n547), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(new_n300), .ZN(new_n557));
  INV_X1    g0357(.A(new_n555), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n558), .A2(new_n553), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n559), .A2(new_n297), .A3(new_n547), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n543), .A2(new_n557), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n556), .A2(G200), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n536), .B1(new_n330), .B2(new_n332), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n541), .B1(new_n563), .B2(G20), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n564), .A2(new_n535), .A3(new_n537), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n531), .B1(new_n565), .B2(new_n254), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n547), .A2(new_n554), .A3(G190), .A4(new_n555), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n533), .A2(G87), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n562), .A2(new_n566), .A3(new_n567), .A4(new_n568), .ZN(new_n569));
  AND2_X1   g0369(.A1(new_n561), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n264), .A2(new_n205), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n571), .B1(new_n485), .B2(new_n205), .ZN(new_n572));
  INV_X1    g0372(.A(new_n572), .ZN(new_n573));
  OAI211_X1 g0373(.A(G107), .B(new_n397), .C1(new_n387), .C2(new_n398), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n259), .A2(G77), .ZN(new_n575));
  NAND2_X1  g0375(.A1(G97), .A2(G107), .ZN(new_n576));
  AOI21_X1  g0376(.A(KEYINPUT6), .B1(new_n207), .B2(new_n576), .ZN(new_n577));
  AND3_X1   g0377(.A1(new_n206), .A2(KEYINPUT6), .A3(G97), .ZN(new_n578));
  OAI21_X1  g0378(.A(G20), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n574), .A2(new_n575), .A3(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT82), .ZN(new_n581));
  AND3_X1   g0381(.A1(new_n580), .A2(new_n581), .A3(new_n254), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n581), .B1(new_n580), .B2(new_n254), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n573), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(new_n473), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n466), .B1(new_n585), .B2(new_n471), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n586), .A2(G257), .A3(new_n279), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n476), .A2(new_n587), .ZN(new_n588));
  OAI211_X1 g0388(.A(G244), .B(new_n272), .C1(new_n317), .C2(new_n318), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT4), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n271), .A2(KEYINPUT4), .A3(G244), .A4(new_n272), .ZN(new_n592));
  NAND2_X1  g0392(.A1(G33), .A2(G283), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n271), .A2(G250), .A3(G1698), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n591), .A2(new_n592), .A3(new_n593), .A4(new_n594), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n588), .B1(new_n595), .B2(new_n280), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n300), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n596), .A2(new_n297), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n584), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n580), .A2(new_n254), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(KEYINPUT82), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n580), .A2(new_n581), .A3(new_n254), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n597), .A2(G200), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n596), .A2(G190), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n604), .A2(new_n605), .A3(new_n573), .A4(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n570), .A2(new_n600), .A3(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT85), .ZN(new_n609));
  OAI211_X1 g0409(.A(G264), .B(G1698), .C1(new_n317), .C2(new_n318), .ZN(new_n610));
  OAI211_X1 g0410(.A(G257), .B(new_n272), .C1(new_n317), .C2(new_n318), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n390), .A2(G303), .A3(new_n391), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n610), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  AND2_X1   g0413(.A1(new_n613), .A2(new_n280), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n586), .A2(new_n279), .ZN(new_n615));
  INV_X1    g0415(.A(G270), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n476), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  OAI21_X1  g0417(.A(KEYINPUT84), .B1(new_n614), .B2(new_n617), .ZN(new_n618));
  AOI22_X1  g0418(.A1(new_n468), .A2(G270), .B1(new_n474), .B2(new_n475), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n613), .A2(new_n280), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT84), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n619), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n593), .B(new_n210), .C1(G33), .C2(new_n205), .ZN(new_n623));
  INV_X1    g0423(.A(G116), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(G20), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n623), .A2(new_n254), .A3(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT20), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n623), .A2(KEYINPUT20), .A3(new_n254), .A4(new_n625), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n263), .A2(G116), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n631), .B1(new_n533), .B2(G116), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n300), .B1(new_n630), .B2(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n618), .A2(new_n622), .A3(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT21), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n618), .A2(KEYINPUT21), .A3(new_n622), .A4(new_n633), .ZN(new_n637));
  AND3_X1   g0437(.A1(new_n619), .A2(G179), .A3(new_n620), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n630), .A2(new_n632), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n636), .A2(new_n637), .A3(new_n640), .ZN(new_n641));
  AND3_X1   g0441(.A1(new_n619), .A2(new_n621), .A3(new_n620), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n621), .B1(new_n619), .B2(new_n620), .ZN(new_n643));
  OAI21_X1  g0443(.A(G190), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n639), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n618), .A2(G200), .A3(new_n622), .ZN(new_n646));
  AND3_X1   g0446(.A1(new_n644), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n609), .B1(new_n641), .B2(new_n647), .ZN(new_n648));
  AOI22_X1  g0448(.A1(new_n634), .A2(new_n635), .B1(new_n639), .B2(new_n638), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n644), .A2(new_n646), .A3(new_n645), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n649), .A2(new_n650), .A3(KEYINPUT85), .A4(new_n637), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n608), .B1(new_n648), .B2(new_n651), .ZN(new_n652));
  AND3_X1   g0452(.A1(new_n458), .A2(new_n530), .A3(new_n652), .ZN(G372));
  NAND2_X1  g0453(.A1(new_n452), .A2(new_n433), .ZN(new_n654));
  INV_X1    g0454(.A(new_n375), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n353), .A2(new_n655), .ZN(new_n656));
  AND4_X1   g0456(.A1(KEYINPUT17), .A2(new_n405), .A3(new_n408), .A4(new_n421), .ZN(new_n657));
  AOI21_X1  g0457(.A(KEYINPUT17), .B1(new_n425), .B2(new_n421), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n358), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n654), .B1(new_n656), .B2(new_n661), .ZN(new_n662));
  AOI22_X1  g0462(.A1(new_n662), .A2(new_n296), .B1(new_n299), .B2(new_n301), .ZN(new_n663));
  INV_X1    g0463(.A(new_n600), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(new_n570), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT89), .ZN(new_n666));
  AND3_X1   g0466(.A1(new_n546), .A2(new_n666), .A3(new_n280), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n666), .B1(new_n546), .B2(new_n280), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n559), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(new_n300), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n670), .A2(new_n560), .A3(new_n543), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n669), .A2(G200), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n672), .A2(new_n566), .A3(new_n567), .A4(new_n568), .ZN(new_n673));
  AND3_X1   g0473(.A1(new_n664), .A2(new_n671), .A3(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT26), .ZN(new_n675));
  MUX2_X1   g0475(.A(new_n665), .B(new_n674), .S(new_n675), .Z(new_n676));
  INV_X1    g0476(.A(new_n527), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n677), .A2(new_n641), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n508), .A2(new_n600), .A3(new_n673), .A4(new_n607), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n671), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n676), .A2(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n663), .B1(new_n457), .B2(new_n681), .ZN(G369));
  NAND3_X1  g0482(.A1(new_n209), .A2(new_n210), .A3(G13), .ZN(new_n683));
  OR2_X1    g0483(.A1(new_n683), .A2(KEYINPUT27), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(KEYINPUT27), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n684), .A2(G213), .A3(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(G343), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n645), .A2(new_n689), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n690), .B1(new_n648), .B2(new_n651), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n641), .A2(new_n690), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(G330), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n525), .A2(new_n688), .ZN(new_n698));
  AOI22_X1  g0498(.A1(new_n530), .A2(new_n698), .B1(new_n677), .B2(new_n688), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n688), .B1(new_n649), .B2(new_n637), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n530), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n677), .A2(new_n689), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n701), .A2(new_n706), .ZN(G399));
  INV_X1    g0507(.A(new_n213), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n708), .A2(G41), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n541), .A2(G116), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n710), .A2(G1), .A3(new_n711), .ZN(new_n712));
  OAI22_X1  g0512(.A1(new_n712), .A2(KEYINPUT90), .B1(new_n219), .B2(new_n710), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n713), .B1(KEYINPUT90), .B2(new_n712), .ZN(new_n714));
  XOR2_X1   g0514(.A(new_n714), .B(KEYINPUT28), .Z(new_n715));
  OAI21_X1  g0515(.A(new_n689), .B1(new_n676), .B2(new_n680), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT29), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n664), .A2(new_n675), .A3(new_n570), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n719), .B1(new_n674), .B2(new_n675), .ZN(new_n720));
  OAI211_X1 g0520(.A(KEYINPUT29), .B(new_n689), .C1(new_n680), .C2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n529), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n528), .B1(new_n527), .B2(new_n508), .ZN(new_n723));
  OAI211_X1 g0523(.A(new_n652), .B(new_n689), .C1(new_n722), .C2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT31), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n689), .A2(new_n725), .ZN(new_n726));
  AND3_X1   g0526(.A1(new_n547), .A2(new_n554), .A3(new_n555), .ZN(new_n727));
  AND2_X1   g0527(.A1(new_n727), .A2(new_n478), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n728), .A2(KEYINPUT30), .A3(new_n638), .A4(new_n596), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n597), .A2(new_n520), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n669), .A2(new_n618), .A3(new_n297), .A4(new_n622), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n730), .B1(new_n731), .B2(KEYINPUT92), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n642), .A2(new_n643), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT92), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n733), .A2(new_n734), .A3(new_n297), .A4(new_n669), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n638), .A2(new_n727), .A3(new_n596), .A4(new_n478), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT91), .ZN(new_n737));
  AOI21_X1  g0537(.A(KEYINPUT30), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n728), .A2(KEYINPUT91), .A3(new_n638), .A4(new_n596), .ZN(new_n739));
  AOI22_X1  g0539(.A1(new_n732), .A2(new_n735), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n729), .B1(new_n740), .B2(KEYINPUT93), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n731), .A2(KEYINPUT92), .ZN(new_n742));
  INV_X1    g0542(.A(new_n730), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n742), .A2(new_n735), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n738), .A2(new_n739), .ZN(new_n745));
  AND3_X1   g0545(.A1(new_n744), .A2(new_n745), .A3(KEYINPUT93), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n726), .B1(new_n741), .B2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT94), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n744), .A2(new_n745), .A3(new_n729), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(new_n688), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n748), .B1(new_n750), .B2(new_n725), .ZN(new_n751));
  AOI211_X1 g0551(.A(KEYINPUT94), .B(KEYINPUT31), .C1(new_n749), .C2(new_n688), .ZN(new_n752));
  OAI211_X1 g0552(.A(new_n724), .B(new_n747), .C1(new_n751), .C2(new_n752), .ZN(new_n753));
  AOI22_X1  g0553(.A1(new_n718), .A2(new_n721), .B1(new_n753), .B2(G330), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n715), .B1(new_n754), .B2(G1), .ZN(G364));
  AND2_X1   g0555(.A1(new_n210), .A2(G13), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n209), .B1(new_n756), .B2(G45), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n709), .A2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n694), .A2(new_n695), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n697), .A2(new_n760), .A3(new_n761), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n216), .B1(G20), .B2(new_n300), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n210), .A2(new_n377), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n297), .A2(G200), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(G58), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n271), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n356), .A2(G179), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n765), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(new_n540), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n297), .A2(new_n356), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n210), .A2(G190), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n772), .B1(G68), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n774), .A2(new_n766), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n774), .A2(new_n770), .ZN(new_n779));
  OAI221_X1 g0579(.A(new_n777), .B1(new_n274), .B2(new_n778), .C1(new_n206), .C2(new_n779), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n297), .A2(new_n356), .A3(G190), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(G20), .ZN(new_n782));
  AOI211_X1 g0582(.A(new_n769), .B(new_n780), .C1(G97), .C2(new_n782), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n774), .A2(new_n297), .A3(new_n356), .ZN(new_n784));
  OR2_X1    g0584(.A1(new_n784), .A2(KEYINPUT96), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n784), .A2(KEYINPUT96), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n787), .A2(new_n381), .ZN(new_n788));
  XNOR2_X1  g0588(.A(KEYINPUT97), .B(KEYINPUT32), .ZN(new_n789));
  XNOR2_X1  g0589(.A(new_n788), .B(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(KEYINPUT95), .ZN(new_n791));
  AND3_X1   g0591(.A1(new_n773), .A2(new_n765), .A3(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n791), .B1(new_n773), .B2(new_n765), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  OAI211_X1 g0594(.A(new_n783), .B(new_n790), .C1(new_n265), .C2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n787), .ZN(new_n796));
  INV_X1    g0596(.A(new_n794), .ZN(new_n797));
  AOI22_X1  g0597(.A1(new_n796), .A2(G329), .B1(G326), .B2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n271), .ZN(new_n799));
  INV_X1    g0599(.A(G283), .ZN(new_n800));
  INV_X1    g0600(.A(new_n782), .ZN(new_n801));
  INV_X1    g0601(.A(G294), .ZN(new_n802));
  OAI221_X1 g0602(.A(new_n799), .B1(new_n779), .B2(new_n800), .C1(new_n801), .C2(new_n802), .ZN(new_n803));
  XOR2_X1   g0603(.A(KEYINPUT33), .B(G317), .Z(new_n804));
  INV_X1    g0604(.A(G303), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n804), .A2(new_n775), .B1(new_n771), .B2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(G322), .ZN(new_n807));
  INV_X1    g0607(.A(G311), .ZN(new_n808));
  OAI22_X1  g0608(.A1(new_n767), .A2(new_n807), .B1(new_n778), .B2(new_n808), .ZN(new_n809));
  NOR3_X1   g0609(.A1(new_n803), .A2(new_n806), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n798), .A2(new_n810), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n764), .B1(new_n795), .B2(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(G13), .A2(G33), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n814), .A2(G20), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n815), .A2(new_n763), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n708), .A2(new_n799), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n817), .A2(G355), .B1(new_n624), .B2(new_n708), .ZN(new_n818));
  AND2_X1   g0618(.A1(new_n251), .A2(G45), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n708), .A2(new_n271), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n820), .B1(G45), .B2(new_n219), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n818), .B1(new_n819), .B2(new_n821), .ZN(new_n822));
  AOI211_X1 g0622(.A(new_n760), .B(new_n812), .C1(new_n816), .C2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n694), .ZN(new_n824));
  INV_X1    g0624(.A(new_n815), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n823), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n762), .A2(new_n826), .ZN(G396));
  NAND2_X1  g0627(.A1(new_n655), .A2(new_n689), .ZN(new_n828));
  OAI22_X1  g0628(.A1(new_n378), .A2(new_n376), .B1(new_n366), .B2(new_n689), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n829), .A2(new_n375), .ZN(new_n830));
  AND2_X1   g0630(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n716), .A2(new_n832), .ZN(new_n833));
  OAI211_X1 g0633(.A(new_n689), .B(new_n831), .C1(new_n676), .C2(new_n680), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n753), .A2(G330), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n759), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n837), .B1(new_n836), .B2(new_n835), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n764), .A2(new_n814), .ZN(new_n839));
  XNOR2_X1  g0639(.A(new_n839), .B(KEYINPUT98), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n760), .B1(new_n841), .B2(new_n274), .ZN(new_n842));
  OAI22_X1  g0642(.A1(new_n787), .A2(new_n808), .B1(new_n805), .B2(new_n794), .ZN(new_n843));
  OAI22_X1  g0643(.A1(new_n767), .A2(new_n802), .B1(new_n778), .B2(new_n624), .ZN(new_n844));
  OAI22_X1  g0644(.A1(new_n771), .A2(new_n206), .B1(new_n779), .B2(new_n540), .ZN(new_n845));
  OAI221_X1 g0645(.A(new_n799), .B1(new_n775), .B2(new_n800), .C1(new_n801), .C2(new_n205), .ZN(new_n846));
  NOR4_X1   g0646(.A1(new_n843), .A2(new_n844), .A3(new_n845), .A4(new_n846), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n271), .B1(new_n779), .B2(new_n304), .ZN(new_n848));
  INV_X1    g0648(.A(new_n771), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n848), .B1(G50), .B2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(G132), .ZN(new_n851));
  OAI221_X1 g0651(.A(new_n850), .B1(new_n768), .B2(new_n801), .C1(new_n851), .C2(new_n787), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT34), .ZN(new_n853));
  INV_X1    g0653(.A(new_n767), .ZN(new_n854));
  INV_X1    g0654(.A(new_n778), .ZN(new_n855));
  AOI22_X1  g0655(.A1(G143), .A2(new_n854), .B1(new_n855), .B2(G159), .ZN(new_n856));
  INV_X1    g0656(.A(G150), .ZN(new_n857));
  INV_X1    g0657(.A(G137), .ZN(new_n858));
  OAI221_X1 g0658(.A(new_n856), .B1(new_n857), .B2(new_n775), .C1(new_n858), .C2(new_n794), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n852), .B1(new_n853), .B2(new_n859), .ZN(new_n860));
  OR2_X1    g0660(.A1(new_n859), .A2(new_n853), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n847), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  OAI221_X1 g0662(.A(new_n842), .B1(new_n764), .B2(new_n862), .C1(new_n831), .C2(new_n814), .ZN(new_n863));
  AND2_X1   g0663(.A1(new_n838), .A2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(G384));
  NOR2_X1   g0665(.A1(new_n577), .A2(new_n578), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  AND2_X1   g0667(.A1(new_n867), .A2(KEYINPUT35), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n867), .A2(KEYINPUT35), .ZN(new_n869));
  NOR4_X1   g0669(.A1(new_n868), .A2(new_n869), .A3(new_n218), .A4(new_n624), .ZN(new_n870));
  XNOR2_X1  g0670(.A(new_n870), .B(KEYINPUT36), .ZN(new_n871));
  OR3_X1    g0671(.A1(new_n219), .A2(new_n439), .A3(new_n274), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n201), .A2(G68), .ZN(new_n873));
  AOI211_X1 g0673(.A(new_n209), .B(G13), .C1(new_n872), .C2(new_n873), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n871), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n315), .A2(new_n689), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n352), .A2(new_n660), .A3(new_n877), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n876), .B1(new_n350), .B2(new_n351), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(new_n831), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n750), .A2(new_n725), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n749), .A2(KEYINPUT31), .A3(new_n688), .ZN(new_n883));
  AND2_X1   g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n881), .B1(new_n724), .B2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n686), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n450), .A2(KEYINPUT100), .A3(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT100), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n889), .B1(new_n425), .B2(new_n686), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT37), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n425), .A2(new_n432), .ZN(new_n893));
  AOI211_X1 g0693(.A(new_n407), .B(new_n420), .C1(new_n401), .C2(new_n404), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  AND3_X1   g0695(.A1(new_n891), .A2(new_n892), .A3(new_n895), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n446), .A2(KEYINPUT16), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n408), .B1(new_n396), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n898), .B1(new_n451), .B2(new_n887), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n892), .B1(new_n899), .B2(new_n422), .ZN(new_n900));
  OR2_X1    g0700(.A1(new_n896), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n898), .A2(new_n887), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n901), .B1(new_n456), .B2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT38), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  OAI211_X1 g0705(.A(new_n901), .B(KEYINPUT38), .C1(new_n456), .C2(new_n902), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n886), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  OR2_X1    g0707(.A1(new_n907), .A2(KEYINPUT40), .ZN(new_n908));
  AND2_X1   g0708(.A1(new_n888), .A2(new_n890), .ZN(new_n909));
  AOI21_X1  g0709(.A(KEYINPUT18), .B1(new_n450), .B2(new_n451), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n910), .A2(new_n434), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n909), .B1(new_n911), .B2(new_n427), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n892), .B1(new_n891), .B2(new_n895), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n912), .B1(new_n896), .B2(new_n913), .ZN(new_n914));
  AND3_X1   g0714(.A1(new_n914), .A2(KEYINPUT101), .A3(new_n904), .ZN(new_n915));
  AOI21_X1  g0715(.A(KEYINPUT101), .B1(new_n914), .B2(new_n904), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n906), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n917), .A2(KEYINPUT40), .A3(new_n885), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n908), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n884), .A2(new_n724), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n458), .A2(new_n920), .ZN(new_n921));
  OR2_X1    g0721(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n919), .A2(new_n921), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n922), .A2(G330), .A3(new_n923), .ZN(new_n924));
  XOR2_X1   g0724(.A(new_n924), .B(KEYINPUT102), .Z(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT99), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n834), .A2(new_n828), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n927), .B1(new_n928), .B2(new_n880), .ZN(new_n929));
  INV_X1    g0729(.A(new_n880), .ZN(new_n930));
  AOI211_X1 g0730(.A(KEYINPUT99), .B(new_n930), .C1(new_n834), .C2(new_n828), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n905), .A2(new_n906), .ZN(new_n933));
  AOI22_X1  g0733(.A1(new_n932), .A2(new_n933), .B1(new_n911), .B2(new_n686), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT39), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n917), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n353), .A2(new_n689), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n905), .A2(KEYINPUT39), .A3(new_n906), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n936), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n934), .A2(new_n940), .ZN(new_n941));
  NAND4_X1  g0741(.A1(new_n718), .A2(new_n456), .A3(new_n380), .A4(new_n721), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(new_n663), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n941), .B(new_n943), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n926), .A2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(new_n944), .ZN(new_n946));
  OAI22_X1  g0746(.A1(new_n925), .A2(new_n946), .B1(new_n209), .B2(new_n756), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n875), .B1(new_n945), .B2(new_n947), .ZN(G367));
  NAND2_X1  g0748(.A1(new_n664), .A2(new_n688), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n584), .A2(new_n688), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n600), .A2(new_n607), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n530), .A2(new_n702), .A3(new_n952), .ZN(new_n953));
  OR2_X1    g0753(.A1(new_n953), .A2(KEYINPUT42), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n953), .A2(KEYINPUT42), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n600), .B1(new_n951), .B2(new_n527), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n956), .A2(new_n689), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n954), .A2(new_n955), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n566), .A2(new_n568), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(new_n688), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n671), .A2(new_n960), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(KEYINPUT103), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n673), .A2(new_n671), .A3(new_n960), .ZN(new_n963));
  OR2_X1    g0763(.A1(new_n963), .A2(KEYINPUT104), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(KEYINPUT104), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n962), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(KEYINPUT43), .ZN(new_n967));
  XNOR2_X1  g0767(.A(KEYINPUT105), .B(KEYINPUT43), .ZN(new_n968));
  NAND4_X1  g0768(.A1(new_n962), .A2(new_n964), .A3(new_n965), .A4(new_n968), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n958), .A2(new_n967), .A3(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n970), .B1(new_n958), .B2(new_n969), .ZN(new_n971));
  INV_X1    g0771(.A(new_n952), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n701), .A2(new_n972), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n971), .B(new_n973), .ZN(new_n974));
  XOR2_X1   g0774(.A(new_n709), .B(KEYINPUT41), .Z(new_n975));
  OR3_X1    g0775(.A1(new_n705), .A2(KEYINPUT106), .A3(new_n972), .ZN(new_n976));
  INV_X1    g0776(.A(KEYINPUT45), .ZN(new_n977));
  OAI21_X1  g0777(.A(KEYINPUT106), .B1(new_n705), .B2(new_n972), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n976), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n979), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n977), .B1(new_n976), .B2(new_n978), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT107), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n705), .A2(new_n972), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT44), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n983), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n705), .A2(KEYINPUT44), .A3(new_n972), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n984), .A2(new_n985), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n988), .B1(KEYINPUT107), .B2(new_n989), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n700), .B1(new_n982), .B2(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(new_n702), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n699), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n993), .A2(new_n703), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n696), .A2(KEYINPUT108), .ZN(new_n995));
  OR2_X1    g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n696), .A2(KEYINPUT108), .ZN(new_n997));
  INV_X1    g0797(.A(new_n997), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n994), .B1(new_n998), .B2(new_n995), .ZN(new_n999));
  AND2_X1   g0799(.A1(new_n996), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n1000), .A2(new_n754), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1001), .A2(KEYINPUT109), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n990), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n981), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1004), .A2(new_n979), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1003), .A2(new_n1005), .A3(new_n701), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT109), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n1000), .A2(new_n1007), .A3(new_n754), .ZN(new_n1008));
  NAND4_X1  g0808(.A1(new_n991), .A2(new_n1002), .A3(new_n1006), .A4(new_n1008), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n975), .B1(new_n1009), .B2(new_n754), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n974), .B1(new_n1010), .B2(new_n758), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n816), .B1(new_n213), .B2(new_n361), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1012), .B1(new_n820), .B2(new_n237), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n796), .A2(G137), .B1(G143), .B2(new_n797), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n779), .A2(new_n274), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n857), .A2(new_n767), .B1(new_n775), .B2(new_n381), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n201), .ZN(new_n1017));
  AOI211_X1 g0817(.A(new_n1015), .B(new_n1016), .C1(new_n1017), .C2(new_n855), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n801), .A2(new_n304), .ZN(new_n1019));
  AOI211_X1 g0819(.A(new_n799), .B(new_n1019), .C1(G58), .C2(new_n849), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1014), .A2(new_n1018), .A3(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(G317), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n799), .B1(new_n205), .B2(new_n779), .C1(new_n787), .C2(new_n1022), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(KEYINPUT111), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n849), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n1025), .A2(KEYINPUT110), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1026), .B1(G311), .B2(new_n797), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n775), .A2(new_n802), .B1(new_n778), .B2(new_n800), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1028), .B1(G303), .B2(new_n854), .ZN(new_n1029));
  AOI21_X1  g0829(.A(KEYINPUT46), .B1(new_n849), .B2(G116), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1030), .B1(G107), .B2(new_n782), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1025), .A2(KEYINPUT110), .ZN(new_n1032));
  NAND4_X1  g0832(.A1(new_n1027), .A2(new_n1029), .A3(new_n1031), .A4(new_n1032), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1021), .B1(new_n1024), .B2(new_n1033), .ZN(new_n1034));
  XOR2_X1   g0834(.A(KEYINPUT112), .B(KEYINPUT47), .Z(new_n1035));
  XNOR2_X1  g0835(.A(new_n1034), .B(new_n1035), .ZN(new_n1036));
  AOI211_X1 g0836(.A(new_n760), .B(new_n1013), .C1(new_n1036), .C2(new_n763), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1037), .B1(new_n966), .B2(new_n825), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1011), .A2(new_n1038), .ZN(G387));
  INV_X1    g0839(.A(new_n711), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n817), .A2(new_n1040), .B1(new_n206), .B2(new_n708), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n242), .A2(new_n465), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n256), .A2(new_n265), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT50), .ZN(new_n1044));
  OAI211_X1 g0844(.A(new_n711), .B(new_n465), .C1(new_n304), .C2(new_n274), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n820), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1041), .B1(new_n1042), .B2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n760), .B1(new_n1047), .B2(new_n816), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n771), .A2(new_n274), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1049), .B1(G50), .B2(new_n854), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n1050), .B1(new_n304), .B2(new_n778), .C1(new_n364), .C2(new_n775), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n787), .A2(new_n857), .B1(new_n381), .B2(new_n794), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n801), .A2(new_n361), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n271), .B1(new_n779), .B2(new_n205), .ZN(new_n1054));
  NOR4_X1   g0854(.A1(new_n1051), .A2(new_n1052), .A3(new_n1053), .A4(new_n1054), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(G311), .A2(new_n776), .B1(new_n855), .B2(G303), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n1056), .B1(new_n1022), .B2(new_n767), .C1(new_n794), .C2(new_n807), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n1057), .ZN(new_n1058));
  OR2_X1    g0858(.A1(new_n1058), .A2(KEYINPUT48), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1058), .A2(KEYINPUT48), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n849), .A2(G294), .B1(G283), .B2(new_n782), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1059), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n1062), .ZN(new_n1063));
  OR2_X1    g0863(.A1(new_n1063), .A2(KEYINPUT49), .ZN(new_n1064));
  INV_X1    g0864(.A(G326), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n799), .B1(new_n624), .B2(new_n779), .C1(new_n787), .C2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1066), .B1(new_n1063), .B2(KEYINPUT49), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1055), .B1(new_n1064), .B2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1048), .B1(new_n1068), .B2(new_n764), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1069), .B1(new_n699), .B2(new_n815), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(new_n1000), .B2(new_n758), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1001), .A2(new_n709), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n1000), .A2(new_n754), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1071), .B1(new_n1072), .B2(new_n1073), .ZN(G393));
  INV_X1    g0874(.A(new_n1006), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n701), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n972), .A2(new_n815), .ZN(new_n1078));
  NOR3_X1   g0878(.A1(new_n247), .A2(new_n708), .A3(new_n271), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n816), .B1(new_n205), .B2(new_n213), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n759), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n797), .A2(G150), .B1(G159), .B2(new_n854), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1082), .ZN(new_n1083));
  XOR2_X1   g0883(.A(KEYINPUT113), .B(KEYINPUT51), .Z(new_n1084));
  NOR2_X1   g0884(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n1017), .A2(new_n776), .B1(new_n855), .B2(new_n256), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1086), .B1(new_n304), .B2(new_n771), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n801), .A2(new_n274), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n271), .B1(new_n779), .B2(new_n540), .ZN(new_n1089));
  OR3_X1    g0889(.A1(new_n1087), .A2(new_n1088), .A3(new_n1089), .ZN(new_n1090));
  AOI211_X1 g0890(.A(new_n1085), .B(new_n1090), .C1(G143), .C2(new_n796), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n794), .A2(new_n1022), .B1(new_n808), .B2(new_n767), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n1093), .B(KEYINPUT52), .ZN(new_n1094));
  OAI221_X1 g0894(.A(new_n799), .B1(new_n779), .B2(new_n206), .C1(new_n801), .C2(new_n624), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(G303), .A2(new_n776), .B1(new_n855), .B2(G294), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1096), .B1(new_n800), .B2(new_n771), .ZN(new_n1097));
  AOI211_X1 g0897(.A(new_n1095), .B(new_n1097), .C1(G322), .C2(new_n796), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n1091), .A2(new_n1092), .B1(new_n1094), .B2(new_n1098), .ZN(new_n1099));
  XOR2_X1   g0899(.A(new_n1099), .B(KEYINPUT114), .Z(new_n1100));
  AOI21_X1  g0900(.A(new_n1081), .B1(new_n1100), .B2(new_n763), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(new_n1077), .A2(new_n758), .B1(new_n1078), .B2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1001), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1103), .A2(new_n1009), .A3(new_n709), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1102), .A2(new_n1104), .ZN(G390));
  INV_X1    g0905(.A(G128), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n794), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n849), .A2(G150), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(new_n1108), .B(KEYINPUT53), .ZN(new_n1109));
  AOI211_X1 g0909(.A(new_n1107), .B(new_n1109), .C1(G125), .C2(new_n796), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(KEYINPUT54), .B(G143), .ZN(new_n1111));
  OAI22_X1  g0911(.A1(new_n767), .A2(new_n851), .B1(new_n778), .B2(new_n1111), .ZN(new_n1112));
  OAI221_X1 g0912(.A(new_n271), .B1(new_n775), .B2(new_n858), .C1(new_n801), .C2(new_n381), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n779), .ZN(new_n1114));
  AOI211_X1 g0914(.A(new_n1112), .B(new_n1113), .C1(new_n1017), .C2(new_n1114), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(G116), .A2(new_n854), .B1(new_n855), .B2(G97), .ZN(new_n1116));
  OAI221_X1 g0916(.A(new_n1116), .B1(new_n304), .B2(new_n779), .C1(new_n206), .C2(new_n775), .ZN(new_n1117));
  NOR4_X1   g0917(.A1(new_n1117), .A2(new_n271), .A3(new_n772), .A4(new_n1088), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n796), .A2(G294), .B1(G283), .B2(new_n797), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n1110), .A2(new_n1115), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  OAI221_X1 g0920(.A(new_n759), .B1(new_n256), .B2(new_n840), .C1(new_n1120), .C2(new_n764), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n896), .A2(new_n900), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n910), .B1(new_n436), .B2(new_n452), .ZN(new_n1123));
  AOI21_X1  g0923(.A(KEYINPUT81), .B1(new_n1123), .B2(new_n454), .ZN(new_n1124));
  NOR3_X1   g0924(.A1(new_n435), .A2(new_n428), .A3(new_n437), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n659), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n902), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1122), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(KEYINPUT101), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n891), .B1(new_n659), .B2(new_n654), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n891), .A2(new_n895), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1131), .A2(KEYINPUT37), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n891), .A2(new_n892), .A3(new_n895), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1130), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1129), .B1(new_n1134), .B2(KEYINPUT38), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n914), .A2(KEYINPUT101), .A3(new_n904), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(new_n1128), .A2(KEYINPUT38), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n939), .B1(new_n1137), .B2(KEYINPUT39), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1121), .B1(new_n1138), .B2(new_n813), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n886), .A2(new_n695), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n938), .B1(new_n928), .B2(new_n880), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1141), .B1(new_n936), .B2(new_n939), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n689), .B(new_n830), .C1(new_n680), .C2(new_n720), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(new_n828), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n938), .B1(new_n1144), .B2(new_n880), .ZN(new_n1145));
  AND2_X1   g0945(.A1(new_n917), .A2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1140), .B1(new_n1142), .B2(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1141), .ZN(new_n1148));
  AND3_X1   g0948(.A1(new_n905), .A2(KEYINPUT39), .A3(new_n906), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1150));
  AOI21_X1  g0950(.A(KEYINPUT39), .B1(new_n1150), .B2(new_n906), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1148), .B1(new_n1149), .B2(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1146), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n753), .A2(G330), .A3(new_n831), .A4(new_n880), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1152), .A2(new_n1153), .A3(new_n1154), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1147), .A2(new_n1155), .A3(KEYINPUT115), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1146), .B1(new_n1138), .B2(new_n1148), .ZN(new_n1157));
  INV_X1    g0957(.A(KEYINPUT115), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1157), .A2(new_n1158), .A3(new_n1154), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1156), .A2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1139), .B1(new_n1160), .B2(new_n758), .ZN(new_n1161));
  INV_X1    g0961(.A(KEYINPUT116), .ZN(new_n1162));
  AND3_X1   g0962(.A1(new_n530), .A2(new_n652), .A3(new_n689), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n882), .A2(new_n883), .ZN(new_n1164));
  OAI211_X1 g0964(.A(G330), .B(new_n831), .C1(new_n1163), .C2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1165), .A2(new_n930), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1144), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1166), .A2(new_n1167), .A3(new_n1154), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n753), .A2(G330), .A3(new_n831), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(new_n1169), .A2(new_n930), .B1(new_n885), .B2(G330), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n928), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1168), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  NAND4_X1  g0972(.A1(new_n920), .A2(new_n380), .A3(G330), .A4(new_n456), .ZN(new_n1173));
  AND3_X1   g0973(.A1(new_n942), .A2(new_n1173), .A3(new_n663), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1162), .B1(new_n1172), .B2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1172), .A2(new_n1162), .A3(new_n1174), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1176), .A2(KEYINPUT117), .A3(new_n1177), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n709), .B1(new_n1160), .B2(new_n1178), .ZN(new_n1179));
  AND3_X1   g0979(.A1(new_n1172), .A2(new_n1162), .A3(new_n1174), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n1180), .A2(new_n1175), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(new_n1156), .A2(new_n1159), .B1(new_n1181), .B2(KEYINPUT117), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1161), .B1(new_n1179), .B2(new_n1182), .ZN(G378));
  OAI21_X1  g0983(.A(new_n759), .B1(new_n1017), .B2(new_n839), .ZN(new_n1184));
  INV_X1    g0984(.A(G41), .ZN(new_n1185));
  AOI21_X1  g0985(.A(G50), .B1(new_n391), .B2(new_n1185), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(new_n796), .A2(G283), .B1(G116), .B2(new_n797), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(G107), .A2(new_n854), .B1(new_n855), .B2(new_n362), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(G97), .A2(new_n776), .B1(new_n1114), .B2(G58), .ZN(new_n1189));
  NOR4_X1   g0989(.A1(new_n1019), .A2(new_n1049), .A3(G41), .A4(new_n271), .ZN(new_n1190));
  NAND4_X1  g0990(.A1(new_n1187), .A2(new_n1188), .A3(new_n1189), .A4(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(KEYINPUT58), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1186), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n775), .A2(new_n851), .B1(new_n778), .B2(new_n858), .ZN(new_n1194));
  OAI22_X1  g0994(.A1(new_n1106), .A2(new_n767), .B1(new_n771), .B2(new_n1111), .ZN(new_n1195));
  AOI211_X1 g0995(.A(new_n1194), .B(new_n1195), .C1(G150), .C2(new_n782), .ZN(new_n1196));
  INV_X1    g0996(.A(G125), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1196), .B1(new_n1197), .B2(new_n794), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1198), .A2(KEYINPUT59), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n796), .A2(G124), .ZN(new_n1200));
  AOI211_X1 g1000(.A(G33), .B(G41), .C1(new_n1114), .C2(G159), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1199), .A2(new_n1200), .A3(new_n1201), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n1198), .A2(KEYINPUT59), .ZN(new_n1203));
  OAI221_X1 g1003(.A(new_n1193), .B1(new_n1192), .B2(new_n1191), .C1(new_n1202), .C2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1184), .B1(new_n1204), .B2(new_n763), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n269), .A2(new_n686), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(new_n303), .B(new_n1206), .ZN(new_n1207));
  XNOR2_X1  g1007(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1208));
  XNOR2_X1  g1008(.A(new_n1207), .B(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1209), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1205), .B1(new_n1210), .B2(new_n814), .ZN(new_n1211));
  XOR2_X1   g1011(.A(new_n1211), .B(KEYINPUT118), .Z(new_n1212));
  OAI211_X1 g1012(.A(new_n918), .B(G330), .C1(new_n907), .C2(KEYINPUT40), .ZN(new_n1213));
  AND2_X1   g1013(.A1(new_n1213), .A2(new_n1209), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n1213), .A2(new_n1209), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n941), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n908), .A2(G330), .A3(new_n918), .A4(new_n1210), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1213), .A2(new_n1209), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1217), .A2(new_n1218), .A3(new_n940), .A4(new_n934), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1216), .A2(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1212), .B1(new_n1220), .B2(new_n758), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1181), .B1(new_n1156), .B2(new_n1159), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1174), .ZN(new_n1223));
  OAI211_X1 g1023(.A(KEYINPUT57), .B(new_n1220), .C1(new_n1222), .C2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1224), .A2(new_n709), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1154), .ZN(new_n1226));
  NOR4_X1   g1026(.A1(new_n1142), .A2(new_n1146), .A3(new_n1226), .A4(KEYINPUT115), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1158), .B1(new_n1157), .B2(new_n1154), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1227), .B1(new_n1228), .B2(new_n1147), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1174), .B1(new_n1229), .B2(new_n1181), .ZN(new_n1230));
  AOI21_X1  g1030(.A(KEYINPUT57), .B1(new_n1230), .B2(new_n1220), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1221), .B1(new_n1225), .B2(new_n1231), .ZN(G375));
  NAND2_X1  g1032(.A1(new_n1172), .A2(new_n758), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n760), .B1(new_n841), .B2(new_n304), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(G97), .A2(new_n849), .B1(new_n855), .B2(G107), .ZN(new_n1235));
  OAI221_X1 g1035(.A(new_n1235), .B1(new_n624), .B2(new_n775), .C1(new_n800), .C2(new_n767), .ZN(new_n1236));
  NOR4_X1   g1036(.A1(new_n1236), .A2(new_n271), .A3(new_n1015), .A4(new_n1053), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n796), .A2(G303), .B1(G294), .B2(new_n797), .ZN(new_n1238));
  OAI221_X1 g1038(.A(new_n271), .B1(new_n779), .B2(new_n768), .C1(new_n801), .C2(new_n265), .ZN(new_n1239));
  OAI22_X1  g1039(.A1(new_n771), .A2(new_n381), .B1(new_n778), .B2(new_n857), .ZN(new_n1240));
  OAI22_X1  g1040(.A1(new_n858), .A2(new_n767), .B1(new_n775), .B2(new_n1111), .ZN(new_n1241));
  NOR3_X1   g1041(.A1(new_n1239), .A2(new_n1240), .A3(new_n1241), .ZN(new_n1242));
  AOI22_X1  g1042(.A1(new_n796), .A2(G128), .B1(G132), .B2(new_n797), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(new_n1237), .A2(new_n1238), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  OAI221_X1 g1044(.A(new_n1234), .B1(new_n764), .B2(new_n1244), .C1(new_n880), .C2(new_n814), .ZN(new_n1245));
  AND2_X1   g1045(.A1(new_n1233), .A2(new_n1245), .ZN(new_n1246));
  OR2_X1    g1046(.A1(new_n1172), .A2(new_n1174), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1181), .A2(new_n1247), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1246), .B1(new_n1248), .B2(new_n975), .ZN(G381));
  NAND2_X1  g1049(.A1(G378), .A2(KEYINPUT119), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT119), .ZN(new_n1251));
  OAI211_X1 g1051(.A(new_n1251), .B(new_n1161), .C1(new_n1179), .C2(new_n1182), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1250), .A2(new_n1252), .ZN(new_n1253));
  OR2_X1    g1053(.A1(new_n1253), .A2(G375), .ZN(new_n1254));
  NOR4_X1   g1054(.A1(G390), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1255), .A2(new_n1011), .A3(new_n1038), .ZN(new_n1256));
  OR3_X1    g1056(.A1(new_n1254), .A2(G381), .A3(new_n1256), .ZN(G407));
  OAI211_X1 g1057(.A(G407), .B(G213), .C1(G343), .C2(new_n1254), .ZN(new_n1258));
  XNOR2_X1  g1058(.A(new_n1258), .B(KEYINPUT120), .ZN(G409));
  INV_X1    g1059(.A(KEYINPUT125), .ZN(new_n1260));
  INV_X1    g1060(.A(G390), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(G387), .A2(new_n1261), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1011), .A2(G390), .A3(new_n1038), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1262), .A2(KEYINPUT123), .A3(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT123), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1011), .A2(G390), .A3(new_n1265), .A4(new_n1038), .ZN(new_n1266));
  XNOR2_X1  g1066(.A(G393), .B(G396), .ZN(new_n1267));
  AND2_X1   g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1264), .A2(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1267), .B1(G387), .B2(new_n1261), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1263), .A2(KEYINPUT122), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT122), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1011), .A2(G390), .A3(new_n1272), .A4(new_n1038), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1270), .A2(new_n1271), .A3(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1269), .A2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT61), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n687), .A2(G213), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n975), .ZN(new_n1280));
  OAI211_X1 g1080(.A(new_n1280), .B(new_n1220), .C1(new_n1222), .C2(new_n1223), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(new_n1221), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1250), .A2(new_n1252), .A3(new_n1282), .ZN(new_n1283));
  OAI211_X1 g1083(.A(G378), .B(new_n1221), .C1(new_n1225), .C2(new_n1231), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1279), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1248), .A2(KEYINPUT60), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT60), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n710), .B1(new_n1247), .B2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1286), .A2(new_n1288), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1289), .A2(G384), .A3(new_n1246), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1288), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1291), .B1(new_n1248), .B2(KEYINPUT60), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1246), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n864), .B1(new_n1292), .B2(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(G2897), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1278), .A2(new_n1295), .ZN(new_n1296));
  AND3_X1   g1096(.A1(new_n1290), .A2(new_n1294), .A3(new_n1296), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1296), .B1(new_n1290), .B2(new_n1294), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1277), .B1(new_n1285), .B2(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1290), .A2(new_n1294), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1302), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1301), .A2(new_n1278), .A3(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT124), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT62), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1300), .B1(new_n1306), .B2(new_n1307), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1304), .A2(new_n1305), .A3(KEYINPUT62), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1276), .B1(new_n1308), .B2(new_n1309), .ZN(new_n1310));
  AOI211_X1 g1110(.A(new_n1279), .B(new_n1302), .C1(new_n1283), .C2(new_n1284), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1311), .A2(KEYINPUT63), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1285), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT121), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1314), .B1(new_n1297), .B2(new_n1298), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1299), .A2(KEYINPUT121), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1313), .A2(new_n1315), .A3(new_n1316), .ZN(new_n1317));
  NOR2_X1   g1117(.A1(new_n1275), .A2(KEYINPUT61), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT63), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1304), .A2(new_n1319), .ZN(new_n1320));
  NAND4_X1  g1120(.A1(new_n1312), .A2(new_n1317), .A3(new_n1318), .A4(new_n1320), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1321), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1260), .B1(new_n1310), .B2(new_n1322), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1307), .B1(new_n1311), .B2(KEYINPUT124), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1300), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1324), .A2(new_n1325), .A3(new_n1309), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1326), .A2(new_n1275), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1327), .A2(KEYINPUT125), .A3(new_n1321), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1323), .A2(new_n1328), .ZN(G405));
  AND3_X1   g1129(.A1(G375), .A2(new_n1250), .A3(new_n1252), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT126), .ZN(new_n1331));
  OAI21_X1  g1131(.A(new_n1284), .B1(new_n1331), .B2(new_n1302), .ZN(new_n1332));
  NOR2_X1   g1132(.A1(new_n1330), .A2(new_n1332), .ZN(new_n1333));
  XNOR2_X1  g1133(.A(new_n1333), .B(new_n1275), .ZN(new_n1334));
  NOR2_X1   g1134(.A1(new_n1303), .A2(KEYINPUT126), .ZN(new_n1335));
  XNOR2_X1  g1135(.A(new_n1334), .B(new_n1335), .ZN(G402));
endmodule


