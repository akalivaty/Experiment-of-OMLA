

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725;

  INV_X1 U373 ( .A(G953), .ZN(n712) );
  XNOR2_X2 U374 ( .A(n529), .B(KEYINPUT1), .ZN(n569) );
  NOR2_X1 U375 ( .A1(n566), .A2(n635), .ZN(n540) );
  XNOR2_X1 U376 ( .A(n539), .B(n372), .ZN(n566) );
  XNOR2_X1 U377 ( .A(n407), .B(n406), .ZN(n493) );
  XNOR2_X1 U378 ( .A(n445), .B(n444), .ZN(n574) );
  XNOR2_X1 U379 ( .A(n376), .B(n460), .ZN(n423) );
  XNOR2_X1 U380 ( .A(n423), .B(KEYINPUT92), .ZN(n709) );
  XNOR2_X1 U381 ( .A(n367), .B(G128), .ZN(n438) );
  INV_X1 U382 ( .A(G143), .ZN(n367) );
  XNOR2_X1 U383 ( .A(KEYINPUT3), .B(G119), .ZN(n417) );
  AND2_X1 U384 ( .A1(n609), .A2(n353), .ZN(n362) );
  NOR2_X1 U385 ( .A1(G953), .A2(G237), .ZN(n466) );
  XNOR2_X1 U386 ( .A(n373), .B(KEYINPUT70), .ZN(n375) );
  XOR2_X1 U387 ( .A(KEYINPUT4), .B(G137), .Z(n373) );
  XOR2_X1 U388 ( .A(G104), .B(G110), .Z(n378) );
  XOR2_X1 U389 ( .A(G146), .B(G140), .Z(n379) );
  INV_X1 U390 ( .A(KEYINPUT78), .ZN(n381) );
  NOR2_X1 U391 ( .A1(n520), .A2(n672), .ZN(n678) );
  INV_X1 U392 ( .A(G469), .ZN(n386) );
  XNOR2_X1 U393 ( .A(KEYINPUT75), .B(KEYINPUT16), .ZN(n428) );
  XNOR2_X1 U394 ( .A(G113), .B(G104), .ZN(n474) );
  XNOR2_X1 U395 ( .A(n393), .B(n392), .ZN(n396) );
  XNOR2_X1 U396 ( .A(n391), .B(n390), .ZN(n393) );
  XNOR2_X1 U397 ( .A(n395), .B(KEYINPUT10), .ZN(n708) );
  XNOR2_X1 U398 ( .A(n370), .B(KEYINPUT100), .ZN(n369) );
  XNOR2_X1 U399 ( .A(KEYINPUT7), .B(KEYINPUT9), .ZN(n370) );
  XNOR2_X1 U400 ( .A(n371), .B(G107), .ZN(n459) );
  XNOR2_X1 U401 ( .A(G122), .B(G116), .ZN(n371) );
  XNOR2_X1 U402 ( .A(n438), .B(n366), .ZN(n460) );
  INV_X1 U403 ( .A(G134), .ZN(n366) );
  INV_X1 U404 ( .A(n582), .ZN(n583) );
  XNOR2_X1 U405 ( .A(n357), .B(n441), .ZN(n586) );
  NAND2_X1 U406 ( .A1(n355), .A2(n519), .ZN(n354) );
  XNOR2_X1 U407 ( .A(n356), .B(n502), .ZN(n355) );
  XNOR2_X1 U408 ( .A(G478), .B(n464), .ZN(n510) );
  XNOR2_X1 U409 ( .A(n359), .B(n491), .ZN(n498) );
  OR2_X1 U410 ( .A1(n507), .A2(n490), .ZN(n359) );
  XNOR2_X1 U411 ( .A(KEYINPUT96), .B(KEYINPUT99), .ZN(n469) );
  NAND2_X1 U412 ( .A1(G234), .A2(G237), .ZN(n449) );
  XOR2_X1 U413 ( .A(G146), .B(KEYINPUT95), .Z(n412) );
  XNOR2_X1 U414 ( .A(G113), .B(G116), .ZN(n414) );
  XNOR2_X1 U415 ( .A(G128), .B(G110), .ZN(n388) );
  XNOR2_X1 U416 ( .A(G131), .B(KEYINPUT69), .ZN(n374) );
  XNOR2_X1 U417 ( .A(G143), .B(G122), .ZN(n473) );
  XNOR2_X1 U418 ( .A(n394), .B(G146), .ZN(n436) );
  INV_X1 U419 ( .A(G125), .ZN(n394) );
  XNOR2_X1 U420 ( .A(KEYINPUT87), .B(KEYINPUT4), .ZN(n437) );
  XNOR2_X1 U421 ( .A(n427), .B(n426), .ZN(n680) );
  INV_X1 U422 ( .A(G237), .ZN(n442) );
  XNOR2_X1 U423 ( .A(n709), .B(n385), .ZN(n694) );
  XNOR2_X1 U424 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U425 ( .A(n380), .B(n379), .ZN(n384) );
  XNOR2_X1 U426 ( .A(n521), .B(n365), .ZN(n670) );
  INV_X1 U427 ( .A(KEYINPUT41), .ZN(n365) );
  OR2_X1 U428 ( .A1(n574), .A2(n676), .ZN(n547) );
  XNOR2_X1 U429 ( .A(n547), .B(KEYINPUT19), .ZN(n554) );
  NOR2_X1 U430 ( .A1(n527), .A2(n544), .ZN(n528) );
  XNOR2_X1 U431 ( .A(n480), .B(n479), .ZN(n511) );
  XNOR2_X1 U432 ( .A(n432), .B(n431), .ZN(n357) );
  XNOR2_X1 U433 ( .A(G119), .B(G137), .ZN(n398) );
  XNOR2_X1 U434 ( .A(n368), .B(n460), .ZN(n463) );
  XNOR2_X1 U435 ( .A(n459), .B(n369), .ZN(n368) );
  NAND2_X2 U436 ( .A1(n361), .A2(n360), .ZN(n703) );
  NAND2_X1 U437 ( .A1(n649), .A2(n351), .ZN(n360) );
  NAND2_X1 U438 ( .A1(n362), .A2(n643), .ZN(n361) );
  AND2_X1 U439 ( .A1(n590), .A2(G953), .ZN(n707) );
  XNOR2_X1 U440 ( .A(n364), .B(n363), .ZN(n725) );
  XNOR2_X1 U441 ( .A(n531), .B(KEYINPUT107), .ZN(n363) );
  NOR2_X1 U442 ( .A1(n670), .A2(n556), .ZN(n364) );
  INV_X1 U443 ( .A(KEYINPUT42), .ZN(n531) );
  NAND2_X1 U444 ( .A1(n498), .A2(n358), .ZN(n496) );
  AND2_X1 U445 ( .A1(n494), .A2(n492), .ZN(n358) );
  AND2_X1 U446 ( .A1(n498), .A2(n492), .ZN(n516) );
  INV_X1 U447 ( .A(n710), .ZN(n643) );
  AND2_X1 U448 ( .A1(n583), .A2(KEYINPUT2), .ZN(n351) );
  NOR2_X1 U449 ( .A1(n357), .A2(n608), .ZN(n352) );
  AND2_X1 U450 ( .A1(n583), .A2(n581), .ZN(n353) );
  XNOR2_X2 U451 ( .A(n354), .B(KEYINPUT45), .ZN(n609) );
  NAND2_X1 U452 ( .A1(n501), .A2(n722), .ZN(n356) );
  XNOR2_X1 U453 ( .A(n396), .B(n708), .ZN(n401) );
  NOR2_X1 U454 ( .A1(G902), .A2(n596), .ZN(n479) );
  XNOR2_X1 U455 ( .A(KEYINPUT83), .B(KEYINPUT39), .ZN(n372) );
  INV_X1 U456 ( .A(KEYINPUT46), .ZN(n541) );
  INV_X1 U457 ( .A(KEYINPUT5), .ZN(n413) );
  XNOR2_X1 U458 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U459 ( .A(n416), .B(n415), .ZN(n421) );
  XNOR2_X1 U460 ( .A(n375), .B(n465), .ZN(n376) );
  XNOR2_X1 U461 ( .A(n405), .B(n404), .ZN(n406) );
  INV_X1 U462 ( .A(KEYINPUT77), .ZN(n392) );
  XNOR2_X1 U463 ( .A(n384), .B(n383), .ZN(n385) );
  BUF_X1 U464 ( .A(n710), .Z(n711) );
  XNOR2_X1 U465 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U466 ( .A(n486), .B(n485), .ZN(n722) );
  XNOR2_X1 U467 ( .A(n374), .B(KEYINPUT68), .ZN(n465) );
  XNOR2_X1 U468 ( .A(G101), .B(G107), .ZN(n377) );
  XNOR2_X1 U469 ( .A(n378), .B(n377), .ZN(n380) );
  NAND2_X1 U470 ( .A1(G227), .A2(n712), .ZN(n382) );
  NOR2_X1 U471 ( .A1(G902), .A2(n694), .ZN(n387) );
  XNOR2_X2 U472 ( .A(n387), .B(n386), .ZN(n529) );
  INV_X1 U473 ( .A(n569), .ZN(n543) );
  XOR2_X1 U474 ( .A(KEYINPUT93), .B(KEYINPUT94), .Z(n389) );
  XNOR2_X1 U475 ( .A(n389), .B(n388), .ZN(n391) );
  XOR2_X1 U476 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n390) );
  XNOR2_X1 U477 ( .A(n436), .B(G140), .ZN(n395) );
  NAND2_X1 U478 ( .A1(G234), .A2(n712), .ZN(n397) );
  XOR2_X1 U479 ( .A(KEYINPUT8), .B(n397), .Z(n461) );
  NAND2_X1 U480 ( .A1(n461), .A2(G221), .ZN(n399) );
  XNOR2_X1 U481 ( .A(n401), .B(n400), .ZN(n705) );
  NOR2_X1 U482 ( .A1(G902), .A2(n705), .ZN(n407) );
  XNOR2_X1 U483 ( .A(KEYINPUT88), .B(KEYINPUT15), .ZN(n402) );
  XNOR2_X1 U484 ( .A(n402), .B(G902), .ZN(n582) );
  NAND2_X1 U485 ( .A1(n582), .A2(G234), .ZN(n403) );
  XNOR2_X1 U486 ( .A(KEYINPUT20), .B(n403), .ZN(n408) );
  NAND2_X1 U487 ( .A1(G217), .A2(n408), .ZN(n405) );
  INV_X1 U488 ( .A(KEYINPUT25), .ZN(n404) );
  AND2_X1 U489 ( .A1(n408), .A2(G221), .ZN(n410) );
  INV_X1 U490 ( .A(KEYINPUT21), .ZN(n409) );
  XNOR2_X1 U491 ( .A(n410), .B(n409), .ZN(n654) );
  NOR2_X2 U492 ( .A1(n493), .A2(n654), .ZN(n506) );
  INV_X1 U493 ( .A(n506), .ZN(n657) );
  NOR2_X2 U494 ( .A1(n543), .A2(n657), .ZN(n503) );
  NAND2_X1 U495 ( .A1(n466), .A2(G210), .ZN(n411) );
  XNOR2_X1 U496 ( .A(n412), .B(n411), .ZN(n416) );
  XNOR2_X1 U497 ( .A(n417), .B(KEYINPUT72), .ZN(n419) );
  XNOR2_X1 U498 ( .A(G101), .B(KEYINPUT71), .ZN(n418) );
  XNOR2_X1 U499 ( .A(n419), .B(n418), .ZN(n431) );
  INV_X1 U500 ( .A(n431), .ZN(n420) );
  XNOR2_X1 U501 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U502 ( .A(n423), .B(n422), .ZN(n602) );
  INV_X1 U503 ( .A(G902), .ZN(n443) );
  NAND2_X1 U504 ( .A1(n602), .A2(n443), .ZN(n424) );
  XNOR2_X2 U505 ( .A(n424), .B(G472), .ZN(n663) );
  INV_X1 U506 ( .A(KEYINPUT6), .ZN(n425) );
  XNOR2_X1 U507 ( .A(n663), .B(n425), .ZN(n545) );
  NAND2_X1 U508 ( .A1(n503), .A2(n545), .ZN(n427) );
  XOR2_X1 U509 ( .A(KEYINPUT86), .B(KEYINPUT33), .Z(n426) );
  XNOR2_X1 U510 ( .A(n428), .B(G110), .ZN(n429) );
  XNOR2_X1 U511 ( .A(n429), .B(n474), .ZN(n430) );
  XNOR2_X1 U512 ( .A(n430), .B(n459), .ZN(n432) );
  XNOR2_X1 U513 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n434) );
  NAND2_X1 U514 ( .A1(n712), .A2(G224), .ZN(n433) );
  XNOR2_X1 U515 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U516 ( .A(n436), .B(n435), .ZN(n440) );
  XNOR2_X1 U517 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U518 ( .A(n440), .B(n439), .ZN(n441) );
  NAND2_X1 U519 ( .A1(n586), .A2(n582), .ZN(n445) );
  NAND2_X1 U520 ( .A1(n443), .A2(n442), .ZN(n446) );
  NAND2_X1 U521 ( .A1(n446), .A2(G210), .ZN(n444) );
  NAND2_X1 U522 ( .A1(n446), .A2(G214), .ZN(n448) );
  INV_X1 U523 ( .A(KEYINPUT89), .ZN(n447) );
  XNOR2_X1 U524 ( .A(n448), .B(n447), .ZN(n570) );
  INV_X1 U525 ( .A(n570), .ZN(n676) );
  XNOR2_X1 U526 ( .A(n449), .B(KEYINPUT14), .ZN(n452) );
  NAND2_X1 U527 ( .A1(G952), .A2(n452), .ZN(n450) );
  XOR2_X1 U528 ( .A(KEYINPUT90), .B(n450), .Z(n684) );
  NAND2_X1 U529 ( .A1(n684), .A2(n712), .ZN(n525) );
  NOR2_X1 U530 ( .A1(G898), .A2(n712), .ZN(n451) );
  XOR2_X1 U531 ( .A(KEYINPUT91), .B(n451), .Z(n608) );
  NAND2_X1 U532 ( .A1(G902), .A2(n452), .ZN(n522) );
  INV_X1 U533 ( .A(n522), .ZN(n453) );
  NAND2_X1 U534 ( .A1(n608), .A2(n453), .ZN(n454) );
  NAND2_X1 U535 ( .A1(n525), .A2(n454), .ZN(n455) );
  NAND2_X1 U536 ( .A1(n554), .A2(n455), .ZN(n456) );
  XNOR2_X1 U537 ( .A(n456), .B(KEYINPUT0), .ZN(n507) );
  NOR2_X1 U538 ( .A1(n680), .A2(n507), .ZN(n458) );
  XNOR2_X1 U539 ( .A(KEYINPUT74), .B(KEYINPUT34), .ZN(n457) );
  XNOR2_X1 U540 ( .A(n458), .B(n457), .ZN(n484) );
  NAND2_X1 U541 ( .A1(G217), .A2(n461), .ZN(n462) );
  XNOR2_X1 U542 ( .A(n463), .B(n462), .ZN(n700) );
  NOR2_X1 U543 ( .A1(G902), .A2(n700), .ZN(n464) );
  INV_X1 U544 ( .A(n510), .ZN(n481) );
  XNOR2_X1 U545 ( .A(KEYINPUT13), .B(G475), .ZN(n480) );
  XNOR2_X1 U546 ( .A(n465), .B(n708), .ZN(n478) );
  XOR2_X1 U547 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n468) );
  NAND2_X1 U548 ( .A1(G214), .A2(n466), .ZN(n467) );
  XNOR2_X1 U549 ( .A(n468), .B(n467), .ZN(n472) );
  XOR2_X1 U550 ( .A(KEYINPUT98), .B(KEYINPUT97), .Z(n470) );
  XNOR2_X1 U551 ( .A(n470), .B(n469), .ZN(n471) );
  XOR2_X1 U552 ( .A(n472), .B(n471), .Z(n476) );
  XNOR2_X1 U553 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X1 U554 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U555 ( .A(n478), .B(n477), .ZN(n596) );
  NAND2_X1 U556 ( .A1(n481), .A2(n511), .ZN(n482) );
  XNOR2_X1 U557 ( .A(n482), .B(KEYINPUT102), .ZN(n553) );
  INV_X1 U558 ( .A(n553), .ZN(n483) );
  NAND2_X1 U559 ( .A1(n484), .A2(n483), .ZN(n486) );
  XNOR2_X1 U560 ( .A(KEYINPUT79), .B(KEYINPUT35), .ZN(n485) );
  INV_X1 U561 ( .A(n511), .ZN(n487) );
  NAND2_X1 U562 ( .A1(n487), .A2(n510), .ZN(n488) );
  XNOR2_X1 U563 ( .A(n488), .B(KEYINPUT101), .ZN(n674) );
  INV_X1 U564 ( .A(n654), .ZN(n489) );
  NAND2_X1 U565 ( .A1(n674), .A2(n489), .ZN(n490) );
  XNOR2_X1 U566 ( .A(KEYINPUT65), .B(KEYINPUT22), .ZN(n491) );
  INV_X1 U567 ( .A(n545), .ZN(n492) );
  AND2_X1 U568 ( .A1(n569), .A2(n493), .ZN(n494) );
  XNOR2_X1 U569 ( .A(KEYINPUT64), .B(KEYINPUT32), .ZN(n495) );
  XNOR2_X1 U570 ( .A(n496), .B(n495), .ZN(n594) );
  INV_X1 U571 ( .A(n663), .ZN(n527) );
  NAND2_X1 U572 ( .A1(n493), .A2(n527), .ZN(n497) );
  NOR2_X1 U573 ( .A1(n569), .A2(n497), .ZN(n499) );
  AND2_X1 U574 ( .A1(n499), .A2(n498), .ZN(n627) );
  INV_X1 U575 ( .A(n627), .ZN(n500) );
  AND2_X1 U576 ( .A1(n594), .A2(n500), .ZN(n501) );
  NOR2_X1 U577 ( .A1(KEYINPUT44), .A2(KEYINPUT73), .ZN(n502) );
  NAND2_X1 U578 ( .A1(n503), .A2(n663), .ZN(n665) );
  OR2_X1 U579 ( .A1(n665), .A2(n507), .ZN(n505) );
  INV_X1 U580 ( .A(KEYINPUT31), .ZN(n504) );
  XNOR2_X1 U581 ( .A(n505), .B(n504), .ZN(n637) );
  NAND2_X1 U582 ( .A1(n506), .A2(n529), .ZN(n534) );
  NOR2_X1 U583 ( .A1(n534), .A2(n663), .ZN(n509) );
  INV_X1 U584 ( .A(n507), .ZN(n508) );
  NAND2_X1 U585 ( .A1(n509), .A2(n508), .ZN(n621) );
  NAND2_X1 U586 ( .A1(n637), .A2(n621), .ZN(n513) );
  NAND2_X1 U587 ( .A1(n511), .A2(n510), .ZN(n635) );
  INV_X1 U588 ( .A(n635), .ZN(n632) );
  NOR2_X1 U589 ( .A1(n511), .A2(n510), .ZN(n628) );
  NOR2_X1 U590 ( .A1(n632), .A2(n628), .ZN(n671) );
  XNOR2_X1 U591 ( .A(KEYINPUT81), .B(n671), .ZN(n512) );
  NAND2_X1 U592 ( .A1(n513), .A2(n512), .ZN(n515) );
  NAND2_X1 U593 ( .A1(KEYINPUT44), .A2(KEYINPUT73), .ZN(n514) );
  NAND2_X1 U594 ( .A1(n515), .A2(n514), .ZN(n518) );
  NOR2_X1 U595 ( .A1(n569), .A2(n493), .ZN(n517) );
  AND2_X1 U596 ( .A1(n517), .A2(n516), .ZN(n617) );
  NOR2_X1 U597 ( .A1(n518), .A2(n617), .ZN(n519) );
  INV_X1 U598 ( .A(n674), .ZN(n520) );
  XOR2_X1 U599 ( .A(KEYINPUT38), .B(n574), .Z(n672) );
  NAND2_X1 U600 ( .A1(n570), .A2(n678), .ZN(n521) );
  AND2_X1 U601 ( .A1(n489), .A2(n493), .ZN(n526) );
  NOR2_X1 U602 ( .A1(G900), .A2(n522), .ZN(n523) );
  NAND2_X1 U603 ( .A1(G953), .A2(n523), .ZN(n524) );
  NAND2_X1 U604 ( .A1(n525), .A2(n524), .ZN(n537) );
  NAND2_X1 U605 ( .A1(n526), .A2(n537), .ZN(n544) );
  XNOR2_X1 U606 ( .A(KEYINPUT28), .B(n528), .ZN(n530) );
  NAND2_X1 U607 ( .A1(n530), .A2(n529), .ZN(n556) );
  XOR2_X1 U608 ( .A(KEYINPUT30), .B(KEYINPUT105), .Z(n533) );
  NAND2_X1 U609 ( .A1(n663), .A2(n570), .ZN(n532) );
  XNOR2_X1 U610 ( .A(n533), .B(n532), .ZN(n535) );
  NOR2_X1 U611 ( .A1(n535), .A2(n534), .ZN(n536) );
  NAND2_X1 U612 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U613 ( .A(n538), .B(KEYINPUT76), .ZN(n550) );
  OR2_X2 U614 ( .A1(n550), .A2(n672), .ZN(n539) );
  XNOR2_X1 U615 ( .A(n540), .B(KEYINPUT40), .ZN(n724) );
  NOR2_X1 U616 ( .A1(n725), .A2(n724), .ZN(n542) );
  XNOR2_X1 U617 ( .A(n542), .B(n541), .ZN(n564) );
  NOR2_X1 U618 ( .A1(n544), .A2(n635), .ZN(n546) );
  NAND2_X1 U619 ( .A1(n546), .A2(n545), .ZN(n568) );
  NOR2_X1 U620 ( .A1(n568), .A2(n547), .ZN(n548) );
  XOR2_X1 U621 ( .A(KEYINPUT36), .B(n548), .Z(n549) );
  NOR2_X1 U622 ( .A1(n543), .A2(n549), .ZN(n641) );
  NOR2_X1 U623 ( .A1(n550), .A2(n574), .ZN(n551) );
  XOR2_X1 U624 ( .A(KEYINPUT106), .B(n551), .Z(n552) );
  NOR2_X1 U625 ( .A1(n553), .A2(n552), .ZN(n631) );
  NOR2_X1 U626 ( .A1(n641), .A2(n631), .ZN(n562) );
  INV_X1 U627 ( .A(n554), .ZN(n555) );
  NOR2_X1 U628 ( .A1(n556), .A2(n555), .ZN(n633) );
  NOR2_X1 U629 ( .A1(KEYINPUT47), .A2(KEYINPUT81), .ZN(n557) );
  XNOR2_X1 U630 ( .A(n557), .B(n671), .ZN(n558) );
  NAND2_X1 U631 ( .A1(n633), .A2(n558), .ZN(n560) );
  OR2_X1 U632 ( .A1(n633), .A2(KEYINPUT47), .ZN(n559) );
  NAND2_X1 U633 ( .A1(n560), .A2(n559), .ZN(n561) );
  NAND2_X1 U634 ( .A1(n562), .A2(n561), .ZN(n563) );
  NOR2_X2 U635 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U636 ( .A(n565), .B(KEYINPUT48), .ZN(n579) );
  INV_X1 U637 ( .A(n628), .ZN(n638) );
  OR2_X1 U638 ( .A1(n638), .A2(n566), .ZN(n567) );
  XNOR2_X1 U639 ( .A(n567), .B(KEYINPUT108), .ZN(n720) );
  XOR2_X1 U640 ( .A(KEYINPUT43), .B(KEYINPUT103), .Z(n573) );
  NOR2_X1 U641 ( .A1(n569), .A2(n568), .ZN(n571) );
  NAND2_X1 U642 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U643 ( .A(n573), .B(n572), .ZN(n575) );
  AND2_X1 U644 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U645 ( .A(n576), .B(KEYINPUT104), .ZN(n723) );
  INV_X1 U646 ( .A(n723), .ZN(n577) );
  AND2_X1 U647 ( .A1(n720), .A2(n577), .ZN(n578) );
  NAND2_X1 U648 ( .A1(n579), .A2(n578), .ZN(n580) );
  INV_X1 U649 ( .A(n580), .ZN(n646) );
  NAND2_X1 U650 ( .A1(n609), .A2(n646), .ZN(n649) );
  XNOR2_X1 U651 ( .A(n580), .B(KEYINPUT82), .ZN(n710) );
  INV_X1 U652 ( .A(KEYINPUT2), .ZN(n581) );
  NAND2_X1 U653 ( .A1(n703), .A2(G210), .ZN(n589) );
  XOR2_X1 U654 ( .A(KEYINPUT55), .B(KEYINPUT85), .Z(n585) );
  XNOR2_X1 U655 ( .A(KEYINPUT54), .B(KEYINPUT121), .ZN(n584) );
  XNOR2_X1 U656 ( .A(n585), .B(n584), .ZN(n587) );
  XOR2_X1 U657 ( .A(n587), .B(n586), .Z(n588) );
  XNOR2_X1 U658 ( .A(n589), .B(n588), .ZN(n591) );
  INV_X1 U659 ( .A(G952), .ZN(n590) );
  NOR2_X2 U660 ( .A1(n591), .A2(n707), .ZN(n593) );
  XNOR2_X1 U661 ( .A(KEYINPUT122), .B(KEYINPUT56), .ZN(n592) );
  XNOR2_X1 U662 ( .A(n593), .B(n592), .ZN(G51) );
  XNOR2_X1 U663 ( .A(n594), .B(G119), .ZN(G21) );
  NAND2_X1 U664 ( .A1(n703), .A2(G475), .ZN(n598) );
  XOR2_X1 U665 ( .A(KEYINPUT66), .B(KEYINPUT59), .Z(n595) );
  XNOR2_X1 U666 ( .A(n596), .B(n595), .ZN(n597) );
  XNOR2_X1 U667 ( .A(n598), .B(n597), .ZN(n599) );
  NOR2_X2 U668 ( .A1(n599), .A2(n707), .ZN(n601) );
  XOR2_X1 U669 ( .A(KEYINPUT67), .B(KEYINPUT60), .Z(n600) );
  XNOR2_X1 U670 ( .A(n601), .B(n600), .ZN(G60) );
  NAND2_X1 U671 ( .A1(n703), .A2(G472), .ZN(n604) );
  XOR2_X1 U672 ( .A(KEYINPUT62), .B(n602), .Z(n603) );
  XNOR2_X1 U673 ( .A(n604), .B(n603), .ZN(n605) );
  NOR2_X2 U674 ( .A1(n605), .A2(n707), .ZN(n607) );
  XOR2_X1 U675 ( .A(KEYINPUT84), .B(KEYINPUT63), .Z(n606) );
  XNOR2_X1 U676 ( .A(n607), .B(n606), .ZN(G57) );
  NAND2_X1 U677 ( .A1(n609), .A2(n712), .ZN(n610) );
  XNOR2_X1 U678 ( .A(n610), .B(KEYINPUT125), .ZN(n615) );
  NAND2_X1 U679 ( .A1(G953), .A2(G224), .ZN(n611) );
  XNOR2_X1 U680 ( .A(KEYINPUT61), .B(n611), .ZN(n612) );
  NAND2_X1 U681 ( .A1(n612), .A2(G898), .ZN(n613) );
  XOR2_X1 U682 ( .A(KEYINPUT124), .B(n613), .Z(n614) );
  NOR2_X1 U683 ( .A1(n615), .A2(n614), .ZN(n616) );
  XOR2_X1 U684 ( .A(n352), .B(n616), .Z(G69) );
  XNOR2_X1 U685 ( .A(G101), .B(n617), .ZN(n618) );
  XNOR2_X1 U686 ( .A(n618), .B(KEYINPUT109), .ZN(G3) );
  NOR2_X1 U687 ( .A1(n635), .A2(n621), .ZN(n619) );
  XOR2_X1 U688 ( .A(KEYINPUT110), .B(n619), .Z(n620) );
  XNOR2_X1 U689 ( .A(G104), .B(n620), .ZN(G6) );
  NOR2_X1 U690 ( .A1(n638), .A2(n621), .ZN(n626) );
  XOR2_X1 U691 ( .A(KEYINPUT27), .B(KEYINPUT112), .Z(n623) );
  XNOR2_X1 U692 ( .A(G107), .B(KEYINPUT111), .ZN(n622) );
  XNOR2_X1 U693 ( .A(n623), .B(n622), .ZN(n624) );
  XNOR2_X1 U694 ( .A(KEYINPUT26), .B(n624), .ZN(n625) );
  XNOR2_X1 U695 ( .A(n626), .B(n625), .ZN(G9) );
  XOR2_X1 U696 ( .A(G110), .B(n627), .Z(G12) );
  XOR2_X1 U697 ( .A(G128), .B(KEYINPUT29), .Z(n630) );
  NAND2_X1 U698 ( .A1(n633), .A2(n628), .ZN(n629) );
  XNOR2_X1 U699 ( .A(n630), .B(n629), .ZN(G30) );
  XOR2_X1 U700 ( .A(G143), .B(n631), .Z(G45) );
  NAND2_X1 U701 ( .A1(n633), .A2(n632), .ZN(n634) );
  XNOR2_X1 U702 ( .A(n634), .B(G146), .ZN(G48) );
  NOR2_X1 U703 ( .A1(n635), .A2(n637), .ZN(n636) );
  XOR2_X1 U704 ( .A(G113), .B(n636), .Z(G15) );
  NOR2_X1 U705 ( .A1(n638), .A2(n637), .ZN(n640) );
  XNOR2_X1 U706 ( .A(G116), .B(KEYINPUT113), .ZN(n639) );
  XNOR2_X1 U707 ( .A(n640), .B(n639), .ZN(G18) );
  XNOR2_X1 U708 ( .A(G125), .B(n641), .ZN(n642) );
  XNOR2_X1 U709 ( .A(n642), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U710 ( .A(KEYINPUT53), .B(KEYINPUT120), .Z(n693) );
  NAND2_X1 U711 ( .A1(n609), .A2(n643), .ZN(n645) );
  OR2_X1 U712 ( .A1(KEYINPUT2), .A2(KEYINPUT80), .ZN(n644) );
  NAND2_X1 U713 ( .A1(n645), .A2(n644), .ZN(n648) );
  NAND2_X1 U714 ( .A1(n646), .A2(KEYINPUT2), .ZN(n647) );
  NAND2_X1 U715 ( .A1(n648), .A2(n647), .ZN(n691) );
  INV_X1 U716 ( .A(n649), .ZN(n651) );
  NAND2_X1 U717 ( .A1(KEYINPUT80), .A2(KEYINPUT2), .ZN(n650) );
  NOR2_X1 U718 ( .A1(n651), .A2(n650), .ZN(n689) );
  NOR2_X1 U719 ( .A1(n670), .A2(n680), .ZN(n652) );
  XOR2_X1 U720 ( .A(KEYINPUT119), .B(n652), .Z(n653) );
  NOR2_X1 U721 ( .A1(G953), .A2(n653), .ZN(n687) );
  NAND2_X1 U722 ( .A1(n654), .A2(n493), .ZN(n655) );
  XNOR2_X1 U723 ( .A(n655), .B(KEYINPUT115), .ZN(n656) );
  XNOR2_X1 U724 ( .A(KEYINPUT49), .B(n656), .ZN(n661) );
  NAND2_X1 U725 ( .A1(n657), .A2(n543), .ZN(n658) );
  XNOR2_X1 U726 ( .A(n658), .B(KEYINPUT50), .ZN(n659) );
  XNOR2_X1 U727 ( .A(KEYINPUT116), .B(n659), .ZN(n660) );
  NAND2_X1 U728 ( .A1(n661), .A2(n660), .ZN(n662) );
  NOR2_X1 U729 ( .A1(n663), .A2(n662), .ZN(n664) );
  XNOR2_X1 U730 ( .A(KEYINPUT117), .B(n664), .ZN(n666) );
  NAND2_X1 U731 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X1 U732 ( .A(n667), .B(KEYINPUT51), .ZN(n668) );
  XNOR2_X1 U733 ( .A(n668), .B(KEYINPUT118), .ZN(n669) );
  NOR2_X1 U734 ( .A1(n670), .A2(n669), .ZN(n682) );
  NOR2_X1 U735 ( .A1(n672), .A2(n671), .ZN(n673) );
  NOR2_X1 U736 ( .A1(n674), .A2(n673), .ZN(n675) );
  NOR2_X1 U737 ( .A1(n676), .A2(n675), .ZN(n677) );
  NOR2_X1 U738 ( .A1(n678), .A2(n677), .ZN(n679) );
  NOR2_X1 U739 ( .A1(n680), .A2(n679), .ZN(n681) );
  NOR2_X1 U740 ( .A1(n682), .A2(n681), .ZN(n683) );
  XOR2_X1 U741 ( .A(KEYINPUT52), .B(n683), .Z(n685) );
  NAND2_X1 U742 ( .A1(n685), .A2(n684), .ZN(n686) );
  NAND2_X1 U743 ( .A1(n687), .A2(n686), .ZN(n688) );
  NOR2_X1 U744 ( .A1(n689), .A2(n688), .ZN(n690) );
  NAND2_X1 U745 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U746 ( .A(n693), .B(n692), .ZN(G75) );
  XOR2_X1 U747 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n696) );
  XNOR2_X1 U748 ( .A(n694), .B(KEYINPUT123), .ZN(n695) );
  XNOR2_X1 U749 ( .A(n696), .B(n695), .ZN(n698) );
  NAND2_X1 U750 ( .A1(n703), .A2(G469), .ZN(n697) );
  XOR2_X1 U751 ( .A(n698), .B(n697), .Z(n699) );
  NOR2_X1 U752 ( .A1(n707), .A2(n699), .ZN(G54) );
  NAND2_X1 U753 ( .A1(n703), .A2(G478), .ZN(n701) );
  XNOR2_X1 U754 ( .A(n701), .B(n700), .ZN(n702) );
  NOR2_X1 U755 ( .A1(n707), .A2(n702), .ZN(G63) );
  NAND2_X1 U756 ( .A1(n703), .A2(G217), .ZN(n704) );
  XNOR2_X1 U757 ( .A(n705), .B(n704), .ZN(n706) );
  NOR2_X1 U758 ( .A1(n707), .A2(n706), .ZN(G66) );
  XNOR2_X1 U759 ( .A(n709), .B(n708), .ZN(n714) );
  XNOR2_X1 U760 ( .A(n714), .B(n711), .ZN(n713) );
  NAND2_X1 U761 ( .A1(n713), .A2(n712), .ZN(n719) );
  XNOR2_X1 U762 ( .A(G227), .B(n714), .ZN(n715) );
  NAND2_X1 U763 ( .A1(n715), .A2(G900), .ZN(n716) );
  XNOR2_X1 U764 ( .A(KEYINPUT126), .B(n716), .ZN(n717) );
  NAND2_X1 U765 ( .A1(n717), .A2(G953), .ZN(n718) );
  NAND2_X1 U766 ( .A1(n719), .A2(n718), .ZN(G72) );
  XNOR2_X1 U767 ( .A(G134), .B(n720), .ZN(n721) );
  XNOR2_X1 U768 ( .A(n721), .B(KEYINPUT114), .ZN(G36) );
  XNOR2_X1 U769 ( .A(G122), .B(n722), .ZN(G24) );
  XOR2_X1 U770 ( .A(G140), .B(n723), .Z(G42) );
  XOR2_X1 U771 ( .A(n724), .B(G131), .Z(G33) );
  XOR2_X1 U772 ( .A(G137), .B(n725), .Z(G39) );
endmodule

