//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 1 1 1 0 1 1 0 1 0 0 1 1 0 1 0 0 0 1 1 0 0 0 1 0 0 1 0 0 1 1 1 0 1 1 1 1 0 0 0 0 1 0 0 1 1 0 1 1 0 0 1 0 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:00 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1263, new_n1264, new_n1265, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT64), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT0), .Z(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  OAI21_X1  g0012(.A(G50), .B1(G58), .B2(G68), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  AOI21_X1  g0014(.A(new_n209), .B1(new_n212), .B2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G68), .A2(G238), .B1(G107), .B2(G264), .ZN(new_n216));
  INV_X1    g0016(.A(G87), .ZN(new_n217));
  INV_X1    g0017(.A(G250), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(G58), .ZN(new_n220));
  INV_X1    g0020(.A(G232), .ZN(new_n221));
  INV_X1    g0021(.A(G97), .ZN(new_n222));
  INV_X1    g0022(.A(G257), .ZN(new_n223));
  OAI22_X1  g0023(.A1(new_n220), .A2(new_n221), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n219), .A2(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(G244), .ZN(new_n226));
  XNOR2_X1  g0026(.A(KEYINPUT66), .B(G77), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n225), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT65), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n206), .B1(new_n228), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n231), .A2(KEYINPUT1), .ZN(new_n232));
  OR2_X1    g0032(.A1(new_n231), .A2(KEYINPUT1), .ZN(new_n233));
  NAND3_X1  g0033(.A1(new_n215), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT67), .ZN(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(new_n221), .ZN(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT2), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G264), .B(G270), .Z(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n239), .B(new_n242), .Z(G358));
  XNOR2_X1  g0043(.A(G50), .B(G68), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G58), .B(G77), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n244), .B(new_n245), .Z(new_n246));
  XOR2_X1   g0046(.A(G87), .B(G97), .Z(new_n247));
  XOR2_X1   g0047(.A(G107), .B(G116), .Z(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(new_n246), .B(new_n249), .Z(G351));
  NAND2_X1  g0050(.A1(G33), .A2(G41), .ZN(new_n251));
  NAND4_X1  g0051(.A1(new_n251), .A2(KEYINPUT68), .A3(G1), .A4(G13), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  AND2_X1   g0053(.A1(G1), .A2(G13), .ZN(new_n254));
  AOI21_X1  g0054(.A(KEYINPUT68), .B1(new_n254), .B2(new_n251), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT69), .ZN(new_n257));
  INV_X1    g0057(.A(G1), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n258), .B1(G41), .B2(G45), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  NAND4_X1  g0060(.A1(new_n256), .A2(new_n257), .A3(G274), .A4(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT68), .ZN(new_n262));
  AND2_X1   g0062(.A1(G33), .A2(G41), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n262), .B1(new_n263), .B2(new_n210), .ZN(new_n264));
  NAND4_X1  g0064(.A1(new_n264), .A2(new_n260), .A3(G274), .A4(new_n252), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(KEYINPUT69), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n261), .A2(new_n266), .ZN(new_n267));
  AND3_X1   g0067(.A1(new_n264), .A2(new_n259), .A3(new_n252), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n254), .A2(new_n251), .ZN(new_n269));
  INV_X1    g0069(.A(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(KEYINPUT3), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT3), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n269), .B1(new_n274), .B2(new_n227), .ZN(new_n275));
  XNOR2_X1  g0075(.A(KEYINPUT3), .B(G33), .ZN(new_n276));
  NOR2_X1   g0076(.A1(G222), .A2(G1698), .ZN(new_n277));
  INV_X1    g0077(.A(G1698), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n278), .A2(G223), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n276), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  AOI22_X1  g0080(.A1(new_n268), .A2(G226), .B1(new_n275), .B2(new_n280), .ZN(new_n281));
  AND2_X1   g0081(.A1(new_n267), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G200), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n284), .B1(G190), .B2(new_n282), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT74), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT10), .ZN(new_n288));
  INV_X1    g0088(.A(new_n285), .ZN(new_n289));
  INV_X1    g0089(.A(G150), .ZN(new_n290));
  NOR2_X1   g0090(.A1(G20), .A2(G33), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  OAI22_X1  g0092(.A1(new_n290), .A2(new_n292), .B1(new_n201), .B2(new_n211), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n220), .A2(KEYINPUT8), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT8), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(G58), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT70), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  XNOR2_X1  g0099(.A(KEYINPUT8), .B(G58), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(KEYINPUT70), .ZN(new_n301));
  AND2_X1   g0101(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n270), .A2(G20), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n293), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND3_X1  g0104(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(new_n210), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n304), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(G50), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n309), .B1(new_n258), .B2(G20), .ZN(new_n310));
  XNOR2_X1  g0110(.A(new_n310), .B(KEYINPUT71), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n258), .A2(G13), .A3(G20), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n311), .A2(new_n307), .A3(new_n312), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n313), .B1(G50), .B2(new_n312), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n308), .A2(new_n314), .ZN(new_n315));
  XNOR2_X1  g0115(.A(new_n315), .B(KEYINPUT9), .ZN(new_n316));
  OAI211_X1 g0116(.A(new_n287), .B(new_n288), .C1(new_n289), .C2(new_n316), .ZN(new_n317));
  XOR2_X1   g0117(.A(new_n315), .B(KEYINPUT9), .Z(new_n318));
  OAI211_X1 g0118(.A(new_n318), .B(new_n285), .C1(new_n286), .C2(KEYINPUT10), .ZN(new_n319));
  INV_X1    g0119(.A(G179), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n282), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT72), .ZN(new_n322));
  XNOR2_X1  g0122(.A(new_n321), .B(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n315), .ZN(new_n324));
  OAI211_X1 g0124(.A(new_n323), .B(new_n324), .C1(G169), .C2(new_n282), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n317), .A2(new_n319), .A3(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT17), .ZN(new_n327));
  INV_X1    g0127(.A(new_n269), .ZN(new_n328));
  NAND2_X1  g0128(.A1(G33), .A2(G87), .ZN(new_n329));
  XNOR2_X1  g0129(.A(new_n329), .B(KEYINPUT79), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT76), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n331), .B1(new_n272), .B2(G33), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n270), .A2(KEYINPUT76), .A3(KEYINPUT3), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n332), .A2(new_n273), .A3(new_n333), .ZN(new_n334));
  OR2_X1    g0134(.A1(G223), .A2(G1698), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n335), .B1(G226), .B2(new_n278), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n330), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  AOI22_X1  g0137(.A1(new_n328), .A2(new_n337), .B1(new_n268), .B2(G232), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n267), .A2(new_n338), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n339), .A2(G190), .ZN(new_n340));
  AND2_X1   g0140(.A1(new_n265), .A2(KEYINPUT69), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n265), .A2(KEYINPUT69), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n337), .A2(new_n328), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n268), .A2(G232), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  OAI21_X1  g0146(.A(KEYINPUT80), .B1(new_n343), .B2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT80), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n267), .A2(new_n338), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n340), .B1(new_n350), .B2(new_n283), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n334), .A2(new_n211), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT7), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n353), .A2(KEYINPUT77), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  XNOR2_X1  g0155(.A(KEYINPUT77), .B(KEYINPUT7), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n334), .A2(new_n211), .A3(new_n356), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n355), .A2(G68), .A3(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(G68), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n220), .A2(new_n359), .ZN(new_n360));
  NOR2_X1   g0160(.A1(G58), .A2(G68), .ZN(new_n361));
  OAI21_X1  g0161(.A(G20), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n291), .A2(G159), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n358), .A2(KEYINPUT16), .A3(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT16), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n353), .B1(new_n276), .B2(G20), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n274), .A2(KEYINPUT7), .A3(new_n211), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n359), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n367), .B1(new_n370), .B2(new_n364), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n366), .A2(new_n306), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n299), .A2(new_n301), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(new_n312), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n307), .B1(G1), .B2(new_n211), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n375), .A2(new_n299), .A3(new_n301), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT78), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n374), .A2(new_n376), .A3(KEYINPUT78), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n372), .A2(new_n381), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n327), .B1(new_n351), .B2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(G169), .ZN(new_n384));
  AND3_X1   g0184(.A1(new_n267), .A2(new_n338), .A3(new_n348), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n348), .B1(new_n267), .B2(new_n338), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n384), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n339), .A2(G179), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n387), .A2(new_n382), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(KEYINPUT18), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT18), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n387), .A2(new_n382), .A3(new_n392), .A4(new_n389), .ZN(new_n393));
  AND2_X1   g0193(.A1(new_n372), .A2(new_n381), .ZN(new_n394));
  AOI21_X1  g0194(.A(G200), .B1(new_n347), .B2(new_n349), .ZN(new_n395));
  OAI211_X1 g0195(.A(new_n394), .B(KEYINPUT17), .C1(new_n395), .C2(new_n340), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n383), .A2(new_n391), .A3(new_n393), .A4(new_n396), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n375), .A2(new_n202), .ZN(new_n398));
  XOR2_X1   g0198(.A(new_n398), .B(KEYINPUT73), .Z(new_n399));
  INV_X1    g0199(.A(new_n227), .ZN(new_n400));
  XNOR2_X1  g0200(.A(KEYINPUT15), .B(G87), .ZN(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  AOI22_X1  g0202(.A1(new_n400), .A2(G20), .B1(new_n402), .B2(new_n303), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n403), .B1(new_n292), .B2(new_n300), .ZN(new_n404));
  INV_X1    g0204(.A(new_n312), .ZN(new_n405));
  AOI22_X1  g0205(.A1(new_n404), .A2(new_n306), .B1(new_n227), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n399), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n276), .A2(G238), .A3(G1698), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n276), .A2(G232), .A3(new_n278), .ZN(new_n409));
  INV_X1    g0209(.A(G107), .ZN(new_n410));
  OAI211_X1 g0210(.A(new_n408), .B(new_n409), .C1(new_n410), .C2(new_n276), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(new_n328), .ZN(new_n412));
  INV_X1    g0212(.A(new_n268), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n412), .B1(new_n413), .B2(new_n226), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n414), .A2(new_n343), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n407), .B1(new_n415), .B2(G190), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n416), .B1(new_n283), .B2(new_n415), .ZN(new_n417));
  INV_X1    g0217(.A(new_n415), .ZN(new_n418));
  AOI22_X1  g0218(.A1(new_n418), .A2(new_n384), .B1(new_n399), .B2(new_n406), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n415), .A2(new_n320), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n417), .A2(new_n421), .ZN(new_n422));
  OR3_X1    g0222(.A1(new_n326), .A2(new_n397), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n303), .A2(G77), .ZN(new_n424));
  OAI221_X1 g0224(.A(new_n424), .B1(new_n211), .B2(G68), .C1(new_n309), .C2(new_n292), .ZN(new_n425));
  AND3_X1   g0225(.A1(new_n425), .A2(KEYINPUT11), .A3(new_n306), .ZN(new_n426));
  AOI21_X1  g0226(.A(KEYINPUT11), .B1(new_n425), .B2(new_n306), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT12), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n428), .B1(new_n405), .B2(new_n359), .ZN(new_n429));
  NOR3_X1   g0229(.A1(new_n312), .A2(KEYINPUT12), .A3(G68), .ZN(new_n430));
  OAI22_X1  g0230(.A1(new_n375), .A2(new_n359), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NOR3_X1   g0231(.A1(new_n426), .A2(new_n427), .A3(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT14), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT13), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT75), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n436), .B1(new_n341), .B2(new_n342), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n261), .A2(KEYINPUT75), .A3(new_n266), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n264), .A2(G238), .A3(new_n259), .A4(new_n252), .ZN(new_n440));
  NOR2_X1   g0240(.A1(G226), .A2(G1698), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n441), .B1(new_n221), .B2(G1698), .ZN(new_n442));
  AOI22_X1  g0242(.A1(new_n442), .A2(new_n276), .B1(G33), .B2(G97), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n440), .B1(new_n443), .B2(new_n269), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n435), .B1(new_n439), .B2(new_n445), .ZN(new_n446));
  AOI211_X1 g0246(.A(KEYINPUT13), .B(new_n444), .C1(new_n437), .C2(new_n438), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n434), .B(G169), .C1(new_n446), .C2(new_n447), .ZN(new_n448));
  NOR3_X1   g0248(.A1(new_n341), .A2(new_n342), .A3(new_n436), .ZN(new_n449));
  AOI21_X1  g0249(.A(KEYINPUT75), .B1(new_n261), .B2(new_n266), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n445), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(KEYINPUT13), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n439), .A2(new_n435), .A3(new_n445), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n452), .A2(G179), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n448), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n452), .A2(new_n453), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n434), .B1(new_n456), .B2(G169), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n433), .B1(new_n455), .B2(new_n457), .ZN(new_n458));
  OAI21_X1  g0258(.A(G200), .B1(new_n446), .B2(new_n447), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n452), .A2(G190), .A3(new_n453), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n459), .A2(new_n460), .A3(new_n432), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n458), .A2(new_n461), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n423), .A2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT83), .ZN(new_n465));
  AND2_X1   g0265(.A1(KEYINPUT5), .A2(G41), .ZN(new_n466));
  NOR2_X1   g0266(.A1(KEYINPUT5), .A2(G41), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n258), .B(G45), .C1(new_n466), .C2(new_n467), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n256), .A2(new_n465), .A3(G257), .A4(new_n468), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n468), .A2(new_n264), .A3(G257), .A4(new_n252), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(KEYINPUT83), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n258), .A2(G45), .ZN(new_n472));
  OR2_X1    g0272(.A1(KEYINPUT5), .A2(G41), .ZN(new_n473));
  NAND2_X1  g0273(.A1(KEYINPUT5), .A2(G41), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n472), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n475), .A2(G274), .A3(new_n264), .A4(new_n252), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n469), .A2(new_n471), .A3(new_n476), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n271), .A2(new_n273), .A3(G250), .A4(G1698), .ZN(new_n478));
  AND2_X1   g0278(.A1(KEYINPUT4), .A2(G244), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n271), .A2(new_n273), .A3(new_n479), .A4(new_n278), .ZN(new_n480));
  NAND2_X1  g0280(.A1(G33), .A2(G283), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n478), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n226), .A2(G1698), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n332), .A2(new_n333), .A3(new_n484), .A4(new_n273), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT4), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n269), .B1(new_n483), .B2(new_n487), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n384), .B1(new_n477), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n291), .A2(G77), .ZN(new_n490));
  NAND2_X1  g0290(.A1(KEYINPUT6), .A2(G97), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n491), .A2(G107), .ZN(new_n492));
  XNOR2_X1  g0292(.A(G97), .B(G107), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT6), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n490), .B1(new_n495), .B2(new_n211), .ZN(new_n496));
  AOI21_X1  g0296(.A(KEYINPUT7), .B1(new_n274), .B2(new_n211), .ZN(new_n497));
  AOI211_X1 g0297(.A(new_n353), .B(G20), .C1(new_n271), .C2(new_n273), .ZN(new_n498));
  OAI21_X1  g0298(.A(G107), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n496), .B1(new_n499), .B2(KEYINPUT81), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n410), .B1(new_n368), .B2(new_n369), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT81), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n307), .B1(new_n500), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n405), .A2(new_n222), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n258), .A2(G33), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n307), .A2(new_n312), .A3(new_n506), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n505), .B1(new_n507), .B2(new_n222), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n489), .B1(new_n504), .B2(new_n508), .ZN(new_n509));
  AND2_X1   g0309(.A1(new_n485), .A2(new_n486), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n328), .B1(new_n510), .B2(new_n482), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(KEYINPUT82), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT82), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n513), .B(new_n328), .C1(new_n510), .C2(new_n482), .ZN(new_n514));
  AOI211_X1 g0314(.A(G179), .B(new_n477), .C1(new_n512), .C2(new_n514), .ZN(new_n515));
  OAI21_X1  g0315(.A(KEYINPUT84), .B1(new_n509), .B2(new_n515), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n504), .A2(new_n508), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n477), .A2(new_n488), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(G190), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n477), .B1(new_n512), .B2(new_n514), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n517), .B(new_n519), .C1(new_n283), .C2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n512), .A2(new_n514), .ZN(new_n522));
  INV_X1    g0322(.A(new_n477), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n522), .A2(new_n320), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n493), .A2(new_n494), .ZN(new_n525));
  INV_X1    g0325(.A(new_n492), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(G20), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n490), .B(new_n528), .C1(new_n501), .C2(new_n502), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n499), .A2(KEYINPUT81), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n306), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(new_n508), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT84), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n524), .A2(new_n533), .A3(new_n534), .A4(new_n489), .ZN(new_n535));
  AND3_X1   g0335(.A1(new_n516), .A2(new_n521), .A3(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT22), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n211), .A2(G87), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n537), .B1(new_n274), .B2(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT23), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n540), .B1(new_n211), .B2(G107), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n410), .A2(KEYINPUT23), .A3(G20), .ZN(new_n542));
  AND2_X1   g0342(.A1(G33), .A2(G116), .ZN(new_n543));
  AOI22_X1  g0343(.A1(new_n541), .A2(new_n542), .B1(new_n211), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n539), .A2(new_n544), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n332), .A2(new_n333), .A3(new_n211), .A4(new_n273), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n537), .A2(new_n217), .ZN(new_n547));
  INV_X1    g0347(.A(new_n547), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  OAI21_X1  g0349(.A(KEYINPUT24), .B1(new_n545), .B2(new_n549), .ZN(new_n550));
  AND3_X1   g0350(.A1(new_n332), .A2(new_n273), .A3(new_n333), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n551), .A2(new_n211), .A3(new_n547), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT24), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n552), .A2(new_n553), .A3(new_n539), .A4(new_n544), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n550), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(new_n306), .ZN(new_n556));
  INV_X1    g0356(.A(new_n507), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT25), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n558), .B1(new_n312), .B2(G107), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n405), .A2(KEYINPUT25), .A3(new_n410), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n557), .A2(G107), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n468), .A2(new_n264), .A3(new_n252), .ZN(new_n562));
  INV_X1    g0362(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n223), .A2(G1698), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n564), .B1(G250), .B2(G1698), .ZN(new_n565));
  INV_X1    g0365(.A(G294), .ZN(new_n566));
  OAI22_X1  g0366(.A1(new_n334), .A2(new_n565), .B1(new_n270), .B2(new_n566), .ZN(new_n567));
  AOI22_X1  g0367(.A1(new_n563), .A2(G264), .B1(new_n567), .B2(new_n328), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n568), .A2(G190), .A3(new_n476), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n567), .A2(new_n328), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n256), .A2(G264), .A3(new_n468), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n570), .A2(new_n476), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(G200), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n556), .A2(new_n561), .A3(new_n569), .A4(new_n573), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n307), .B1(new_n550), .B2(new_n554), .ZN(new_n575));
  INV_X1    g0375(.A(new_n561), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n570), .A2(new_n571), .A3(G179), .A4(new_n476), .ZN(new_n577));
  OAI22_X1  g0377(.A1(new_n575), .A2(new_n576), .B1(KEYINPUT91), .B2(new_n577), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n384), .B1(new_n568), .B2(new_n476), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n577), .A2(KEYINPUT91), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n574), .B1(new_n578), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(KEYINPUT92), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT92), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n574), .B(new_n584), .C1(new_n581), .C2(new_n578), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(G270), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n476), .B1(new_n562), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n223), .A2(new_n278), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n589), .B1(G264), .B2(new_n278), .ZN(new_n590));
  XNOR2_X1  g0390(.A(KEYINPUT88), .B(G303), .ZN(new_n591));
  OAI22_X1  g0391(.A1(new_n334), .A2(new_n590), .B1(new_n276), .B2(new_n591), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n588), .B1(new_n328), .B2(new_n592), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n593), .A2(new_n384), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT90), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n312), .A2(G116), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(G116), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n597), .B1(new_n507), .B2(new_n598), .ZN(new_n599));
  AOI22_X1  g0399(.A1(new_n305), .A2(new_n210), .B1(G20), .B2(new_n598), .ZN(new_n600));
  AOI21_X1  g0400(.A(G20), .B1(G33), .B2(G283), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n270), .A2(G97), .ZN(new_n602));
  AND3_X1   g0402(.A1(new_n601), .A2(new_n602), .A3(KEYINPUT89), .ZN(new_n603));
  AOI21_X1  g0403(.A(KEYINPUT89), .B1(new_n601), .B2(new_n602), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n600), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT20), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  OAI211_X1 g0407(.A(KEYINPUT20), .B(new_n600), .C1(new_n603), .C2(new_n604), .ZN(new_n608));
  AOI211_X1 g0408(.A(new_n595), .B(new_n599), .C1(new_n607), .C2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n607), .A2(new_n608), .ZN(new_n610));
  INV_X1    g0410(.A(new_n599), .ZN(new_n611));
  AOI21_X1  g0411(.A(KEYINPUT90), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n594), .B1(new_n609), .B2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT21), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n592), .A2(new_n328), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n616), .B(new_n476), .C1(new_n587), .C2(new_n562), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n617), .A2(new_n320), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n618), .B1(new_n609), .B2(new_n612), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n594), .B(KEYINPUT21), .C1(new_n612), .C2(new_n609), .ZN(new_n620));
  INV_X1    g0420(.A(new_n609), .ZN(new_n621));
  INV_X1    g0421(.A(new_n612), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n617), .A2(G200), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n593), .A2(G190), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n621), .A2(new_n622), .A3(new_n623), .A4(new_n624), .ZN(new_n625));
  AND4_X1   g0425(.A1(new_n615), .A2(new_n619), .A3(new_n620), .A4(new_n625), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n402), .A2(new_n312), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n551), .A2(KEYINPUT86), .A3(new_n211), .A4(G68), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT86), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n629), .B1(new_n546), .B2(new_n359), .ZN(new_n630));
  AOI21_X1  g0430(.A(G20), .B1(G33), .B2(G97), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT19), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(KEYINPUT85), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT85), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(KEYINPUT19), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n631), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n217), .A2(new_n222), .A3(new_n410), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n303), .A2(G97), .ZN(new_n638));
  XNOR2_X1  g0438(.A(KEYINPUT85), .B(KEYINPUT19), .ZN(new_n639));
  AOI22_X1  g0439(.A1(new_n636), .A2(new_n637), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n628), .A2(new_n630), .A3(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n627), .B1(new_n641), .B2(new_n306), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n557), .A2(G87), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n226), .A2(G1698), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n645), .B1(G238), .B2(G1698), .ZN(new_n646));
  OAI22_X1  g0446(.A1(new_n334), .A2(new_n646), .B1(new_n270), .B2(new_n598), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(new_n328), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n472), .A2(G274), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n649), .B1(new_n218), .B2(new_n472), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(new_n256), .ZN(new_n651));
  AOI21_X1  g0451(.A(G200), .B1(new_n648), .B2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(G190), .ZN(new_n653));
  AOI22_X1  g0453(.A1(new_n647), .A2(new_n328), .B1(new_n650), .B2(new_n256), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n652), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n507), .A2(new_n401), .ZN(new_n656));
  AOI211_X1 g0456(.A(new_n627), .B(new_n656), .C1(new_n641), .C2(new_n306), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n654), .A2(new_n320), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n658), .B1(new_n654), .B2(G169), .ZN(new_n659));
  OAI22_X1  g0459(.A1(new_n644), .A2(new_n655), .B1(new_n657), .B2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT87), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  AOI21_X1  g0462(.A(G169), .B1(new_n648), .B2(new_n651), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n663), .B1(new_n320), .B2(new_n654), .ZN(new_n664));
  INV_X1    g0464(.A(new_n656), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n642), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n648), .A2(new_n651), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n668), .A2(G190), .ZN(new_n669));
  OAI211_X1 g0469(.A(new_n642), .B(new_n643), .C1(new_n669), .C2(new_n652), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n667), .A2(KEYINPUT87), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n662), .A2(new_n671), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n536), .A2(new_n586), .A3(new_n626), .A4(new_n672), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n464), .A2(new_n673), .ZN(G372));
  NAND2_X1  g0474(.A1(new_n383), .A2(new_n396), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n461), .A2(new_n420), .A3(new_n419), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n675), .B1(new_n458), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n391), .A2(new_n393), .ZN(new_n678));
  OAI211_X1 g0478(.A(new_n319), .B(new_n317), .C1(new_n677), .C2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT93), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT26), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n516), .A2(new_n535), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n681), .B1(new_n672), .B2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n660), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n509), .A2(new_n515), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n667), .B1(new_n686), .B2(KEYINPUT26), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n680), .B1(new_n683), .B2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n667), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n524), .A2(new_n533), .A3(new_n489), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n690), .A2(new_n660), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n689), .B1(new_n691), .B2(new_n681), .ZN(new_n692));
  AOI22_X1  g0492(.A1(new_n662), .A2(new_n671), .B1(new_n516), .B2(new_n535), .ZN(new_n693));
  OAI211_X1 g0493(.A(new_n692), .B(KEYINPUT93), .C1(new_n693), .C2(new_n681), .ZN(new_n694));
  OR2_X1    g0494(.A1(new_n578), .A2(new_n581), .ZN(new_n695));
  AND4_X1   g0495(.A1(new_n695), .A2(new_n615), .A3(new_n619), .A4(new_n620), .ZN(new_n696));
  AND3_X1   g0496(.A1(new_n667), .A2(new_n574), .A3(new_n670), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n697), .A2(new_n516), .A3(new_n535), .A4(new_n521), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n688), .A2(new_n694), .A3(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  OAI211_X1 g0502(.A(new_n325), .B(new_n679), .C1(new_n464), .C2(new_n702), .ZN(G369));
  INV_X1    g0503(.A(G13), .ZN(new_n704));
  NOR3_X1   g0504(.A1(new_n704), .A2(G1), .A3(G20), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT27), .ZN(new_n707));
  OAI21_X1  g0507(.A(KEYINPUT94), .B1(new_n705), .B2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NOR3_X1   g0509(.A1(new_n705), .A2(KEYINPUT94), .A3(new_n707), .ZN(new_n710));
  OAI221_X1 g0510(.A(G213), .B1(KEYINPUT27), .B2(new_n706), .C1(new_n709), .C2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(G343), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n713), .B1(new_n609), .B2(new_n612), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n626), .A2(new_n714), .ZN(new_n715));
  AND2_X1   g0515(.A1(new_n620), .A2(new_n619), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(new_n615), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n715), .B1(new_n718), .B2(new_n714), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(G330), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n713), .B1(new_n575), .B2(new_n576), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n586), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n713), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n722), .B1(new_n695), .B2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n720), .A2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n586), .A2(new_n717), .A3(new_n723), .ZN(new_n728));
  INV_X1    g0528(.A(new_n695), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(new_n723), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n727), .A2(new_n732), .ZN(G399));
  INV_X1    g0533(.A(new_n207), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n734), .A2(G41), .ZN(new_n735));
  NOR4_X1   g0535(.A1(new_n735), .A2(new_n258), .A3(G116), .A4(new_n637), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n736), .B1(new_n214), .B2(new_n735), .ZN(new_n737));
  XOR2_X1   g0537(.A(new_n737), .B(KEYINPUT28), .Z(new_n738));
  OAI221_X1 g0538(.A(new_n667), .B1(new_n681), .B2(new_n691), .C1(new_n696), .C2(new_n698), .ZN(new_n739));
  AND2_X1   g0539(.A1(new_n693), .A2(new_n681), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n723), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(KEYINPUT29), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT29), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n701), .A2(new_n743), .A3(new_n723), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n617), .A2(new_n320), .A3(new_n668), .A4(new_n572), .ZN(new_n745));
  OR2_X1    g0545(.A1(new_n520), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(KEYINPUT30), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n593), .A2(G179), .A3(new_n654), .A4(new_n568), .ZN(new_n748));
  INV_X1    g0548(.A(new_n518), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n747), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  AND2_X1   g0550(.A1(new_n568), .A2(new_n654), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n618), .A2(new_n751), .A3(KEYINPUT30), .A4(new_n518), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n746), .A2(new_n750), .A3(new_n752), .ZN(new_n753));
  AND3_X1   g0553(.A1(new_n753), .A2(KEYINPUT31), .A3(new_n713), .ZN(new_n754));
  AOI21_X1  g0554(.A(KEYINPUT31), .B1(new_n753), .B2(new_n713), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n756), .B1(new_n673), .B2(new_n713), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(G330), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n742), .A2(new_n744), .A3(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n738), .B1(new_n760), .B2(G1), .ZN(G364));
  NOR2_X1   g0561(.A1(new_n704), .A2(G20), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n258), .B1(new_n762), .B2(G45), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n735), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n207), .A2(new_n276), .ZN(new_n766));
  INV_X1    g0566(.A(G355), .ZN(new_n767));
  OAI22_X1  g0567(.A1(new_n766), .A2(new_n767), .B1(G116), .B2(new_n207), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n734), .A2(new_n551), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(G45), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n770), .B1(new_n771), .B2(new_n214), .ZN(new_n772));
  OR2_X1    g0572(.A1(new_n246), .A2(new_n771), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n768), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(G13), .A2(G33), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(G20), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n210), .B1(G20), .B2(new_n384), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n765), .B1(new_n774), .B2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(KEYINPUT95), .ZN(new_n782));
  AND2_X1   g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n211), .A2(G190), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NOR3_X1   g0585(.A1(new_n785), .A2(G179), .A3(new_n283), .ZN(new_n786));
  XNOR2_X1  g0586(.A(new_n786), .B(KEYINPUT97), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(G283), .ZN(new_n788));
  NOR2_X1   g0588(.A1(G179), .A2(G200), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n211), .B1(new_n789), .B2(G190), .ZN(new_n790));
  OR2_X1    g0590(.A1(new_n790), .A2(KEYINPUT98), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n790), .A2(KEYINPUT98), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(G294), .ZN(new_n795));
  NAND3_X1  g0595(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(G190), .ZN(new_n797));
  INV_X1    g0597(.A(G317), .ZN(new_n798));
  OR2_X1    g0598(.A1(new_n798), .A2(KEYINPUT33), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n798), .A2(KEYINPUT33), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n797), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(G311), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n320), .A2(G200), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n803), .A2(new_n784), .ZN(new_n804));
  OAI211_X1 g0604(.A(new_n801), .B(new_n274), .C1(new_n802), .C2(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n796), .A2(new_n653), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n805), .B1(G326), .B2(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n211), .A2(new_n653), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n808), .A2(new_n803), .ZN(new_n809));
  INV_X1    g0609(.A(G322), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n784), .A2(new_n789), .ZN(new_n811));
  INV_X1    g0611(.A(G329), .ZN(new_n812));
  OAI22_X1  g0612(.A1(new_n809), .A2(new_n810), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n808), .A2(new_n320), .A3(G200), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n813), .B1(G303), .B2(new_n815), .ZN(new_n816));
  NAND4_X1  g0616(.A1(new_n788), .A2(new_n795), .A3(new_n807), .A4(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(G159), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n811), .A2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n820), .A2(KEYINPUT32), .ZN(new_n821));
  AOI211_X1 g0621(.A(new_n274), .B(new_n821), .C1(G87), .C2(new_n815), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n794), .A2(G97), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n787), .A2(G107), .ZN(new_n824));
  AOI22_X1  g0624(.A1(new_n820), .A2(KEYINPUT32), .B1(new_n797), .B2(G68), .ZN(new_n825));
  NAND4_X1  g0625(.A1(new_n822), .A2(new_n823), .A3(new_n824), .A4(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n809), .ZN(new_n827));
  INV_X1    g0627(.A(new_n804), .ZN(new_n828));
  AOI22_X1  g0628(.A1(new_n827), .A2(G58), .B1(new_n828), .B2(new_n400), .ZN(new_n829));
  INV_X1    g0629(.A(new_n806), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n829), .B1(new_n309), .B2(new_n830), .ZN(new_n831));
  XOR2_X1   g0631(.A(new_n831), .B(KEYINPUT96), .Z(new_n832));
  OAI21_X1  g0632(.A(new_n817), .B1(new_n826), .B2(new_n832), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n783), .B1(new_n778), .B2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n777), .ZN(new_n835));
  OAI221_X1 g0635(.A(new_n834), .B1(new_n782), .B2(new_n781), .C1(new_n719), .C2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n765), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n720), .A2(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n719), .A2(G330), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n836), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  XOR2_X1   g0640(.A(new_n840), .B(KEYINPUT99), .Z(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(G396));
  NOR2_X1   g0642(.A1(new_n421), .A2(new_n713), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n407), .A2(new_n713), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n417), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n843), .B1(new_n845), .B2(new_n421), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n846), .B1(new_n701), .B2(new_n723), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n417), .A2(new_n421), .A3(new_n723), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n692), .B1(new_n693), .B2(new_n681), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n699), .B1(new_n849), .B2(new_n680), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n848), .B1(new_n850), .B2(new_n694), .ZN(new_n851));
  OR2_X1    g0651(.A1(new_n847), .A2(new_n851), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n765), .B1(new_n852), .B2(new_n758), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n853), .B1(new_n758), .B2(new_n852), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n778), .A2(new_n775), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n837), .B1(new_n202), .B2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n778), .ZN(new_n857));
  INV_X1    g0657(.A(new_n797), .ZN(new_n858));
  INV_X1    g0658(.A(G283), .ZN(new_n859));
  OAI221_X1 g0659(.A(new_n274), .B1(new_n811), .B2(new_n802), .C1(new_n858), .C2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n787), .A2(G87), .ZN(new_n861));
  OAI22_X1  g0661(.A1(new_n814), .A2(new_n410), .B1(new_n809), .B2(new_n566), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n862), .B1(G116), .B2(new_n828), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  AOI211_X1 g0664(.A(new_n860), .B(new_n864), .C1(G303), .C2(new_n806), .ZN(new_n865));
  AOI22_X1  g0665(.A1(G143), .A2(new_n827), .B1(new_n828), .B2(G159), .ZN(new_n866));
  INV_X1    g0666(.A(G137), .ZN(new_n867));
  OAI221_X1 g0667(.A(new_n866), .B1(new_n830), .B2(new_n867), .C1(new_n290), .C2(new_n858), .ZN(new_n868));
  XNOR2_X1  g0668(.A(KEYINPUT100), .B(KEYINPUT34), .ZN(new_n869));
  OR2_X1    g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n787), .A2(G68), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n794), .A2(G58), .ZN(new_n872));
  INV_X1    g0672(.A(new_n811), .ZN(new_n873));
  AOI22_X1  g0673(.A1(new_n815), .A2(G50), .B1(new_n873), .B2(G132), .ZN(new_n874));
  NAND4_X1  g0674(.A1(new_n871), .A2(new_n551), .A3(new_n872), .A4(new_n874), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n875), .B1(new_n868), .B2(new_n869), .ZN(new_n876));
  AOI22_X1  g0676(.A1(new_n865), .A2(new_n823), .B1(new_n870), .B2(new_n876), .ZN(new_n877));
  OAI221_X1 g0677(.A(new_n856), .B1(new_n857), .B2(new_n877), .C1(new_n846), .C2(new_n776), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n854), .A2(new_n878), .ZN(G384));
  OR2_X1    g0679(.A1(new_n527), .A2(KEYINPUT35), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n527), .A2(KEYINPUT35), .ZN(new_n881));
  NAND4_X1  g0681(.A1(new_n880), .A2(G116), .A3(new_n212), .A4(new_n881), .ZN(new_n882));
  XOR2_X1   g0682(.A(new_n882), .B(KEYINPUT36), .Z(new_n883));
  OR3_X1    g0683(.A1(new_n227), .A2(new_n213), .A3(new_n360), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n309), .A2(G68), .ZN(new_n885));
  AOI211_X1 g0685(.A(new_n258), .B(G13), .C1(new_n884), .C2(new_n885), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n883), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n366), .A2(new_n306), .ZN(new_n888));
  AOI21_X1  g0688(.A(KEYINPUT16), .B1(new_n358), .B2(new_n365), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n377), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n711), .ZN(new_n891));
  AND2_X1   g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n397), .A2(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n394), .B1(new_n395), .B2(new_n340), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT37), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n382), .A2(new_n891), .ZN(new_n896));
  NAND4_X1  g0696(.A1(new_n894), .A2(new_n895), .A3(new_n390), .A4(new_n896), .ZN(new_n897));
  AOI21_X1  g0697(.A(G169), .B1(new_n347), .B2(new_n349), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n711), .B1(new_n898), .B2(new_n388), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n283), .B1(new_n385), .B2(new_n386), .ZN(new_n900));
  INV_X1    g0700(.A(new_n340), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  AOI22_X1  g0702(.A1(new_n899), .A2(new_n890), .B1(new_n902), .B2(new_n394), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n897), .B1(new_n903), .B2(new_n895), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n893), .A2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT38), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n893), .A2(KEYINPUT38), .A3(new_n904), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  OAI21_X1  g0709(.A(G169), .B1(new_n446), .B2(new_n447), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(KEYINPUT14), .ZN(new_n911));
  NAND4_X1  g0711(.A1(new_n461), .A2(new_n911), .A3(new_n454), .A4(new_n448), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n723), .A2(new_n432), .ZN(new_n913));
  AOI21_X1  g0713(.A(KEYINPUT102), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(new_n913), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n458), .A2(new_n461), .A3(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n912), .A2(KEYINPUT102), .A3(new_n913), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n915), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n843), .B(KEYINPUT101), .ZN(new_n920));
  OAI211_X1 g0720(.A(new_n909), .B(new_n919), .C1(new_n851), .C2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n678), .A2(new_n711), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(KEYINPUT103), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT103), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n921), .A2(new_n925), .A3(new_n922), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT39), .ZN(new_n927));
  AND3_X1   g0727(.A1(new_n893), .A2(KEYINPUT38), .A3(new_n904), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n894), .A2(new_n390), .A3(new_n896), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(KEYINPUT37), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n897), .ZN(new_n931));
  INV_X1    g0731(.A(new_n896), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n397), .A2(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(KEYINPUT38), .B1(new_n931), .B2(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n927), .B1(new_n928), .B2(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n907), .A2(KEYINPUT39), .A3(new_n908), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  OR2_X1    g0737(.A1(new_n458), .A2(new_n713), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(new_n939), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n924), .A2(new_n926), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n679), .A2(new_n325), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n742), .A2(new_n744), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n942), .B1(new_n943), .B2(new_n463), .ZN(new_n944));
  XOR2_X1   g0744(.A(new_n941), .B(new_n944), .Z(new_n945));
  NAND2_X1  g0745(.A1(new_n917), .A2(new_n918), .ZN(new_n946));
  OAI211_X1 g0746(.A(new_n757), .B(new_n846), .C1(new_n946), .C2(new_n914), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT40), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT104), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(new_n928), .B2(new_n934), .ZN(new_n951));
  AND2_X1   g0751(.A1(new_n931), .A2(new_n933), .ZN(new_n952));
  OAI211_X1 g0752(.A(new_n908), .B(KEYINPUT104), .C1(new_n952), .C2(KEYINPUT38), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n949), .A2(new_n951), .A3(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(KEYINPUT38), .B1(new_n893), .B2(new_n904), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n928), .A2(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n948), .B1(new_n947), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n954), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n463), .A2(new_n757), .ZN(new_n959));
  OR2_X1    g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n958), .A2(new_n959), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n960), .A2(G330), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n945), .A2(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n963), .B1(new_n258), .B2(new_n762), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n945), .A2(new_n962), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n887), .B1(new_n964), .B2(new_n965), .ZN(G367));
  NAND2_X1  g0766(.A1(new_n644), .A2(new_n713), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n684), .A2(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n667), .B2(new_n967), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(KEYINPUT43), .ZN(new_n970));
  XOR2_X1   g0770(.A(new_n970), .B(KEYINPUT105), .Z(new_n971));
  OAI21_X1  g0771(.A(new_n536), .B1(new_n517), .B2(new_n723), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n685), .A2(new_n713), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n728), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(KEYINPUT42), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n682), .B1(new_n974), .B2(new_n729), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n978), .A2(new_n713), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n971), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  OR2_X1    g0780(.A1(new_n969), .A2(KEYINPUT43), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(KEYINPUT106), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n726), .A2(new_n974), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n983), .A2(new_n984), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n981), .A2(KEYINPUT106), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n988), .B(new_n989), .ZN(new_n990));
  XOR2_X1   g0790(.A(new_n735), .B(KEYINPUT41), .Z(new_n991));
  OAI21_X1  g0791(.A(new_n725), .B1(new_n718), .B2(new_n713), .ZN(new_n992));
  OR2_X1    g0792(.A1(new_n728), .A2(KEYINPUT107), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n728), .A2(KEYINPUT107), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n992), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(new_n720), .ZN(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(new_n760), .ZN(new_n998));
  INV_X1    g0798(.A(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(new_n974), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n1000), .A2(new_n731), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1001), .B(KEYINPUT45), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n732), .A2(new_n974), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT44), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1005), .B(new_n727), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n999), .A2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n991), .B1(new_n1007), .B2(new_n760), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n990), .B1(new_n764), .B2(new_n1008), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n779), .B1(new_n207), .B2(new_n401), .C1(new_n770), .C2(new_n242), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n276), .B1(new_n811), .B2(new_n867), .C1(new_n858), .C2(new_n818), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n1011), .B1(G143), .B2(new_n806), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n794), .A2(G68), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n400), .A2(new_n786), .B1(new_n815), .B2(G58), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(G150), .A2(new_n827), .B1(new_n828), .B2(G50), .ZN(new_n1015));
  NAND4_X1  g0815(.A1(new_n1012), .A2(new_n1013), .A3(new_n1014), .A4(new_n1015), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n814), .A2(new_n598), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1017), .B(KEYINPUT46), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1018), .B1(G294), .B2(new_n797), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n804), .A2(new_n859), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n809), .A2(new_n591), .B1(new_n811), .B2(new_n798), .ZN(new_n1021));
  AOI211_X1 g0821(.A(new_n1020), .B(new_n1021), .C1(G97), .C2(new_n786), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n551), .B1(new_n806), .B2(G311), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1019), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n793), .A2(new_n410), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1016), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  XOR2_X1   g0826(.A(new_n1026), .B(KEYINPUT47), .Z(new_n1027));
  OAI211_X1 g0827(.A(new_n765), .B(new_n1010), .C1(new_n1027), .C2(new_n857), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(KEYINPUT108), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(new_n835), .B2(new_n969), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1009), .A2(new_n1030), .ZN(G387));
  NOR2_X1   g0831(.A1(new_n724), .A2(new_n835), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n637), .A2(G116), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n766), .A2(new_n1033), .B1(G107), .B2(new_n207), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n239), .A2(G45), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n1035), .B(KEYINPUT109), .ZN(new_n1036));
  OAI211_X1 g0836(.A(new_n1033), .B(new_n771), .C1(new_n359), .C2(new_n202), .ZN(new_n1037));
  XOR2_X1   g0837(.A(KEYINPUT110), .B(KEYINPUT50), .Z(new_n1038));
  NOR3_X1   g0838(.A1(new_n1038), .A2(G50), .A3(new_n300), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1038), .B1(G50), .B2(new_n300), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n770), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1034), .B1(new_n1036), .B2(new_n1042), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n765), .B1(new_n1043), .B2(new_n780), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n787), .A2(G97), .B1(new_n302), .B2(new_n797), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n815), .A2(new_n400), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1046), .B1(new_n309), .B2(new_n809), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n804), .A2(new_n359), .B1(new_n811), .B2(new_n290), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n551), .B1(new_n830), .B2(new_n818), .ZN(new_n1049));
  NOR3_X1   g0849(.A1(new_n1047), .A2(new_n1048), .A3(new_n1049), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n794), .A2(new_n402), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1045), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n591), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n827), .A2(G317), .B1(new_n828), .B2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1054), .B1(new_n810), .B2(new_n830), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1055), .B1(G311), .B2(new_n797), .ZN(new_n1056));
  OR2_X1    g0856(.A1(new_n1056), .A2(KEYINPUT48), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1056), .A2(KEYINPUT48), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n794), .A2(G283), .B1(G294), .B2(new_n815), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1057), .A2(new_n1058), .A3(new_n1059), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT111), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1061), .A2(KEYINPUT49), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n786), .A2(G116), .B1(G326), .B2(new_n873), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1062), .A2(new_n334), .A3(new_n1063), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n1061), .A2(KEYINPUT49), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1052), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  AOI211_X1 g0866(.A(new_n1032), .B(new_n1044), .C1(new_n1066), .C2(new_n778), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1067), .B1(new_n997), .B2(new_n764), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n998), .A2(new_n735), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n997), .A2(new_n760), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1068), .B1(new_n1069), .B2(new_n1070), .ZN(G393));
  INV_X1    g0871(.A(new_n735), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1072), .B1(new_n999), .B2(new_n1006), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1073), .B1(new_n999), .B2(new_n1006), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1000), .A2(new_n777), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(new_n1075), .B(KEYINPUT112), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n794), .A2(G116), .B1(new_n1053), .B2(new_n797), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1077), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n1078), .A2(KEYINPUT113), .B1(G294), .B2(new_n828), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1079), .B1(KEYINPUT113), .B2(new_n1078), .ZN(new_n1080));
  XOR2_X1   g0880(.A(new_n1080), .B(KEYINPUT114), .Z(new_n1081));
  INV_X1    g0881(.A(new_n824), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n827), .A2(G311), .B1(G317), .B2(new_n806), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(new_n1083), .B(KEYINPUT52), .ZN(new_n1084));
  OAI221_X1 g0884(.A(new_n274), .B1(new_n811), .B2(new_n810), .C1(new_n814), .C2(new_n859), .ZN(new_n1085));
  NOR4_X1   g0885(.A1(new_n1081), .A2(new_n1082), .A3(new_n1084), .A4(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n828), .A2(new_n297), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n815), .A2(G68), .B1(new_n873), .B2(G143), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n334), .B1(new_n797), .B2(G50), .ZN(new_n1089));
  NAND4_X1  g0889(.A1(new_n861), .A2(new_n1087), .A3(new_n1088), .A4(new_n1089), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n830), .A2(new_n290), .B1(new_n809), .B2(new_n818), .ZN(new_n1091));
  INV_X1    g0891(.A(KEYINPUT51), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n794), .A2(G77), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NOR3_X1   g0896(.A1(new_n1090), .A2(new_n1093), .A3(new_n1096), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n778), .B1(new_n1086), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n769), .A2(new_n249), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n780), .B1(new_n734), .B2(G97), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n837), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  AND3_X1   g0901(.A1(new_n1076), .A2(new_n1098), .A3(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1102), .B1(new_n1006), .B2(new_n764), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1074), .A2(new_n1103), .ZN(new_n1104));
  OR2_X1    g0904(.A1(new_n1104), .A2(KEYINPUT115), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1104), .A2(KEYINPUT115), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1105), .A2(new_n1106), .ZN(G390));
  INV_X1    g0907(.A(new_n846), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n758), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1109), .A2(new_n919), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n848), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n920), .B1(new_n701), .B2(new_n1111), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n946), .A2(new_n914), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n938), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(KEYINPUT116), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  OAI211_X1 g0916(.A(KEYINPUT116), .B(new_n938), .C1(new_n1112), .C2(new_n1113), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1116), .A2(new_n937), .A3(new_n1117), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n723), .B(new_n846), .C1(new_n739), .C2(new_n740), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1119), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n919), .B1(new_n1120), .B2(new_n920), .ZN(new_n1121));
  NAND4_X1  g0921(.A1(new_n1121), .A2(new_n938), .A3(new_n951), .A4(new_n953), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1110), .B1(new_n1118), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1118), .A2(new_n1110), .A3(new_n1122), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n1120), .A2(new_n920), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1113), .B1(new_n758), .B2(new_n1108), .ZN(new_n1127));
  AND3_X1   g0927(.A1(new_n1110), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1112), .B1(new_n1110), .B2(new_n1127), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n463), .A2(G330), .A3(new_n757), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n944), .A2(new_n1131), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1124), .A2(new_n1125), .A3(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1110), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1135));
  AND2_X1   g0935(.A1(new_n1110), .A2(new_n1127), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1135), .B1(new_n1136), .B2(new_n1112), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1132), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  AND3_X1   g0939(.A1(new_n1118), .A2(new_n1110), .A3(new_n1122), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1139), .B1(new_n1140), .B2(new_n1123), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1134), .A2(new_n1141), .A3(new_n735), .ZN(new_n1142));
  OAI221_X1 g0942(.A(new_n274), .B1(new_n814), .B2(new_n217), .C1(new_n859), .C2(new_n830), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1143), .B1(G107), .B2(new_n797), .ZN(new_n1144));
  OAI22_X1  g0944(.A1(new_n809), .A2(new_n598), .B1(new_n804), .B2(new_n222), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1145), .B1(G294), .B2(new_n873), .ZN(new_n1146));
  NAND4_X1  g0946(.A1(new_n1144), .A2(new_n871), .A3(new_n1094), .A4(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n786), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n276), .B1(new_n1148), .B2(new_n309), .ZN(new_n1149));
  INV_X1    g0949(.A(KEYINPUT117), .ZN(new_n1150));
  OR2_X1    g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n814), .A2(new_n290), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(new_n1152), .B(KEYINPUT53), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1151), .A2(new_n1153), .A3(new_n1154), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(KEYINPUT54), .B(G143), .ZN(new_n1156));
  INV_X1    g0956(.A(G125), .ZN(new_n1157));
  OAI22_X1  g0957(.A1(new_n804), .A2(new_n1156), .B1(new_n811), .B2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1158), .B1(G132), .B2(new_n827), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n797), .A2(G137), .B1(new_n806), .B2(G128), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n1159), .B(new_n1160), .C1(new_n818), .C2(new_n793), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1147), .B1(new_n1155), .B2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1162), .A2(new_n778), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n855), .ZN(new_n1164));
  OAI211_X1 g0964(.A(new_n1163), .B(new_n765), .C1(new_n302), .C2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1165), .B1(new_n937), .B2(new_n775), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n1140), .A2(new_n1123), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1166), .B1(new_n1167), .B2(new_n764), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1142), .A2(new_n1168), .ZN(G378));
  INV_X1    g0969(.A(KEYINPUT121), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n951), .A2(new_n953), .ZN(new_n1171));
  NAND4_X1  g0971(.A1(new_n919), .A2(KEYINPUT40), .A3(new_n757), .A4(new_n846), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n957), .B(G330), .C1(new_n1171), .C2(new_n1172), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n315), .A2(new_n711), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(new_n326), .B(new_n1174), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1176), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(new_n1175), .B(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1173), .A2(new_n1179), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n954), .A2(G330), .A3(new_n957), .A4(new_n1178), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n1182), .A2(new_n941), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n939), .B1(new_n923), .B2(KEYINPUT103), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(new_n1181), .A2(new_n1180), .B1(new_n1184), .B2(new_n926), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1170), .B1(new_n1183), .B2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1182), .A2(new_n941), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n1180), .A2(new_n1184), .A3(new_n1181), .A4(new_n926), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1187), .A2(KEYINPUT121), .A3(new_n1188), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1186), .A2(new_n764), .A3(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n837), .B1(new_n309), .B2(new_n855), .ZN(new_n1191));
  OAI221_X1 g0991(.A(new_n1046), .B1(new_n401), .B2(new_n804), .C1(new_n830), .C2(new_n598), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1192), .B1(G97), .B2(new_n797), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n1148), .A2(new_n220), .ZN(new_n1194));
  OAI22_X1  g0994(.A1(new_n809), .A2(new_n410), .B1(new_n811), .B2(new_n859), .ZN(new_n1195));
  NOR4_X1   g0995(.A1(new_n1194), .A2(G41), .A3(new_n551), .A4(new_n1195), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1193), .A2(new_n1013), .A3(new_n1196), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(new_n1197), .B(KEYINPUT58), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(G33), .A2(G41), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n1199), .A2(G50), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1200), .B1(new_n551), .B2(G41), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n793), .A2(new_n290), .B1(new_n830), .B2(new_n1157), .ZN(new_n1202));
  XNOR2_X1  g1002(.A(new_n1202), .B(KEYINPUT118), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n797), .A2(G132), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n827), .A2(G128), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1156), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(new_n815), .A2(new_n1206), .B1(new_n828), .B2(G137), .ZN(new_n1207));
  NAND4_X1  g1007(.A1(new_n1203), .A2(new_n1204), .A3(new_n1205), .A4(new_n1207), .ZN(new_n1208));
  XOR2_X1   g1008(.A(new_n1208), .B(KEYINPUT119), .Z(new_n1209));
  INV_X1    g1009(.A(new_n1209), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n1210), .A2(KEYINPUT59), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1199), .B1(new_n1148), .B2(new_n818), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1212), .B1(G124), .B2(new_n873), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT59), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1213), .B1(new_n1209), .B2(new_n1214), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n1198), .B(new_n1201), .C1(new_n1211), .C2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1216), .A2(KEYINPUT120), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1217), .A2(new_n778), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1216), .A2(KEYINPUT120), .ZN(new_n1219));
  OAI221_X1 g1019(.A(new_n1191), .B1(new_n1218), .B2(new_n1219), .C1(new_n1178), .C2(new_n776), .ZN(new_n1220));
  AND3_X1   g1020(.A1(new_n1190), .A2(KEYINPUT122), .A3(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(KEYINPUT122), .B1(new_n1190), .B2(new_n1220), .ZN(new_n1222));
  OR2_X1    g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(KEYINPUT57), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1186), .A2(new_n1189), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1132), .B1(new_n1167), .B2(new_n1133), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1224), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  OAI21_X1  g1027(.A(KEYINPUT123), .B1(new_n1183), .B2(new_n1185), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT123), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1188), .A2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1228), .A2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1134), .A2(new_n1138), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1231), .A2(KEYINPUT57), .A3(new_n1232), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1227), .A2(new_n735), .A3(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1223), .A2(new_n1234), .ZN(G375));
  NAND2_X1  g1035(.A1(new_n1113), .A2(new_n775), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n765), .B1(G68), .B2(new_n1164), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n276), .B1(new_n873), .B2(G303), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1238), .B1(new_n858), .B2(new_n598), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1239), .B1(G294), .B2(new_n806), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n787), .A2(G77), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n809), .A2(new_n859), .B1(new_n804), .B2(new_n410), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1242), .B1(G97), .B2(new_n815), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1240), .A2(new_n1051), .A3(new_n1241), .A4(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1194), .B1(G137), .B2(new_n827), .ZN(new_n1245));
  OAI22_X1  g1045(.A1(new_n814), .A2(new_n818), .B1(new_n804), .B2(new_n290), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1246), .B1(G128), .B2(new_n873), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(new_n1206), .A2(new_n797), .B1(G132), .B2(new_n806), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1245), .A2(new_n551), .A3(new_n1247), .A4(new_n1248), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n793), .A2(new_n309), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1244), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1237), .B1(new_n1251), .B2(new_n778), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(new_n1137), .A2(new_n764), .B1(new_n1236), .B2(new_n1252), .ZN(new_n1253));
  OR2_X1    g1053(.A1(new_n1133), .A2(new_n991), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1253), .B1(new_n1254), .B2(new_n1255), .ZN(G381));
  INV_X1    g1056(.A(G375), .ZN(new_n1257));
  INV_X1    g1057(.A(G390), .ZN(new_n1258));
  INV_X1    g1058(.A(G378), .ZN(new_n1259));
  OR2_X1    g1059(.A1(G393), .A2(G396), .ZN(new_n1260));
  NOR4_X1   g1060(.A1(G387), .A2(G384), .A3(G381), .A4(new_n1260), .ZN(new_n1261));
  NAND4_X1  g1061(.A1(new_n1257), .A2(new_n1258), .A3(new_n1259), .A4(new_n1261), .ZN(G407));
  NAND2_X1  g1062(.A1(new_n712), .A2(G213), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1263), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1257), .A2(new_n1259), .A3(new_n1264), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(G407), .A2(new_n1265), .A3(G213), .ZN(G409));
  OAI211_X1 g1066(.A(new_n1234), .B(G378), .C1(new_n1222), .C2(new_n1221), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1231), .A2(new_n764), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(new_n1220), .ZN(new_n1269));
  NOR3_X1   g1069(.A1(new_n1225), .A2(new_n1226), .A3(new_n991), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1259), .B1(new_n1269), .B2(new_n1270), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1264), .B1(new_n1267), .B2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT125), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT124), .ZN(new_n1275));
  OAI211_X1 g1075(.A(new_n1275), .B(new_n1139), .C1(new_n1255), .C2(KEYINPUT60), .ZN(new_n1276));
  AOI21_X1  g1076(.A(KEYINPUT60), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1277));
  OAI21_X1  g1077(.A(KEYINPUT124), .B1(new_n1277), .B2(new_n1133), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1072), .B1(new_n1255), .B2(KEYINPUT60), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1276), .A2(new_n1278), .A3(new_n1279), .ZN(new_n1280));
  AND3_X1   g1080(.A1(new_n1280), .A2(G384), .A3(new_n1253), .ZN(new_n1281));
  AOI21_X1  g1081(.A(G384), .B1(new_n1280), .B2(new_n1253), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1274), .B1(new_n1281), .B2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1280), .A2(new_n1253), .ZN(new_n1284));
  INV_X1    g1084(.A(G384), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1280), .A2(G384), .A3(new_n1253), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1286), .A2(KEYINPUT125), .A3(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1264), .A2(G2897), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1283), .A2(new_n1288), .A3(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1291), .A2(G2897), .A3(new_n1264), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1290), .A2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1293), .ZN(new_n1294));
  AOI21_X1  g1094(.A(KEYINPUT61), .B1(new_n1273), .B2(new_n1294), .ZN(new_n1295));
  AND2_X1   g1095(.A1(new_n1283), .A2(new_n1288), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1272), .A2(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT63), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(G387), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1258), .A2(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(G390), .A2(G387), .ZN(new_n1302));
  XNOR2_X1  g1102(.A(G393), .B(new_n841), .ZN(new_n1303));
  NAND4_X1  g1103(.A1(new_n1301), .A2(new_n1302), .A3(KEYINPUT126), .A4(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1303), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1300), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1306));
  OAI21_X1  g1106(.A(KEYINPUT126), .B1(G390), .B2(G387), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1305), .B1(new_n1306), .B2(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1304), .A2(new_n1308), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1272), .A2(KEYINPUT63), .A3(new_n1296), .ZN(new_n1310));
  NAND4_X1  g1110(.A1(new_n1295), .A2(new_n1299), .A3(new_n1309), .A4(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT62), .ZN(new_n1312));
  AND3_X1   g1112(.A1(new_n1272), .A2(new_n1312), .A3(new_n1296), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT61), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1314), .B1(new_n1272), .B2(new_n1293), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1312), .B1(new_n1272), .B2(new_n1296), .ZN(new_n1316));
  NOR3_X1   g1116(.A1(new_n1313), .A2(new_n1315), .A3(new_n1316), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1311), .B1(new_n1317), .B2(new_n1309), .ZN(G405));
  NAND2_X1  g1118(.A1(G375), .A2(new_n1259), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1319), .A2(new_n1267), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1291), .B1(new_n1274), .B2(KEYINPUT127), .ZN(new_n1321));
  NOR2_X1   g1121(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT127), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1296), .A2(new_n1323), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n1324), .B1(new_n1267), .B2(new_n1319), .ZN(new_n1325));
  OAI211_X1 g1125(.A(new_n1304), .B(new_n1308), .C1(new_n1322), .C2(new_n1325), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1320), .A2(new_n1323), .A3(new_n1296), .ZN(new_n1327));
  OAI211_X1 g1127(.A(new_n1327), .B(new_n1309), .C1(new_n1320), .C2(new_n1321), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1326), .A2(new_n1328), .ZN(G402));
endmodule


