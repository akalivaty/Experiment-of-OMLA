

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595;

  XNOR2_X1 U326 ( .A(n449), .B(n294), .ZN(n342) );
  XNOR2_X1 U327 ( .A(n307), .B(KEYINPUT89), .ZN(n308) );
  NOR2_X1 U328 ( .A1(n548), .A2(n297), .ZN(n571) );
  XNOR2_X1 U329 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U330 ( .A(n309), .B(n308), .ZN(n312) );
  AND2_X1 U331 ( .A1(G232GAT), .A2(G233GAT), .ZN(n294) );
  XNOR2_X1 U332 ( .A(n356), .B(n355), .ZN(n401) );
  XOR2_X1 U333 ( .A(n359), .B(n358), .Z(n295) );
  XOR2_X1 U334 ( .A(KEYINPUT102), .B(n478), .Z(n296) );
  XOR2_X1 U335 ( .A(KEYINPUT55), .B(n465), .Z(n297) );
  INV_X1 U336 ( .A(n560), .ZN(n399) );
  NOR2_X1 U337 ( .A1(n404), .A2(n403), .ZN(n405) );
  XNOR2_X1 U338 ( .A(n341), .B(n340), .ZN(n361) );
  XNOR2_X1 U339 ( .A(n368), .B(n367), .ZN(n369) );
  XNOR2_X1 U340 ( .A(n342), .B(n361), .ZN(n343) );
  XNOR2_X1 U341 ( .A(KEYINPUT37), .B(KEYINPUT106), .ZN(n485) );
  XNOR2_X1 U342 ( .A(n370), .B(n369), .ZN(n374) );
  XNOR2_X1 U343 ( .A(n486), .B(n485), .ZN(n509) );
  XNOR2_X1 U344 ( .A(n585), .B(KEYINPUT41), .ZN(n562) );
  XNOR2_X1 U345 ( .A(n378), .B(n377), .ZN(n585) );
  INV_X1 U346 ( .A(G85GAT), .ZN(n489) );
  XNOR2_X1 U347 ( .A(n423), .B(n313), .ZN(n548) );
  XNOR2_X1 U348 ( .A(n492), .B(G176GAT), .ZN(n493) );
  XNOR2_X1 U349 ( .A(n489), .B(KEYINPUT116), .ZN(n490) );
  XNOR2_X1 U350 ( .A(n494), .B(n493), .ZN(G1349GAT) );
  XNOR2_X1 U351 ( .A(n491), .B(n490), .ZN(G1336GAT) );
  XOR2_X1 U352 ( .A(KEYINPUT18), .B(KEYINPUT91), .Z(n299) );
  XNOR2_X1 U353 ( .A(KEYINPUT19), .B(KEYINPUT17), .ZN(n298) );
  XNOR2_X1 U354 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U355 ( .A(G169GAT), .B(n300), .Z(n423) );
  XOR2_X1 U356 ( .A(KEYINPUT90), .B(G176GAT), .Z(n302) );
  XNOR2_X1 U357 ( .A(G43GAT), .B(G183GAT), .ZN(n301) );
  XOR2_X1 U358 ( .A(n302), .B(n301), .Z(n306) );
  XOR2_X1 U359 ( .A(G15GAT), .B(G127GAT), .Z(n318) );
  XOR2_X1 U360 ( .A(G190GAT), .B(G99GAT), .Z(n303) );
  XNOR2_X1 U361 ( .A(n318), .B(n303), .ZN(n304) );
  XOR2_X1 U362 ( .A(G120GAT), .B(G71GAT), .Z(n367) );
  XNOR2_X1 U363 ( .A(n304), .B(n367), .ZN(n305) );
  XNOR2_X1 U364 ( .A(n306), .B(n305), .ZN(n309) );
  NAND2_X1 U365 ( .A1(G227GAT), .A2(G233GAT), .ZN(n307) );
  XNOR2_X1 U366 ( .A(G113GAT), .B(G134GAT), .ZN(n310) );
  XNOR2_X1 U367 ( .A(n310), .B(KEYINPUT0), .ZN(n441) );
  XOR2_X1 U368 ( .A(n441), .B(KEYINPUT20), .Z(n311) );
  XNOR2_X1 U369 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U370 ( .A(KEYINPUT45), .B(KEYINPUT117), .Z(n359) );
  INV_X1 U371 ( .A(G155GAT), .ZN(n314) );
  NAND2_X1 U372 ( .A1(G22GAT), .A2(n314), .ZN(n317) );
  INV_X1 U373 ( .A(G22GAT), .ZN(n315) );
  NAND2_X1 U374 ( .A1(n315), .A2(G155GAT), .ZN(n316) );
  NAND2_X1 U375 ( .A1(n317), .A2(n316), .ZN(n448) );
  XOR2_X1 U376 ( .A(n448), .B(n318), .Z(n320) );
  NAND2_X1 U377 ( .A1(G231GAT), .A2(G233GAT), .ZN(n319) );
  XNOR2_X1 U378 ( .A(n320), .B(n319), .ZN(n331) );
  XOR2_X1 U379 ( .A(KEYINPUT15), .B(KEYINPUT87), .Z(n326) );
  XNOR2_X1 U380 ( .A(G57GAT), .B(KEYINPUT75), .ZN(n321) );
  XNOR2_X1 U381 ( .A(n321), .B(KEYINPUT13), .ZN(n376) );
  XOR2_X1 U382 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n323) );
  XNOR2_X1 U383 ( .A(G78GAT), .B(G64GAT), .ZN(n322) );
  XNOR2_X1 U384 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U385 ( .A(n376), .B(n324), .ZN(n325) );
  XNOR2_X1 U386 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U387 ( .A(G8GAT), .B(G183GAT), .Z(n413) );
  XOR2_X1 U388 ( .A(n327), .B(n413), .Z(n329) );
  XNOR2_X1 U389 ( .A(G71GAT), .B(G211GAT), .ZN(n328) );
  XNOR2_X1 U390 ( .A(n329), .B(n328), .ZN(n330) );
  XNOR2_X1 U391 ( .A(n331), .B(n330), .ZN(n333) );
  XOR2_X1 U392 ( .A(KEYINPUT73), .B(G1GAT), .Z(n390) );
  INV_X1 U393 ( .A(n390), .ZN(n332) );
  XOR2_X1 U394 ( .A(n333), .B(n332), .Z(n588) );
  XOR2_X1 U395 ( .A(KEYINPUT85), .B(G92GAT), .Z(n335) );
  XNOR2_X1 U396 ( .A(G190GAT), .B(G218GAT), .ZN(n334) );
  XNOR2_X1 U397 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U398 ( .A(G36GAT), .B(n336), .Z(n419) );
  XOR2_X1 U399 ( .A(G50GAT), .B(G162GAT), .Z(n449) );
  NAND2_X1 U400 ( .A1(KEYINPUT79), .A2(n489), .ZN(n339) );
  INV_X1 U401 ( .A(KEYINPUT79), .ZN(n337) );
  NAND2_X1 U402 ( .A1(n337), .A2(G85GAT), .ZN(n338) );
  NAND2_X1 U403 ( .A1(n339), .A2(n338), .ZN(n341) );
  XNOR2_X1 U404 ( .A(G99GAT), .B(G106GAT), .ZN(n340) );
  XNOR2_X1 U405 ( .A(n419), .B(n343), .ZN(n356) );
  XOR2_X1 U406 ( .A(KEYINPUT82), .B(KEYINPUT66), .Z(n345) );
  XNOR2_X1 U407 ( .A(KEYINPUT9), .B(KEYINPUT11), .ZN(n344) );
  XNOR2_X1 U408 ( .A(n345), .B(n344), .ZN(n349) );
  XOR2_X1 U409 ( .A(KEYINPUT10), .B(KEYINPUT84), .Z(n347) );
  XNOR2_X1 U410 ( .A(G134GAT), .B(KEYINPUT83), .ZN(n346) );
  XNOR2_X1 U411 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U412 ( .A(n349), .B(n348), .Z(n354) );
  XOR2_X1 U413 ( .A(KEYINPUT8), .B(KEYINPUT72), .Z(n351) );
  XNOR2_X1 U414 ( .A(G43GAT), .B(G29GAT), .ZN(n350) );
  XNOR2_X1 U415 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U416 ( .A(KEYINPUT7), .B(n352), .ZN(n398) );
  INV_X1 U417 ( .A(n398), .ZN(n353) );
  XOR2_X1 U418 ( .A(KEYINPUT86), .B(n401), .Z(n572) );
  XNOR2_X1 U419 ( .A(KEYINPUT36), .B(KEYINPUT105), .ZN(n357) );
  XOR2_X1 U420 ( .A(n572), .B(n357), .Z(n591) );
  NAND2_X1 U421 ( .A1(n588), .A2(n591), .ZN(n358) );
  INV_X1 U422 ( .A(KEYINPUT81), .ZN(n360) );
  XNOR2_X1 U423 ( .A(n361), .B(n360), .ZN(n363) );
  NAND2_X1 U424 ( .A1(G230GAT), .A2(G233GAT), .ZN(n362) );
  XNOR2_X1 U425 ( .A(n363), .B(n362), .ZN(n370) );
  XOR2_X1 U426 ( .A(KEYINPUT76), .B(KEYINPUT31), .Z(n365) );
  XNOR2_X1 U427 ( .A(G204GAT), .B(G92GAT), .ZN(n364) );
  XNOR2_X1 U428 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U429 ( .A(G176GAT), .B(G64GAT), .Z(n412) );
  XOR2_X1 U430 ( .A(n366), .B(n412), .Z(n368) );
  XOR2_X1 U431 ( .A(KEYINPUT80), .B(KEYINPUT32), .Z(n372) );
  XNOR2_X1 U432 ( .A(KEYINPUT33), .B(KEYINPUT77), .ZN(n371) );
  XNOR2_X1 U433 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U434 ( .A(n374), .B(n373), .Z(n378) );
  XNOR2_X1 U435 ( .A(G78GAT), .B(KEYINPUT78), .ZN(n375) );
  XNOR2_X1 U436 ( .A(n375), .B(G148GAT), .ZN(n462) );
  XNOR2_X1 U437 ( .A(n462), .B(n376), .ZN(n377) );
  XOR2_X1 U438 ( .A(G197GAT), .B(G22GAT), .Z(n380) );
  XNOR2_X1 U439 ( .A(G169GAT), .B(G141GAT), .ZN(n379) );
  XNOR2_X1 U440 ( .A(n380), .B(n379), .ZN(n384) );
  XOR2_X1 U441 ( .A(G8GAT), .B(KEYINPUT69), .Z(n382) );
  XNOR2_X1 U442 ( .A(KEYINPUT68), .B(KEYINPUT29), .ZN(n381) );
  XNOR2_X1 U443 ( .A(n382), .B(n381), .ZN(n383) );
  XOR2_X1 U444 ( .A(n384), .B(n383), .Z(n396) );
  XOR2_X1 U445 ( .A(KEYINPUT74), .B(KEYINPUT71), .Z(n386) );
  XNOR2_X1 U446 ( .A(KEYINPUT70), .B(KEYINPUT30), .ZN(n385) );
  XNOR2_X1 U447 ( .A(n386), .B(n385), .ZN(n394) );
  XOR2_X1 U448 ( .A(G15GAT), .B(G113GAT), .Z(n388) );
  XNOR2_X1 U449 ( .A(G50GAT), .B(G36GAT), .ZN(n387) );
  XNOR2_X1 U450 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U451 ( .A(n390), .B(n389), .Z(n392) );
  NAND2_X1 U452 ( .A1(G229GAT), .A2(G233GAT), .ZN(n391) );
  XNOR2_X1 U453 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U454 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U455 ( .A(n396), .B(n395), .ZN(n397) );
  XOR2_X1 U456 ( .A(n398), .B(n397), .Z(n560) );
  NOR2_X1 U457 ( .A1(n585), .A2(n399), .ZN(n400) );
  NAND2_X1 U458 ( .A1(n295), .A2(n400), .ZN(n407) );
  INV_X1 U459 ( .A(n588), .ZN(n566) );
  NAND2_X1 U460 ( .A1(n401), .A2(n566), .ZN(n404) );
  NOR2_X1 U461 ( .A1(n560), .A2(n562), .ZN(n402) );
  XNOR2_X1 U462 ( .A(n402), .B(KEYINPUT46), .ZN(n403) );
  XNOR2_X1 U463 ( .A(n405), .B(KEYINPUT47), .ZN(n406) );
  NAND2_X1 U464 ( .A1(n407), .A2(n406), .ZN(n409) );
  XOR2_X1 U465 ( .A(KEYINPUT48), .B(KEYINPUT64), .Z(n408) );
  XNOR2_X1 U466 ( .A(n409), .B(n408), .ZN(n544) );
  XOR2_X1 U467 ( .A(G204GAT), .B(G211GAT), .Z(n411) );
  XNOR2_X1 U468 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n410) );
  XNOR2_X1 U469 ( .A(n411), .B(n410), .ZN(n461) );
  XNOR2_X1 U470 ( .A(n461), .B(n412), .ZN(n414) );
  XNOR2_X1 U471 ( .A(n414), .B(n413), .ZN(n418) );
  XOR2_X1 U472 ( .A(KEYINPUT99), .B(KEYINPUT97), .Z(n416) );
  NAND2_X1 U473 ( .A1(G226GAT), .A2(G233GAT), .ZN(n415) );
  XNOR2_X1 U474 ( .A(n416), .B(n415), .ZN(n417) );
  XOR2_X1 U475 ( .A(n418), .B(n417), .Z(n421) );
  XNOR2_X1 U476 ( .A(n419), .B(KEYINPUT98), .ZN(n420) );
  XNOR2_X1 U477 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U478 ( .A(n423), .B(n422), .ZN(n535) );
  NOR2_X1 U479 ( .A1(n544), .A2(n535), .ZN(n424) );
  XNOR2_X1 U480 ( .A(n424), .B(KEYINPUT54), .ZN(n444) );
  XOR2_X1 U481 ( .A(G85GAT), .B(G162GAT), .Z(n426) );
  XNOR2_X1 U482 ( .A(G29GAT), .B(G127GAT), .ZN(n425) );
  XNOR2_X1 U483 ( .A(n426), .B(n425), .ZN(n430) );
  XOR2_X1 U484 ( .A(G57GAT), .B(G155GAT), .Z(n428) );
  XNOR2_X1 U485 ( .A(G120GAT), .B(G148GAT), .ZN(n427) );
  XNOR2_X1 U486 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U487 ( .A(n430), .B(n429), .Z(n435) );
  XOR2_X1 U488 ( .A(KEYINPUT95), .B(KEYINPUT6), .Z(n432) );
  NAND2_X1 U489 ( .A1(G225GAT), .A2(G233GAT), .ZN(n431) );
  XNOR2_X1 U490 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U491 ( .A(KEYINPUT1), .B(n433), .ZN(n434) );
  XNOR2_X1 U492 ( .A(n435), .B(n434), .ZN(n439) );
  XOR2_X1 U493 ( .A(KEYINPUT96), .B(KEYINPUT5), .Z(n437) );
  XNOR2_X1 U494 ( .A(G1GAT), .B(KEYINPUT4), .ZN(n436) );
  XNOR2_X1 U495 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U496 ( .A(n439), .B(n438), .Z(n443) );
  XNOR2_X1 U497 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n440) );
  XNOR2_X1 U498 ( .A(n440), .B(KEYINPUT2), .ZN(n457) );
  XNOR2_X1 U499 ( .A(n441), .B(n457), .ZN(n442) );
  XNOR2_X1 U500 ( .A(n443), .B(n442), .ZN(n523) );
  NAND2_X1 U501 ( .A1(n444), .A2(n523), .ZN(n445) );
  XNOR2_X1 U502 ( .A(n445), .B(KEYINPUT65), .ZN(n580) );
  XOR2_X1 U503 ( .A(KEYINPUT94), .B(KEYINPUT24), .Z(n447) );
  XNOR2_X1 U504 ( .A(KEYINPUT93), .B(KEYINPUT22), .ZN(n446) );
  XNOR2_X1 U505 ( .A(n447), .B(n446), .ZN(n453) );
  XNOR2_X1 U506 ( .A(n449), .B(n448), .ZN(n451) );
  XOR2_X1 U507 ( .A(G106GAT), .B(G218GAT), .Z(n450) );
  XNOR2_X1 U508 ( .A(n451), .B(n450), .ZN(n452) );
  XOR2_X1 U509 ( .A(n453), .B(n452), .Z(n455) );
  NAND2_X1 U510 ( .A1(G228GAT), .A2(G233GAT), .ZN(n454) );
  XNOR2_X1 U511 ( .A(n455), .B(n454), .ZN(n456) );
  XOR2_X1 U512 ( .A(n456), .B(KEYINPUT23), .Z(n459) );
  XNOR2_X1 U513 ( .A(n457), .B(KEYINPUT92), .ZN(n458) );
  XNOR2_X1 U514 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U515 ( .A(n461), .B(n460), .ZN(n464) );
  INV_X1 U516 ( .A(n462), .ZN(n463) );
  XNOR2_X1 U517 ( .A(n464), .B(n463), .ZN(n471) );
  NAND2_X1 U518 ( .A1(n580), .A2(n471), .ZN(n465) );
  NAND2_X1 U519 ( .A1(n571), .A2(n399), .ZN(n467) );
  XNOR2_X1 U520 ( .A(G169GAT), .B(KEYINPUT120), .ZN(n466) );
  XNOR2_X1 U521 ( .A(n467), .B(n466), .ZN(G1348GAT) );
  OR2_X1 U522 ( .A1(n535), .A2(n548), .ZN(n468) );
  NAND2_X1 U523 ( .A1(n468), .A2(n471), .ZN(n469) );
  XNOR2_X1 U524 ( .A(n469), .B(KEYINPUT25), .ZN(n470) );
  XNOR2_X1 U525 ( .A(n470), .B(KEYINPUT101), .ZN(n476) );
  INV_X1 U526 ( .A(n548), .ZN(n482) );
  NOR2_X1 U527 ( .A1(n482), .A2(n471), .ZN(n472) );
  XNOR2_X1 U528 ( .A(n472), .B(KEYINPUT26), .ZN(n581) );
  XOR2_X1 U529 ( .A(KEYINPUT27), .B(KEYINPUT100), .Z(n473) );
  XOR2_X1 U530 ( .A(n535), .B(n473), .Z(n479) );
  INV_X1 U531 ( .A(n479), .ZN(n474) );
  NAND2_X1 U532 ( .A1(n581), .A2(n474), .ZN(n475) );
  NAND2_X1 U533 ( .A1(n476), .A2(n475), .ZN(n477) );
  NAND2_X1 U534 ( .A1(n477), .A2(n523), .ZN(n478) );
  NOR2_X1 U535 ( .A1(n523), .A2(n479), .ZN(n542) );
  XOR2_X1 U536 ( .A(KEYINPUT28), .B(KEYINPUT67), .Z(n480) );
  XNOR2_X1 U537 ( .A(n471), .B(n480), .ZN(n546) );
  NAND2_X1 U538 ( .A1(n542), .A2(n546), .ZN(n481) );
  NOR2_X1 U539 ( .A1(n482), .A2(n481), .ZN(n483) );
  NOR2_X1 U540 ( .A1(n296), .A2(n483), .ZN(n498) );
  NOR2_X1 U541 ( .A1(n588), .A2(n498), .ZN(n484) );
  NAND2_X1 U542 ( .A1(n591), .A2(n484), .ZN(n486) );
  INV_X1 U543 ( .A(n562), .ZN(n550) );
  NAND2_X1 U544 ( .A1(n560), .A2(n550), .ZN(n487) );
  XNOR2_X1 U545 ( .A(n487), .B(KEYINPUT109), .ZN(n520) );
  NAND2_X1 U546 ( .A1(n509), .A2(n520), .ZN(n488) );
  XOR2_X1 U547 ( .A(KEYINPUT115), .B(n488), .Z(n538) );
  NOR2_X1 U548 ( .A1(n523), .A2(n538), .ZN(n491) );
  NAND2_X1 U549 ( .A1(n571), .A2(n550), .ZN(n494) );
  XOR2_X1 U550 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n492) );
  NOR2_X1 U551 ( .A1(n585), .A2(n560), .ZN(n508) );
  OR2_X1 U552 ( .A1(n566), .A2(n572), .ZN(n495) );
  XNOR2_X1 U553 ( .A(n495), .B(KEYINPUT16), .ZN(n496) );
  XNOR2_X1 U554 ( .A(n496), .B(KEYINPUT88), .ZN(n497) );
  NOR2_X1 U555 ( .A1(n498), .A2(n497), .ZN(n521) );
  NAND2_X1 U556 ( .A1(n508), .A2(n521), .ZN(n506) );
  NOR2_X1 U557 ( .A1(n523), .A2(n506), .ZN(n499) );
  XOR2_X1 U558 ( .A(G1GAT), .B(n499), .Z(n500) );
  XNOR2_X1 U559 ( .A(KEYINPUT34), .B(n500), .ZN(G1324GAT) );
  NOR2_X1 U560 ( .A1(n535), .A2(n506), .ZN(n502) );
  XNOR2_X1 U561 ( .A(KEYINPUT103), .B(KEYINPUT104), .ZN(n501) );
  XNOR2_X1 U562 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U563 ( .A(G8GAT), .B(n503), .ZN(G1325GAT) );
  NOR2_X1 U564 ( .A1(n548), .A2(n506), .ZN(n505) );
  XNOR2_X1 U565 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n504) );
  XNOR2_X1 U566 ( .A(n505), .B(n504), .ZN(G1326GAT) );
  NOR2_X1 U567 ( .A1(n546), .A2(n506), .ZN(n507) );
  XOR2_X1 U568 ( .A(G22GAT), .B(n507), .Z(G1327GAT) );
  XNOR2_X1 U569 ( .A(KEYINPUT39), .B(KEYINPUT107), .ZN(n512) );
  NAND2_X1 U570 ( .A1(n509), .A2(n508), .ZN(n510) );
  XNOR2_X1 U571 ( .A(n510), .B(KEYINPUT38), .ZN(n518) );
  NOR2_X1 U572 ( .A1(n523), .A2(n518), .ZN(n511) );
  XNOR2_X1 U573 ( .A(n512), .B(n511), .ZN(n513) );
  XOR2_X1 U574 ( .A(G29GAT), .B(n513), .Z(G1328GAT) );
  NOR2_X1 U575 ( .A1(n518), .A2(n535), .ZN(n514) );
  XOR2_X1 U576 ( .A(KEYINPUT108), .B(n514), .Z(n515) );
  XNOR2_X1 U577 ( .A(G36GAT), .B(n515), .ZN(G1329GAT) );
  NOR2_X1 U578 ( .A1(n518), .A2(n548), .ZN(n516) );
  XOR2_X1 U579 ( .A(KEYINPUT40), .B(n516), .Z(n517) );
  XNOR2_X1 U580 ( .A(G43GAT), .B(n517), .ZN(G1330GAT) );
  NOR2_X1 U581 ( .A1(n546), .A2(n518), .ZN(n519) );
  XOR2_X1 U582 ( .A(G50GAT), .B(n519), .Z(G1331GAT) );
  XNOR2_X1 U583 ( .A(KEYINPUT42), .B(KEYINPUT111), .ZN(n525) );
  NAND2_X1 U584 ( .A1(n521), .A2(n520), .ZN(n522) );
  XNOR2_X1 U585 ( .A(n522), .B(KEYINPUT110), .ZN(n530) );
  NOR2_X1 U586 ( .A1(n523), .A2(n530), .ZN(n524) );
  XNOR2_X1 U587 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U588 ( .A(G57GAT), .B(n526), .ZN(G1332GAT) );
  NOR2_X1 U589 ( .A1(n530), .A2(n535), .ZN(n527) );
  XOR2_X1 U590 ( .A(KEYINPUT112), .B(n527), .Z(n528) );
  XNOR2_X1 U591 ( .A(G64GAT), .B(n528), .ZN(G1333GAT) );
  NOR2_X1 U592 ( .A1(n530), .A2(n548), .ZN(n529) );
  XOR2_X1 U593 ( .A(G71GAT), .B(n529), .Z(G1334GAT) );
  NOR2_X1 U594 ( .A1(n530), .A2(n546), .ZN(n534) );
  XOR2_X1 U595 ( .A(KEYINPUT113), .B(KEYINPUT43), .Z(n532) );
  XNOR2_X1 U596 ( .A(G78GAT), .B(KEYINPUT114), .ZN(n531) );
  XNOR2_X1 U597 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U598 ( .A(n534), .B(n533), .ZN(G1335GAT) );
  NOR2_X1 U599 ( .A1(n535), .A2(n538), .ZN(n536) );
  XOR2_X1 U600 ( .A(G92GAT), .B(n536), .Z(G1337GAT) );
  NOR2_X1 U601 ( .A1(n548), .A2(n538), .ZN(n537) );
  XOR2_X1 U602 ( .A(G99GAT), .B(n537), .Z(G1338GAT) );
  INV_X1 U603 ( .A(KEYINPUT44), .ZN(n540) );
  NOR2_X1 U604 ( .A1(n546), .A2(n538), .ZN(n539) );
  XNOR2_X1 U605 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U606 ( .A(G106GAT), .B(n541), .ZN(G1339GAT) );
  INV_X1 U607 ( .A(n542), .ZN(n543) );
  NOR2_X1 U608 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U609 ( .A(KEYINPUT118), .B(n545), .ZN(n559) );
  NAND2_X1 U610 ( .A1(n546), .A2(n559), .ZN(n547) );
  NOR2_X1 U611 ( .A1(n548), .A2(n547), .ZN(n556) );
  NAND2_X1 U612 ( .A1(n399), .A2(n556), .ZN(n549) );
  XNOR2_X1 U613 ( .A(G113GAT), .B(n549), .ZN(G1340GAT) );
  XOR2_X1 U614 ( .A(KEYINPUT49), .B(KEYINPUT119), .Z(n552) );
  NAND2_X1 U615 ( .A1(n556), .A2(n550), .ZN(n551) );
  XNOR2_X1 U616 ( .A(n552), .B(n551), .ZN(n553) );
  XOR2_X1 U617 ( .A(G120GAT), .B(n553), .Z(G1341GAT) );
  NAND2_X1 U618 ( .A1(n556), .A2(n588), .ZN(n554) );
  XNOR2_X1 U619 ( .A(n554), .B(KEYINPUT50), .ZN(n555) );
  XNOR2_X1 U620 ( .A(G127GAT), .B(n555), .ZN(G1342GAT) );
  XOR2_X1 U621 ( .A(G134GAT), .B(KEYINPUT51), .Z(n558) );
  NAND2_X1 U622 ( .A1(n556), .A2(n572), .ZN(n557) );
  XNOR2_X1 U623 ( .A(n558), .B(n557), .ZN(G1343GAT) );
  NAND2_X1 U624 ( .A1(n581), .A2(n559), .ZN(n568) );
  NOR2_X1 U625 ( .A1(n560), .A2(n568), .ZN(n561) );
  XOR2_X1 U626 ( .A(G141GAT), .B(n561), .Z(G1344GAT) );
  NOR2_X1 U627 ( .A1(n562), .A2(n568), .ZN(n564) );
  XNOR2_X1 U628 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n564), .B(n563), .ZN(n565) );
  XNOR2_X1 U630 ( .A(G148GAT), .B(n565), .ZN(G1345GAT) );
  NOR2_X1 U631 ( .A1(n566), .A2(n568), .ZN(n567) );
  XOR2_X1 U632 ( .A(G155GAT), .B(n567), .Z(G1346GAT) );
  NOR2_X1 U633 ( .A1(n401), .A2(n568), .ZN(n569) );
  XOR2_X1 U634 ( .A(G162GAT), .B(n569), .Z(G1347GAT) );
  NAND2_X1 U635 ( .A1(n571), .A2(n588), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n570), .B(G183GAT), .ZN(G1350GAT) );
  AND2_X1 U637 ( .A1(n572), .A2(n571), .ZN(n576) );
  XNOR2_X1 U638 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n573), .B(KEYINPUT121), .ZN(n574) );
  XNOR2_X1 U640 ( .A(KEYINPUT122), .B(n574), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(G1351GAT) );
  XOR2_X1 U642 ( .A(KEYINPUT125), .B(KEYINPUT60), .Z(n578) );
  XNOR2_X1 U643 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n577) );
  XNOR2_X1 U644 ( .A(n578), .B(n577), .ZN(n579) );
  XOR2_X1 U645 ( .A(KEYINPUT124), .B(n579), .Z(n584) );
  NAND2_X1 U646 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n582), .B(KEYINPUT123), .ZN(n592) );
  NAND2_X1 U648 ( .A1(n592), .A2(n399), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(G1352GAT) );
  XOR2_X1 U650 ( .A(G204GAT), .B(KEYINPUT61), .Z(n587) );
  NAND2_X1 U651 ( .A1(n592), .A2(n585), .ZN(n586) );
  XNOR2_X1 U652 ( .A(n587), .B(n586), .ZN(G1353GAT) );
  NAND2_X1 U653 ( .A1(n592), .A2(n588), .ZN(n589) );
  XNOR2_X1 U654 ( .A(n589), .B(KEYINPUT126), .ZN(n590) );
  XNOR2_X1 U655 ( .A(G211GAT), .B(n590), .ZN(G1354GAT) );
  XOR2_X1 U656 ( .A(KEYINPUT127), .B(KEYINPUT62), .Z(n594) );
  NAND2_X1 U657 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U658 ( .A(n594), .B(n593), .ZN(n595) );
  XNOR2_X1 U659 ( .A(G218GAT), .B(n595), .ZN(G1355GAT) );
endmodule

