

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U550 ( .A(KEYINPUT17), .ZN(n533) );
  XNOR2_X1 U551 ( .A(n723), .B(n722), .ZN(n724) );
  INV_X1 U552 ( .A(KEYINPUT29), .ZN(n722) );
  XNOR2_X1 U553 ( .A(n744), .B(KEYINPUT97), .ZN(n739) );
  NOR2_X1 U554 ( .A1(n782), .A2(n781), .ZN(n784) );
  INV_X1 U555 ( .A(KEYINPUT103), .ZN(n783) );
  NOR2_X1 U556 ( .A1(G651), .A2(G543), .ZN(n661) );
  NAND2_X1 U557 ( .A1(n888), .A2(G138), .ZN(n536) );
  XOR2_X1 U558 ( .A(KEYINPUT30), .B(n729), .Z(n515) );
  AND2_X1 U559 ( .A1(n814), .A2(n826), .ZN(n516) );
  AND2_X1 U560 ( .A1(n707), .A2(G1996), .ZN(n702) );
  NOR2_X1 U561 ( .A1(n945), .A2(n705), .ZN(n706) );
  INV_X1 U562 ( .A(KEYINPUT31), .ZN(n733) );
  XNOR2_X1 U563 ( .A(n733), .B(KEYINPUT96), .ZN(n734) );
  BUF_X1 U564 ( .A(n726), .Z(n746) );
  NOR2_X1 U565 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U566 ( .A1(n803), .A2(n693), .ZN(n726) );
  XNOR2_X1 U567 ( .A(n554), .B(KEYINPUT66), .ZN(n555) );
  NOR2_X1 U568 ( .A1(G164), .A2(G1384), .ZN(n803) );
  XNOR2_X1 U569 ( .A(G2104), .B(KEYINPUT65), .ZN(n538) );
  XNOR2_X1 U570 ( .A(n556), .B(n555), .ZN(n558) );
  NAND2_X1 U571 ( .A1(n516), .A2(n815), .ZN(n816) );
  XNOR2_X1 U572 ( .A(n784), .B(n783), .ZN(n817) );
  NOR2_X1 U573 ( .A1(G651), .A2(n644), .ZN(n652) );
  XNOR2_X1 U574 ( .A(KEYINPUT1), .B(n518), .ZN(n653) );
  NOR2_X1 U575 ( .A1(n542), .A2(n541), .ZN(G164) );
  XOR2_X1 U576 ( .A(KEYINPUT0), .B(G543), .Z(n644) );
  NAND2_X1 U577 ( .A1(n652), .A2(G51), .ZN(n520) );
  INV_X1 U578 ( .A(G651), .ZN(n523) );
  NOR2_X1 U579 ( .A1(G543), .A2(n523), .ZN(n517) );
  XOR2_X1 U580 ( .A(KEYINPUT70), .B(n517), .Z(n518) );
  NAND2_X1 U581 ( .A1(G63), .A2(n653), .ZN(n519) );
  NAND2_X1 U582 ( .A1(n520), .A2(n519), .ZN(n521) );
  XNOR2_X1 U583 ( .A(KEYINPUT6), .B(n521), .ZN(n530) );
  NAND2_X1 U584 ( .A1(n661), .A2(G89), .ZN(n522) );
  XNOR2_X1 U585 ( .A(n522), .B(KEYINPUT4), .ZN(n526) );
  OR2_X1 U586 ( .A1(n523), .A2(n644), .ZN(n524) );
  XOR2_X1 U587 ( .A(KEYINPUT68), .B(n524), .Z(n657) );
  NAND2_X1 U588 ( .A1(G76), .A2(n657), .ZN(n525) );
  NAND2_X1 U589 ( .A1(n526), .A2(n525), .ZN(n527) );
  XOR2_X1 U590 ( .A(KEYINPUT5), .B(n527), .Z(n528) );
  XNOR2_X1 U591 ( .A(KEYINPUT78), .B(n528), .ZN(n529) );
  NOR2_X1 U592 ( .A1(n530), .A2(n529), .ZN(n531) );
  XOR2_X1 U593 ( .A(KEYINPUT7), .B(n531), .Z(G168) );
  XNOR2_X1 U594 ( .A(G168), .B(KEYINPUT8), .ZN(n532) );
  XNOR2_X1 U595 ( .A(n532), .B(KEYINPUT79), .ZN(G286) );
  NOR2_X1 U596 ( .A1(G2104), .A2(G2105), .ZN(n534) );
  XNOR2_X2 U597 ( .A(n534), .B(n533), .ZN(n888) );
  INV_X1 U598 ( .A(G2105), .ZN(n551) );
  INV_X1 U599 ( .A(n538), .ZN(n553) );
  AND2_X1 U600 ( .A1(n551), .A2(n553), .ZN(n887) );
  NAND2_X1 U601 ( .A1(n887), .A2(G102), .ZN(n535) );
  NAND2_X1 U602 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U603 ( .A(KEYINPUT88), .B(n537), .ZN(n542) );
  AND2_X1 U604 ( .A1(n538), .A2(G2105), .ZN(n883) );
  NAND2_X1 U605 ( .A1(G126), .A2(n883), .ZN(n540) );
  AND2_X1 U606 ( .A1(G2104), .A2(G2105), .ZN(n884) );
  NAND2_X1 U607 ( .A1(G114), .A2(n884), .ZN(n539) );
  NAND2_X1 U608 ( .A1(n540), .A2(n539), .ZN(n541) );
  NAND2_X1 U609 ( .A1(n661), .A2(G91), .ZN(n544) );
  NAND2_X1 U610 ( .A1(G78), .A2(n657), .ZN(n543) );
  NAND2_X1 U611 ( .A1(n544), .A2(n543), .ZN(n548) );
  NAND2_X1 U612 ( .A1(n652), .A2(G53), .ZN(n546) );
  NAND2_X1 U613 ( .A1(G65), .A2(n653), .ZN(n545) );
  NAND2_X1 U614 ( .A1(n546), .A2(n545), .ZN(n547) );
  OR2_X1 U615 ( .A1(n548), .A2(n547), .ZN(G299) );
  NAND2_X1 U616 ( .A1(G137), .A2(n888), .ZN(n550) );
  NAND2_X1 U617 ( .A1(G113), .A2(n884), .ZN(n549) );
  AND2_X1 U618 ( .A1(n550), .A2(n549), .ZN(n690) );
  AND2_X1 U619 ( .A1(n551), .A2(G101), .ZN(n552) );
  NAND2_X1 U620 ( .A1(n553), .A2(n552), .ZN(n556) );
  INV_X1 U621 ( .A(KEYINPUT23), .ZN(n554) );
  NAND2_X1 U622 ( .A1(G125), .A2(n883), .ZN(n557) );
  NAND2_X1 U623 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U624 ( .A(KEYINPUT67), .B(n559), .ZN(n691) );
  AND2_X1 U625 ( .A1(n690), .A2(n691), .ZN(G160) );
  XOR2_X1 U626 ( .A(G2446), .B(G2430), .Z(n561) );
  XNOR2_X1 U627 ( .A(G2451), .B(KEYINPUT108), .ZN(n560) );
  XNOR2_X1 U628 ( .A(n561), .B(n560), .ZN(n562) );
  XOR2_X1 U629 ( .A(n562), .B(G2427), .Z(n564) );
  XNOR2_X1 U630 ( .A(G1348), .B(G1341), .ZN(n563) );
  XNOR2_X1 U631 ( .A(n564), .B(n563), .ZN(n568) );
  XOR2_X1 U632 ( .A(G2443), .B(G2435), .Z(n566) );
  XNOR2_X1 U633 ( .A(G2438), .B(G2454), .ZN(n565) );
  XNOR2_X1 U634 ( .A(n566), .B(n565), .ZN(n567) );
  XOR2_X1 U635 ( .A(n568), .B(n567), .Z(n569) );
  AND2_X1 U636 ( .A1(G14), .A2(n569), .ZN(G401) );
  AND2_X1 U637 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U638 ( .A(G132), .ZN(G219) );
  INV_X1 U639 ( .A(G57), .ZN(G237) );
  NAND2_X1 U640 ( .A1(n661), .A2(G88), .ZN(n571) );
  NAND2_X1 U641 ( .A1(G75), .A2(n657), .ZN(n570) );
  NAND2_X1 U642 ( .A1(n571), .A2(n570), .ZN(n575) );
  NAND2_X1 U643 ( .A1(n652), .A2(G50), .ZN(n573) );
  NAND2_X1 U644 ( .A1(G62), .A2(n653), .ZN(n572) );
  NAND2_X1 U645 ( .A1(n573), .A2(n572), .ZN(n574) );
  NOR2_X1 U646 ( .A1(n575), .A2(n574), .ZN(G166) );
  NAND2_X1 U647 ( .A1(G7), .A2(G661), .ZN(n576) );
  XNOR2_X1 U648 ( .A(n576), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U649 ( .A(G223), .ZN(n836) );
  NAND2_X1 U650 ( .A1(n836), .A2(G567), .ZN(n577) );
  XNOR2_X1 U651 ( .A(n577), .B(KEYINPUT11), .ZN(n578) );
  XNOR2_X1 U652 ( .A(KEYINPUT75), .B(n578), .ZN(G234) );
  NAND2_X1 U653 ( .A1(n661), .A2(G81), .ZN(n579) );
  XNOR2_X1 U654 ( .A(n579), .B(KEYINPUT12), .ZN(n581) );
  NAND2_X1 U655 ( .A1(G68), .A2(n657), .ZN(n580) );
  NAND2_X1 U656 ( .A1(n581), .A2(n580), .ZN(n583) );
  XOR2_X1 U657 ( .A(KEYINPUT76), .B(KEYINPUT13), .Z(n582) );
  XNOR2_X1 U658 ( .A(n583), .B(n582), .ZN(n586) );
  NAND2_X1 U659 ( .A1(G56), .A2(n653), .ZN(n584) );
  XOR2_X1 U660 ( .A(KEYINPUT14), .B(n584), .Z(n585) );
  NOR2_X1 U661 ( .A1(n586), .A2(n585), .ZN(n588) );
  NAND2_X1 U662 ( .A1(n652), .A2(G43), .ZN(n587) );
  NAND2_X1 U663 ( .A1(n588), .A2(n587), .ZN(n945) );
  INV_X1 U664 ( .A(G860), .ZN(n610) );
  OR2_X1 U665 ( .A1(n945), .A2(n610), .ZN(G153) );
  NAND2_X1 U666 ( .A1(G52), .A2(n652), .ZN(n589) );
  XOR2_X1 U667 ( .A(KEYINPUT72), .B(n589), .Z(n595) );
  NAND2_X1 U668 ( .A1(G77), .A2(n657), .ZN(n590) );
  XOR2_X1 U669 ( .A(KEYINPUT73), .B(n590), .Z(n592) );
  NAND2_X1 U670 ( .A1(n661), .A2(G90), .ZN(n591) );
  NAND2_X1 U671 ( .A1(n592), .A2(n591), .ZN(n593) );
  XOR2_X1 U672 ( .A(KEYINPUT9), .B(n593), .Z(n594) );
  NOR2_X1 U673 ( .A1(n595), .A2(n594), .ZN(n597) );
  NAND2_X1 U674 ( .A1(G64), .A2(n653), .ZN(n596) );
  NAND2_X1 U675 ( .A1(n597), .A2(n596), .ZN(G301) );
  NAND2_X1 U676 ( .A1(G868), .A2(G301), .ZN(n607) );
  NAND2_X1 U677 ( .A1(n652), .A2(G54), .ZN(n599) );
  NAND2_X1 U678 ( .A1(G79), .A2(n657), .ZN(n598) );
  NAND2_X1 U679 ( .A1(n599), .A2(n598), .ZN(n604) );
  NAND2_X1 U680 ( .A1(n661), .A2(G92), .ZN(n601) );
  NAND2_X1 U681 ( .A1(G66), .A2(n653), .ZN(n600) );
  NAND2_X1 U682 ( .A1(n601), .A2(n600), .ZN(n602) );
  XOR2_X1 U683 ( .A(KEYINPUT77), .B(n602), .Z(n603) );
  NOR2_X1 U684 ( .A1(n604), .A2(n603), .ZN(n605) );
  XOR2_X2 U685 ( .A(KEYINPUT15), .B(n605), .Z(n954) );
  OR2_X1 U686 ( .A1(n954), .A2(G868), .ZN(n606) );
  NAND2_X1 U687 ( .A1(n607), .A2(n606), .ZN(G284) );
  INV_X1 U688 ( .A(G868), .ZN(n672) );
  NOR2_X1 U689 ( .A1(G286), .A2(n672), .ZN(n609) );
  NOR2_X1 U690 ( .A1(G868), .A2(G299), .ZN(n608) );
  NOR2_X1 U691 ( .A1(n609), .A2(n608), .ZN(G297) );
  NAND2_X1 U692 ( .A1(n610), .A2(G559), .ZN(n611) );
  NAND2_X1 U693 ( .A1(n611), .A2(n954), .ZN(n612) );
  XNOR2_X1 U694 ( .A(n612), .B(KEYINPUT80), .ZN(n613) );
  XNOR2_X1 U695 ( .A(KEYINPUT16), .B(n613), .ZN(G148) );
  NOR2_X1 U696 ( .A1(G868), .A2(n945), .ZN(n616) );
  NAND2_X1 U697 ( .A1(G868), .A2(n954), .ZN(n614) );
  NOR2_X1 U698 ( .A1(G559), .A2(n614), .ZN(n615) );
  NOR2_X1 U699 ( .A1(n616), .A2(n615), .ZN(G282) );
  NAND2_X1 U700 ( .A1(G123), .A2(n883), .ZN(n617) );
  XOR2_X1 U701 ( .A(KEYINPUT81), .B(n617), .Z(n618) );
  XNOR2_X1 U702 ( .A(n618), .B(KEYINPUT18), .ZN(n620) );
  NAND2_X1 U703 ( .A1(G111), .A2(n884), .ZN(n619) );
  NAND2_X1 U704 ( .A1(n620), .A2(n619), .ZN(n624) );
  NAND2_X1 U705 ( .A1(G99), .A2(n887), .ZN(n622) );
  NAND2_X1 U706 ( .A1(G135), .A2(n888), .ZN(n621) );
  NAND2_X1 U707 ( .A1(n622), .A2(n621), .ZN(n623) );
  NOR2_X1 U708 ( .A1(n624), .A2(n623), .ZN(n625) );
  XNOR2_X1 U709 ( .A(KEYINPUT82), .B(n625), .ZN(n966) );
  XNOR2_X1 U710 ( .A(n966), .B(G2096), .ZN(n627) );
  INV_X1 U711 ( .A(G2100), .ZN(n626) );
  NAND2_X1 U712 ( .A1(n627), .A2(n626), .ZN(G156) );
  NAND2_X1 U713 ( .A1(n661), .A2(G93), .ZN(n629) );
  NAND2_X1 U714 ( .A1(G67), .A2(n653), .ZN(n628) );
  NAND2_X1 U715 ( .A1(n629), .A2(n628), .ZN(n632) );
  NAND2_X1 U716 ( .A1(G80), .A2(n657), .ZN(n630) );
  XNOR2_X1 U717 ( .A(KEYINPUT83), .B(n630), .ZN(n631) );
  NOR2_X1 U718 ( .A1(n632), .A2(n631), .ZN(n634) );
  NAND2_X1 U719 ( .A1(n652), .A2(G55), .ZN(n633) );
  NAND2_X1 U720 ( .A1(n634), .A2(n633), .ZN(n673) );
  NAND2_X1 U721 ( .A1(n954), .A2(G559), .ZN(n670) );
  XNOR2_X1 U722 ( .A(n945), .B(n670), .ZN(n635) );
  NOR2_X1 U723 ( .A1(G860), .A2(n635), .ZN(n636) );
  XOR2_X1 U724 ( .A(n673), .B(n636), .Z(G145) );
  NAND2_X1 U725 ( .A1(n652), .A2(G48), .ZN(n638) );
  NAND2_X1 U726 ( .A1(G61), .A2(n653), .ZN(n637) );
  NAND2_X1 U727 ( .A1(n638), .A2(n637), .ZN(n641) );
  NAND2_X1 U728 ( .A1(n657), .A2(G73), .ZN(n639) );
  XOR2_X1 U729 ( .A(KEYINPUT2), .B(n639), .Z(n640) );
  NOR2_X1 U730 ( .A1(n641), .A2(n640), .ZN(n643) );
  NAND2_X1 U731 ( .A1(n661), .A2(G86), .ZN(n642) );
  NAND2_X1 U732 ( .A1(n643), .A2(n642), .ZN(G305) );
  NAND2_X1 U733 ( .A1(G87), .A2(n644), .ZN(n645) );
  XNOR2_X1 U734 ( .A(n645), .B(KEYINPUT84), .ZN(n650) );
  NAND2_X1 U735 ( .A1(G49), .A2(n652), .ZN(n647) );
  NAND2_X1 U736 ( .A1(G74), .A2(G651), .ZN(n646) );
  NAND2_X1 U737 ( .A1(n647), .A2(n646), .ZN(n648) );
  NOR2_X1 U738 ( .A1(n653), .A2(n648), .ZN(n649) );
  NAND2_X1 U739 ( .A1(n650), .A2(n649), .ZN(n651) );
  XOR2_X1 U740 ( .A(KEYINPUT85), .B(n651), .Z(G288) );
  NAND2_X1 U741 ( .A1(n652), .A2(G47), .ZN(n656) );
  NAND2_X1 U742 ( .A1(G60), .A2(n653), .ZN(n654) );
  XOR2_X1 U743 ( .A(KEYINPUT71), .B(n654), .Z(n655) );
  NAND2_X1 U744 ( .A1(n656), .A2(n655), .ZN(n660) );
  NAND2_X1 U745 ( .A1(G72), .A2(n657), .ZN(n658) );
  XNOR2_X1 U746 ( .A(KEYINPUT69), .B(n658), .ZN(n659) );
  NOR2_X1 U747 ( .A1(n660), .A2(n659), .ZN(n663) );
  NAND2_X1 U748 ( .A1(n661), .A2(G85), .ZN(n662) );
  NAND2_X1 U749 ( .A1(n663), .A2(n662), .ZN(G290) );
  XOR2_X1 U750 ( .A(G305), .B(G288), .Z(n664) );
  XNOR2_X1 U751 ( .A(n945), .B(n664), .ZN(n665) );
  XNOR2_X1 U752 ( .A(n665), .B(G290), .ZN(n666) );
  XNOR2_X1 U753 ( .A(n666), .B(G299), .ZN(n667) );
  XNOR2_X1 U754 ( .A(n673), .B(n667), .ZN(n669) );
  XNOR2_X1 U755 ( .A(G166), .B(KEYINPUT19), .ZN(n668) );
  XNOR2_X1 U756 ( .A(n669), .B(n668), .ZN(n904) );
  XOR2_X1 U757 ( .A(n904), .B(n670), .Z(n671) );
  NAND2_X1 U758 ( .A1(G868), .A2(n671), .ZN(n675) );
  NAND2_X1 U759 ( .A1(n673), .A2(n672), .ZN(n674) );
  NAND2_X1 U760 ( .A1(n675), .A2(n674), .ZN(G295) );
  NAND2_X1 U761 ( .A1(G2084), .A2(G2078), .ZN(n676) );
  XOR2_X1 U762 ( .A(KEYINPUT20), .B(n676), .Z(n677) );
  NAND2_X1 U763 ( .A1(G2090), .A2(n677), .ZN(n678) );
  XNOR2_X1 U764 ( .A(KEYINPUT21), .B(n678), .ZN(n679) );
  NAND2_X1 U765 ( .A1(n679), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U766 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U767 ( .A(KEYINPUT74), .B(G82), .Z(G220) );
  NAND2_X1 U768 ( .A1(G108), .A2(G120), .ZN(n680) );
  NOR2_X1 U769 ( .A1(G237), .A2(n680), .ZN(n681) );
  NAND2_X1 U770 ( .A1(G69), .A2(n681), .ZN(n840) );
  NAND2_X1 U771 ( .A1(n840), .A2(G567), .ZN(n687) );
  NOR2_X1 U772 ( .A1(G220), .A2(G219), .ZN(n682) );
  XNOR2_X1 U773 ( .A(KEYINPUT22), .B(n682), .ZN(n683) );
  NAND2_X1 U774 ( .A1(n683), .A2(G96), .ZN(n684) );
  NOR2_X1 U775 ( .A1(G218), .A2(n684), .ZN(n685) );
  XOR2_X1 U776 ( .A(KEYINPUT86), .B(n685), .Z(n841) );
  NAND2_X1 U777 ( .A1(G2106), .A2(n841), .ZN(n686) );
  NAND2_X1 U778 ( .A1(n687), .A2(n686), .ZN(n842) );
  NAND2_X1 U779 ( .A1(G483), .A2(G661), .ZN(n688) );
  NOR2_X1 U780 ( .A1(n842), .A2(n688), .ZN(n689) );
  XOR2_X1 U781 ( .A(KEYINPUT87), .B(n689), .Z(n839) );
  NAND2_X1 U782 ( .A1(n839), .A2(G36), .ZN(G176) );
  INV_X1 U783 ( .A(G301), .ZN(G171) );
  INV_X1 U784 ( .A(G166), .ZN(G303) );
  XOR2_X1 U785 ( .A(G2078), .B(KEYINPUT25), .Z(n999) );
  AND2_X1 U786 ( .A1(n690), .A2(G40), .ZN(n692) );
  NAND2_X1 U787 ( .A1(n692), .A2(n691), .ZN(n802) );
  INV_X1 U788 ( .A(n802), .ZN(n693) );
  NOR2_X1 U789 ( .A1(n999), .A2(n746), .ZN(n694) );
  XNOR2_X1 U790 ( .A(n694), .B(KEYINPUT91), .ZN(n696) );
  INV_X1 U791 ( .A(n726), .ZN(n707) );
  OR2_X1 U792 ( .A1(G1961), .A2(n707), .ZN(n695) );
  NAND2_X1 U793 ( .A1(n696), .A2(n695), .ZN(n730) );
  NAND2_X1 U794 ( .A1(n730), .A2(G171), .ZN(n725) );
  NAND2_X1 U795 ( .A1(n707), .A2(G2072), .ZN(n697) );
  XOR2_X1 U796 ( .A(KEYINPUT27), .B(n697), .Z(n699) );
  NAND2_X1 U797 ( .A1(G1956), .A2(n746), .ZN(n698) );
  NAND2_X1 U798 ( .A1(n699), .A2(n698), .ZN(n717) );
  NOR2_X1 U799 ( .A1(G299), .A2(n717), .ZN(n700) );
  XOR2_X1 U800 ( .A(KEYINPUT94), .B(n700), .Z(n716) );
  XOR2_X1 U801 ( .A(KEYINPUT64), .B(KEYINPUT26), .Z(n701) );
  XNOR2_X1 U802 ( .A(n702), .B(n701), .ZN(n704) );
  NAND2_X1 U803 ( .A1(n746), .A2(G1341), .ZN(n703) );
  NAND2_X1 U804 ( .A1(n704), .A2(n703), .ZN(n705) );
  OR2_X1 U805 ( .A1(n954), .A2(n706), .ZN(n714) );
  NAND2_X1 U806 ( .A1(n954), .A2(n706), .ZN(n712) );
  AND2_X1 U807 ( .A1(n707), .A2(G2067), .ZN(n708) );
  XNOR2_X1 U808 ( .A(n708), .B(KEYINPUT93), .ZN(n710) );
  NAND2_X1 U809 ( .A1(n746), .A2(G1348), .ZN(n709) );
  NAND2_X1 U810 ( .A1(n710), .A2(n709), .ZN(n711) );
  NAND2_X1 U811 ( .A1(n712), .A2(n711), .ZN(n713) );
  NAND2_X1 U812 ( .A1(n714), .A2(n713), .ZN(n715) );
  NAND2_X1 U813 ( .A1(n716), .A2(n715), .ZN(n721) );
  NAND2_X1 U814 ( .A1(n717), .A2(G299), .ZN(n718) );
  XNOR2_X1 U815 ( .A(n718), .B(KEYINPUT92), .ZN(n719) );
  XNOR2_X1 U816 ( .A(KEYINPUT28), .B(n719), .ZN(n720) );
  NAND2_X1 U817 ( .A1(n721), .A2(n720), .ZN(n723) );
  NAND2_X1 U818 ( .A1(n725), .A2(n724), .ZN(n737) );
  NOR2_X1 U819 ( .A1(G2084), .A2(n746), .ZN(n741) );
  NAND2_X1 U820 ( .A1(G8), .A2(n726), .ZN(n780) );
  NOR2_X1 U821 ( .A1(G1966), .A2(n780), .ZN(n738) );
  NOR2_X1 U822 ( .A1(n741), .A2(n738), .ZN(n727) );
  NAND2_X1 U823 ( .A1(G8), .A2(n727), .ZN(n728) );
  XNOR2_X1 U824 ( .A(n728), .B(KEYINPUT95), .ZN(n729) );
  NOR2_X1 U825 ( .A1(G168), .A2(n515), .ZN(n732) );
  NOR2_X1 U826 ( .A1(G171), .A2(n730), .ZN(n731) );
  NOR2_X1 U827 ( .A1(n732), .A2(n731), .ZN(n735) );
  XNOR2_X1 U828 ( .A(n735), .B(n734), .ZN(n736) );
  NAND2_X1 U829 ( .A1(n737), .A2(n736), .ZN(n744) );
  XNOR2_X1 U830 ( .A(n740), .B(KEYINPUT98), .ZN(n743) );
  NAND2_X1 U831 ( .A1(n741), .A2(G8), .ZN(n742) );
  NAND2_X1 U832 ( .A1(n743), .A2(n742), .ZN(n770) );
  XOR2_X1 U833 ( .A(KEYINPUT32), .B(KEYINPUT101), .Z(n755) );
  NAND2_X1 U834 ( .A1(n744), .A2(G286), .ZN(n752) );
  NOR2_X1 U835 ( .A1(G1971), .A2(n780), .ZN(n745) );
  XNOR2_X1 U836 ( .A(KEYINPUT99), .B(n745), .ZN(n749) );
  NOR2_X1 U837 ( .A1(G2090), .A2(n746), .ZN(n747) );
  NOR2_X1 U838 ( .A1(G166), .A2(n747), .ZN(n748) );
  NAND2_X1 U839 ( .A1(n749), .A2(n748), .ZN(n750) );
  XNOR2_X1 U840 ( .A(n750), .B(KEYINPUT100), .ZN(n751) );
  NAND2_X1 U841 ( .A1(n752), .A2(n751), .ZN(n753) );
  NAND2_X1 U842 ( .A1(G8), .A2(n753), .ZN(n754) );
  XNOR2_X1 U843 ( .A(n755), .B(n754), .ZN(n769) );
  NAND2_X1 U844 ( .A1(G1976), .A2(G288), .ZN(n948) );
  INV_X1 U845 ( .A(n948), .ZN(n756) );
  OR2_X1 U846 ( .A1(n780), .A2(n756), .ZN(n760) );
  INV_X1 U847 ( .A(n760), .ZN(n757) );
  AND2_X1 U848 ( .A1(n769), .A2(n757), .ZN(n758) );
  NAND2_X1 U849 ( .A1(n770), .A2(n758), .ZN(n762) );
  NOR2_X1 U850 ( .A1(G1976), .A2(G288), .ZN(n764) );
  NOR2_X1 U851 ( .A1(G1971), .A2(G303), .ZN(n759) );
  NOR2_X1 U852 ( .A1(n764), .A2(n759), .ZN(n957) );
  OR2_X1 U853 ( .A1(n760), .A2(n957), .ZN(n761) );
  NAND2_X1 U854 ( .A1(n762), .A2(n761), .ZN(n763) );
  NOR2_X1 U855 ( .A1(KEYINPUT33), .A2(n763), .ZN(n767) );
  NAND2_X1 U856 ( .A1(n764), .A2(KEYINPUT33), .ZN(n765) );
  NOR2_X1 U857 ( .A1(n765), .A2(n780), .ZN(n766) );
  NOR2_X1 U858 ( .A1(n767), .A2(n766), .ZN(n768) );
  XOR2_X1 U859 ( .A(G1981), .B(G305), .Z(n940) );
  NAND2_X1 U860 ( .A1(n768), .A2(n940), .ZN(n777) );
  NAND2_X1 U861 ( .A1(n770), .A2(n769), .ZN(n773) );
  NOR2_X1 U862 ( .A1(G2090), .A2(G303), .ZN(n771) );
  NAND2_X1 U863 ( .A1(G8), .A2(n771), .ZN(n772) );
  NAND2_X1 U864 ( .A1(n773), .A2(n772), .ZN(n774) );
  NAND2_X1 U865 ( .A1(n780), .A2(n774), .ZN(n775) );
  XNOR2_X1 U866 ( .A(n775), .B(KEYINPUT102), .ZN(n776) );
  NAND2_X1 U867 ( .A1(n777), .A2(n776), .ZN(n782) );
  NOR2_X1 U868 ( .A1(G1981), .A2(G305), .ZN(n778) );
  XOR2_X1 U869 ( .A(n778), .B(KEYINPUT24), .Z(n779) );
  NOR2_X1 U870 ( .A1(n780), .A2(n779), .ZN(n781) );
  NAND2_X1 U871 ( .A1(n883), .A2(G129), .ZN(n791) );
  NAND2_X1 U872 ( .A1(G141), .A2(n888), .ZN(n786) );
  NAND2_X1 U873 ( .A1(G117), .A2(n884), .ZN(n785) );
  NAND2_X1 U874 ( .A1(n786), .A2(n785), .ZN(n789) );
  NAND2_X1 U875 ( .A1(n887), .A2(G105), .ZN(n787) );
  XOR2_X1 U876 ( .A(KEYINPUT38), .B(n787), .Z(n788) );
  NOR2_X1 U877 ( .A1(n789), .A2(n788), .ZN(n790) );
  NAND2_X1 U878 ( .A1(n791), .A2(n790), .ZN(n792) );
  XOR2_X1 U879 ( .A(KEYINPUT89), .B(n792), .Z(n871) );
  NAND2_X1 U880 ( .A1(G1996), .A2(n871), .ZN(n793) );
  XOR2_X1 U881 ( .A(KEYINPUT90), .B(n793), .Z(n801) );
  NAND2_X1 U882 ( .A1(G95), .A2(n887), .ZN(n795) );
  NAND2_X1 U883 ( .A1(G131), .A2(n888), .ZN(n794) );
  NAND2_X1 U884 ( .A1(n795), .A2(n794), .ZN(n799) );
  NAND2_X1 U885 ( .A1(G119), .A2(n883), .ZN(n797) );
  NAND2_X1 U886 ( .A1(G107), .A2(n884), .ZN(n796) );
  NAND2_X1 U887 ( .A1(n797), .A2(n796), .ZN(n798) );
  NOR2_X1 U888 ( .A1(n799), .A2(n798), .ZN(n896) );
  INV_X1 U889 ( .A(G1991), .ZN(n994) );
  NOR2_X1 U890 ( .A1(n896), .A2(n994), .ZN(n800) );
  NOR2_X1 U891 ( .A1(n801), .A2(n800), .ZN(n982) );
  NOR2_X1 U892 ( .A1(n803), .A2(n802), .ZN(n830) );
  INV_X1 U893 ( .A(n830), .ZN(n804) );
  NOR2_X1 U894 ( .A1(n982), .A2(n804), .ZN(n821) );
  INV_X1 U895 ( .A(n821), .ZN(n814) );
  NAND2_X1 U896 ( .A1(G104), .A2(n887), .ZN(n806) );
  NAND2_X1 U897 ( .A1(G140), .A2(n888), .ZN(n805) );
  NAND2_X1 U898 ( .A1(n806), .A2(n805), .ZN(n807) );
  XNOR2_X1 U899 ( .A(KEYINPUT34), .B(n807), .ZN(n812) );
  NAND2_X1 U900 ( .A1(G128), .A2(n883), .ZN(n809) );
  NAND2_X1 U901 ( .A1(G116), .A2(n884), .ZN(n808) );
  NAND2_X1 U902 ( .A1(n809), .A2(n808), .ZN(n810) );
  XOR2_X1 U903 ( .A(KEYINPUT35), .B(n810), .Z(n811) );
  NOR2_X1 U904 ( .A1(n812), .A2(n811), .ZN(n813) );
  XNOR2_X1 U905 ( .A(KEYINPUT36), .B(n813), .ZN(n900) );
  XNOR2_X1 U906 ( .A(KEYINPUT37), .B(G2067), .ZN(n828) );
  NOR2_X1 U907 ( .A1(n900), .A2(n828), .ZN(n971) );
  NAND2_X1 U908 ( .A1(n830), .A2(n971), .ZN(n826) );
  XNOR2_X1 U909 ( .A(G1986), .B(G290), .ZN(n956) );
  NAND2_X1 U910 ( .A1(n956), .A2(n830), .ZN(n815) );
  OR2_X1 U911 ( .A1(n817), .A2(n816), .ZN(n833) );
  XNOR2_X1 U912 ( .A(KEYINPUT39), .B(KEYINPUT105), .ZN(n824) );
  NOR2_X1 U913 ( .A1(G1986), .A2(G290), .ZN(n818) );
  AND2_X1 U914 ( .A1(n994), .A2(n896), .ZN(n967) );
  NOR2_X1 U915 ( .A1(n818), .A2(n967), .ZN(n819) );
  XNOR2_X1 U916 ( .A(n819), .B(KEYINPUT104), .ZN(n820) );
  NOR2_X1 U917 ( .A1(n821), .A2(n820), .ZN(n822) );
  NOR2_X1 U918 ( .A1(G1996), .A2(n871), .ZN(n984) );
  NOR2_X1 U919 ( .A1(n822), .A2(n984), .ZN(n823) );
  XOR2_X1 U920 ( .A(n824), .B(n823), .Z(n825) );
  NAND2_X1 U921 ( .A1(n826), .A2(n825), .ZN(n827) );
  XNOR2_X1 U922 ( .A(n827), .B(KEYINPUT106), .ZN(n829) );
  NAND2_X1 U923 ( .A1(n900), .A2(n828), .ZN(n968) );
  NAND2_X1 U924 ( .A1(n829), .A2(n968), .ZN(n831) );
  NAND2_X1 U925 ( .A1(n831), .A2(n830), .ZN(n832) );
  NAND2_X1 U926 ( .A1(n833), .A2(n832), .ZN(n835) );
  XOR2_X1 U927 ( .A(KEYINPUT40), .B(KEYINPUT107), .Z(n834) );
  XNOR2_X1 U928 ( .A(n835), .B(n834), .ZN(G329) );
  NAND2_X1 U929 ( .A1(G2106), .A2(n836), .ZN(G217) );
  AND2_X1 U930 ( .A1(G15), .A2(G2), .ZN(n837) );
  NAND2_X1 U931 ( .A1(G661), .A2(n837), .ZN(G259) );
  NAND2_X1 U932 ( .A1(G3), .A2(G1), .ZN(n838) );
  NAND2_X1 U933 ( .A1(n839), .A2(n838), .ZN(G188) );
  XNOR2_X1 U934 ( .A(G120), .B(KEYINPUT109), .ZN(G236) );
  INV_X1 U936 ( .A(G108), .ZN(G238) );
  INV_X1 U937 ( .A(G96), .ZN(G221) );
  NOR2_X1 U938 ( .A1(n841), .A2(n840), .ZN(G325) );
  INV_X1 U939 ( .A(G325), .ZN(G261) );
  INV_X1 U940 ( .A(n842), .ZN(G319) );
  XOR2_X1 U941 ( .A(G2100), .B(G2096), .Z(n844) );
  XNOR2_X1 U942 ( .A(KEYINPUT42), .B(G2678), .ZN(n843) );
  XNOR2_X1 U943 ( .A(n844), .B(n843), .ZN(n848) );
  XOR2_X1 U944 ( .A(KEYINPUT43), .B(G2090), .Z(n846) );
  XNOR2_X1 U945 ( .A(G2067), .B(G2072), .ZN(n845) );
  XNOR2_X1 U946 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U947 ( .A(n848), .B(n847), .Z(n850) );
  XNOR2_X1 U948 ( .A(G2084), .B(G2078), .ZN(n849) );
  XNOR2_X1 U949 ( .A(n850), .B(n849), .ZN(G227) );
  XNOR2_X1 U950 ( .A(G1996), .B(KEYINPUT110), .ZN(n860) );
  XOR2_X1 U951 ( .A(G1956), .B(G1961), .Z(n852) );
  XNOR2_X1 U952 ( .A(G1991), .B(G1981), .ZN(n851) );
  XNOR2_X1 U953 ( .A(n852), .B(n851), .ZN(n856) );
  XOR2_X1 U954 ( .A(G1966), .B(G1971), .Z(n854) );
  XNOR2_X1 U955 ( .A(G1986), .B(G1976), .ZN(n853) );
  XNOR2_X1 U956 ( .A(n854), .B(n853), .ZN(n855) );
  XOR2_X1 U957 ( .A(n856), .B(n855), .Z(n858) );
  XNOR2_X1 U958 ( .A(G2474), .B(KEYINPUT41), .ZN(n857) );
  XNOR2_X1 U959 ( .A(n858), .B(n857), .ZN(n859) );
  XNOR2_X1 U960 ( .A(n860), .B(n859), .ZN(G229) );
  NAND2_X1 U961 ( .A1(G100), .A2(n887), .ZN(n862) );
  NAND2_X1 U962 ( .A1(G112), .A2(n884), .ZN(n861) );
  NAND2_X1 U963 ( .A1(n862), .A2(n861), .ZN(n870) );
  NAND2_X1 U964 ( .A1(n888), .A2(G136), .ZN(n863) );
  XNOR2_X1 U965 ( .A(KEYINPUT112), .B(n863), .ZN(n867) );
  XOR2_X1 U966 ( .A(KEYINPUT111), .B(KEYINPUT44), .Z(n865) );
  NAND2_X1 U967 ( .A1(G124), .A2(n883), .ZN(n864) );
  XNOR2_X1 U968 ( .A(n865), .B(n864), .ZN(n866) );
  NAND2_X1 U969 ( .A1(n867), .A2(n866), .ZN(n868) );
  XOR2_X1 U970 ( .A(KEYINPUT113), .B(n868), .Z(n869) );
  NOR2_X1 U971 ( .A1(n870), .A2(n869), .ZN(G162) );
  XNOR2_X1 U972 ( .A(G162), .B(n871), .ZN(n872) );
  XNOR2_X1 U973 ( .A(n872), .B(n966), .ZN(n880) );
  NAND2_X1 U974 ( .A1(G103), .A2(n887), .ZN(n874) );
  NAND2_X1 U975 ( .A1(G139), .A2(n888), .ZN(n873) );
  NAND2_X1 U976 ( .A1(n874), .A2(n873), .ZN(n879) );
  NAND2_X1 U977 ( .A1(G127), .A2(n883), .ZN(n876) );
  NAND2_X1 U978 ( .A1(G115), .A2(n884), .ZN(n875) );
  NAND2_X1 U979 ( .A1(n876), .A2(n875), .ZN(n877) );
  XOR2_X1 U980 ( .A(KEYINPUT47), .B(n877), .Z(n878) );
  NOR2_X1 U981 ( .A1(n879), .A2(n878), .ZN(n974) );
  XOR2_X1 U982 ( .A(n880), .B(n974), .Z(n882) );
  XNOR2_X1 U983 ( .A(G164), .B(G160), .ZN(n881) );
  XNOR2_X1 U984 ( .A(n882), .B(n881), .ZN(n902) );
  XOR2_X1 U985 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n898) );
  NAND2_X1 U986 ( .A1(G130), .A2(n883), .ZN(n886) );
  NAND2_X1 U987 ( .A1(G118), .A2(n884), .ZN(n885) );
  NAND2_X1 U988 ( .A1(n886), .A2(n885), .ZN(n894) );
  NAND2_X1 U989 ( .A1(G106), .A2(n887), .ZN(n890) );
  NAND2_X1 U990 ( .A1(G142), .A2(n888), .ZN(n889) );
  NAND2_X1 U991 ( .A1(n890), .A2(n889), .ZN(n891) );
  XOR2_X1 U992 ( .A(KEYINPUT45), .B(n891), .Z(n892) );
  XNOR2_X1 U993 ( .A(KEYINPUT114), .B(n892), .ZN(n893) );
  NOR2_X1 U994 ( .A1(n894), .A2(n893), .ZN(n895) );
  XNOR2_X1 U995 ( .A(n896), .B(n895), .ZN(n897) );
  XNOR2_X1 U996 ( .A(n898), .B(n897), .ZN(n899) );
  XOR2_X1 U997 ( .A(n900), .B(n899), .Z(n901) );
  XNOR2_X1 U998 ( .A(n902), .B(n901), .ZN(n903) );
  NOR2_X1 U999 ( .A1(G37), .A2(n903), .ZN(G395) );
  XNOR2_X1 U1000 ( .A(n954), .B(G286), .ZN(n905) );
  XNOR2_X1 U1001 ( .A(n905), .B(n904), .ZN(n906) );
  XNOR2_X1 U1002 ( .A(n906), .B(G171), .ZN(n907) );
  NOR2_X1 U1003 ( .A1(G37), .A2(n907), .ZN(G397) );
  NOR2_X1 U1004 ( .A1(G227), .A2(G229), .ZN(n908) );
  XOR2_X1 U1005 ( .A(KEYINPUT49), .B(n908), .Z(n909) );
  NAND2_X1 U1006 ( .A1(G319), .A2(n909), .ZN(n910) );
  NOR2_X1 U1007 ( .A1(G401), .A2(n910), .ZN(n911) );
  XOR2_X1 U1008 ( .A(KEYINPUT115), .B(n911), .Z(n914) );
  NOR2_X1 U1009 ( .A1(G395), .A2(G397), .ZN(n912) );
  XNOR2_X1 U1010 ( .A(KEYINPUT116), .B(n912), .ZN(n913) );
  NAND2_X1 U1011 ( .A1(n914), .A2(n913), .ZN(G225) );
  INV_X1 U1012 ( .A(G225), .ZN(G308) );
  INV_X1 U1013 ( .A(G69), .ZN(G235) );
  XOR2_X1 U1014 ( .A(KEYINPUT123), .B(G4), .Z(n916) );
  XNOR2_X1 U1015 ( .A(G1348), .B(KEYINPUT59), .ZN(n915) );
  XNOR2_X1 U1016 ( .A(n916), .B(n915), .ZN(n920) );
  XNOR2_X1 U1017 ( .A(G1981), .B(G6), .ZN(n918) );
  XNOR2_X1 U1018 ( .A(G19), .B(G1341), .ZN(n917) );
  NOR2_X1 U1019 ( .A1(n918), .A2(n917), .ZN(n919) );
  NAND2_X1 U1020 ( .A1(n920), .A2(n919), .ZN(n923) );
  XNOR2_X1 U1021 ( .A(KEYINPUT122), .B(G1956), .ZN(n921) );
  XNOR2_X1 U1022 ( .A(G20), .B(n921), .ZN(n922) );
  NOR2_X1 U1023 ( .A1(n923), .A2(n922), .ZN(n924) );
  XNOR2_X1 U1024 ( .A(KEYINPUT60), .B(n924), .ZN(n925) );
  XNOR2_X1 U1025 ( .A(n925), .B(KEYINPUT124), .ZN(n929) );
  XNOR2_X1 U1026 ( .A(G1966), .B(G21), .ZN(n927) );
  XNOR2_X1 U1027 ( .A(G1961), .B(G5), .ZN(n926) );
  NOR2_X1 U1028 ( .A1(n927), .A2(n926), .ZN(n928) );
  NAND2_X1 U1029 ( .A1(n929), .A2(n928), .ZN(n937) );
  XNOR2_X1 U1030 ( .A(G1986), .B(G24), .ZN(n931) );
  XNOR2_X1 U1031 ( .A(G22), .B(G1971), .ZN(n930) );
  NOR2_X1 U1032 ( .A1(n931), .A2(n930), .ZN(n934) );
  XNOR2_X1 U1033 ( .A(G1976), .B(KEYINPUT125), .ZN(n932) );
  XNOR2_X1 U1034 ( .A(n932), .B(G23), .ZN(n933) );
  NAND2_X1 U1035 ( .A1(n934), .A2(n933), .ZN(n935) );
  XNOR2_X1 U1036 ( .A(KEYINPUT58), .B(n935), .ZN(n936) );
  NOR2_X1 U1037 ( .A1(n937), .A2(n936), .ZN(n938) );
  XOR2_X1 U1038 ( .A(KEYINPUT61), .B(n938), .Z(n939) );
  NOR2_X1 U1039 ( .A1(G16), .A2(n939), .ZN(n964) );
  XOR2_X1 U1040 ( .A(G16), .B(KEYINPUT56), .Z(n962) );
  XNOR2_X1 U1041 ( .A(G1966), .B(G168), .ZN(n941) );
  NAND2_X1 U1042 ( .A1(n941), .A2(n940), .ZN(n942) );
  XNOR2_X1 U1043 ( .A(n942), .B(KEYINPUT57), .ZN(n953) );
  NAND2_X1 U1044 ( .A1(G1971), .A2(G303), .ZN(n944) );
  XOR2_X1 U1045 ( .A(G1956), .B(G299), .Z(n943) );
  NAND2_X1 U1046 ( .A1(n944), .A2(n943), .ZN(n947) );
  XNOR2_X1 U1047 ( .A(G1341), .B(n945), .ZN(n946) );
  NOR2_X1 U1048 ( .A1(n947), .A2(n946), .ZN(n949) );
  NAND2_X1 U1049 ( .A1(n949), .A2(n948), .ZN(n951) );
  XNOR2_X1 U1050 ( .A(G1961), .B(G301), .ZN(n950) );
  NOR2_X1 U1051 ( .A1(n951), .A2(n950), .ZN(n952) );
  NAND2_X1 U1052 ( .A1(n953), .A2(n952), .ZN(n960) );
  XOR2_X1 U1053 ( .A(G1348), .B(n954), .Z(n955) );
  NOR2_X1 U1054 ( .A1(n956), .A2(n955), .ZN(n958) );
  NAND2_X1 U1055 ( .A1(n958), .A2(n957), .ZN(n959) );
  NOR2_X1 U1056 ( .A1(n960), .A2(n959), .ZN(n961) );
  NOR2_X1 U1057 ( .A1(n962), .A2(n961), .ZN(n963) );
  NOR2_X1 U1058 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1059 ( .A(n965), .B(KEYINPUT126), .ZN(n993) );
  NOR2_X1 U1060 ( .A1(n967), .A2(n966), .ZN(n973) );
  XNOR2_X1 U1061 ( .A(G2084), .B(G160), .ZN(n969) );
  NAND2_X1 U1062 ( .A1(n969), .A2(n968), .ZN(n970) );
  NOR2_X1 U1063 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1064 ( .A1(n973), .A2(n972), .ZN(n980) );
  XNOR2_X1 U1065 ( .A(G2072), .B(n974), .ZN(n976) );
  XNOR2_X1 U1066 ( .A(G164), .B(G2078), .ZN(n975) );
  NAND2_X1 U1067 ( .A1(n976), .A2(n975), .ZN(n977) );
  XOR2_X1 U1068 ( .A(KEYINPUT50), .B(n977), .Z(n978) );
  XNOR2_X1 U1069 ( .A(KEYINPUT117), .B(n978), .ZN(n979) );
  NOR2_X1 U1070 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1071 ( .A1(n982), .A2(n981), .ZN(n987) );
  XOR2_X1 U1072 ( .A(G2090), .B(G162), .Z(n983) );
  NOR2_X1 U1073 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1074 ( .A(n985), .B(KEYINPUT51), .ZN(n986) );
  NOR2_X1 U1075 ( .A1(n987), .A2(n986), .ZN(n988) );
  XNOR2_X1 U1076 ( .A(KEYINPUT52), .B(n988), .ZN(n990) );
  INV_X1 U1077 ( .A(KEYINPUT55), .ZN(n989) );
  NAND2_X1 U1078 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1079 ( .A1(n991), .A2(G29), .ZN(n992) );
  NAND2_X1 U1080 ( .A1(n993), .A2(n992), .ZN(n1020) );
  XOR2_X1 U1081 ( .A(G2090), .B(G35), .Z(n1010) );
  XNOR2_X1 U1082 ( .A(G25), .B(n994), .ZN(n995) );
  NAND2_X1 U1083 ( .A1(n995), .A2(G28), .ZN(n996) );
  XNOR2_X1 U1084 ( .A(KEYINPUT118), .B(n996), .ZN(n1006) );
  XNOR2_X1 U1085 ( .A(G2067), .B(G26), .ZN(n998) );
  XNOR2_X1 U1086 ( .A(G1996), .B(G32), .ZN(n997) );
  NOR2_X1 U1087 ( .A1(n998), .A2(n997), .ZN(n1003) );
  XNOR2_X1 U1088 ( .A(n999), .B(G27), .ZN(n1001) );
  XNOR2_X1 U1089 ( .A(G33), .B(G2072), .ZN(n1000) );
  NOR2_X1 U1090 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1091 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XOR2_X1 U1092 ( .A(n1004), .B(KEYINPUT119), .Z(n1005) );
  NOR2_X1 U1093 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XOR2_X1 U1094 ( .A(KEYINPUT53), .B(n1007), .Z(n1008) );
  XNOR2_X1 U1095 ( .A(n1008), .B(KEYINPUT120), .ZN(n1009) );
  NAND2_X1 U1096 ( .A1(n1010), .A2(n1009), .ZN(n1013) );
  XNOR2_X1 U1097 ( .A(G34), .B(G2084), .ZN(n1011) );
  XNOR2_X1 U1098 ( .A(KEYINPUT54), .B(n1011), .ZN(n1012) );
  NOR2_X1 U1099 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1100 ( .A(KEYINPUT55), .B(n1014), .ZN(n1016) );
  INV_X1 U1101 ( .A(G29), .ZN(n1015) );
  NAND2_X1 U1102 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1103 ( .A1(n1017), .A2(G11), .ZN(n1018) );
  XOR2_X1 U1104 ( .A(KEYINPUT121), .B(n1018), .Z(n1019) );
  NOR2_X1 U1105 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1106 ( .A(KEYINPUT62), .B(n1021), .ZN(G311) );
  INV_X1 U1107 ( .A(G311), .ZN(G150) );
endmodule

