//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 0 1 1 1 1 0 0 1 0 0 1 1 1 0 0 1 1 0 0 0 0 0 1 0 0 1 0 0 0 1 1 1 1 0 1 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:29 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n766,
    new_n767, new_n768, new_n769, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n786, new_n787, new_n789, new_n790,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n803, new_n804, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n819, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1040, new_n1041,
    new_n1042, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1061, new_n1062, new_n1063, new_n1064, new_n1065, new_n1066,
    new_n1067, new_n1068, new_n1069, new_n1070, new_n1071, new_n1072,
    new_n1073, new_n1074, new_n1075, new_n1076, new_n1077, new_n1078,
    new_n1080, new_n1081, new_n1082, new_n1083, new_n1084, new_n1085,
    new_n1086, new_n1087, new_n1088, new_n1089, new_n1090, new_n1091,
    new_n1092;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT76), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G469), .ZN(new_n191));
  INV_X1    g005(.A(G902), .ZN(new_n192));
  XNOR2_X1  g006(.A(G110), .B(G140), .ZN(new_n193));
  INV_X1    g007(.A(G953), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G227), .ZN(new_n195));
  XOR2_X1   g009(.A(new_n193), .B(new_n195), .Z(new_n196));
  INV_X1    g010(.A(KEYINPUT64), .ZN(new_n197));
  INV_X1    g011(.A(G143), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(KEYINPUT64), .A2(G143), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n199), .A2(G146), .A3(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G146), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G143), .ZN(new_n203));
  INV_X1    g017(.A(G128), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n204), .A2(KEYINPUT1), .ZN(new_n205));
  AND3_X1   g019(.A1(new_n201), .A2(new_n203), .A3(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(new_n203), .ZN(new_n207));
  AND2_X1   g021(.A1(KEYINPUT64), .A2(G143), .ZN(new_n208));
  NOR2_X1   g022(.A1(KEYINPUT64), .A2(G143), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n207), .B1(new_n210), .B2(G146), .ZN(new_n211));
  INV_X1    g025(.A(new_n211), .ZN(new_n212));
  AOI21_X1  g026(.A(G146), .B1(new_n199), .B2(new_n200), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT1), .ZN(new_n214));
  OAI21_X1  g028(.A(G128), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n206), .B1(new_n212), .B2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G107), .ZN(new_n217));
  OAI21_X1  g031(.A(KEYINPUT77), .B1(new_n217), .B2(G104), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT77), .ZN(new_n219));
  INV_X1    g033(.A(G104), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n219), .A2(new_n220), .A3(G107), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n217), .A2(G104), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n218), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(G101), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n217), .A2(G104), .ZN(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G101), .ZN(new_n227));
  AND3_X1   g041(.A1(new_n217), .A2(KEYINPUT3), .A3(G104), .ZN(new_n228));
  AOI21_X1  g042(.A(KEYINPUT3), .B1(new_n217), .B2(G104), .ZN(new_n229));
  OAI211_X1 g043(.A(new_n226), .B(new_n227), .C1(new_n228), .C2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n224), .A2(new_n230), .ZN(new_n231));
  OAI21_X1  g045(.A(KEYINPUT78), .B1(new_n216), .B2(new_n231), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n201), .A2(new_n203), .A3(new_n205), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n202), .B1(new_n208), .B2(new_n209), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n204), .B1(new_n234), .B2(KEYINPUT1), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n233), .B1(new_n235), .B2(new_n211), .ZN(new_n236));
  AND2_X1   g050(.A1(new_n224), .A2(new_n230), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT78), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n236), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  AOI21_X1  g053(.A(KEYINPUT10), .B1(new_n232), .B2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(G137), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n241), .A2(KEYINPUT11), .A3(G134), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT11), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G137), .ZN(new_n244));
  AND2_X1   g058(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(G131), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n241), .A2(KEYINPUT11), .ZN(new_n247));
  INV_X1    g061(.A(G134), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(KEYINPUT65), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT65), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(G134), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n247), .A2(new_n249), .A3(new_n251), .ZN(new_n252));
  AND3_X1   g066(.A1(new_n245), .A2(new_n246), .A3(new_n252), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n246), .B1(new_n245), .B2(new_n252), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  XNOR2_X1  g070(.A(KEYINPUT0), .B(G128), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n198), .A2(G146), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n257), .B1(new_n234), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(KEYINPUT0), .A2(G128), .ZN(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n259), .B1(new_n211), .B2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT4), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT3), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n264), .B1(new_n220), .B2(G107), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n217), .A2(KEYINPUT3), .A3(G104), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n225), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n263), .B1(new_n267), .B2(new_n227), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n226), .B1(new_n228), .B2(new_n229), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(G101), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n269), .A2(new_n263), .A3(G101), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n262), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n234), .A2(new_n258), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n204), .B1(new_n203), .B2(KEYINPUT1), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(new_n233), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n278), .A2(new_n237), .A3(KEYINPUT10), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n273), .A2(new_n279), .ZN(new_n280));
  NOR3_X1   g094(.A1(new_n240), .A2(new_n256), .A3(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT10), .ZN(new_n282));
  AND3_X1   g096(.A1(new_n236), .A2(new_n237), .A3(new_n238), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n238), .B1(new_n236), .B2(new_n237), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n282), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(new_n280), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n255), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  OAI211_X1 g101(.A(KEYINPUT81), .B(new_n196), .C1(new_n281), .C2(new_n287), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n278), .A2(new_n237), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n289), .B1(new_n232), .B2(new_n239), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n255), .A2(KEYINPUT79), .ZN(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(KEYINPUT12), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT12), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n283), .A2(new_n284), .ZN(new_n295));
  OAI211_X1 g109(.A(new_n294), .B(new_n291), .C1(new_n295), .C2(new_n289), .ZN(new_n296));
  INV_X1    g110(.A(new_n196), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n285), .A2(new_n286), .A3(new_n255), .ZN(new_n298));
  NAND4_X1  g112(.A1(new_n293), .A2(new_n296), .A3(new_n297), .A4(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n288), .A2(new_n299), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n256), .B1(new_n240), .B2(new_n280), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(new_n298), .ZN(new_n302));
  AOI21_X1  g116(.A(KEYINPUT81), .B1(new_n302), .B2(new_n196), .ZN(new_n303));
  OAI211_X1 g117(.A(new_n191), .B(new_n192), .C1(new_n300), .C2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n293), .A2(new_n296), .A3(new_n298), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(new_n196), .ZN(new_n307));
  AOI21_X1  g121(.A(KEYINPUT80), .B1(new_n298), .B2(new_n297), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n298), .A2(KEYINPUT80), .A3(new_n297), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(new_n301), .ZN(new_n310));
  OAI211_X1 g124(.A(new_n307), .B(G469), .C1(new_n308), .C2(new_n310), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n191), .A2(new_n192), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n190), .B1(new_n305), .B2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT82), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n304), .A2(new_n313), .A3(new_n311), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n318), .A2(KEYINPUT82), .A3(new_n190), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  XNOR2_X1  g134(.A(G110), .B(G122), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(G119), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G116), .ZN(new_n324));
  INV_X1    g138(.A(G116), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(G119), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  XNOR2_X1  g141(.A(KEYINPUT2), .B(G113), .ZN(new_n328));
  OR2_X1    g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n329), .A2(new_n224), .A3(new_n230), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT5), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT66), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n325), .A2(G119), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n323), .A2(G116), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n332), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n324), .A2(new_n326), .A3(KEYINPUT66), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n331), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  OAI21_X1  g151(.A(G113), .B1(new_n324), .B2(KEYINPUT5), .ZN(new_n338));
  OAI21_X1  g152(.A(KEYINPUT84), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  AND3_X1   g153(.A1(new_n324), .A2(new_n326), .A3(KEYINPUT66), .ZN(new_n340));
  AOI21_X1  g154(.A(KEYINPUT66), .B1(new_n324), .B2(new_n326), .ZN(new_n341));
  OAI21_X1  g155(.A(KEYINPUT5), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT84), .ZN(new_n343));
  INV_X1    g157(.A(new_n338), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n342), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n330), .B1(new_n339), .B2(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n335), .A2(new_n328), .A3(new_n336), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(new_n329), .ZN(new_n348));
  AND3_X1   g162(.A1(new_n271), .A2(new_n348), .A3(new_n272), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n322), .B1(new_n346), .B2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n330), .ZN(new_n351));
  NOR3_X1   g165(.A1(new_n337), .A2(KEYINPUT84), .A3(new_n338), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n343), .B1(new_n342), .B2(new_n344), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n351), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n271), .A2(new_n348), .A3(new_n272), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n354), .A2(new_n355), .A3(new_n321), .ZN(new_n356));
  NAND4_X1  g170(.A1(new_n350), .A2(new_n356), .A3(KEYINPUT85), .A4(KEYINPUT6), .ZN(new_n357));
  AND3_X1   g171(.A1(new_n350), .A2(new_n356), .A3(KEYINPUT6), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT6), .ZN(new_n359));
  OAI211_X1 g173(.A(new_n359), .B(new_n322), .C1(new_n346), .C2(new_n349), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT85), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n357), .B1(new_n358), .B2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n259), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n211), .A2(new_n261), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(G125), .ZN(new_n367));
  INV_X1    g181(.A(G125), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n277), .A2(new_n368), .A3(new_n233), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(G224), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n371), .A2(G953), .ZN(new_n372));
  XNOR2_X1  g186(.A(new_n372), .B(KEYINPUT86), .ZN(new_n373));
  XNOR2_X1  g187(.A(new_n370), .B(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n363), .A2(new_n375), .ZN(new_n376));
  OAI21_X1  g190(.A(G210), .B1(G237), .B2(G902), .ZN(new_n377));
  OAI21_X1  g191(.A(KEYINPUT7), .B1(new_n371), .B2(G953), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  OAI211_X1 g193(.A(new_n369), .B(new_n379), .C1(new_n262), .C2(new_n368), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(KEYINPUT89), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT89), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n367), .A2(new_n382), .A3(new_n369), .A4(new_n379), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  OAI211_X1 g198(.A(KEYINPUT88), .B(new_n369), .C1(new_n262), .C2(new_n368), .ZN(new_n385));
  OAI211_X1 g199(.A(new_n385), .B(new_n378), .C1(KEYINPUT88), .C2(new_n369), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n384), .A2(new_n356), .A3(new_n386), .ZN(new_n387));
  XNOR2_X1  g201(.A(new_n321), .B(KEYINPUT8), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n329), .B1(new_n352), .B2(new_n353), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(new_n231), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT87), .ZN(new_n392));
  NOR3_X1   g206(.A1(new_n327), .A2(new_n392), .A3(new_n331), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n392), .B1(new_n327), .B2(new_n331), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(new_n344), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n351), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n389), .B1(new_n391), .B2(new_n396), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n192), .B1(new_n387), .B2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n376), .A2(new_n377), .A3(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(new_n377), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n350), .A2(new_n356), .A3(KEYINPUT6), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n402), .A2(new_n361), .A3(new_n360), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n374), .B1(new_n403), .B2(new_n357), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n401), .B1(new_n404), .B2(new_n398), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n400), .A2(new_n405), .A3(KEYINPUT90), .ZN(new_n406));
  OAI21_X1  g220(.A(G214), .B1(G237), .B2(G902), .ZN(new_n407));
  XNOR2_X1  g221(.A(new_n407), .B(KEYINPUT83), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n398), .B1(new_n363), .B2(new_n375), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT90), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n410), .A2(new_n411), .A3(new_n377), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n406), .A2(new_n409), .A3(new_n412), .ZN(new_n413));
  XNOR2_X1  g227(.A(G113), .B(G122), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n414), .B(new_n220), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(G237), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n417), .A2(new_n194), .A3(G214), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT91), .ZN(new_n419));
  NAND4_X1  g233(.A1(new_n418), .A2(new_n199), .A3(new_n419), .A4(new_n200), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n417), .A2(new_n194), .A3(G143), .A4(G214), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n419), .B1(new_n210), .B2(new_n418), .ZN(new_n423));
  OAI21_X1  g237(.A(G131), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT92), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n199), .A2(new_n200), .ZN(new_n426));
  AND3_X1   g240(.A1(new_n417), .A2(new_n194), .A3(G214), .ZN(new_n427));
  OAI21_X1  g241(.A(KEYINPUT91), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND4_X1  g242(.A1(new_n428), .A2(new_n246), .A3(new_n421), .A4(new_n420), .ZN(new_n429));
  AND3_X1   g243(.A1(new_n424), .A2(new_n425), .A3(new_n429), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n425), .B1(new_n424), .B2(new_n429), .ZN(new_n431));
  INV_X1    g245(.A(G140), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(G125), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n368), .A2(G140), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n433), .A2(new_n434), .A3(KEYINPUT16), .ZN(new_n435));
  OR3_X1    g249(.A1(new_n368), .A2(KEYINPUT16), .A3(G140), .ZN(new_n436));
  AND3_X1   g250(.A1(new_n435), .A2(G146), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(KEYINPUT73), .ZN(new_n438));
  XNOR2_X1  g252(.A(G125), .B(G140), .ZN(new_n439));
  AND2_X1   g253(.A1(new_n439), .A2(KEYINPUT19), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n439), .A2(KEYINPUT19), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n202), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n435), .A2(new_n436), .A3(G146), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT73), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n438), .A2(new_n442), .A3(new_n445), .ZN(new_n446));
  NOR3_X1   g260(.A1(new_n430), .A2(new_n431), .A3(new_n446), .ZN(new_n447));
  OAI211_X1 g261(.A(KEYINPUT18), .B(G131), .C1(new_n422), .C2(new_n423), .ZN(new_n448));
  NAND2_X1  g262(.A1(KEYINPUT18), .A2(G131), .ZN(new_n449));
  NAND4_X1  g263(.A1(new_n428), .A2(new_n421), .A3(new_n420), .A4(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n433), .A2(new_n434), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(G146), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n439), .A2(new_n202), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n448), .A2(new_n450), .A3(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n416), .B1(new_n447), .B2(new_n456), .ZN(new_n457));
  OAI211_X1 g271(.A(KEYINPUT17), .B(G131), .C1(new_n422), .C2(new_n423), .ZN(new_n458));
  AOI21_X1  g272(.A(G146), .B1(new_n435), .B2(new_n436), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n437), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(KEYINPUT93), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT93), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n458), .A2(new_n460), .A3(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT17), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n424), .A2(new_n465), .A3(new_n429), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n462), .A2(new_n464), .A3(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n467), .A2(new_n455), .A3(new_n415), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n457), .A2(new_n468), .ZN(new_n469));
  NOR2_X1   g283(.A1(G475), .A2(G902), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(KEYINPUT20), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT20), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n469), .A2(new_n473), .A3(new_n470), .ZN(new_n474));
  AND3_X1   g288(.A1(new_n467), .A2(new_n455), .A3(new_n415), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n415), .B1(new_n467), .B2(new_n455), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n192), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  AOI22_X1  g291(.A1(new_n472), .A2(new_n474), .B1(G475), .B2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT95), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n479), .B1(new_n198), .B2(G128), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n204), .A2(KEYINPUT95), .A3(G143), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n199), .A2(G128), .A3(new_n200), .ZN(new_n483));
  XNOR2_X1  g297(.A(KEYINPUT65), .B(G134), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n482), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  XNOR2_X1  g299(.A(G116), .B(G122), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(new_n217), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n486), .A2(new_n217), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT13), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n482), .B1(new_n483), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n483), .A2(new_n490), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT94), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n483), .A2(KEYINPUT94), .A3(new_n490), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n491), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  OAI221_X1 g310(.A(new_n485), .B1(new_n488), .B2(new_n489), .C1(new_n496), .C2(new_n248), .ZN(new_n497));
  XOR2_X1   g311(.A(KEYINPUT70), .B(G217), .Z(new_n498));
  NOR3_X1   g312(.A1(new_n498), .A2(G953), .A3(new_n187), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT98), .ZN(new_n500));
  AND3_X1   g314(.A1(new_n482), .A2(new_n483), .A3(new_n484), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n484), .B1(new_n482), .B2(new_n483), .ZN(new_n502));
  OAI21_X1  g316(.A(KEYINPUT96), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n482), .A2(new_n483), .ZN(new_n504));
  INV_X1    g318(.A(new_n484), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT96), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n506), .A2(new_n507), .A3(new_n485), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n503), .A2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(G122), .ZN(new_n510));
  OAI21_X1  g324(.A(KEYINPUT14), .B1(new_n510), .B2(G116), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT14), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n512), .A2(new_n325), .A3(G122), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n510), .A2(G116), .ZN(new_n514));
  AND4_X1   g328(.A1(KEYINPUT97), .A2(new_n511), .A3(new_n513), .A4(new_n514), .ZN(new_n515));
  OAI21_X1  g329(.A(G107), .B1(new_n513), .B2(KEYINPUT97), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n487), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n500), .B1(new_n509), .B2(new_n518), .ZN(new_n519));
  AOI211_X1 g333(.A(KEYINPUT98), .B(new_n517), .C1(new_n503), .C2(new_n508), .ZN(new_n520));
  OAI211_X1 g334(.A(new_n497), .B(new_n499), .C1(new_n519), .C2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(KEYINPUT99), .ZN(new_n522));
  NOR3_X1   g336(.A1(new_n501), .A2(new_n502), .A3(KEYINPUT96), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n507), .B1(new_n506), .B2(new_n485), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n518), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(KEYINPUT98), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n509), .A2(new_n500), .A3(new_n518), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT99), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n528), .A2(new_n529), .A3(new_n497), .A4(new_n499), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n497), .B1(new_n519), .B2(new_n520), .ZN(new_n531));
  INV_X1    g345(.A(new_n499), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n522), .A2(new_n530), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(new_n192), .ZN(new_n535));
  INV_X1    g349(.A(G478), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n536), .A2(KEYINPUT15), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(G952), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n539), .A2(G953), .ZN(new_n540));
  NAND2_X1  g354(.A1(G234), .A2(G237), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n541), .A2(G902), .A3(G953), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  XNOR2_X1  g359(.A(KEYINPUT21), .B(G898), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n543), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(new_n537), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n534), .A2(new_n192), .A3(new_n549), .ZN(new_n550));
  NAND4_X1  g364(.A1(new_n478), .A2(new_n538), .A3(new_n548), .A4(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(KEYINPUT100), .ZN(new_n552));
  AND3_X1   g366(.A1(new_n534), .A2(new_n192), .A3(new_n549), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n549), .B1(new_n534), .B2(new_n192), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT100), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n555), .A2(new_n556), .A3(new_n478), .A4(new_n548), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n413), .B1(new_n552), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n320), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(KEYINPUT74), .A2(KEYINPUT25), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  OAI21_X1  g375(.A(KEYINPUT23), .B1(new_n204), .B2(G119), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n204), .A2(G119), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n562), .A2(KEYINPUT72), .A3(new_n563), .ZN(new_n564));
  OAI21_X1  g378(.A(KEYINPUT72), .B1(new_n323), .B2(G128), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n323), .A2(G128), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n565), .A2(KEYINPUT23), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n564), .A2(new_n567), .ZN(new_n568));
  XNOR2_X1  g382(.A(G119), .B(G128), .ZN(new_n569));
  XNOR2_X1  g383(.A(KEYINPUT24), .B(G110), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  OAI22_X1  g385(.A1(new_n568), .A2(G110), .B1(new_n569), .B2(new_n571), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n572), .A2(new_n438), .A3(new_n445), .A4(new_n453), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n571), .A2(KEYINPUT71), .A3(new_n569), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT71), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n566), .A2(new_n563), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n575), .B1(new_n576), .B2(new_n570), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n574), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n568), .A2(G110), .ZN(new_n579));
  OAI211_X1 g393(.A(new_n578), .B(new_n579), .C1(new_n459), .C2(new_n437), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n573), .A2(new_n580), .ZN(new_n581));
  XNOR2_X1  g395(.A(KEYINPUT22), .B(G137), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n194), .A2(G221), .A3(G234), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n582), .B(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n581), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n573), .A2(new_n580), .A3(new_n584), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n586), .A2(new_n192), .A3(new_n587), .ZN(new_n588));
  NOR2_X1   g402(.A1(KEYINPUT74), .A2(KEYINPUT25), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n561), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n589), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n586), .A2(new_n192), .A3(new_n587), .A4(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n498), .B1(G234), .B2(new_n192), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT75), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n586), .A2(new_n587), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n594), .A2(G902), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n595), .A2(new_n596), .A3(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n594), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n603), .B1(new_n590), .B2(new_n592), .ZN(new_n604));
  OAI21_X1  g418(.A(KEYINPUT75), .B1(new_n604), .B2(new_n600), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT32), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT31), .ZN(new_n608));
  OAI211_X1 g422(.A(new_n365), .B(new_n364), .C1(new_n253), .C2(new_n254), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n245), .A2(new_n246), .A3(new_n252), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n246), .B1(G134), .B2(G137), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n611), .B1(new_n505), .B2(G137), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n275), .B1(new_n234), .B2(new_n258), .ZN(new_n613));
  OAI211_X1 g427(.A(new_n610), .B(new_n612), .C1(new_n613), .C2(new_n206), .ZN(new_n614));
  INV_X1    g428(.A(new_n348), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n609), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT28), .ZN(new_n617));
  AND2_X1   g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n615), .B1(new_n609), .B2(new_n614), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(new_n616), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n618), .B1(new_n621), .B2(KEYINPUT28), .ZN(new_n622));
  XNOR2_X1  g436(.A(KEYINPUT67), .B(KEYINPUT27), .ZN(new_n623));
  INV_X1    g437(.A(G210), .ZN(new_n624));
  NOR3_X1   g438(.A1(new_n624), .A2(G237), .A3(G953), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n623), .B(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(KEYINPUT26), .B(G101), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n626), .B(new_n627), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n608), .B1(new_n622), .B2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT30), .ZN(new_n630));
  AND3_X1   g444(.A1(new_n609), .A2(new_n630), .A3(new_n614), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n630), .B1(new_n609), .B2(new_n614), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n348), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n633), .A2(new_n616), .A3(new_n628), .ZN(new_n634));
  AND3_X1   g448(.A1(new_n609), .A2(new_n615), .A3(new_n614), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n609), .A2(new_n614), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(KEYINPUT30), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n609), .A2(new_n614), .A3(new_n630), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n635), .B1(new_n639), .B2(new_n348), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT68), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n640), .A2(new_n641), .A3(new_n608), .A4(new_n628), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n633), .A2(new_n608), .A3(new_n616), .A4(new_n628), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(KEYINPUT68), .ZN(new_n644));
  AOI22_X1  g458(.A1(new_n629), .A2(new_n634), .B1(new_n642), .B2(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(G472), .A2(G902), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(KEYINPUT69), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n607), .B1(new_n645), .B2(new_n647), .ZN(new_n648));
  OAI21_X1  g462(.A(KEYINPUT28), .B1(new_n635), .B2(new_n619), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n616), .A2(new_n617), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n628), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n634), .B1(new_n651), .B2(KEYINPUT31), .ZN(new_n652));
  AND2_X1   g466(.A1(new_n643), .A2(KEYINPUT68), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n643), .A2(KEYINPUT68), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n652), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n647), .A2(new_n607), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n649), .A2(KEYINPUT29), .A3(new_n628), .A4(new_n650), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n649), .A2(new_n628), .A3(new_n650), .ZN(new_n658));
  INV_X1    g472(.A(KEYINPUT29), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n628), .B1(new_n633), .B2(new_n616), .ZN(new_n661));
  OAI211_X1 g475(.A(new_n192), .B(new_n657), .C1(new_n660), .C2(new_n661), .ZN(new_n662));
  AOI22_X1  g476(.A1(new_n655), .A2(new_n656), .B1(new_n662), .B2(G472), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n606), .B1(new_n648), .B2(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n559), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(new_n227), .ZN(G3));
  INV_X1    g481(.A(G472), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n668), .B1(new_n655), .B2(new_n192), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n642), .A2(new_n644), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n647), .B1(new_n671), .B2(new_n652), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n674), .A2(new_n606), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n320), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n477), .A2(G475), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n473), .B1(new_n469), .B2(new_n470), .ZN(new_n678));
  INV_X1    g492(.A(new_n470), .ZN(new_n679));
  AOI211_X1 g493(.A(KEYINPUT20), .B(new_n679), .C1(new_n457), .C2(new_n468), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n677), .B1(new_n678), .B2(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT33), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n534), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n531), .A2(KEYINPUT102), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(new_n499), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n531), .A2(KEYINPUT102), .A3(new_n532), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n685), .A2(KEYINPUT33), .A3(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT103), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n536), .A2(G902), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n683), .A2(new_n687), .A3(new_n688), .A4(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n535), .A2(new_n536), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n682), .B1(new_n684), .B2(new_n499), .ZN(new_n693));
  AOI22_X1  g507(.A1(new_n682), .A2(new_n534), .B1(new_n693), .B2(new_n686), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n688), .B1(new_n694), .B2(new_n689), .ZN(new_n695));
  OAI21_X1  g509(.A(new_n681), .B1(new_n692), .B2(new_n695), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n400), .A2(new_n405), .A3(KEYINPUT101), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT101), .ZN(new_n698));
  OAI211_X1 g512(.A(new_n698), .B(new_n401), .C1(new_n404), .C2(new_n398), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n697), .A2(new_n407), .A3(new_n699), .ZN(new_n700));
  NOR4_X1   g514(.A1(new_n676), .A2(new_n547), .A3(new_n696), .A4(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(KEYINPUT34), .B(G104), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n701), .B(new_n702), .ZN(G6));
  INV_X1    g517(.A(KEYINPUT104), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n472), .A2(new_n704), .A3(new_n474), .ZN(new_n705));
  AOI22_X1  g519(.A1(new_n678), .A2(KEYINPUT104), .B1(G475), .B2(new_n477), .ZN(new_n706));
  OAI211_X1 g520(.A(new_n705), .B(new_n706), .C1(new_n553), .C2(new_n554), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n547), .B(KEYINPUT105), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  NOR4_X1   g523(.A1(new_n676), .A2(new_n700), .A3(new_n707), .A4(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(KEYINPUT35), .B(G107), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n710), .B(new_n711), .ZN(G9));
  XNOR2_X1  g526(.A(new_n581), .B(KEYINPUT106), .ZN(new_n713));
  OR2_X1    g527(.A1(new_n585), .A2(KEYINPUT36), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n713), .B(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(new_n715), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n595), .B1(new_n716), .B2(new_n599), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n670), .A2(new_n673), .A3(new_n717), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n559), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(KEYINPUT37), .B(G110), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n719), .B(new_n720), .ZN(G12));
  INV_X1    g535(.A(new_n656), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n657), .A2(new_n192), .ZN(new_n723));
  AND2_X1   g537(.A1(new_n658), .A2(new_n659), .ZN(new_n724));
  INV_X1    g538(.A(new_n661), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n723), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  OAI22_X1  g540(.A1(new_n645), .A2(new_n722), .B1(new_n726), .B2(new_n668), .ZN(new_n727));
  INV_X1    g541(.A(new_n647), .ZN(new_n728));
  AOI21_X1  g542(.A(KEYINPUT32), .B1(new_n655), .B2(new_n728), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n717), .B1(new_n727), .B2(new_n729), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n730), .A2(new_n700), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n194), .A2(G900), .ZN(new_n732));
  INV_X1    g546(.A(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n541), .A2(G902), .ZN(new_n734));
  OR3_X1    g548(.A1(new_n733), .A2(KEYINPUT107), .A3(new_n734), .ZN(new_n735));
  OAI21_X1  g549(.A(KEYINPUT107), .B1(new_n733), .B2(new_n734), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n735), .A2(new_n542), .A3(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n707), .A2(new_n738), .ZN(new_n739));
  AOI21_X1  g553(.A(KEYINPUT82), .B1(new_n318), .B2(new_n190), .ZN(new_n740));
  AND3_X1   g554(.A1(new_n318), .A2(KEYINPUT82), .A3(new_n190), .ZN(new_n741));
  OAI211_X1 g555(.A(new_n731), .B(new_n739), .C1(new_n740), .C2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G128), .ZN(G30));
  XNOR2_X1  g557(.A(new_n737), .B(KEYINPUT39), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n320), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n745), .A2(KEYINPUT40), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n406), .A2(new_n412), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT38), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n406), .A2(KEYINPUT38), .A3(new_n412), .ZN(new_n750));
  AND2_X1   g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(new_n628), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n620), .A2(new_n616), .A3(new_n752), .ZN(new_n753));
  OAI211_X1 g567(.A(new_n192), .B(new_n753), .C1(new_n640), .C2(new_n752), .ZN(new_n754));
  AOI22_X1  g568(.A1(new_n655), .A2(new_n656), .B1(G472), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n648), .A2(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n555), .A2(new_n478), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n604), .B1(new_n598), .B2(new_n715), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n758), .A2(new_n407), .A3(new_n759), .ZN(new_n760));
  NOR3_X1   g574(.A1(new_n751), .A2(new_n757), .A3(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT40), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n320), .A2(new_n762), .A3(new_n744), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n746), .A2(new_n761), .A3(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(new_n426), .ZN(G45));
  OAI211_X1 g579(.A(new_n681), .B(new_n737), .C1(new_n692), .C2(new_n695), .ZN(new_n766));
  INV_X1    g580(.A(new_n766), .ZN(new_n767));
  OAI211_X1 g581(.A(new_n767), .B(new_n731), .C1(new_n740), .C2(new_n741), .ZN(new_n768));
  XNOR2_X1  g582(.A(KEYINPUT108), .B(G146), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n768), .B(new_n769), .ZN(G48));
  NOR2_X1   g584(.A1(new_n700), .A2(new_n547), .ZN(new_n771));
  AND2_X1   g585(.A1(new_n690), .A2(new_n691), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n683), .A2(new_n687), .ZN(new_n773));
  INV_X1    g587(.A(new_n689), .ZN(new_n774));
  OAI21_X1  g588(.A(KEYINPUT103), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n478), .B1(new_n772), .B2(new_n775), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n192), .B1(new_n300), .B2(new_n303), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(G469), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n778), .A2(new_n188), .A3(new_n304), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n771), .A2(new_n664), .A3(new_n776), .A4(new_n780), .ZN(new_n781));
  XOR2_X1   g595(.A(KEYINPUT41), .B(G113), .Z(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(KEYINPUT109), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n781), .B(new_n783), .ZN(G15));
  INV_X1    g598(.A(new_n700), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n707), .A2(new_n709), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n785), .A2(new_n780), .A3(new_n664), .A4(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G116), .ZN(G18));
  NAND2_X1  g602(.A1(new_n552), .A2(new_n557), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n731), .A2(new_n789), .A3(new_n780), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G119), .ZN(G21));
  NOR2_X1   g605(.A1(new_n700), .A2(new_n779), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n538), .A2(new_n550), .ZN(new_n793));
  AOI21_X1  g607(.A(KEYINPUT110), .B1(new_n793), .B2(new_n681), .ZN(new_n794));
  OAI211_X1 g608(.A(new_n681), .B(KEYINPUT110), .C1(new_n553), .C2(new_n554), .ZN(new_n795));
  INV_X1    g609(.A(new_n795), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n604), .A2(new_n600), .ZN(new_n798));
  INV_X1    g612(.A(new_n798), .ZN(new_n799));
  NOR4_X1   g613(.A1(new_n669), .A2(new_n799), .A3(new_n672), .A4(new_n709), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n792), .A2(new_n797), .A3(new_n800), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(G122), .ZN(G24));
  NOR2_X1   g616(.A1(new_n766), .A2(new_n718), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n803), .A2(new_n792), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(G125), .ZN(G27));
  INV_X1    g619(.A(new_n188), .ZN(new_n806));
  INV_X1    g620(.A(new_n314), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n806), .B1(new_n807), .B2(new_n304), .ZN(new_n808));
  INV_X1    g622(.A(new_n407), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n809), .B1(new_n406), .B2(new_n412), .ZN(new_n810));
  AND3_X1   g624(.A1(new_n664), .A2(new_n808), .A3(new_n810), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n766), .A2(KEYINPUT42), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n799), .B1(new_n648), .B2(new_n663), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n808), .A2(new_n814), .A3(new_n810), .ZN(new_n815));
  OAI21_X1  g629(.A(KEYINPUT42), .B1(new_n815), .B2(new_n766), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n813), .A2(new_n816), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(new_n246), .ZN(G33));
  NAND4_X1  g632(.A1(new_n664), .A2(new_n808), .A3(new_n739), .A4(new_n810), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(G134), .ZN(G36));
  AOI21_X1  g634(.A(new_n681), .B1(new_n772), .B2(new_n775), .ZN(new_n821));
  OAI21_X1  g635(.A(KEYINPUT112), .B1(new_n821), .B2(KEYINPUT43), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n478), .B1(new_n692), .B2(new_n695), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT112), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT43), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n823), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n775), .A2(new_n691), .A3(new_n690), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n681), .B(KEYINPUT113), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n827), .A2(KEYINPUT43), .A3(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n822), .A2(new_n826), .A3(new_n829), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n759), .B1(new_n670), .B2(new_n673), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT44), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n307), .B1(new_n310), .B2(new_n308), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT45), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n191), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  OAI211_X1 g651(.A(new_n307), .B(KEYINPUT45), .C1(new_n308), .C2(new_n310), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n312), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  OR2_X1    g653(.A1(new_n839), .A2(KEYINPUT46), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT46), .ZN(new_n841));
  AOI211_X1 g655(.A(new_n841), .B(new_n312), .C1(new_n837), .C2(new_n838), .ZN(new_n842));
  INV_X1    g656(.A(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n840), .A2(new_n843), .A3(new_n304), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n844), .A2(KEYINPUT111), .A3(new_n188), .A4(new_n744), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT111), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n304), .B1(new_n839), .B2(KEYINPUT46), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n188), .B1(new_n847), .B2(new_n842), .ZN(new_n848));
  INV_X1    g662(.A(new_n744), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n846), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n845), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n830), .A2(KEYINPUT44), .A3(new_n831), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n834), .A2(new_n851), .A3(new_n810), .A4(new_n852), .ZN(new_n853));
  XNOR2_X1  g667(.A(new_n853), .B(G137), .ZN(G39));
  NAND3_X1  g668(.A1(new_n844), .A2(KEYINPUT47), .A3(new_n188), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT47), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n848), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(new_n810), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n648), .A2(new_n663), .ZN(new_n860));
  INV_X1    g674(.A(new_n606), .ZN(new_n861));
  NOR3_X1   g675(.A1(new_n859), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n858), .A2(new_n767), .A3(new_n862), .ZN(new_n863));
  XNOR2_X1  g677(.A(new_n863), .B(G140), .ZN(G42));
  INV_X1    g678(.A(KEYINPUT115), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n669), .A2(new_n672), .A3(new_n759), .ZN(new_n866));
  OAI211_X1 g680(.A(new_n320), .B(new_n558), .C1(new_n664), .C2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT114), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n868), .B1(new_n553), .B2(new_n554), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n538), .A2(KEYINPUT114), .A3(new_n550), .ZN(new_n870));
  AND2_X1   g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n696), .B1(new_n871), .B2(new_n681), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n413), .A2(new_n709), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n320), .A2(new_n872), .A3(new_n675), .A4(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n867), .A2(new_n874), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n790), .A2(new_n781), .A3(new_n801), .A4(new_n787), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  AND2_X1   g691(.A1(new_n742), .A2(new_n804), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT110), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n879), .B1(new_n555), .B2(new_n478), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n698), .B1(new_n410), .B2(new_n377), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n809), .B1(new_n881), .B2(new_n405), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n880), .A2(new_n882), .A3(new_n699), .A4(new_n795), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n717), .A2(new_n738), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n756), .A2(new_n188), .A3(new_n318), .A4(new_n884), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n860), .A2(new_n882), .A3(new_n699), .A4(new_n717), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n887), .B1(new_n317), .B2(new_n319), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n886), .B1(new_n888), .B2(new_n767), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT52), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n878), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n866), .A2(new_n827), .A3(new_n681), .A4(new_n737), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n808), .A2(new_n810), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n741), .A2(new_n740), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n759), .B1(new_n648), .B2(new_n663), .ZN(new_n895));
  AND3_X1   g709(.A1(new_n705), .A2(new_n706), .A3(new_n737), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n895), .A2(new_n871), .A3(new_n810), .A4(new_n896), .ZN(new_n897));
  OAI221_X1 g711(.A(new_n819), .B1(new_n892), .B2(new_n893), .C1(new_n894), .C2(new_n897), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n898), .A2(new_n817), .ZN(new_n899));
  AND2_X1   g713(.A1(new_n756), .A2(new_n884), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n900), .A2(new_n797), .A3(new_n785), .A4(new_n808), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n768), .A2(new_n742), .A3(new_n804), .A4(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(KEYINPUT52), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n877), .A2(new_n891), .A3(new_n899), .A4(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT53), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n865), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n891), .A2(new_n903), .ZN(new_n907));
  AND2_X1   g721(.A1(new_n867), .A2(new_n874), .ZN(new_n908));
  INV_X1    g722(.A(new_n817), .ZN(new_n909));
  AND4_X1   g723(.A1(new_n781), .A2(new_n790), .A3(new_n787), .A4(new_n801), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n819), .B1(new_n894), .B2(new_n897), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n892), .A2(new_n893), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n908), .A2(new_n909), .A3(new_n910), .A4(new_n913), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n905), .B1(new_n907), .B2(new_n914), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n902), .B(new_n890), .ZN(new_n916));
  AND3_X1   g730(.A1(new_n781), .A2(new_n801), .A3(new_n787), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n917), .A2(new_n790), .A3(new_n874), .A4(new_n867), .ZN(new_n918));
  AND4_X1   g732(.A1(new_n895), .A2(new_n871), .A3(new_n810), .A4(new_n896), .ZN(new_n919));
  AOI22_X1  g733(.A1(new_n919), .A2(new_n320), .B1(new_n811), .B2(new_n739), .ZN(new_n920));
  INV_X1    g734(.A(new_n912), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n920), .A2(new_n816), .A3(new_n813), .A4(new_n921), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n918), .A2(new_n922), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n916), .A2(new_n923), .A3(KEYINPUT115), .A4(KEYINPUT53), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n906), .A2(new_n915), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n925), .A2(KEYINPUT54), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n674), .A2(new_n799), .ZN(new_n927));
  AND4_X1   g741(.A1(new_n809), .A2(new_n749), .A3(new_n750), .A4(new_n780), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n830), .A2(new_n543), .A3(new_n927), .A4(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT116), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n930), .A2(KEYINPUT50), .ZN(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n929), .B(new_n932), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n859), .A2(new_n779), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n830), .A2(new_n543), .A3(new_n866), .A4(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT117), .ZN(new_n936));
  NOR3_X1   g750(.A1(new_n756), .A2(new_n606), .A3(new_n542), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n934), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n606), .A2(new_n542), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n780), .A2(new_n757), .A3(new_n810), .A4(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n940), .A2(KEYINPUT117), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n827), .A2(new_n681), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n938), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n778), .A2(new_n189), .A3(new_n304), .ZN(new_n944));
  AND3_X1   g758(.A1(new_n855), .A2(new_n857), .A3(new_n944), .ZN(new_n945));
  NAND4_X1  g759(.A1(new_n830), .A2(new_n543), .A3(new_n927), .A4(new_n810), .ZN(new_n946));
  OAI211_X1 g760(.A(new_n935), .B(new_n943), .C1(new_n945), .C2(new_n946), .ZN(new_n947));
  OAI21_X1  g761(.A(KEYINPUT51), .B1(new_n933), .B2(new_n947), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n929), .B(new_n931), .ZN(new_n949));
  OR2_X1    g763(.A1(new_n945), .A2(new_n946), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT51), .ZN(new_n951));
  AND2_X1   g765(.A1(new_n935), .A2(new_n943), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n949), .A2(new_n950), .A3(new_n951), .A4(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT118), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n830), .A2(new_n543), .A3(new_n814), .A4(new_n934), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT48), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n955), .B(new_n956), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n938), .A2(new_n776), .A3(new_n941), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n830), .A2(new_n543), .A3(new_n927), .ZN(new_n959));
  INV_X1    g773(.A(new_n792), .ZN(new_n960));
  OAI211_X1 g774(.A(new_n540), .B(new_n958), .C1(new_n959), .C2(new_n960), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n954), .B1(new_n957), .B2(new_n961), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n955), .B(KEYINPUT48), .ZN(new_n963));
  INV_X1    g777(.A(new_n961), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n963), .A2(new_n964), .A3(KEYINPUT118), .ZN(new_n965));
  AOI22_X1  g779(.A1(new_n948), .A2(new_n953), .B1(new_n962), .B2(new_n965), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n916), .A2(new_n923), .A3(KEYINPUT53), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT54), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n967), .A2(new_n915), .A3(new_n968), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n926), .A2(new_n966), .A3(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n970), .A2(KEYINPUT119), .ZN(new_n971));
  AND3_X1   g785(.A1(new_n967), .A2(new_n915), .A3(new_n968), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n972), .B1(KEYINPUT54), .B2(new_n925), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT119), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n973), .A2(new_n974), .A3(new_n966), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n539), .A2(new_n194), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n971), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  AND3_X1   g791(.A1(new_n751), .A2(new_n827), .A3(new_n828), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n798), .A2(new_n190), .A3(new_n409), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n778), .A2(new_n304), .ZN(new_n980));
  AOI211_X1 g794(.A(new_n979), .B(new_n756), .C1(KEYINPUT49), .C2(new_n980), .ZN(new_n981));
  OAI211_X1 g795(.A(new_n978), .B(new_n981), .C1(KEYINPUT49), .C2(new_n980), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n977), .A2(new_n982), .ZN(G75));
  NOR2_X1   g797(.A1(new_n194), .A2(G952), .ZN(new_n984));
  INV_X1    g798(.A(new_n984), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n967), .A2(new_n915), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n986), .A2(G902), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n987), .A2(new_n624), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n363), .B(new_n375), .ZN(new_n989));
  XNOR2_X1  g803(.A(new_n989), .B(KEYINPUT55), .ZN(new_n990));
  XOR2_X1   g804(.A(KEYINPUT121), .B(KEYINPUT56), .Z(new_n991));
  OR2_X1    g805(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n985), .B1(new_n988), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n988), .A2(KEYINPUT120), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT56), .ZN(new_n995));
  INV_X1    g809(.A(KEYINPUT120), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n996), .B1(new_n987), .B2(new_n624), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n994), .A2(new_n995), .A3(new_n997), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n993), .B1(new_n998), .B2(new_n990), .ZN(G51));
  INV_X1    g813(.A(KEYINPUT122), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n837), .A2(new_n838), .ZN(new_n1001));
  AOI211_X1 g815(.A(new_n192), .B(new_n1001), .C1(new_n967), .C2(new_n915), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n312), .B(KEYINPUT57), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n968), .B1(new_n967), .B2(new_n915), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n1003), .B1(new_n972), .B2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g819(.A1(new_n300), .A2(new_n303), .ZN(new_n1006));
  INV_X1    g820(.A(new_n1006), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n1002), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n1000), .B1(new_n1008), .B2(new_n984), .ZN(new_n1009));
  AOI21_X1  g823(.A(KEYINPUT53), .B1(new_n916), .B2(new_n923), .ZN(new_n1010));
  NOR3_X1   g824(.A1(new_n907), .A2(new_n914), .A3(new_n905), .ZN(new_n1011));
  OAI21_X1  g825(.A(KEYINPUT54), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1012), .A2(new_n969), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n1006), .B1(new_n1013), .B2(new_n1003), .ZN(new_n1014));
  OAI211_X1 g828(.A(KEYINPUT122), .B(new_n985), .C1(new_n1014), .C2(new_n1002), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1009), .A2(new_n1015), .ZN(G54));
  NAND4_X1  g830(.A1(new_n986), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n1017));
  INV_X1    g831(.A(new_n469), .ZN(new_n1018));
  AND2_X1   g832(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NOR2_X1   g833(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1020));
  NOR3_X1   g834(.A1(new_n1019), .A2(new_n1020), .A3(new_n984), .ZN(G60));
  NAND2_X1  g835(.A1(G478), .A2(G902), .ZN(new_n1022));
  XOR2_X1   g836(.A(new_n1022), .B(KEYINPUT59), .Z(new_n1023));
  NOR2_X1   g837(.A1(new_n773), .A2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g838(.A(new_n1024), .B1(new_n972), .B2(new_n1004), .ZN(new_n1025));
  INV_X1    g839(.A(KEYINPUT123), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g841(.A1(new_n1013), .A2(KEYINPUT123), .A3(new_n1024), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g843(.A(new_n773), .B1(new_n973), .B2(new_n1023), .ZN(new_n1030));
  AND3_X1   g844(.A1(new_n1029), .A2(new_n985), .A3(new_n1030), .ZN(G63));
  XOR2_X1   g845(.A(KEYINPUT124), .B(KEYINPUT60), .Z(new_n1032));
  NAND2_X1  g846(.A1(G217), .A2(G902), .ZN(new_n1033));
  XNOR2_X1  g847(.A(new_n1032), .B(new_n1033), .ZN(new_n1034));
  NAND2_X1  g848(.A1(new_n986), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g849(.A1(new_n1035), .A2(new_n597), .ZN(new_n1036));
  OAI211_X1 g850(.A(new_n1036), .B(new_n985), .C1(new_n716), .C2(new_n1035), .ZN(new_n1037));
  INV_X1    g851(.A(KEYINPUT61), .ZN(new_n1038));
  XNOR2_X1  g852(.A(new_n1037), .B(new_n1038), .ZN(G66));
  OAI21_X1  g853(.A(G953), .B1(new_n546), .B2(new_n371), .ZN(new_n1040));
  OAI21_X1  g854(.A(new_n1040), .B1(new_n877), .B2(G953), .ZN(new_n1041));
  OAI211_X1 g855(.A(new_n403), .B(new_n357), .C1(G898), .C2(new_n194), .ZN(new_n1042));
  XNOR2_X1  g856(.A(new_n1041), .B(new_n1042), .ZN(G69));
  AOI21_X1  g857(.A(new_n194), .B1(G227), .B2(G900), .ZN(new_n1044));
  AOI21_X1  g858(.A(new_n817), .B1(new_n739), .B2(new_n811), .ZN(new_n1045));
  INV_X1    g859(.A(new_n851), .ZN(new_n1046));
  NAND3_X1  g860(.A1(new_n797), .A2(new_n785), .A3(new_n814), .ZN(new_n1047));
  OAI211_X1 g861(.A(new_n863), .B(new_n1045), .C1(new_n1046), .C2(new_n1047), .ZN(new_n1048));
  AND3_X1   g862(.A1(new_n768), .A2(new_n742), .A3(new_n804), .ZN(new_n1049));
  NAND2_X1  g863(.A1(new_n853), .A2(new_n1049), .ZN(new_n1050));
  INV_X1    g864(.A(KEYINPUT126), .ZN(new_n1051));
  NAND2_X1  g865(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g866(.A1(new_n853), .A2(KEYINPUT126), .A3(new_n1049), .ZN(new_n1053));
  AOI21_X1  g867(.A(new_n1048), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g868(.A(new_n733), .B1(new_n1054), .B2(G953), .ZN(new_n1055));
  NOR2_X1   g869(.A1(new_n440), .A2(new_n441), .ZN(new_n1056));
  XNOR2_X1  g870(.A(new_n639), .B(new_n1056), .ZN(new_n1057));
  INV_X1    g871(.A(new_n1057), .ZN(new_n1058));
  NAND2_X1  g872(.A1(new_n1055), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g873(.A(KEYINPUT62), .ZN(new_n1060));
  NAND3_X1  g874(.A1(new_n764), .A2(new_n1060), .A3(new_n1049), .ZN(new_n1061));
  INV_X1    g875(.A(KEYINPUT125), .ZN(new_n1062));
  XNOR2_X1  g876(.A(new_n1061), .B(new_n1062), .ZN(new_n1063));
  NAND2_X1  g877(.A1(new_n764), .A2(new_n1049), .ZN(new_n1064));
  NAND2_X1  g878(.A1(new_n1064), .A2(KEYINPUT62), .ZN(new_n1065));
  INV_X1    g879(.A(new_n745), .ZN(new_n1066));
  NAND4_X1  g880(.A1(new_n1066), .A2(new_n664), .A3(new_n810), .A4(new_n872), .ZN(new_n1067));
  NAND4_X1  g881(.A1(new_n1065), .A2(new_n853), .A3(new_n863), .A4(new_n1067), .ZN(new_n1068));
  OAI21_X1  g882(.A(new_n194), .B1(new_n1063), .B2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g883(.A1(new_n1069), .A2(new_n1057), .ZN(new_n1070));
  AOI21_X1  g884(.A(new_n1044), .B1(new_n1059), .B2(new_n1070), .ZN(new_n1071));
  INV_X1    g885(.A(new_n1048), .ZN(new_n1072));
  AND3_X1   g886(.A1(new_n853), .A2(KEYINPUT126), .A3(new_n1049), .ZN(new_n1073));
  AOI21_X1  g887(.A(KEYINPUT126), .B1(new_n853), .B2(new_n1049), .ZN(new_n1074));
  OAI21_X1  g888(.A(new_n1072), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g889(.A(new_n732), .B1(new_n1075), .B2(new_n194), .ZN(new_n1076));
  OAI211_X1 g890(.A(new_n1070), .B(new_n1044), .C1(new_n1076), .C2(new_n1057), .ZN(new_n1077));
  INV_X1    g891(.A(new_n1077), .ZN(new_n1078));
  NOR2_X1   g892(.A1(new_n1071), .A2(new_n1078), .ZN(G72));
  NAND2_X1  g893(.A1(G472), .A2(G902), .ZN(new_n1080));
  XOR2_X1   g894(.A(new_n1080), .B(KEYINPUT63), .Z(new_n1081));
  OR2_X1    g895(.A1(new_n1063), .A2(new_n1068), .ZN(new_n1082));
  OAI21_X1  g896(.A(new_n1081), .B1(new_n1082), .B2(new_n918), .ZN(new_n1083));
  OR2_X1    g897(.A1(new_n640), .A2(new_n752), .ZN(new_n1084));
  INV_X1    g898(.A(new_n1084), .ZN(new_n1085));
  AOI21_X1  g899(.A(new_n984), .B1(new_n1083), .B2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g900(.A(new_n1081), .B1(new_n1075), .B2(new_n918), .ZN(new_n1087));
  NAND3_X1  g901(.A1(new_n1087), .A2(new_n640), .A3(new_n752), .ZN(new_n1088));
  NAND2_X1  g902(.A1(new_n725), .A2(new_n634), .ZN(new_n1089));
  NAND2_X1  g903(.A1(new_n1089), .A2(new_n1081), .ZN(new_n1090));
  XNOR2_X1  g904(.A(new_n1090), .B(KEYINPUT127), .ZN(new_n1091));
  NAND2_X1  g905(.A1(new_n925), .A2(new_n1091), .ZN(new_n1092));
  AND3_X1   g906(.A1(new_n1086), .A2(new_n1088), .A3(new_n1092), .ZN(G57));
endmodule


