//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 0 1 0 0 0 0 0 0 0 1 0 1 0 1 1 0 1 1 1 1 1 1 0 1 0 0 1 0 0 1 1 0 0 1 1 1 0 1 0 0 1 0 0 0 1 1 1 1 0 1 0 1 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:52 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1278,
    new_n1279, new_n1281, new_n1282, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1351, new_n1352, new_n1353;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G13), .ZN(new_n204));
  INV_X1    g0004(.A(new_n204), .ZN(new_n205));
  OAI21_X1  g0005(.A(G250), .B1(G257), .B2(G264), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  AND2_X1   g0007(.A1(G1), .A2(G13), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  OAI21_X1  g0011(.A(G50), .B1(G58), .B2(G68), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  AOI22_X1  g0013(.A1(new_n207), .A2(KEYINPUT0), .B1(new_n211), .B2(new_n213), .ZN(new_n214));
  OAI21_X1  g0014(.A(new_n214), .B1(KEYINPUT0), .B2(new_n207), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT64), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n217));
  XOR2_X1   g0017(.A(new_n217), .B(KEYINPUT65), .Z(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G116), .B2(G270), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n221));
  NAND3_X1  g0021(.A1(new_n219), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n203), .B1(new_n218), .B2(new_n222), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT1), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n216), .A2(new_n224), .ZN(G361));
  XOR2_X1   g0025(.A(G238), .B(G244), .Z(new_n226));
  XNOR2_X1  g0026(.A(G226), .B(G232), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G250), .B(G257), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT67), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G264), .B(G270), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n230), .B(new_n234), .ZN(G358));
  XOR2_X1   g0035(.A(G68), .B(G77), .Z(new_n236));
  XNOR2_X1  g0036(.A(G50), .B(G58), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT68), .B(KEYINPUT69), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XOR2_X1   g0041(.A(G107), .B(G116), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G351));
  INV_X1    g0044(.A(G33), .ZN(new_n245));
  OAI21_X1  g0045(.A(KEYINPUT72), .B1(new_n203), .B2(new_n245), .ZN(new_n246));
  INV_X1    g0046(.A(KEYINPUT72), .ZN(new_n247));
  NAND4_X1  g0047(.A1(new_n247), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n248));
  INV_X1    g0048(.A(G1), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n249), .A2(G13), .A3(G20), .ZN(new_n250));
  NAND4_X1  g0050(.A1(new_n246), .A2(new_n209), .A3(new_n248), .A4(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n249), .A2(G20), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n252), .A2(G68), .A3(new_n253), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n246), .A2(new_n209), .A3(new_n248), .ZN(new_n255));
  NOR2_X1   g0055(.A1(G20), .A2(G33), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G50), .ZN(new_n258));
  OAI22_X1  g0058(.A1(new_n257), .A2(new_n258), .B1(new_n210), .B2(G68), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n210), .A2(G33), .ZN(new_n260));
  INV_X1    g0060(.A(G77), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n255), .B1(new_n259), .B2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT11), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n254), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n250), .ZN(new_n266));
  INV_X1    g0066(.A(G68), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  XNOR2_X1  g0068(.A(new_n268), .B(KEYINPUT12), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n263), .A2(new_n264), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n265), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G169), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT13), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT3), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(new_n245), .ZN(new_n276));
  NAND2_X1  g0076(.A1(KEYINPUT3), .A2(G33), .ZN(new_n277));
  AOI21_X1  g0077(.A(G1698), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G226), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n276), .A2(new_n277), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n280), .A2(G232), .A3(G1698), .ZN(new_n281));
  NAND2_X1  g0081(.A1(G33), .A2(G97), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n279), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(G33), .A2(G41), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n208), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n283), .A2(new_n286), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n249), .B1(G41), .B2(G45), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT70), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  OAI211_X1 g0090(.A(new_n249), .B(KEYINPUT70), .C1(G41), .C2(G45), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G274), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n293), .B1(new_n208), .B2(new_n284), .ZN(new_n294));
  OR2_X1    g0094(.A1(G41), .A2(G45), .ZN(new_n295));
  AOI22_X1  g0095(.A1(new_n295), .A2(new_n249), .B1(new_n208), .B2(new_n284), .ZN(new_n296));
  AOI22_X1  g0096(.A1(new_n292), .A2(new_n294), .B1(new_n296), .B2(G238), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n274), .B1(new_n287), .B2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n287), .A2(new_n274), .A3(new_n297), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n273), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT14), .ZN(new_n302));
  INV_X1    g0102(.A(new_n300), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n303), .A2(new_n298), .ZN(new_n304));
  AOI22_X1  g0104(.A1(new_n301), .A2(new_n302), .B1(new_n304), .B2(G179), .ZN(new_n305));
  OAI21_X1  g0105(.A(G169), .B1(new_n303), .B2(new_n298), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(KEYINPUT14), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n272), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  OAI21_X1  g0108(.A(G200), .B1(new_n303), .B2(new_n298), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n299), .A2(G190), .A3(new_n300), .ZN(new_n310));
  AND3_X1   g0110(.A1(new_n309), .A2(new_n310), .A3(new_n272), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n308), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n292), .A2(new_n294), .ZN(new_n313));
  INV_X1    g0113(.A(G226), .ZN(new_n314));
  INV_X1    g0114(.A(new_n296), .ZN(new_n315));
  OAI211_X1 g0115(.A(new_n313), .B(KEYINPUT71), .C1(new_n314), .C2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT71), .ZN(new_n317));
  INV_X1    g0117(.A(new_n313), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n315), .A2(new_n314), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n317), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n280), .A2(G1698), .ZN(new_n321));
  INV_X1    g0121(.A(G223), .ZN(new_n322));
  OAI22_X1  g0122(.A1(new_n321), .A2(new_n322), .B1(new_n261), .B2(new_n280), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n323), .B1(G222), .B2(new_n278), .ZN(new_n324));
  OAI211_X1 g0124(.A(new_n316), .B(new_n320), .C1(new_n324), .C2(new_n285), .ZN(new_n325));
  OR2_X1    g0125(.A1(new_n325), .A2(G179), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n252), .A2(G50), .A3(new_n253), .ZN(new_n327));
  XNOR2_X1  g0127(.A(KEYINPUT8), .B(G58), .ZN(new_n328));
  INV_X1    g0128(.A(G150), .ZN(new_n329));
  OAI22_X1  g0129(.A1(new_n328), .A2(new_n260), .B1(new_n329), .B2(new_n257), .ZN(new_n330));
  NOR2_X1   g0130(.A1(G50), .A2(G58), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n210), .B1(new_n331), .B2(new_n267), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n255), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  OAI211_X1 g0133(.A(new_n327), .B(new_n333), .C1(G50), .C2(new_n250), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n325), .A2(new_n273), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n326), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(G190), .ZN(new_n338));
  OR2_X1    g0138(.A1(new_n325), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n325), .A2(G200), .ZN(new_n340));
  XNOR2_X1  g0140(.A(new_n334), .B(KEYINPUT9), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n339), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(KEYINPUT10), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT10), .ZN(new_n344));
  NAND4_X1  g0144(.A1(new_n339), .A2(new_n344), .A3(new_n340), .A4(new_n341), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n337), .B1(new_n343), .B2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT17), .ZN(new_n347));
  INV_X1    g0147(.A(G1698), .ZN(new_n348));
  AND2_X1   g0148(.A1(KEYINPUT3), .A2(G33), .ZN(new_n349));
  NOR2_X1   g0149(.A1(KEYINPUT3), .A2(G33), .ZN(new_n350));
  OAI211_X1 g0150(.A(G223), .B(new_n348), .C1(new_n349), .C2(new_n350), .ZN(new_n351));
  OAI211_X1 g0151(.A(G226), .B(G1698), .C1(new_n349), .C2(new_n350), .ZN(new_n352));
  NAND2_X1  g0152(.A1(G33), .A2(G87), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n351), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(new_n286), .ZN(new_n355));
  AOI22_X1  g0155(.A1(new_n292), .A2(new_n294), .B1(new_n296), .B2(G232), .ZN(new_n356));
  AOI21_X1  g0156(.A(G200), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  AND2_X1   g0157(.A1(new_n355), .A2(new_n356), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n357), .B1(new_n338), .B2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(new_n328), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(new_n253), .ZN(new_n361));
  OAI22_X1  g0161(.A1(new_n361), .A2(new_n251), .B1(new_n250), .B2(new_n360), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  XNOR2_X1  g0163(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n349), .A2(new_n350), .ZN(new_n366));
  AOI21_X1  g0166(.A(KEYINPUT7), .B1(new_n366), .B2(new_n210), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n276), .A2(KEYINPUT7), .A3(new_n210), .A4(new_n277), .ZN(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  OAI21_X1  g0169(.A(G68), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(G58), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n371), .A2(new_n267), .ZN(new_n372));
  NOR2_X1   g0172(.A1(G58), .A2(G68), .ZN(new_n373));
  OAI21_X1  g0173(.A(G20), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n256), .A2(G159), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n365), .B1(new_n370), .B2(new_n377), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n276), .A2(new_n210), .A3(new_n277), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT7), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n267), .B1(new_n381), .B2(new_n368), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n374), .A2(KEYINPUT16), .A3(new_n375), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n255), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n363), .B1(new_n378), .B2(new_n384), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n347), .B1(new_n359), .B2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(G179), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n355), .A2(new_n356), .A3(new_n387), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n388), .B1(new_n358), .B2(G169), .ZN(new_n389));
  AND3_X1   g0189(.A1(new_n246), .A2(new_n209), .A3(new_n248), .ZN(new_n390));
  AND3_X1   g0190(.A1(new_n374), .A2(KEYINPUT16), .A3(new_n375), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n390), .B1(new_n370), .B2(new_n391), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n364), .B1(new_n382), .B2(new_n376), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n362), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  OAI21_X1  g0194(.A(KEYINPUT18), .B1(new_n389), .B2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(new_n388), .ZN(new_n396));
  AOI21_X1  g0196(.A(G169), .B1(new_n355), .B2(new_n356), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT18), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n398), .A2(new_n385), .A3(new_n399), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n355), .A2(new_n356), .A3(new_n338), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n401), .B1(new_n358), .B2(G200), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n402), .A2(new_n394), .A3(KEYINPUT17), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n386), .A2(new_n395), .A3(new_n400), .A4(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT73), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n328), .B1(new_n406), .B2(new_n257), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n407), .B1(new_n406), .B2(new_n257), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n408), .B1(new_n210), .B2(new_n261), .ZN(new_n409));
  XNOR2_X1  g0209(.A(KEYINPUT15), .B(G87), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT74), .ZN(new_n411));
  XNOR2_X1  g0211(.A(new_n410), .B(new_n411), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n412), .A2(new_n260), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n255), .B1(new_n409), .B2(new_n413), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n252), .A2(G77), .A3(new_n253), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n266), .A2(new_n261), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n414), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n318), .B1(G244), .B2(new_n296), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n280), .A2(G232), .A3(new_n348), .ZN(new_n419));
  INV_X1    g0219(.A(G107), .ZN(new_n420));
  INV_X1    g0220(.A(G238), .ZN(new_n421));
  OAI221_X1 g0221(.A(new_n419), .B1(new_n420), .B2(new_n280), .C1(new_n321), .C2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(new_n286), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n418), .A2(new_n387), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n418), .A2(new_n423), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(new_n273), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n417), .A2(new_n424), .A3(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n425), .A2(G200), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n425), .A2(new_n338), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n417), .A2(new_n430), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n428), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n312), .A2(new_n346), .A3(new_n405), .A4(new_n432), .ZN(new_n433));
  OAI211_X1 g0233(.A(G264), .B(G1698), .C1(new_n349), .C2(new_n350), .ZN(new_n434));
  OAI211_X1 g0234(.A(G257), .B(new_n348), .C1(new_n349), .C2(new_n350), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n276), .A2(G303), .A3(new_n277), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n434), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(KEYINPUT80), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT80), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n434), .A2(new_n435), .A3(new_n439), .A4(new_n436), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n285), .B1(new_n438), .B2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(G45), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n442), .A2(G1), .ZN(new_n443));
  AND2_X1   g0243(.A1(KEYINPUT5), .A2(G41), .ZN(new_n444));
  NOR2_X1   g0244(.A1(KEYINPUT5), .A2(G41), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n443), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n446), .A2(G270), .A3(new_n285), .ZN(new_n447));
  XNOR2_X1  g0247(.A(KEYINPUT5), .B(G41), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n294), .A2(new_n443), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  OAI21_X1  g0250(.A(G200), .B1(new_n441), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n249), .A2(G33), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n390), .A2(G116), .A3(new_n250), .A4(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(G116), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n266), .A2(new_n454), .ZN(new_n455));
  AOI21_X1  g0255(.A(G20), .B1(G33), .B2(G283), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n245), .A2(G97), .ZN(new_n457));
  AOI22_X1  g0257(.A1(new_n456), .A2(new_n457), .B1(G20), .B2(new_n454), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n255), .A2(KEYINPUT20), .A3(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  AOI21_X1  g0260(.A(KEYINPUT20), .B1(new_n255), .B2(new_n458), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n453), .B(new_n455), .C1(new_n460), .C2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT81), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n255), .A2(new_n458), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT20), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(new_n459), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n468), .A2(KEYINPUT81), .A3(new_n453), .A4(new_n455), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n451), .A2(new_n464), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(KEYINPUT82), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n438), .A2(new_n440), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(new_n286), .ZN(new_n473));
  AND2_X1   g0273(.A1(new_n447), .A2(new_n449), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n473), .A2(G190), .A3(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT82), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n451), .A2(new_n464), .A3(new_n476), .A4(new_n469), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n471), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  OAI21_X1  g0278(.A(G169), .B1(new_n441), .B2(new_n450), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n479), .B1(new_n464), .B2(new_n469), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n464), .A2(new_n469), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n474), .A2(G179), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n441), .A2(new_n482), .ZN(new_n483));
  AOI22_X1  g0283(.A1(new_n480), .A2(KEYINPUT21), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n273), .B1(new_n473), .B2(new_n474), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n481), .A2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT21), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n478), .A2(new_n484), .A3(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n446), .A2(G264), .A3(new_n285), .ZN(new_n490));
  AND2_X1   g0290(.A1(new_n490), .A2(new_n449), .ZN(new_n491));
  OAI211_X1 g0291(.A(G257), .B(G1698), .C1(new_n349), .C2(new_n350), .ZN(new_n492));
  OAI211_X1 g0292(.A(G250), .B(new_n348), .C1(new_n349), .C2(new_n350), .ZN(new_n493));
  NAND2_X1  g0293(.A1(G33), .A2(G294), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n492), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(new_n286), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n491), .A2(new_n338), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n490), .A2(new_n449), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n498), .B1(new_n286), .B2(new_n495), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n497), .B1(new_n499), .B2(G200), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n210), .B(G87), .C1(new_n349), .C2(new_n350), .ZN(new_n501));
  AND2_X1   g0301(.A1(KEYINPUT83), .A2(KEYINPUT22), .ZN(new_n502));
  NOR2_X1   g0302(.A1(KEYINPUT83), .A2(KEYINPUT22), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n501), .A2(new_n504), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n280), .A2(new_n210), .A3(G87), .A4(new_n502), .ZN(new_n506));
  NAND2_X1  g0306(.A1(G33), .A2(G116), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n507), .A2(G20), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT23), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n509), .B1(new_n210), .B2(G107), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n420), .A2(KEYINPUT23), .A3(G20), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n508), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n505), .A2(new_n506), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(KEYINPUT24), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT24), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n505), .A2(new_n506), .A3(new_n512), .A4(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n255), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n266), .A2(new_n420), .ZN(new_n519));
  NOR2_X1   g0319(.A1(KEYINPUT84), .A2(KEYINPUT25), .ZN(new_n520));
  OR2_X1    g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  AND2_X1   g0321(.A1(KEYINPUT84), .A2(KEYINPUT25), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n522), .B1(new_n519), .B2(new_n520), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n252), .A2(new_n452), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n524), .B1(new_n525), .B2(new_n420), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n500), .A2(new_n518), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n491), .A2(new_n496), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n529), .A2(new_n387), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n273), .B1(new_n491), .B2(new_n496), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n390), .B1(new_n514), .B2(new_n516), .ZN(new_n532));
  OAI22_X1  g0332(.A1(new_n530), .A2(new_n531), .B1(new_n532), .B2(new_n526), .ZN(new_n533));
  AND2_X1   g0333(.A1(new_n528), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n446), .A2(G257), .A3(new_n285), .ZN(new_n535));
  INV_X1    g0335(.A(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n278), .A2(KEYINPUT4), .A3(G244), .ZN(new_n537));
  OAI211_X1 g0337(.A(G244), .B(new_n348), .C1(new_n349), .C2(new_n350), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT4), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(G33), .A2(G283), .ZN(new_n541));
  OAI211_X1 g0341(.A(G250), .B(G1698), .C1(new_n349), .C2(new_n350), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n537), .A2(new_n540), .A3(new_n541), .A4(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n536), .B1(new_n543), .B2(new_n286), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n544), .A2(new_n338), .A3(new_n449), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n541), .B(new_n542), .C1(new_n538), .C2(new_n539), .ZN(new_n546));
  AOI21_X1  g0346(.A(KEYINPUT4), .B1(new_n278), .B2(G244), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n286), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  AND3_X1   g0348(.A1(new_n548), .A2(new_n449), .A3(new_n535), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n545), .B1(new_n549), .B2(G200), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n250), .A2(G97), .ZN(new_n551));
  INV_X1    g0351(.A(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(G97), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n552), .B1(new_n525), .B2(new_n553), .ZN(new_n554));
  OAI21_X1  g0354(.A(G107), .B1(new_n367), .B2(new_n369), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(KEYINPUT77), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n420), .B1(new_n381), .B2(new_n368), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT77), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT76), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n560), .A2(new_n420), .A3(KEYINPUT6), .A4(G97), .ZN(new_n561));
  NAND2_X1  g0361(.A1(KEYINPUT6), .A2(G97), .ZN(new_n562));
  OAI21_X1  g0362(.A(KEYINPUT76), .B1(new_n562), .B2(G107), .ZN(new_n563));
  AND2_X1   g0363(.A1(G97), .A2(G107), .ZN(new_n564));
  NOR2_X1   g0364(.A1(G97), .A2(G107), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n561), .B(new_n563), .C1(new_n566), .C2(KEYINPUT6), .ZN(new_n567));
  AOI22_X1  g0367(.A1(new_n567), .A2(G20), .B1(G77), .B2(new_n256), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n556), .A2(new_n559), .A3(new_n568), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n554), .B1(new_n569), .B2(new_n255), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n550), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n569), .A2(new_n255), .ZN(new_n572));
  INV_X1    g0372(.A(new_n554), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g0374(.A(G169), .B1(new_n544), .B2(new_n449), .ZN(new_n575));
  INV_X1    g0375(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n549), .A2(new_n387), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n574), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  OAI211_X1 g0378(.A(G244), .B(G1698), .C1(new_n349), .C2(new_n350), .ZN(new_n579));
  OAI211_X1 g0379(.A(G238), .B(new_n348), .C1(new_n349), .C2(new_n350), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n579), .A2(new_n580), .A3(new_n507), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(new_n286), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n249), .A2(G45), .ZN(new_n583));
  AND2_X1   g0383(.A1(new_n583), .A2(G250), .ZN(new_n584));
  AOI22_X1  g0384(.A1(new_n285), .A2(new_n584), .B1(new_n294), .B2(new_n443), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(G200), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n582), .A2(new_n585), .A3(G190), .ZN(new_n588));
  AND2_X1   g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n590));
  AND3_X1   g0390(.A1(new_n590), .A2(KEYINPUT78), .A3(new_n210), .ZN(new_n591));
  AOI21_X1  g0391(.A(KEYINPUT78), .B1(new_n590), .B2(new_n210), .ZN(new_n592));
  NOR3_X1   g0392(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n593));
  NOR3_X1   g0393(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n210), .B(G68), .C1(new_n349), .C2(new_n350), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n260), .A2(new_n553), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n595), .B1(KEYINPUT19), .B2(new_n596), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n255), .B1(new_n594), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n412), .A2(new_n266), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n252), .A2(G87), .A3(new_n452), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n598), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT79), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n412), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n251), .B1(new_n249), .B2(G33), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n410), .A2(new_n411), .ZN(new_n606));
  INV_X1    g0406(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n410), .A2(new_n411), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n607), .A2(KEYINPUT79), .A3(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n604), .A2(new_n605), .A3(new_n609), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n610), .A2(new_n599), .A3(new_n598), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n586), .A2(G169), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n582), .A2(new_n585), .A3(G179), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  AOI22_X1  g0414(.A1(new_n589), .A2(new_n602), .B1(new_n611), .B2(new_n614), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n534), .A2(new_n571), .A3(new_n578), .A4(new_n615), .ZN(new_n616));
  NOR3_X1   g0416(.A1(new_n433), .A2(new_n489), .A3(new_n616), .ZN(G372));
  INV_X1    g0417(.A(new_n433), .ZN(new_n618));
  AND3_X1   g0418(.A1(new_n582), .A2(new_n585), .A3(G179), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n273), .B1(new_n582), .B2(new_n585), .ZN(new_n620));
  OAI21_X1  g0420(.A(KEYINPUT85), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT85), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n612), .A2(new_n622), .A3(new_n613), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT86), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n601), .A2(new_n625), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n598), .A2(new_n599), .A3(KEYINPUT86), .A4(new_n600), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  AOI22_X1  g0428(.A1(new_n624), .A2(new_n611), .B1(new_n628), .B2(new_n589), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT26), .ZN(new_n630));
  AND3_X1   g0430(.A1(new_n544), .A2(new_n387), .A3(new_n449), .ZN(new_n631));
  NOR3_X1   g0431(.A1(new_n570), .A2(new_n631), .A3(new_n575), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n629), .A2(new_n630), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n624), .A2(new_n611), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n611), .A2(new_n614), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n602), .A2(new_n587), .A3(new_n588), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  OAI21_X1  g0437(.A(KEYINPUT26), .B1(new_n578), .B2(new_n637), .ZN(new_n638));
  AND3_X1   g0438(.A1(new_n633), .A2(new_n634), .A3(new_n638), .ZN(new_n639));
  AND3_X1   g0439(.A1(new_n578), .A2(new_n571), .A3(new_n528), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n481), .A2(new_n483), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n481), .A2(KEYINPUT21), .A3(new_n485), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n488), .A2(new_n641), .A3(new_n642), .A4(new_n533), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n640), .A2(new_n643), .A3(new_n629), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n639), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n618), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g0446(.A(new_n646), .B(KEYINPUT87), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n343), .A2(new_n345), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n386), .A2(new_n403), .ZN(new_n649));
  INV_X1    g0449(.A(new_n272), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n299), .A2(G179), .A3(new_n300), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n651), .B1(new_n306), .B2(KEYINPUT14), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n299), .A2(new_n300), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n302), .B1(new_n653), .B2(G169), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n650), .B1(new_n652), .B2(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n309), .A2(new_n310), .A3(new_n272), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n428), .A2(new_n656), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n649), .B1(new_n655), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n395), .A2(new_n400), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n648), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(new_n336), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT88), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n660), .A2(KEYINPUT88), .A3(new_n336), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n647), .A2(new_n665), .ZN(G369));
  INV_X1    g0466(.A(G330), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n642), .A2(new_n641), .ZN(new_n668));
  AOI21_X1  g0468(.A(KEYINPUT21), .B1(new_n481), .B2(new_n485), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n249), .A2(new_n210), .A3(G13), .ZN(new_n671));
  OR2_X1    g0471(.A1(new_n671), .A2(KEYINPUT27), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(KEYINPUT27), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n672), .A2(G213), .A3(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(G343), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n481), .A2(new_n676), .ZN(new_n677));
  OR2_X1    g0477(.A1(new_n670), .A2(new_n677), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n670), .A2(new_n478), .A3(new_n677), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n667), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n533), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(new_n676), .ZN(new_n682));
  XNOR2_X1  g0482(.A(new_n682), .B(KEYINPUT89), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n676), .B1(new_n532), .B2(new_n526), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n534), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n680), .A2(new_n686), .ZN(new_n687));
  AND2_X1   g0487(.A1(new_n687), .A2(KEYINPUT90), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n687), .A2(KEYINPUT90), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n670), .A2(new_n676), .ZN(new_n692));
  INV_X1    g0492(.A(new_n676), .ZN(new_n693));
  AOI22_X1  g0493(.A1(new_n686), .A2(new_n692), .B1(new_n681), .B2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n691), .A2(new_n694), .ZN(G399));
  NOR2_X1   g0495(.A1(new_n205), .A2(G41), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n696), .A2(new_n249), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n593), .A2(new_n454), .ZN(new_n699));
  INV_X1    g0499(.A(new_n696), .ZN(new_n700));
  OAI22_X1  g0500(.A1(new_n698), .A2(new_n699), .B1(new_n212), .B2(new_n700), .ZN(new_n701));
  XNOR2_X1  g0501(.A(new_n701), .B(KEYINPUT28), .ZN(new_n702));
  AOI211_X1 g0502(.A(KEYINPUT29), .B(new_n676), .C1(new_n639), .C2(new_n644), .ZN(new_n703));
  NOR3_X1   g0503(.A1(new_n668), .A2(new_n669), .A3(new_n681), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n629), .A2(new_n571), .A3(new_n578), .A4(new_n528), .ZN(new_n705));
  OAI21_X1  g0505(.A(KEYINPUT93), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n632), .A2(new_n630), .A3(new_n615), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(new_n634), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n630), .B1(new_n629), .B2(new_n632), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT93), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n640), .A2(new_n643), .A3(new_n711), .A4(new_n629), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n706), .A2(new_n710), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(new_n693), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n703), .B1(new_n714), .B2(KEYINPUT29), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n450), .A2(new_n387), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n473), .A2(KEYINPUT91), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n548), .A2(new_n535), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n491), .A2(new_n496), .A3(new_n582), .A4(new_n585), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT91), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n721), .B1(new_n441), .B2(new_n482), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n717), .A2(new_n720), .A3(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT30), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT92), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n717), .A2(new_n720), .A3(KEYINPUT30), .A4(new_n722), .ZN(new_n728));
  AND3_X1   g0528(.A1(new_n529), .A2(new_n387), .A3(new_n586), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n544), .A2(new_n449), .ZN(new_n730));
  OAI211_X1 g0530(.A(new_n729), .B(new_n730), .C1(new_n450), .C2(new_n441), .ZN(new_n731));
  AND2_X1   g0531(.A1(new_n728), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n723), .A2(KEYINPUT92), .A3(new_n724), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n727), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(new_n676), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT31), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n616), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n738), .A2(new_n670), .A3(new_n478), .A4(new_n693), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n732), .A2(new_n725), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n740), .A2(KEYINPUT31), .A3(new_n676), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n737), .A2(new_n739), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(G330), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n715), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n702), .B1(new_n745), .B2(G1), .ZN(G364));
  NAND2_X1  g0546(.A1(new_n210), .A2(G13), .ZN(new_n747));
  XNOR2_X1  g0547(.A(new_n747), .B(KEYINPUT94), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(G45), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n697), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n205), .A2(new_n366), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(G355), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n753), .B1(G116), .B2(new_n204), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n240), .A2(G45), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n205), .A2(new_n280), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n757), .B1(new_n442), .B2(new_n213), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n754), .B1(new_n755), .B2(new_n758), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n209), .B1(G20), .B2(new_n273), .ZN(new_n760));
  NOR2_X1   g0560(.A1(G13), .A2(G33), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(G20), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n760), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n751), .B1(new_n759), .B2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n210), .A2(G190), .ZN(new_n767));
  OAI21_X1  g0567(.A(KEYINPUT96), .B1(G179), .B2(G200), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR3_X1   g0569(.A1(KEYINPUT96), .A2(G179), .A3(G200), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n767), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(KEYINPUT97), .ZN(new_n772));
  OR2_X1    g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n771), .A2(new_n772), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(G329), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n210), .A2(new_n338), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n778), .A2(new_n387), .A3(G200), .ZN(new_n779));
  XOR2_X1   g0579(.A(new_n779), .B(KEYINPUT98), .Z(new_n780));
  XNOR2_X1  g0580(.A(KEYINPUT33), .B(G317), .ZN(new_n781));
  INV_X1    g0581(.A(KEYINPUT99), .ZN(new_n782));
  OR2_X1    g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g0583(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n784), .A2(G190), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n786), .B1(new_n781), .B2(new_n782), .ZN(new_n787));
  AOI22_X1  g0587(.A1(new_n780), .A2(G303), .B1(new_n783), .B2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n770), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n338), .B1(new_n789), .B2(new_n768), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(new_n210), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(G294), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n387), .A2(G200), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n778), .A2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(G322), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n366), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n767), .A2(new_n387), .A3(G200), .ZN(new_n798));
  INV_X1    g0598(.A(G283), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n767), .A2(new_n794), .ZN(new_n800));
  INV_X1    g0600(.A(G311), .ZN(new_n801));
  OAI22_X1  g0601(.A1(new_n798), .A2(new_n799), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n784), .A2(new_n338), .ZN(new_n803));
  AOI211_X1 g0603(.A(new_n797), .B(new_n802), .C1(G326), .C2(new_n803), .ZN(new_n804));
  NAND4_X1  g0604(.A1(new_n777), .A2(new_n788), .A3(new_n793), .A4(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n776), .A2(G159), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n806), .B(KEYINPUT32), .ZN(new_n807));
  INV_X1    g0607(.A(G87), .ZN(new_n808));
  OAI22_X1  g0608(.A1(new_n779), .A2(new_n808), .B1(new_n800), .B2(new_n261), .ZN(new_n809));
  INV_X1    g0609(.A(new_n798), .ZN(new_n810));
  AOI211_X1 g0610(.A(new_n366), .B(new_n809), .C1(G107), .C2(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n792), .A2(G97), .ZN(new_n812));
  XNOR2_X1  g0612(.A(new_n795), .B(KEYINPUT95), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n814), .A2(G58), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n785), .A2(G68), .B1(new_n803), .B2(G50), .ZN(new_n816));
  NAND4_X1  g0616(.A1(new_n811), .A2(new_n812), .A3(new_n815), .A4(new_n816), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n805), .B1(new_n807), .B2(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n766), .B1(new_n818), .B2(new_n760), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n678), .A2(new_n679), .ZN(new_n820));
  INV_X1    g0620(.A(new_n763), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n819), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n680), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(new_n750), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n820), .A2(G330), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n822), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  XNOR2_X1  g0626(.A(new_n826), .B(KEYINPUT100), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(G396));
  NAND2_X1  g0628(.A1(new_n645), .A2(new_n693), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n427), .A2(new_n676), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  AOI22_X1  g0631(.A1(new_n431), .A2(new_n429), .B1(new_n417), .B2(new_n676), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n831), .B1(new_n832), .B2(new_n428), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n829), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n431), .A2(new_n429), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n417), .A2(new_n676), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n830), .B1(new_n837), .B2(new_n427), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n704), .A2(new_n705), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n633), .A2(new_n634), .A3(new_n638), .ZN(new_n840));
  OAI211_X1 g0640(.A(new_n693), .B(new_n838), .C1(new_n839), .C2(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n834), .A2(new_n841), .ZN(new_n842));
  OR2_X1    g0642(.A1(new_n842), .A2(new_n743), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n751), .B1(new_n842), .B2(new_n743), .ZN(new_n844));
  AND2_X1   g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n776), .A2(G311), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n780), .A2(G107), .ZN(new_n847));
  INV_X1    g0647(.A(new_n803), .ZN(new_n848));
  INV_X1    g0648(.A(G303), .ZN(new_n849));
  OAI22_X1  g0649(.A1(new_n786), .A2(new_n799), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(G294), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n366), .B1(new_n795), .B2(new_n851), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n798), .A2(new_n808), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n800), .A2(new_n454), .ZN(new_n854));
  NOR4_X1   g0654(.A1(new_n850), .A2(new_n852), .A3(new_n853), .A4(new_n854), .ZN(new_n855));
  NAND4_X1  g0655(.A1(new_n846), .A2(new_n812), .A3(new_n847), .A4(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n800), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n857), .A2(G159), .B1(G137), .B2(new_n803), .ZN(new_n858));
  INV_X1    g0658(.A(G143), .ZN(new_n859));
  OAI221_X1 g0659(.A(new_n858), .B1(new_n329), .B2(new_n786), .C1(new_n813), .C2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT34), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n280), .B1(new_n798), .B2(new_n267), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n863), .B1(new_n780), .B2(G50), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n776), .A2(G132), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n792), .A2(G58), .ZN(new_n866));
  NAND4_X1  g0666(.A1(new_n862), .A2(new_n864), .A3(new_n865), .A4(new_n866), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n860), .A2(new_n861), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n856), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n869), .A2(new_n760), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n760), .A2(new_n761), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n750), .B1(new_n261), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n873), .B1(new_n761), .B2(new_n833), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n845), .A2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(G384));
  OR2_X1    g0676(.A1(new_n567), .A2(KEYINPUT35), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n567), .A2(KEYINPUT35), .ZN(new_n878));
  NAND4_X1  g0678(.A1(new_n877), .A2(G116), .A3(new_n211), .A4(new_n878), .ZN(new_n879));
  XOR2_X1   g0679(.A(new_n879), .B(KEYINPUT36), .Z(new_n880));
  OAI211_X1 g0680(.A(new_n213), .B(G77), .C1(new_n371), .C2(new_n267), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n258), .A2(G68), .ZN(new_n882));
  AOI211_X1 g0682(.A(new_n249), .B(G13), .C1(new_n881), .C2(new_n882), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT40), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n398), .A2(new_n385), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n402), .A2(new_n394), .ZN(new_n887));
  INV_X1    g0687(.A(new_n674), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n385), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n886), .A2(new_n887), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(KEYINPUT37), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT101), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT37), .ZN(new_n893));
  NAND4_X1  g0693(.A1(new_n886), .A2(new_n887), .A3(new_n889), .A4(new_n893), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n891), .A2(new_n892), .A3(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n889), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n404), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n890), .A2(KEYINPUT101), .A3(KEYINPUT37), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n895), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT38), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND4_X1  g0701(.A1(new_n895), .A2(KEYINPUT38), .A3(new_n897), .A4(new_n898), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n901), .A2(KEYINPUT102), .A3(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT102), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n899), .A2(new_n904), .A3(new_n900), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n734), .A2(KEYINPUT31), .A3(new_n676), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n737), .A2(new_n739), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n650), .A2(new_n676), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n655), .A2(new_n656), .A3(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n653), .A2(new_n302), .A3(G169), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n307), .A2(new_n911), .A3(new_n651), .ZN(new_n912));
  OAI211_X1 g0712(.A(new_n650), .B(new_n676), .C1(new_n912), .C2(new_n311), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n833), .B1(new_n910), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n908), .A2(new_n914), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n885), .B1(new_n906), .B2(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n891), .A2(KEYINPUT103), .A3(new_n894), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n897), .ZN(new_n918));
  AOI21_X1  g0718(.A(KEYINPUT103), .B1(new_n891), .B2(new_n894), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n900), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n885), .B1(new_n920), .B2(new_n902), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n921), .A2(new_n908), .A3(new_n914), .ZN(new_n922));
  AND2_X1   g0722(.A1(new_n916), .A2(new_n922), .ZN(new_n923));
  NOR3_X1   g0723(.A1(new_n489), .A2(new_n616), .A3(new_n676), .ZN(new_n924));
  AOI21_X1  g0724(.A(KEYINPUT31), .B1(new_n734), .B2(new_n676), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n433), .B1(new_n926), .B2(new_n907), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n667), .B1(new_n923), .B2(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n928), .B1(new_n923), .B2(new_n927), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n902), .A2(KEYINPUT102), .ZN(new_n930));
  AND2_X1   g0730(.A1(new_n890), .A2(KEYINPUT37), .ZN(new_n931));
  AOI22_X1  g0731(.A1(new_n931), .A2(KEYINPUT101), .B1(new_n404), .B2(new_n896), .ZN(new_n932));
  AOI21_X1  g0732(.A(KEYINPUT38), .B1(new_n932), .B2(new_n895), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n930), .A2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(new_n905), .ZN(new_n935));
  OAI21_X1  g0735(.A(KEYINPUT39), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n308), .A2(new_n693), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  AOI21_X1  g0738(.A(KEYINPUT39), .B1(new_n920), .B2(new_n902), .ZN(new_n939));
  INV_X1    g0739(.A(new_n939), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n936), .A2(new_n938), .A3(new_n940), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n930), .B(new_n901), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n910), .A2(new_n913), .ZN(new_n943));
  INV_X1    g0743(.A(new_n943), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n944), .B1(new_n841), .B2(new_n831), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n942), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n659), .A2(new_n674), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n941), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n665), .B1(new_n715), .B2(new_n433), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n948), .B(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n929), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n951), .B1(new_n249), .B2(new_n748), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n929), .A2(new_n950), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n884), .B1(new_n952), .B2(new_n953), .ZN(G367));
  NAND2_X1  g0754(.A1(new_n749), .A2(G1), .ZN(new_n955));
  INV_X1    g0755(.A(new_n955), .ZN(new_n956));
  NOR2_X1   g0756(.A1(KEYINPUT105), .A2(KEYINPUT44), .ZN(new_n957));
  XOR2_X1   g0757(.A(new_n957), .B(KEYINPUT106), .Z(new_n958));
  INV_X1    g0758(.A(new_n958), .ZN(new_n959));
  OAI211_X1 g0759(.A(new_n578), .B(new_n571), .C1(new_n570), .C2(new_n693), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n632), .A2(new_n676), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n694), .A2(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT105), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT44), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n959), .B1(new_n963), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n686), .A2(new_n692), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n681), .A2(new_n693), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n968), .A2(new_n969), .A3(new_n962), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT45), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n694), .A2(KEYINPUT45), .A3(new_n962), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  OAI221_X1 g0774(.A(new_n958), .B1(new_n964), .B2(new_n965), .C1(new_n694), .C2(new_n962), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n967), .A2(new_n974), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(new_n691), .ZN(new_n977));
  NAND4_X1  g0777(.A1(new_n690), .A2(new_n967), .A3(new_n974), .A4(new_n975), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  AOI21_X1  g0779(.A(KEYINPUT107), .B1(new_n686), .B2(new_n692), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n980), .B1(new_n686), .B2(new_n692), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n680), .A2(KEYINPUT108), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT107), .ZN(new_n983));
  OR3_X1    g0783(.A1(new_n686), .A2(new_n983), .A3(new_n692), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n981), .A2(new_n982), .A3(new_n984), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n680), .A2(KEYINPUT108), .ZN(new_n986));
  AND2_X1   g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n985), .A2(new_n986), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(new_n989), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n744), .B1(new_n979), .B2(new_n990), .ZN(new_n991));
  XOR2_X1   g0791(.A(new_n696), .B(KEYINPUT41), .Z(new_n992));
  OAI21_X1  g0792(.A(new_n956), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n578), .B1(new_n960), .B2(new_n533), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT104), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n996), .A2(new_n676), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n994), .A2(new_n995), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n686), .A2(new_n692), .A3(new_n962), .ZN(new_n999));
  AOI22_X1  g0799(.A1(new_n997), .A2(new_n998), .B1(KEYINPUT42), .B2(new_n999), .ZN(new_n1000));
  OR2_X1    g0800(.A1(new_n999), .A2(KEYINPUT42), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  OR3_X1    g0802(.A1(new_n634), .A2(new_n628), .A3(new_n693), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n629), .B1(new_n628), .B2(new_n693), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT43), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1005), .A2(KEYINPUT43), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1002), .A2(new_n1008), .A3(new_n1009), .ZN(new_n1010));
  NAND4_X1  g0810(.A1(new_n1000), .A2(new_n1007), .A3(new_n1006), .A4(new_n1001), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n690), .A2(new_n962), .ZN(new_n1013));
  XOR2_X1   g0813(.A(new_n1012), .B(new_n1013), .Z(new_n1014));
  NAND2_X1  g0814(.A1(new_n993), .A2(new_n1014), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n234), .A2(new_n757), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n764), .B1(new_n412), .B2(new_n204), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n751), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(G159), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n280), .B1(new_n779), .B2(new_n371), .C1(new_n1019), .C2(new_n786), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n798), .A2(new_n261), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1021), .B1(G50), .B2(new_n857), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1022), .B1(new_n329), .B2(new_n795), .ZN(new_n1023));
  AOI211_X1 g0823(.A(new_n1020), .B(new_n1023), .C1(G143), .C2(new_n803), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1024), .B1(new_n267), .B2(new_n791), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1025), .B1(G137), .B2(new_n776), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n780), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n366), .B1(new_n800), .B2(new_n799), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1028), .B1(G97), .B2(new_n810), .ZN(new_n1029));
  OAI211_X1 g0829(.A(new_n1027), .B(new_n1029), .C1(new_n849), .C2(new_n813), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n779), .ZN(new_n1031));
  AOI21_X1  g0831(.A(KEYINPUT46), .B1(new_n1031), .B2(G116), .ZN(new_n1032));
  XOR2_X1   g0832(.A(KEYINPUT109), .B(G311), .Z(new_n1033));
  INV_X1    g0833(.A(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1032), .B1(new_n803), .B2(new_n1034), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n1035), .B1(new_n851), .B2(new_n786), .C1(new_n791), .C2(new_n420), .ZN(new_n1036));
  AOI211_X1 g0836(.A(new_n1030), .B(new_n1036), .C1(G317), .C2(new_n776), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n1026), .A2(new_n1037), .ZN(new_n1038));
  XOR2_X1   g0838(.A(new_n1038), .B(KEYINPUT47), .Z(new_n1039));
  AOI21_X1  g0839(.A(new_n1018), .B1(new_n1039), .B2(new_n760), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1006), .A2(new_n763), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1015), .A2(new_n1042), .ZN(G387));
  NAND2_X1  g0843(.A1(new_n989), .A2(new_n744), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n745), .B1(new_n987), .B2(new_n988), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1044), .A2(new_n696), .A3(new_n1045), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n752), .A2(new_n699), .B1(new_n420), .B2(new_n205), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n230), .A2(new_n442), .ZN(new_n1048));
  AOI211_X1 g0848(.A(G45), .B(new_n699), .C1(G68), .C2(G77), .ZN(new_n1049));
  XOR2_X1   g0849(.A(KEYINPUT110), .B(KEYINPUT50), .Z(new_n1050));
  OAI21_X1  g0850(.A(new_n1050), .B1(G50), .B2(new_n328), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1049), .A2(new_n1051), .ZN(new_n1052));
  NOR3_X1   g0852(.A1(new_n1050), .A2(G50), .A3(new_n328), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n756), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1047), .B1(new_n1048), .B2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n750), .B1(new_n1055), .B2(new_n764), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n280), .B1(new_n798), .B2(new_n553), .C1(new_n328), .C2(new_n786), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1057), .B1(G159), .B2(new_n803), .ZN(new_n1058));
  AND2_X1   g0858(.A1(new_n604), .A2(new_n609), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1059), .A2(new_n792), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1031), .A2(G77), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n795), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(G50), .A2(new_n1062), .B1(new_n857), .B2(G68), .ZN(new_n1063));
  NAND4_X1  g0863(.A1(new_n1058), .A2(new_n1060), .A3(new_n1061), .A4(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1064), .B1(G150), .B2(new_n776), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n366), .B1(new_n798), .B2(new_n454), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n857), .A2(G303), .B1(G322), .B2(new_n803), .ZN(new_n1067));
  INV_X1    g0867(.A(G317), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n1067), .B1(new_n786), .B2(new_n1033), .C1(new_n813), .C2(new_n1068), .ZN(new_n1069));
  INV_X1    g0869(.A(KEYINPUT48), .ZN(new_n1070));
  OR2_X1    g0870(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n792), .A2(G283), .B1(G294), .B2(new_n1031), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1071), .A2(new_n1072), .A3(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(KEYINPUT49), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  AOI211_X1 g0876(.A(new_n1066), .B(new_n1076), .C1(G326), .C2(new_n776), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1065), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n760), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1056), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n686), .A2(new_n821), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(new_n990), .B2(new_n955), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1046), .A2(new_n1084), .ZN(G393));
  INV_X1    g0885(.A(new_n979), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n696), .B1(new_n1086), .B2(new_n1045), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1087), .B1(new_n1045), .B2(new_n1086), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n962), .A2(new_n821), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n1089), .B(KEYINPUT111), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n776), .A2(G322), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n792), .A2(G116), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n366), .B1(new_n798), .B2(new_n420), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n779), .A2(new_n799), .B1(new_n800), .B2(new_n851), .ZN(new_n1094));
  AOI211_X1 g0894(.A(new_n1093), .B(new_n1094), .C1(G303), .C2(new_n785), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n848), .A2(new_n1068), .B1(new_n795), .B2(new_n801), .ZN(new_n1096));
  XNOR2_X1  g0896(.A(new_n1096), .B(KEYINPUT52), .ZN(new_n1097));
  NAND4_X1  g0897(.A1(new_n1091), .A2(new_n1092), .A3(new_n1095), .A4(new_n1097), .ZN(new_n1098));
  AOI211_X1 g0898(.A(new_n366), .B(new_n853), .C1(G68), .C2(new_n1031), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1099), .B1(new_n859), .B2(new_n775), .ZN(new_n1100));
  XOR2_X1   g0900(.A(new_n1100), .B(KEYINPUT112), .Z(new_n1101));
  NAND2_X1  g0901(.A1(new_n792), .A2(G77), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n857), .A2(new_n360), .B1(G50), .B2(new_n785), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n848), .A2(new_n329), .B1(new_n795), .B2(new_n1019), .ZN(new_n1104));
  AND2_X1   g0904(.A1(new_n1104), .A2(KEYINPUT51), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n1104), .A2(KEYINPUT51), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n1102), .B(new_n1103), .C1(new_n1105), .C2(new_n1106), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1098), .B1(new_n1101), .B2(new_n1107), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(new_n1108), .B(KEYINPUT113), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1109), .A2(new_n760), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n243), .A2(new_n756), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n1111), .B(new_n764), .C1(new_n553), .C2(new_n204), .ZN(new_n1112));
  NAND4_X1  g0912(.A1(new_n1090), .A2(new_n751), .A3(new_n1110), .A4(new_n1112), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1113), .B1(new_n1086), .B2(new_n956), .ZN(new_n1114));
  OR2_X1    g0914(.A1(new_n1088), .A2(new_n1114), .ZN(G390));
  NAND3_X1  g0915(.A1(new_n618), .A2(new_n908), .A3(G330), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(KEYINPUT114), .ZN(new_n1117));
  INV_X1    g0917(.A(KEYINPUT114), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n927), .A2(new_n1118), .A3(G330), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n949), .B1(new_n1117), .B2(new_n1119), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n833), .A2(new_n667), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n742), .A2(new_n943), .A3(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n943), .B1(new_n908), .B2(new_n1121), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n837), .A2(new_n427), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n713), .A2(new_n693), .A3(new_n1126), .ZN(new_n1127));
  AND2_X1   g0927(.A1(new_n1127), .A2(new_n831), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1125), .A2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n908), .A2(new_n943), .A3(new_n1121), .ZN(new_n1130));
  AND2_X1   g0930(.A1(new_n742), .A2(new_n1121), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1130), .B1(new_n1131), .B2(new_n943), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n841), .A2(new_n831), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1129), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1120), .A2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n938), .B1(new_n920), .B2(new_n902), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1137), .B1(new_n1128), .B2(new_n944), .ZN(new_n1138));
  INV_X1    g0938(.A(KEYINPUT39), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1139), .B1(new_n903), .B2(new_n905), .ZN(new_n1140));
  OAI22_X1  g0940(.A1(new_n1140), .A2(new_n939), .B1(new_n945), .B2(new_n938), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1138), .A2(new_n1141), .A3(new_n1122), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1133), .A2(new_n943), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n936), .A2(new_n940), .B1(new_n1143), .B2(new_n937), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1137), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1127), .A2(new_n831), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1145), .B1(new_n1146), .B2(new_n943), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n1144), .A2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1142), .B1(new_n1148), .B2(new_n1130), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n700), .B1(new_n1136), .B2(new_n1149), .ZN(new_n1150));
  NOR3_X1   g0950(.A1(new_n1144), .A2(new_n1147), .A3(new_n1123), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1130), .B1(new_n1138), .B2(new_n1141), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1153), .A2(new_n1120), .A3(new_n1135), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1150), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1153), .A2(new_n955), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n761), .B1(new_n1140), .B2(new_n939), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n871), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n751), .B1(new_n360), .B2(new_n1158), .ZN(new_n1159));
  XNOR2_X1  g0959(.A(KEYINPUT54), .B(G143), .ZN(new_n1160));
  OAI22_X1  g0960(.A1(new_n798), .A2(new_n258), .B1(new_n800), .B2(new_n1160), .ZN(new_n1161));
  AOI211_X1 g0961(.A(new_n366), .B(new_n1161), .C1(G132), .C2(new_n1062), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n792), .A2(G159), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n779), .A2(new_n329), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT53), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(new_n1164), .A2(new_n1165), .B1(new_n803), .B2(G128), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1164), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n1167), .A2(KEYINPUT53), .B1(new_n785), .B2(G137), .ZN(new_n1168));
  NAND4_X1  g0968(.A1(new_n1162), .A2(new_n1163), .A3(new_n1166), .A4(new_n1168), .ZN(new_n1169));
  AND2_X1   g0969(.A1(new_n776), .A2(G125), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(new_n857), .A2(G97), .B1(G283), .B2(new_n803), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1171), .B1(new_n420), .B2(new_n786), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1172), .A2(KEYINPUT115), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n780), .A2(G87), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n366), .B1(new_n798), .B2(new_n267), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1175), .B1(G116), .B2(new_n1062), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n1173), .A2(new_n1174), .A3(new_n1102), .A4(new_n1176), .ZN(new_n1177));
  OAI22_X1  g0977(.A1(new_n1172), .A2(KEYINPUT115), .B1(new_n775), .B2(new_n851), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n1169), .A2(new_n1170), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1159), .B1(new_n1179), .B2(new_n760), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1157), .A2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1155), .A2(new_n1156), .A3(new_n1181), .ZN(G378));
  NOR3_X1   g0982(.A1(new_n1140), .A2(new_n937), .A3(new_n939), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n947), .B1(new_n1143), .B2(new_n906), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n943), .A2(new_n838), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1186), .B1(new_n926), .B2(new_n907), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n667), .B1(new_n1187), .B2(new_n921), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n334), .A2(new_n888), .ZN(new_n1189));
  XNOR2_X1  g0989(.A(new_n1189), .B(KEYINPUT55), .ZN(new_n1190));
  OR2_X1    g0990(.A1(new_n346), .A2(new_n1190), .ZN(new_n1191));
  XOR2_X1   g0991(.A(KEYINPUT119), .B(KEYINPUT56), .Z(new_n1192));
  NAND2_X1  g0992(.A1(new_n346), .A2(new_n1190), .ZN(new_n1193));
  AND3_X1   g0993(.A1(new_n1191), .A2(new_n1192), .A3(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1192), .B1(new_n1191), .B2(new_n1193), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  AND3_X1   g0996(.A1(new_n916), .A2(new_n1188), .A3(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1196), .B1(new_n916), .B2(new_n1188), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1185), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1196), .ZN(new_n1200));
  AOI21_X1  g1000(.A(KEYINPUT40), .B1(new_n942), .B2(new_n1187), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n922), .A2(G330), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1200), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n916), .A2(new_n1188), .A3(new_n1196), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1203), .A2(new_n948), .A3(new_n1204), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1199), .A2(new_n1205), .A3(KEYINPUT120), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT120), .ZN(new_n1207));
  NAND4_X1  g1007(.A1(new_n1203), .A2(new_n948), .A3(new_n1207), .A4(new_n1204), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1206), .A2(new_n955), .A3(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1196), .A2(new_n761), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n751), .B1(G50), .B2(new_n1158), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n280), .A2(G41), .ZN(new_n1212));
  AND2_X1   g1012(.A1(new_n1061), .A2(new_n1212), .ZN(new_n1213));
  OAI221_X1 g1013(.A(new_n1213), .B1(new_n371), .B2(new_n798), .C1(new_n775), .C2(new_n799), .ZN(new_n1214));
  XOR2_X1   g1014(.A(new_n1214), .B(KEYINPUT116), .Z(new_n1215));
  NOR2_X1   g1015(.A1(new_n795), .A2(new_n420), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1216), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(new_n1217), .A2(KEYINPUT117), .B1(new_n803), .B2(G116), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT117), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n1216), .A2(new_n1219), .B1(G97), .B2(new_n785), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1218), .B(new_n1220), .C1(new_n791), .C2(new_n267), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1221), .B1(new_n1059), .B2(new_n857), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1215), .A2(KEYINPUT58), .A3(new_n1222), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(G33), .A2(G41), .ZN(new_n1224));
  NOR3_X1   g1024(.A1(new_n1212), .A2(G50), .A3(new_n1224), .ZN(new_n1225));
  XOR2_X1   g1025(.A(KEYINPUT118), .B(G124), .Z(new_n1226));
  OAI221_X1 g1026(.A(new_n1224), .B1(new_n1019), .B2(new_n798), .C1(new_n775), .C2(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(G128), .ZN(new_n1228));
  OAI22_X1  g1028(.A1(new_n779), .A2(new_n1160), .B1(new_n795), .B2(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1229), .B1(G137), .B2(new_n857), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(new_n785), .A2(G132), .B1(new_n803), .B2(G125), .ZN(new_n1231));
  OAI211_X1 g1031(.A(new_n1230), .B(new_n1231), .C1(new_n329), .C2(new_n791), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1227), .B1(new_n1232), .B2(KEYINPUT59), .ZN(new_n1233));
  OR2_X1    g1033(.A1(new_n1232), .A2(KEYINPUT59), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1225), .B1(new_n1233), .B2(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1223), .A2(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(KEYINPUT58), .B1(new_n1215), .B2(new_n1222), .ZN(new_n1237));
  OR2_X1    g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1211), .B1(new_n1238), .B2(new_n760), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1210), .A2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1209), .A2(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT57), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1206), .A2(new_n1208), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1119), .A2(new_n1117), .ZN(new_n1244));
  OAI211_X1 g1044(.A(new_n1244), .B(new_n665), .C1(new_n433), .C2(new_n715), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1245), .B1(new_n1153), .B2(new_n1135), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1242), .B1(new_n1243), .B2(new_n1246), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(new_n1125), .A2(new_n1128), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1120), .B1(new_n1149), .B2(new_n1248), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1242), .B1(new_n1199), .B2(new_n1205), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n700), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1241), .B1(new_n1247), .B2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT121), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  AOI211_X1 g1054(.A(KEYINPUT121), .B(new_n1241), .C1(new_n1247), .C2(new_n1251), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n1254), .A2(new_n1255), .ZN(G375));
  NAND2_X1  g1056(.A1(new_n1245), .A2(new_n1248), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n992), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1136), .A2(new_n1257), .A3(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n944), .A2(new_n761), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n786), .A2(new_n1160), .ZN(new_n1261));
  OAI221_X1 g1061(.A(new_n280), .B1(new_n800), .B2(new_n329), .C1(new_n371), .C2(new_n798), .ZN(new_n1262));
  AOI211_X1 g1062(.A(new_n1261), .B(new_n1262), .C1(G132), .C2(new_n803), .ZN(new_n1263));
  AOI22_X1  g1063(.A1(new_n780), .A2(G159), .B1(new_n814), .B2(G137), .ZN(new_n1264));
  AND2_X1   g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  OAI221_X1 g1065(.A(new_n1265), .B1(new_n258), .B2(new_n791), .C1(new_n1228), .C2(new_n775), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n776), .A2(G303), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n780), .A2(G97), .ZN(new_n1268));
  OAI22_X1  g1068(.A1(new_n786), .A2(new_n454), .B1(new_n848), .B2(new_n851), .ZN(new_n1269));
  OAI22_X1  g1069(.A1(new_n795), .A2(new_n799), .B1(new_n800), .B2(new_n420), .ZN(new_n1270));
  NOR4_X1   g1070(.A1(new_n1269), .A2(new_n1270), .A3(new_n280), .A4(new_n1021), .ZN(new_n1271));
  NAND4_X1  g1071(.A1(new_n1060), .A2(new_n1267), .A3(new_n1268), .A4(new_n1271), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1080), .B1(new_n1266), .B2(new_n1272), .ZN(new_n1273));
  AOI211_X1 g1073(.A(new_n750), .B(new_n1273), .C1(new_n267), .C2(new_n871), .ZN(new_n1274));
  XNOR2_X1  g1074(.A(new_n1274), .B(KEYINPUT122), .ZN(new_n1275));
  AOI22_X1  g1075(.A1(new_n1135), .A2(new_n955), .B1(new_n1260), .B2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1259), .A2(new_n1276), .ZN(G381));
  NAND3_X1  g1077(.A1(new_n1046), .A2(new_n1084), .A3(new_n827), .ZN(new_n1278));
  OR4_X1    g1078(.A1(G384), .A2(G390), .A3(G381), .A4(new_n1278), .ZN(new_n1279));
  OR4_X1    g1079(.A1(G387), .A2(new_n1279), .A3(G378), .A4(G375), .ZN(G407));
  INV_X1    g1080(.A(G378), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1281), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1282));
  OAI211_X1 g1082(.A(G407), .B(G213), .C1(G343), .C2(new_n1282), .ZN(G409));
  AOI21_X1  g1083(.A(new_n827), .B1(new_n1046), .B2(new_n1084), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1284), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(G387), .A2(new_n1278), .A3(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1285), .A2(new_n1278), .ZN(new_n1287));
  AOI22_X1  g1087(.A1(new_n993), .A2(new_n1014), .B1(new_n1041), .B2(new_n1040), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1287), .B1(new_n1288), .B2(KEYINPUT126), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1286), .A2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(G390), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1286), .A2(new_n1289), .A3(G390), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1294), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n956), .B1(new_n1199), .B2(new_n1205), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1296), .B1(new_n1210), .B2(new_n1239), .ZN(new_n1297));
  NAND4_X1  g1097(.A1(new_n1249), .A2(new_n1258), .A3(new_n1208), .A4(new_n1206), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1281), .A2(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1247), .A2(new_n1251), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1241), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1300), .B1(new_n1303), .B2(new_n1281), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n675), .A2(G213), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1245), .A2(new_n1248), .A3(KEYINPUT60), .ZN(new_n1306));
  AND2_X1   g1106(.A1(new_n1306), .A2(new_n696), .ZN(new_n1307));
  OAI21_X1  g1107(.A(KEYINPUT60), .B1(new_n1245), .B2(new_n1248), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1308), .A2(new_n1257), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1307), .A2(new_n1309), .ZN(new_n1310));
  AOI21_X1  g1110(.A(G384), .B1(new_n1310), .B2(new_n1276), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1276), .ZN(new_n1312));
  AOI211_X1 g1112(.A(new_n875), .B(new_n1312), .C1(new_n1307), .C2(new_n1309), .ZN(new_n1313));
  NOR2_X1   g1113(.A1(new_n1311), .A2(new_n1313), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1304), .A2(new_n1305), .A3(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT63), .ZN(new_n1316));
  NOR2_X1   g1116(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1317));
  NOR2_X1   g1117(.A1(new_n1295), .A2(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT61), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1305), .ZN(new_n1321));
  AND2_X1   g1121(.A1(new_n1321), .A2(G2897), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1322), .B1(new_n1311), .B2(new_n1313), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1321), .B1(KEYINPUT124), .B2(G2897), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n1324), .B1(KEYINPUT124), .B2(G2897), .ZN(new_n1325));
  NOR3_X1   g1125(.A1(new_n1311), .A2(new_n1313), .A3(new_n1325), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT125), .ZN(new_n1327));
  OAI21_X1  g1127(.A(new_n1323), .B1(new_n1326), .B2(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1314), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1329), .A2(KEYINPUT125), .A3(new_n1322), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1320), .A2(new_n1328), .A3(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1315), .A2(KEYINPUT123), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT123), .ZN(new_n1333));
  NAND4_X1  g1133(.A1(new_n1304), .A2(new_n1333), .A3(new_n1305), .A4(new_n1314), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1332), .A2(new_n1316), .A3(new_n1334), .ZN(new_n1335));
  NAND4_X1  g1135(.A1(new_n1318), .A2(new_n1319), .A3(new_n1331), .A4(new_n1335), .ZN(new_n1336));
  AOI21_X1  g1136(.A(KEYINPUT62), .B1(new_n1332), .B2(new_n1334), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1315), .A2(KEYINPUT62), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1338), .A2(new_n1331), .A3(new_n1319), .ZN(new_n1339));
  OAI21_X1  g1139(.A(new_n1295), .B1(new_n1337), .B2(new_n1339), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1336), .A2(new_n1340), .ZN(G405));
  NAND2_X1  g1141(.A1(new_n1303), .A2(KEYINPUT121), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1343));
  AOI21_X1  g1143(.A(G378), .B1(new_n1342), .B2(new_n1343), .ZN(new_n1344));
  NOR2_X1   g1144(.A1(new_n1252), .A2(new_n1281), .ZN(new_n1345));
  OAI21_X1  g1145(.A(new_n1314), .B1(new_n1344), .B2(new_n1345), .ZN(new_n1346));
  INV_X1    g1146(.A(new_n1345), .ZN(new_n1347));
  NAND3_X1  g1147(.A1(new_n1282), .A2(new_n1329), .A3(new_n1347), .ZN(new_n1348));
  NAND3_X1  g1148(.A1(new_n1346), .A2(new_n1294), .A3(new_n1348), .ZN(new_n1349));
  AOI21_X1  g1149(.A(new_n1294), .B1(new_n1346), .B2(new_n1348), .ZN(new_n1350));
  INV_X1    g1150(.A(KEYINPUT127), .ZN(new_n1351));
  OAI21_X1  g1151(.A(new_n1349), .B1(new_n1350), .B2(new_n1351), .ZN(new_n1352));
  AOI211_X1 g1152(.A(KEYINPUT127), .B(new_n1294), .C1(new_n1346), .C2(new_n1348), .ZN(new_n1353));
  NOR2_X1   g1153(.A1(new_n1352), .A2(new_n1353), .ZN(G402));
endmodule


