//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0 1 0 1 0 1 1 1 0 0 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 0 1 0 1 0 0 1 0 1 1 1 0 1 1 0 0 1 0 1 0 1 1 0 0 1 0 1 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:07 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1256, new_n1257, new_n1258, new_n1260, new_n1261,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1324, new_n1325, new_n1326;
  INV_X1    g0000(.A(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G58), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NOR2_X1   g0005(.A1(G58), .A2(G68), .ZN(new_n206));
  INV_X1    g0006(.A(KEYINPUT64), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  OAI21_X1  g0008(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n209));
  NAND3_X1  g0009(.A1(new_n208), .A2(G50), .A3(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  INV_X1    g0012(.A(G20), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n211), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G20), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n216), .A2(G13), .ZN(new_n217));
  OAI211_X1 g0017(.A(new_n217), .B(G250), .C1(G257), .C2(G264), .ZN(new_n218));
  XNOR2_X1  g0018(.A(new_n218), .B(KEYINPUT0), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n220));
  INV_X1    g0020(.A(G58), .ZN(new_n221));
  INV_X1    g0021(.A(G232), .ZN(new_n222));
  INV_X1    g0022(.A(G107), .ZN(new_n223));
  INV_X1    g0023(.A(G264), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n220), .B1(new_n221), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(KEYINPUT65), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n229));
  NAND3_X1  g0029(.A1(new_n227), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n225), .A2(new_n226), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n216), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  OAI211_X1 g0032(.A(new_n215), .B(new_n219), .C1(new_n232), .C2(KEYINPUT1), .ZN(new_n233));
  AOI21_X1  g0033(.A(new_n233), .B1(KEYINPUT1), .B2(new_n232), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(new_n222), .ZN(new_n236));
  XOR2_X1   g0036(.A(KEYINPUT2), .B(G226), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT66), .ZN(new_n240));
  XOR2_X1   g0040(.A(G264), .B(G270), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n238), .B(new_n242), .Z(G358));
  NAND2_X1  g0043(.A1(G68), .A2(G77), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n203), .A2(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n245), .B(KEYINPUT67), .Z(new_n246));
  XNOR2_X1  g0046(.A(G50), .B(G58), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(G87), .B(G97), .Z(new_n249));
  XNOR2_X1  g0049(.A(G107), .B(G116), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(new_n248), .B(new_n251), .Z(G351));
  INV_X1    g0052(.A(G13), .ZN(new_n253));
  NOR3_X1   g0053(.A1(new_n253), .A2(new_n213), .A3(G1), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n255), .A2(G50), .ZN(new_n256));
  NAND3_X1  g0056(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(new_n212), .ZN(new_n258));
  INV_X1    g0058(.A(G1), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n258), .B1(new_n259), .B2(G20), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n256), .B1(new_n260), .B2(G50), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  NOR2_X1   g0062(.A1(G50), .A2(G58), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n213), .B1(new_n263), .B2(new_n201), .ZN(new_n264));
  XNOR2_X1  g0064(.A(KEYINPUT8), .B(G58), .ZN(new_n265));
  XNOR2_X1  g0065(.A(new_n265), .B(KEYINPUT70), .ZN(new_n266));
  INV_X1    g0066(.A(G33), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n267), .A2(G20), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G150), .ZN(new_n270));
  NOR2_X1   g0070(.A1(G20), .A2(G33), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n269), .B1(new_n270), .B2(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n264), .B1(new_n273), .B2(KEYINPUT71), .ZN(new_n274));
  AOI22_X1  g0074(.A1(new_n266), .A2(new_n268), .B1(G150), .B2(new_n271), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT71), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n274), .A2(new_n277), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n262), .B1(new_n278), .B2(new_n258), .ZN(new_n279));
  INV_X1    g0079(.A(G274), .ZN(new_n280));
  AND2_X1   g0080(.A1(G1), .A2(G13), .ZN(new_n281));
  NAND2_X1  g0081(.A1(G33), .A2(G41), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n280), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G41), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(KEYINPUT68), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT68), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(G41), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  OAI211_X1 g0088(.A(new_n283), .B(new_n259), .C1(new_n288), .C2(G45), .ZN(new_n289));
  INV_X1    g0089(.A(G45), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n284), .A2(new_n290), .ZN(new_n291));
  AOI22_X1  g0091(.A1(new_n259), .A2(new_n291), .B1(new_n281), .B2(new_n282), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(G226), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n289), .A2(new_n293), .ZN(new_n294));
  OR2_X1    g0094(.A1(G222), .A2(G1698), .ZN(new_n295));
  XNOR2_X1  g0095(.A(KEYINPUT69), .B(G223), .ZN(new_n296));
  INV_X1    g0096(.A(G1698), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n295), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  XNOR2_X1  g0098(.A(KEYINPUT3), .B(G33), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n281), .A2(new_n282), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT3), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(G33), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n267), .A2(KEYINPUT3), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n301), .B1(new_n305), .B2(new_n202), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n294), .B1(new_n300), .B2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G179), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n309), .B1(G169), .B2(new_n307), .ZN(new_n310));
  OR2_X1    g0110(.A1(new_n279), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT10), .ZN(new_n312));
  XOR2_X1   g0112(.A(KEYINPUT73), .B(G200), .Z(new_n313));
  NOR2_X1   g0113(.A1(new_n307), .A2(new_n313), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n314), .B1(G190), .B2(new_n307), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n277), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n275), .A2(new_n276), .ZN(new_n318));
  NOR3_X1   g0118(.A1(new_n317), .A2(new_n264), .A3(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n258), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n261), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT9), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n316), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n320), .B1(new_n274), .B2(new_n277), .ZN(new_n324));
  NOR3_X1   g0124(.A1(new_n324), .A2(new_n322), .A3(new_n262), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n312), .B1(new_n323), .B2(new_n326), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n322), .B1(new_n324), .B2(new_n262), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(new_n315), .ZN(new_n329));
  NOR3_X1   g0129(.A1(new_n329), .A2(KEYINPUT10), .A3(new_n325), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n311), .B1(new_n327), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n292), .A2(G232), .ZN(new_n332));
  AND2_X1   g0132(.A1(new_n289), .A2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(new_n301), .ZN(new_n334));
  INV_X1    g0134(.A(G226), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(G1698), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n336), .B1(G223), .B2(G1698), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n302), .A2(KEYINPUT76), .A3(G33), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT76), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n303), .A2(new_n304), .A3(new_n339), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n337), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(G87), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n267), .A2(new_n342), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n334), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  AND3_X1   g0144(.A1(new_n333), .A2(new_n344), .A3(G179), .ZN(new_n345));
  INV_X1    g0145(.A(G169), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n346), .B1(new_n333), .B2(new_n344), .ZN(new_n347));
  OR2_X1    g0147(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n221), .A2(new_n201), .ZN(new_n349));
  OAI21_X1  g0149(.A(G20), .B1(new_n349), .B2(new_n206), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n271), .A2(G159), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT7), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n353), .B1(new_n299), .B2(G20), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n305), .A2(KEYINPUT7), .A3(new_n213), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n352), .B1(new_n356), .B2(G68), .ZN(new_n357));
  XOR2_X1   g0157(.A(KEYINPUT78), .B(KEYINPUT16), .Z(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n258), .B1(new_n357), .B2(new_n359), .ZN(new_n360));
  AND3_X1   g0160(.A1(new_n350), .A2(KEYINPUT16), .A3(new_n351), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n340), .A2(new_n213), .A3(new_n338), .ZN(new_n362));
  AND2_X1   g0162(.A1(new_n362), .A2(KEYINPUT7), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n340), .A2(new_n353), .A3(new_n213), .A4(new_n338), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(G68), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n361), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT77), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  OAI211_X1 g0168(.A(KEYINPUT77), .B(new_n361), .C1(new_n363), .C2(new_n365), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n360), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n266), .A2(new_n254), .ZN(new_n371));
  INV_X1    g0171(.A(new_n260), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n371), .B1(new_n266), .B2(new_n372), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n348), .B1(new_n370), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(KEYINPUT18), .ZN(new_n375));
  NOR3_X1   g0175(.A1(new_n299), .A2(new_n353), .A3(G20), .ZN(new_n376));
  AOI21_X1  g0176(.A(KEYINPUT7), .B1(new_n305), .B2(new_n213), .ZN(new_n377));
  OAI21_X1  g0177(.A(G68), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(new_n352), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n320), .B1(new_n380), .B2(new_n358), .ZN(new_n381));
  INV_X1    g0181(.A(new_n369), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n362), .A2(KEYINPUT7), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n383), .A2(G68), .A3(new_n364), .ZN(new_n384));
  AOI21_X1  g0184(.A(KEYINPUT77), .B1(new_n384), .B2(new_n361), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n381), .B1(new_n382), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n333), .A2(new_n344), .ZN(new_n387));
  INV_X1    g0187(.A(G200), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n389), .B1(G190), .B2(new_n387), .ZN(new_n390));
  INV_X1    g0190(.A(new_n373), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n386), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT17), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT18), .ZN(new_n395));
  OAI211_X1 g0195(.A(new_n348), .B(new_n395), .C1(new_n370), .C2(new_n373), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n386), .A2(new_n390), .A3(KEYINPUT17), .A4(new_n391), .ZN(new_n397));
  NAND4_X1  g0197(.A1(new_n375), .A2(new_n394), .A3(new_n396), .A4(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n292), .A2(G238), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n289), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n335), .A2(new_n297), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n222), .A2(G1698), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n299), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(G33), .A2(G97), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n301), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT74), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT13), .ZN(new_n407));
  NOR4_X1   g0207(.A1(new_n400), .A2(new_n405), .A3(new_n406), .A4(new_n407), .ZN(new_n408));
  AND2_X1   g0208(.A1(new_n289), .A2(new_n399), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n403), .A2(new_n404), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(new_n334), .ZN(new_n411));
  AOI22_X1  g0211(.A1(new_n409), .A2(new_n411), .B1(KEYINPUT74), .B2(KEYINPUT13), .ZN(new_n412));
  OAI21_X1  g0212(.A(G179), .B1(new_n408), .B2(new_n412), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n411), .A2(KEYINPUT13), .A3(new_n289), .A4(new_n399), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n407), .B1(new_n400), .B2(new_n405), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT14), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n414), .A2(new_n415), .A3(new_n416), .A4(G169), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n413), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n414), .A2(G169), .A3(new_n415), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT75), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n419), .A2(new_n420), .A3(KEYINPUT14), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n419), .A2(KEYINPUT14), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(KEYINPUT75), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n418), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  NOR3_X1   g0224(.A1(new_n255), .A2(KEYINPUT12), .A3(G68), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT12), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n426), .B1(new_n254), .B2(new_n201), .ZN(new_n427));
  OAI22_X1  g0227(.A1(new_n425), .A2(new_n427), .B1(new_n372), .B2(new_n201), .ZN(new_n428));
  AOI22_X1  g0228(.A1(new_n271), .A2(G50), .B1(G20), .B2(new_n201), .ZN(new_n429));
  INV_X1    g0229(.A(new_n268), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n429), .B1(new_n430), .B2(new_n202), .ZN(new_n431));
  AND3_X1   g0231(.A1(new_n431), .A2(KEYINPUT11), .A3(new_n258), .ZN(new_n432));
  AOI21_X1  g0232(.A(KEYINPUT11), .B1(new_n431), .B2(new_n258), .ZN(new_n433));
  NOR3_X1   g0233(.A1(new_n428), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n424), .A2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n408), .A2(new_n412), .ZN(new_n437));
  INV_X1    g0237(.A(G190), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n414), .A2(G200), .A3(new_n415), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(new_n434), .ZN(new_n441));
  OR2_X1    g0241(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  XNOR2_X1  g0242(.A(KEYINPUT15), .B(G87), .ZN(new_n443));
  OAI21_X1  g0243(.A(KEYINPUT72), .B1(new_n443), .B2(new_n430), .ZN(new_n444));
  NAND2_X1  g0244(.A1(G20), .A2(G77), .ZN(new_n445));
  OAI211_X1 g0245(.A(new_n444), .B(new_n445), .C1(new_n265), .C2(new_n272), .ZN(new_n446));
  NOR3_X1   g0246(.A1(new_n443), .A2(new_n430), .A3(KEYINPUT72), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n258), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n255), .A2(G77), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n449), .B1(new_n260), .B2(G77), .ZN(new_n450));
  AND2_X1   g0250(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n299), .A2(G232), .A3(new_n297), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n299), .A2(G1698), .ZN(new_n453));
  INV_X1    g0253(.A(G238), .ZN(new_n454));
  OAI221_X1 g0254(.A(new_n452), .B1(new_n223), .B2(new_n299), .C1(new_n453), .C2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(new_n334), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n292), .A2(G244), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n456), .A2(new_n289), .A3(new_n457), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n451), .B1(new_n458), .B2(new_n438), .ZN(new_n459));
  INV_X1    g0259(.A(new_n313), .ZN(new_n460));
  AND2_X1   g0260(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n451), .B1(new_n458), .B2(new_n346), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n464), .B1(G179), .B2(new_n458), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n436), .A2(new_n442), .A3(new_n463), .A4(new_n465), .ZN(new_n466));
  NOR3_X1   g0266(.A1(new_n331), .A2(new_n398), .A3(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  AOI21_X1  g0268(.A(KEYINPUT5), .B1(new_n285), .B2(new_n287), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n259), .A2(G45), .ZN(new_n470));
  OAI21_X1  g0270(.A(KEYINPUT80), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n284), .A2(KEYINPUT5), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT80), .ZN(new_n473));
  INV_X1    g0273(.A(new_n470), .ZN(new_n474));
  XNOR2_X1  g0274(.A(KEYINPUT68), .B(G41), .ZN(new_n475));
  OAI211_X1 g0275(.A(new_n473), .B(new_n474), .C1(new_n475), .C2(KEYINPUT5), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n471), .A2(new_n283), .A3(new_n472), .A4(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n224), .A2(G1698), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n478), .B1(G257), .B2(G1698), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n479), .B1(new_n338), .B2(new_n340), .ZN(new_n480));
  INV_X1    g0280(.A(G303), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n299), .A2(new_n481), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n334), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  AND2_X1   g0283(.A1(new_n477), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n476), .A2(new_n472), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT5), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n288), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n473), .B1(new_n487), .B2(new_n474), .ZN(new_n488));
  OAI211_X1 g0288(.A(G270), .B(new_n301), .C1(new_n485), .C2(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n484), .A2(G190), .A3(new_n489), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n255), .B(new_n320), .C1(G1), .C2(new_n267), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(G116), .ZN(new_n492));
  INV_X1    g0292(.A(G116), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n255), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(G33), .A2(G283), .ZN(new_n496));
  INV_X1    g0296(.A(G97), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n496), .B(new_n213), .C1(G33), .C2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n493), .A2(G20), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n498), .A2(new_n258), .A3(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT20), .ZN(new_n501));
  OR2_X1    g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n500), .A2(new_n501), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n502), .A2(KEYINPUT84), .A3(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT84), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n500), .A2(new_n505), .A3(new_n501), .ZN(new_n506));
  AND3_X1   g0306(.A1(new_n495), .A2(new_n504), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n490), .A2(new_n507), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n388), .B1(new_n484), .B2(new_n489), .ZN(new_n509));
  OAI21_X1  g0309(.A(KEYINPUT85), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n489), .A2(new_n477), .A3(new_n483), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(G200), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT85), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n512), .A2(new_n513), .A3(new_n507), .A4(new_n490), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n510), .A2(new_n514), .ZN(new_n515));
  NOR3_X1   g0315(.A1(new_n507), .A2(new_n511), .A3(new_n308), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n495), .A2(new_n504), .A3(new_n506), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n511), .A2(new_n517), .A3(G169), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(KEYINPUT21), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n346), .B1(new_n484), .B2(new_n489), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT21), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n520), .A2(new_n521), .A3(new_n517), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n516), .B1(new_n519), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n515), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n271), .A2(G77), .ZN(new_n525));
  XNOR2_X1  g0325(.A(G97), .B(G107), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT79), .ZN(new_n527));
  OR2_X1    g0327(.A1(new_n527), .A2(KEYINPUT6), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  MUX2_X1   g0329(.A(new_n527), .B(G97), .S(KEYINPUT6), .Z(new_n530));
  OAI21_X1  g0330(.A(new_n529), .B1(new_n530), .B2(new_n526), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n525), .B1(new_n531), .B2(new_n213), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n223), .B1(new_n354), .B2(new_n355), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n258), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n255), .A2(G97), .ZN(new_n535));
  INV_X1    g0335(.A(new_n491), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n535), .B1(new_n536), .B2(G97), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n534), .A2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(G244), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n539), .B1(new_n340), .B2(new_n338), .ZN(new_n540));
  AOI21_X1  g0340(.A(KEYINPUT4), .B1(new_n540), .B2(new_n297), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n299), .A2(KEYINPUT4), .A3(G244), .A4(new_n297), .ZN(new_n542));
  INV_X1    g0342(.A(G250), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n542), .B(new_n496), .C1(new_n543), .C2(new_n453), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n334), .B1(new_n541), .B2(new_n544), .ZN(new_n545));
  OAI211_X1 g0345(.A(G257), .B(new_n301), .C1(new_n485), .C2(new_n488), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n545), .A2(new_n477), .A3(new_n546), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n538), .B1(G200), .B2(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(new_n547), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(G190), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  AOI22_X1  g0351(.A1(new_n547), .A2(new_n346), .B1(new_n534), .B2(new_n537), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n545), .A2(new_n308), .A3(new_n546), .A4(new_n477), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n340), .A2(new_n338), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT22), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n557), .A2(new_n342), .ZN(new_n558));
  AND3_X1   g0358(.A1(new_n556), .A2(new_n213), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(G33), .A2(G116), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n560), .A2(G20), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT23), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n562), .B1(new_n213), .B2(G107), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n223), .A2(KEYINPUT23), .A3(G20), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n561), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n342), .A2(G20), .ZN(new_n566));
  AND2_X1   g0366(.A1(new_n299), .A2(new_n566), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n565), .B1(new_n567), .B2(KEYINPUT22), .ZN(new_n568));
  NOR3_X1   g0368(.A1(new_n559), .A2(new_n568), .A3(KEYINPUT24), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT24), .ZN(new_n570));
  INV_X1    g0370(.A(new_n565), .ZN(new_n571));
  AOI21_X1  g0371(.A(KEYINPUT22), .B1(new_n299), .B2(new_n566), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n556), .A2(new_n213), .A3(new_n558), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n570), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n258), .B1(new_n569), .B2(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT25), .ZN(new_n577));
  NOR3_X1   g0377(.A1(new_n255), .A2(new_n577), .A3(G107), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n577), .B1(new_n255), .B2(G107), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n581), .B1(new_n223), .B2(new_n491), .ZN(new_n582));
  INV_X1    g0382(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n576), .A2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(new_n338), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n585), .B1(new_n339), .B2(new_n299), .ZN(new_n586));
  NOR3_X1   g0386(.A1(new_n586), .A2(new_n543), .A3(G1698), .ZN(new_n587));
  NAND2_X1  g0387(.A1(G257), .A2(G1698), .ZN(new_n588));
  INV_X1    g0388(.A(G294), .ZN(new_n589));
  OAI22_X1  g0389(.A1(new_n586), .A2(new_n588), .B1(new_n267), .B2(new_n589), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n334), .B1(new_n587), .B2(new_n590), .ZN(new_n591));
  OAI211_X1 g0391(.A(G264), .B(new_n301), .C1(new_n485), .C2(new_n488), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n591), .A2(new_n477), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(new_n346), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n591), .A2(new_n308), .A3(new_n477), .A4(new_n592), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n584), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n593), .A2(G200), .ZN(new_n597));
  OAI21_X1  g0397(.A(KEYINPUT24), .B1(new_n559), .B2(new_n568), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n573), .A2(new_n574), .A3(new_n570), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n582), .B1(new_n600), .B2(new_n258), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n591), .A2(G190), .A3(new_n477), .A4(new_n592), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n597), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT19), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n268), .A2(new_n604), .A3(G97), .ZN(new_n605));
  NOR3_X1   g0405(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n606), .B1(new_n213), .B2(new_n404), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n605), .B1(new_n607), .B2(new_n604), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n556), .A2(new_n213), .A3(G68), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n258), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n443), .A2(new_n254), .ZN(new_n612));
  OR2_X1    g0412(.A1(new_n491), .A2(new_n443), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n611), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT83), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n320), .B1(new_n608), .B2(new_n609), .ZN(new_n617));
  INV_X1    g0417(.A(new_n612), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n619), .A2(KEYINPUT83), .A3(new_n613), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n540), .A2(G1698), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n556), .A2(G238), .A3(new_n297), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n621), .A2(new_n560), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(new_n334), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT82), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT81), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n470), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n259), .A2(KEYINPUT81), .A3(G45), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(new_n282), .ZN(new_n630));
  OAI21_X1  g0430(.A(G250), .B1(new_n630), .B2(new_n212), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n625), .B1(new_n629), .B2(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n543), .B1(new_n281), .B2(new_n282), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n633), .A2(KEYINPUT82), .A3(new_n628), .A4(new_n627), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n283), .A2(new_n474), .ZN(new_n636));
  AND2_X1   g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n346), .B1(new_n624), .B2(new_n637), .ZN(new_n638));
  AOI22_X1  g0438(.A1(new_n540), .A2(G1698), .B1(G33), .B2(G116), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n301), .B1(new_n639), .B2(new_n622), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n635), .A2(new_n636), .ZN(new_n641));
  NOR3_X1   g0441(.A1(new_n640), .A2(new_n308), .A3(new_n641), .ZN(new_n642));
  OAI211_X1 g0442(.A(new_n616), .B(new_n620), .C1(new_n638), .C2(new_n642), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n460), .B1(new_n640), .B2(new_n641), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n491), .A2(new_n342), .ZN(new_n645));
  NOR3_X1   g0445(.A1(new_n617), .A2(new_n618), .A3(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n624), .A2(new_n637), .ZN(new_n647));
  OAI211_X1 g0447(.A(new_n644), .B(new_n646), .C1(new_n647), .C2(new_n438), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n596), .A2(new_n603), .A3(new_n643), .A4(new_n648), .ZN(new_n649));
  NOR4_X1   g0449(.A1(new_n468), .A2(new_n524), .A3(new_n555), .A4(new_n649), .ZN(G372));
  INV_X1    g0450(.A(new_n311), .ZN(new_n651));
  INV_X1    g0451(.A(new_n465), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n435), .B1(new_n442), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n394), .A2(new_n397), .ZN(new_n654));
  OAI211_X1 g0454(.A(new_n375), .B(new_n396), .C1(new_n653), .C2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT88), .ZN(new_n656));
  OR2_X1    g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  OAI21_X1  g0457(.A(KEYINPUT10), .B1(new_n329), .B2(new_n325), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n323), .A2(new_n312), .A3(new_n326), .ZN(new_n659));
  AOI22_X1  g0459(.A1(new_n655), .A2(new_n656), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n651), .B1(new_n657), .B2(new_n660), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n643), .A2(new_n553), .A3(new_n552), .A4(new_n648), .ZN(new_n662));
  OAI21_X1  g0462(.A(G169), .B1(new_n640), .B2(new_n641), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n624), .A2(new_n637), .A3(G179), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT86), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n663), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n663), .A2(new_n664), .ZN(new_n667));
  AOI22_X1  g0467(.A1(new_n667), .A2(KEYINPUT86), .B1(new_n619), .B2(new_n613), .ZN(new_n668));
  AOI22_X1  g0468(.A1(new_n662), .A2(KEYINPUT26), .B1(new_n666), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n667), .A2(KEYINPUT86), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n670), .A2(new_n614), .A3(new_n666), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT26), .ZN(new_n672));
  AND2_X1   g0472(.A1(new_n552), .A2(new_n553), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n671), .A2(new_n672), .A3(new_n673), .A4(new_n648), .ZN(new_n674));
  INV_X1    g0474(.A(new_n516), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n521), .B1(new_n520), .B2(new_n517), .ZN(new_n676));
  AND4_X1   g0476(.A1(new_n521), .A2(new_n511), .A3(G169), .A4(new_n517), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n675), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT87), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n596), .A2(new_n679), .ZN(new_n680));
  NAND4_X1  g0480(.A1(new_n584), .A2(new_n594), .A3(KEYINPUT87), .A4(new_n595), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n678), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  AOI22_X1  g0482(.A1(new_n548), .A2(new_n550), .B1(new_n552), .B2(new_n553), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n671), .A2(new_n683), .A3(new_n603), .A4(new_n648), .ZN(new_n684));
  OAI211_X1 g0484(.A(new_n669), .B(new_n674), .C1(new_n682), .C2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n661), .B1(new_n468), .B2(new_n686), .ZN(G369));
  NAND3_X1  g0487(.A1(new_n259), .A2(new_n213), .A3(G13), .ZN(new_n688));
  OR2_X1    g0488(.A1(new_n688), .A2(KEYINPUT27), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(KEYINPUT27), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n689), .A2(G213), .A3(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(G343), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n507), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n678), .A2(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n696), .B1(new_n524), .B2(new_n695), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(G330), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  AND2_X1   g0499(.A1(new_n596), .A2(new_n603), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n700), .B1(new_n601), .B2(new_n694), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n701), .B1(new_n596), .B2(new_n694), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n699), .A2(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n523), .A2(new_n693), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(new_n700), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n680), .A2(new_n681), .A3(new_n694), .ZN(new_n706));
  AND2_X1   g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n703), .A2(new_n707), .ZN(G399));
  INV_X1    g0508(.A(new_n217), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n709), .A2(new_n288), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n606), .A2(new_n493), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n711), .A2(G1), .A3(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n714), .B1(new_n210), .B2(new_n711), .ZN(new_n715));
  XNOR2_X1  g0515(.A(new_n715), .B(KEYINPUT28), .ZN(new_n716));
  OR4_X1    g0516(.A1(new_n524), .A2(new_n649), .A3(new_n555), .A4(new_n693), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n484), .A2(new_n591), .A3(new_n489), .A4(new_n592), .ZN(new_n718));
  NOR3_X1   g0518(.A1(new_n718), .A2(new_n664), .A3(new_n547), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n647), .A2(new_n308), .A3(new_n511), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n593), .A2(new_n547), .ZN(new_n721));
  OAI22_X1  g0521(.A1(new_n719), .A2(KEYINPUT30), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  AND2_X1   g0522(.A1(new_n591), .A2(new_n592), .ZN(new_n723));
  INV_X1    g0523(.A(new_n511), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n549), .A2(new_n723), .A3(new_n642), .A4(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT30), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n693), .B1(new_n722), .B2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT31), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n720), .ZN(new_n731));
  INV_X1    g0531(.A(new_n721), .ZN(new_n732));
  AOI22_X1  g0532(.A1(new_n725), .A2(new_n726), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n719), .A2(KEYINPUT30), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n694), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  XNOR2_X1  g0535(.A(KEYINPUT89), .B(KEYINPUT31), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n717), .A2(new_n730), .A3(new_n738), .ZN(new_n739));
  AND2_X1   g0539(.A1(new_n739), .A2(G330), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n685), .A2(new_n694), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT29), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n673), .A2(new_n643), .A3(new_n672), .A4(new_n648), .ZN(new_n744));
  AND2_X1   g0544(.A1(new_n744), .A2(new_n671), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n671), .A2(new_n648), .ZN(new_n746));
  OAI21_X1  g0546(.A(KEYINPUT26), .B1(new_n746), .B2(new_n554), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n523), .A2(new_n596), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  OAI211_X1 g0549(.A(new_n745), .B(new_n747), .C1(new_n684), .C2(new_n749), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n750), .A2(KEYINPUT29), .A3(new_n694), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n740), .B1(new_n743), .B2(new_n751), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n716), .B1(new_n752), .B2(G1), .ZN(G364));
  NOR2_X1   g0553(.A1(new_n253), .A2(G20), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n259), .B1(new_n754), .B2(G45), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n710), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n699), .A2(new_n757), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n758), .B1(G330), .B2(new_n697), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n709), .A2(new_n305), .ZN(new_n760));
  NAND2_X1  g0560(.A1(G355), .A2(KEYINPUT90), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(G355), .A2(KEYINPUT90), .ZN(new_n763));
  OAI22_X1  g0563(.A1(new_n762), .A2(new_n763), .B1(G116), .B2(new_n217), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n248), .A2(G45), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n556), .A2(new_n709), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n767), .B1(new_n290), .B2(new_n211), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n764), .B1(new_n765), .B2(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(G13), .A2(G33), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(G20), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n212), .B1(G20), .B2(new_n346), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n757), .B1(new_n769), .B2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n213), .A2(new_n308), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(G200), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(G190), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(new_n201), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n388), .A2(G190), .ZN(new_n782));
  NOR3_X1   g0582(.A1(new_n782), .A2(new_n213), .A3(new_n308), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n778), .A2(new_n438), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(G50), .ZN(new_n787));
  OAI221_X1 g0587(.A(new_n299), .B1(new_n221), .B2(new_n784), .C1(new_n786), .C2(new_n787), .ZN(new_n788));
  OAI21_X1  g0588(.A(G20), .B1(new_n782), .B2(G179), .ZN(new_n789));
  INV_X1    g0589(.A(KEYINPUT93), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n789), .A2(new_n790), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  AOI211_X1 g0595(.A(new_n781), .B(new_n788), .C1(G97), .C2(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n213), .A2(G179), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n460), .A2(G190), .A3(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(new_n342), .ZN(new_n799));
  NOR2_X1   g0599(.A1(G190), .A2(G200), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n777), .A2(KEYINPUT91), .A3(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(KEYINPUT91), .B1(new_n777), .B2(new_n800), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n799), .B1(G77), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n797), .A2(new_n800), .ZN(new_n807));
  XNOR2_X1  g0607(.A(KEYINPUT92), .B(G159), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  XNOR2_X1  g0609(.A(new_n809), .B(KEYINPUT32), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n460), .A2(new_n438), .A3(new_n797), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(G107), .ZN(new_n813));
  NAND4_X1  g0613(.A1(new_n796), .A2(new_n806), .A3(new_n810), .A4(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n785), .A2(G326), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n299), .B1(new_n783), .B2(G322), .ZN(new_n816));
  XOR2_X1   g0616(.A(KEYINPUT33), .B(G317), .Z(new_n817));
  OAI211_X1 g0617(.A(new_n815), .B(new_n816), .C1(new_n780), .C2(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n818), .B1(G294), .B2(new_n795), .ZN(new_n819));
  XNOR2_X1  g0619(.A(new_n807), .B(KEYINPUT94), .ZN(new_n820));
  AOI22_X1  g0620(.A1(new_n812), .A2(G283), .B1(new_n820), .B2(G329), .ZN(new_n821));
  INV_X1    g0621(.A(new_n798), .ZN(new_n822));
  AOI22_X1  g0622(.A1(new_n805), .A2(G311), .B1(new_n822), .B2(G303), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n819), .A2(new_n821), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n814), .A2(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n776), .B1(new_n825), .B2(new_n773), .ZN(new_n826));
  INV_X1    g0626(.A(new_n772), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n826), .B1(new_n697), .B2(new_n827), .ZN(new_n828));
  AND2_X1   g0628(.A1(new_n759), .A2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(G396));
  INV_X1    g0630(.A(new_n757), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n465), .A2(KEYINPUT96), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT96), .ZN(new_n833));
  OAI211_X1 g0633(.A(new_n464), .B(new_n833), .C1(G179), .C2(new_n458), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n835), .A2(new_n462), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n685), .A2(new_n694), .A3(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n832), .A2(new_n463), .A3(new_n834), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n451), .A2(new_n694), .ZN(new_n840));
  OAI22_X1  g0640(.A1(new_n839), .A2(new_n840), .B1(new_n465), .B2(new_n694), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n841), .B1(new_n685), .B2(new_n694), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n838), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(new_n740), .ZN(new_n844));
  AND2_X1   g0644(.A1(new_n844), .A2(KEYINPUT97), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n844), .A2(KEYINPUT97), .ZN(new_n846));
  OAI221_X1 g0646(.A(new_n831), .B1(new_n740), .B2(new_n843), .C1(new_n845), .C2(new_n846), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n773), .A2(new_n770), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n757), .B1(G77), .B2(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n299), .B1(new_n783), .B2(G294), .ZN(new_n851));
  INV_X1    g0651(.A(G283), .ZN(new_n852));
  OAI221_X1 g0652(.A(new_n851), .B1(new_n780), .B2(new_n852), .C1(new_n481), .C2(new_n786), .ZN(new_n853));
  AOI22_X1  g0653(.A1(new_n805), .A2(G116), .B1(G311), .B2(new_n820), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n812), .A2(G87), .ZN(new_n855));
  OAI211_X1 g0655(.A(new_n854), .B(new_n855), .C1(new_n223), .C2(new_n798), .ZN(new_n856));
  AOI211_X1 g0656(.A(new_n853), .B(new_n856), .C1(G97), .C2(new_n795), .ZN(new_n857));
  XOR2_X1   g0657(.A(new_n857), .B(KEYINPUT95), .Z(new_n858));
  AOI22_X1  g0658(.A1(new_n785), .A2(G137), .B1(G143), .B2(new_n783), .ZN(new_n859));
  OAI221_X1 g0659(.A(new_n859), .B1(new_n270), .B2(new_n780), .C1(new_n804), .C2(new_n808), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n861), .A2(KEYINPUT34), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n812), .A2(G68), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n863), .B1(new_n787), .B2(new_n798), .ZN(new_n864));
  AOI211_X1 g0664(.A(new_n586), .B(new_n864), .C1(G132), .C2(new_n820), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n861), .A2(KEYINPUT34), .ZN(new_n866));
  OAI211_X1 g0666(.A(new_n865), .B(new_n866), .C1(new_n221), .C2(new_n794), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n858), .B1(new_n862), .B2(new_n867), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n850), .B1(new_n868), .B2(new_n773), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n869), .B1(new_n771), .B2(new_n841), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n847), .A2(new_n870), .ZN(G384));
  INV_X1    g0671(.A(KEYINPUT35), .ZN(new_n872));
  OAI211_X1 g0672(.A(G116), .B(new_n214), .C1(new_n531), .C2(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n873), .B1(new_n872), .B2(new_n531), .ZN(new_n874));
  XNOR2_X1  g0674(.A(new_n874), .B(KEYINPUT36), .ZN(new_n875));
  OR3_X1    g0675(.A1(new_n210), .A2(new_n202), .A3(new_n349), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n787), .A2(G68), .ZN(new_n877));
  AOI211_X1 g0677(.A(new_n259), .B(G13), .C1(new_n876), .C2(new_n877), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n875), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n743), .A2(new_n467), .A3(new_n751), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n661), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g0681(.A(new_n881), .B(KEYINPUT101), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n835), .A2(new_n694), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n837), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n368), .A2(new_n369), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n384), .A2(new_n379), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n320), .B1(new_n886), .B2(new_n358), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n373), .B1(new_n885), .B2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n348), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n392), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n888), .A2(new_n691), .ZN(new_n891));
  OAI21_X1  g0691(.A(KEYINPUT37), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(new_n691), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n893), .B1(new_n370), .B2(new_n373), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT37), .ZN(new_n895));
  NAND4_X1  g0695(.A1(new_n374), .A2(new_n894), .A3(new_n895), .A4(new_n392), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n892), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n398), .A2(new_n891), .ZN(new_n898));
  AOI21_X1  g0698(.A(KEYINPUT38), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n897), .A2(new_n898), .A3(KEYINPUT38), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n434), .A2(new_n694), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT98), .ZN(new_n905));
  OAI211_X1 g0705(.A(new_n905), .B(new_n442), .C1(new_n424), .C2(new_n434), .ZN(new_n906));
  OAI211_X1 g0706(.A(KEYINPUT98), .B(new_n442), .C1(new_n424), .C2(new_n434), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n423), .A2(new_n421), .ZN(new_n908));
  NAND4_X1  g0708(.A1(new_n908), .A2(new_n417), .A3(new_n413), .A4(new_n903), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  AOI22_X1  g0710(.A1(new_n904), .A2(new_n906), .B1(new_n907), .B2(new_n910), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n884), .A2(new_n902), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n375), .A2(new_n396), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n691), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n374), .A2(new_n894), .A3(new_n392), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(KEYINPUT37), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n896), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(KEYINPUT99), .ZN(new_n919));
  INV_X1    g0719(.A(new_n894), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n398), .A2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT99), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n917), .A2(new_n922), .A3(new_n896), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n919), .A2(new_n921), .A3(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT38), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT39), .ZN(new_n927));
  NAND4_X1  g0727(.A1(new_n926), .A2(KEYINPUT100), .A3(new_n927), .A4(new_n901), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT100), .ZN(new_n929));
  AOI22_X1  g0729(.A1(new_n918), .A2(KEYINPUT99), .B1(new_n398), .B2(new_n920), .ZN(new_n930));
  AOI21_X1  g0730(.A(KEYINPUT38), .B1(new_n930), .B2(new_n923), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n901), .A2(new_n927), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n929), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n902), .A2(KEYINPUT39), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n928), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n436), .A2(new_n693), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n915), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n882), .B(new_n937), .ZN(new_n938));
  AND2_X1   g0738(.A1(new_n911), .A2(new_n841), .ZN(new_n939));
  OAI211_X1 g0739(.A(KEYINPUT31), .B(new_n693), .C1(new_n722), .C2(new_n727), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n735), .B2(new_n737), .ZN(new_n941));
  NOR4_X1   g0741(.A1(new_n524), .A2(new_n649), .A3(new_n555), .A4(new_n693), .ZN(new_n942));
  OR2_X1    g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n939), .A2(new_n943), .A3(KEYINPUT40), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  AND3_X1   g0745(.A1(new_n897), .A2(new_n898), .A3(KEYINPUT38), .ZN(new_n946));
  NOR3_X1   g0746(.A1(new_n931), .A2(KEYINPUT102), .A3(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT102), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n948), .B1(new_n926), .B2(new_n901), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n945), .B1(new_n947), .B2(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT40), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n946), .A2(new_n899), .ZN(new_n952));
  OAI211_X1 g0752(.A(new_n911), .B(new_n841), .C1(new_n941), .C2(new_n942), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n951), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  AND2_X1   g0754(.A1(new_n950), .A2(new_n954), .ZN(new_n955));
  AND2_X1   g0755(.A1(new_n467), .A2(new_n943), .ZN(new_n956));
  OR2_X1    g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n955), .A2(new_n956), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n957), .A2(G330), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n938), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n960), .B1(new_n259), .B2(new_n754), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n938), .A2(new_n959), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n879), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(KEYINPUT103), .ZN(G367));
  NOR2_X1   g0764(.A1(new_n646), .A2(new_n694), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n668), .A2(new_n666), .A3(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n966), .B1(new_n746), .B2(new_n965), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n967), .A2(KEYINPUT43), .ZN(new_n968));
  XOR2_X1   g0768(.A(new_n968), .B(KEYINPUT104), .Z(new_n969));
  NAND2_X1  g0769(.A1(new_n967), .A2(KEYINPUT43), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n538), .A2(new_n693), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n683), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n673), .A2(new_n693), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n974), .A2(new_n700), .A3(new_n704), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(KEYINPUT42), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n554), .B1(new_n972), .B2(new_n596), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n977), .A2(new_n694), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n975), .A2(KEYINPUT42), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n970), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n969), .B(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(new_n703), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(new_n974), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n982), .B(new_n984), .ZN(new_n985));
  XOR2_X1   g0785(.A(new_n710), .B(KEYINPUT41), .Z(new_n986));
  NAND2_X1  g0786(.A1(new_n707), .A2(new_n974), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n987), .B(KEYINPUT45), .Z(new_n988));
  NOR2_X1   g0788(.A1(new_n707), .A2(new_n974), .ZN(new_n989));
  OR2_X1    g0789(.A1(KEYINPUT105), .A2(KEYINPUT44), .ZN(new_n990));
  AND2_X1   g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(KEYINPUT105), .A2(KEYINPUT44), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n992), .B1(new_n989), .B2(new_n990), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n988), .B1(new_n991), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(new_n983), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n705), .B1(new_n702), .B2(new_n704), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(new_n699), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n752), .A2(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(new_n998), .ZN(new_n999));
  OAI211_X1 g0799(.A(new_n988), .B(new_n703), .C1(new_n991), .C2(new_n993), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n995), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n986), .B1(new_n1001), .B2(new_n752), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n985), .B1(new_n1002), .B2(new_n756), .ZN(new_n1003));
  AND2_X1   g0803(.A1(new_n242), .A2(new_n766), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n774), .B1(new_n217), .B2(new_n443), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n757), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(new_n805), .A2(G50), .B1(new_n812), .B2(G77), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1007), .B1(new_n221), .B2(new_n798), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n794), .A2(new_n201), .ZN(new_n1009));
  XOR2_X1   g0809(.A(KEYINPUT107), .B(G137), .Z(new_n1010));
  OAI221_X1 g0810(.A(new_n299), .B1(new_n807), .B2(new_n1010), .C1(new_n784), .C2(new_n270), .ZN(new_n1011));
  INV_X1    g0811(.A(G143), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n1012), .A2(new_n786), .B1(new_n780), .B2(new_n808), .ZN(new_n1013));
  NOR4_X1   g0813(.A1(new_n1008), .A2(new_n1009), .A3(new_n1011), .A4(new_n1013), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n822), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT46), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1016), .B1(new_n798), .B2(new_n493), .ZN(new_n1017));
  OAI211_X1 g0817(.A(new_n1015), .B(new_n1017), .C1(new_n589), .C2(new_n780), .ZN(new_n1018));
  XOR2_X1   g0818(.A(new_n1018), .B(KEYINPUT106), .Z(new_n1019));
  NOR2_X1   g0819(.A1(new_n794), .A2(new_n223), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n804), .A2(new_n852), .B1(new_n811), .B2(new_n497), .ZN(new_n1021));
  INV_X1    g0821(.A(G317), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n586), .B1(new_n1022), .B2(new_n807), .C1(new_n784), .C2(new_n481), .ZN(new_n1023));
  INV_X1    g0823(.A(G311), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n786), .A2(new_n1024), .ZN(new_n1025));
  NOR4_X1   g0825(.A1(new_n1020), .A2(new_n1021), .A3(new_n1023), .A4(new_n1025), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1014), .B1(new_n1019), .B2(new_n1026), .ZN(new_n1027));
  XOR2_X1   g0827(.A(new_n1027), .B(KEYINPUT47), .Z(new_n1028));
  AOI21_X1  g0828(.A(new_n1006), .B1(new_n1028), .B2(new_n773), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(new_n967), .B2(new_n827), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1003), .A2(new_n1030), .ZN(G387));
  NOR2_X1   g0831(.A1(new_n702), .A2(new_n827), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n760), .A2(new_n712), .B1(new_n223), .B2(new_n709), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n238), .A2(new_n290), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n265), .A2(G50), .ZN(new_n1035));
  XOR2_X1   g0835(.A(new_n1035), .B(KEYINPUT50), .Z(new_n1036));
  NAND3_X1  g0836(.A1(new_n713), .A2(new_n290), .A3(new_n244), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n766), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1033), .B1(new_n1034), .B2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1039), .A2(new_n774), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1040), .A2(new_n757), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n784), .A2(new_n787), .B1(new_n807), .B2(new_n270), .ZN(new_n1042));
  AOI211_X1 g0842(.A(new_n586), .B(new_n1042), .C1(G159), .C2(new_n785), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(G77), .A2(new_n822), .B1(new_n812), .B2(G97), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n805), .A2(G68), .B1(new_n266), .B2(new_n779), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n794), .A2(new_n443), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n1046), .ZN(new_n1047));
  NAND4_X1  g0847(.A1(new_n1043), .A2(new_n1044), .A3(new_n1045), .A4(new_n1047), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n779), .A2(G311), .B1(G317), .B2(new_n783), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(KEYINPUT108), .B(G322), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n1049), .B1(new_n786), .B2(new_n1050), .C1(new_n481), .C2(new_n804), .ZN(new_n1051));
  INV_X1    g0851(.A(KEYINPUT48), .ZN(new_n1052));
  OR2_X1    g0852(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n795), .A2(G283), .B1(new_n822), .B2(G294), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1053), .A2(new_n1054), .A3(new_n1055), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1056), .B(KEYINPUT109), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1057), .A2(KEYINPUT49), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n807), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n556), .B1(G326), .B2(new_n1059), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n1058), .B(new_n1060), .C1(new_n493), .C2(new_n811), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n1057), .A2(KEYINPUT49), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1048), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  AOI211_X1 g0863(.A(new_n1032), .B(new_n1041), .C1(new_n1063), .C2(new_n773), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1064), .B1(new_n997), .B2(new_n756), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n710), .B(KEYINPUT110), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n998), .A2(new_n1066), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n752), .A2(new_n997), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1065), .B1(new_n1067), .B2(new_n1068), .ZN(G393));
  INV_X1    g0869(.A(KEYINPUT111), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n995), .A2(new_n1070), .A3(new_n1000), .ZN(new_n1071));
  OR3_X1    g0871(.A1(new_n994), .A2(new_n1070), .A3(new_n983), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  OAI211_X1 g0873(.A(new_n1001), .B(new_n1066), .C1(new_n1073), .C2(new_n999), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n972), .A2(new_n772), .A3(new_n973), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n767), .A2(new_n251), .ZN(new_n1076));
  AOI211_X1 g0876(.A(new_n775), .B(new_n1076), .C1(G97), .C2(new_n709), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n785), .A2(G150), .B1(G159), .B2(new_n783), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(new_n1078), .B(KEYINPUT51), .ZN(new_n1079));
  OAI221_X1 g0879(.A(new_n855), .B1(new_n201), .B2(new_n798), .C1(new_n265), .C2(new_n804), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n794), .A2(new_n202), .ZN(new_n1081));
  OAI221_X1 g0881(.A(new_n556), .B1(new_n1012), .B2(new_n807), .C1(new_n780), .C2(new_n787), .ZN(new_n1082));
  OR4_X1    g0882(.A1(new_n1079), .A2(new_n1080), .A3(new_n1081), .A4(new_n1082), .ZN(new_n1083));
  OAI221_X1 g0883(.A(new_n305), .B1(new_n807), .B2(new_n1050), .C1(new_n780), .C2(new_n481), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1084), .B1(G107), .B2(new_n812), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n805), .A2(G294), .B1(new_n822), .B2(G283), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n786), .A2(new_n1022), .B1(new_n1024), .B2(new_n784), .ZN(new_n1087));
  INV_X1    g0887(.A(KEYINPUT52), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(G116), .A2(new_n795), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  OR2_X1    g0889(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1090));
  NAND4_X1  g0890(.A1(new_n1085), .A2(new_n1086), .A3(new_n1089), .A4(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1083), .A2(new_n1091), .ZN(new_n1092));
  AOI211_X1 g0892(.A(new_n831), .B(new_n1077), .C1(new_n1092), .C2(new_n773), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n1073), .A2(new_n756), .B1(new_n1075), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1074), .A2(new_n1094), .ZN(G390));
  AOI21_X1  g0895(.A(new_n927), .B1(new_n900), .B2(new_n901), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n932), .B1(new_n925), .B2(new_n924), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1096), .B1(new_n1097), .B2(KEYINPUT100), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n884), .A2(new_n911), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n936), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1098), .A2(new_n1101), .A3(new_n933), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(new_n936), .B(KEYINPUT112), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n750), .A2(new_n694), .A3(new_n836), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(new_n883), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1103), .B1(new_n1105), .B2(new_n911), .ZN(new_n1106));
  OAI21_X1  g0906(.A(KEYINPUT102), .B1(new_n931), .B2(new_n946), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n923), .ZN(new_n1108));
  AND2_X1   g0908(.A1(new_n398), .A2(new_n920), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n922), .B1(new_n917), .B2(new_n896), .ZN(new_n1110));
  NOR3_X1   g0910(.A1(new_n1108), .A2(new_n1109), .A3(new_n1110), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n948), .B(new_n901), .C1(new_n1111), .C2(KEYINPUT38), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1107), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1106), .A2(new_n1113), .ZN(new_n1114));
  NAND4_X1  g0914(.A1(new_n739), .A2(G330), .A3(new_n841), .A4(new_n911), .ZN(new_n1115));
  AND3_X1   g0915(.A1(new_n1102), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1116));
  AND2_X1   g0916(.A1(new_n943), .A2(G330), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1117), .A2(new_n939), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1118), .B1(new_n1102), .B2(new_n1114), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1116), .A2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n739), .A2(G330), .A3(new_n841), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n911), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(new_n1117), .A2(new_n939), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n884), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n943), .A2(G330), .A3(new_n841), .ZN(new_n1125));
  AND2_X1   g0925(.A1(new_n1125), .A2(new_n1122), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1115), .A2(new_n883), .A3(new_n1104), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n1123), .A2(new_n1124), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1117), .A2(new_n467), .ZN(new_n1129));
  AND3_X1   g0929(.A1(new_n661), .A2(new_n1129), .A3(new_n880), .ZN(new_n1130));
  AOI21_X1  g0930(.A(KEYINPUT113), .B1(new_n1128), .B2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1120), .A2(new_n1131), .ZN(new_n1132));
  AND2_X1   g0932(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1133));
  OAI22_X1  g0933(.A1(new_n1133), .A2(KEYINPUT113), .B1(new_n1116), .B2(new_n1119), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1135), .A2(new_n1066), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1102), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1137));
  AND3_X1   g0937(.A1(new_n928), .A2(new_n933), .A3(new_n934), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n1138), .A2(new_n1101), .B1(new_n1113), .B2(new_n1106), .ZN(new_n1139));
  OAI211_X1 g0939(.A(new_n1137), .B(new_n756), .C1(new_n1139), .C2(new_n1118), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1138), .A2(new_n770), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n757), .B1(new_n266), .B2(new_n849), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n299), .B1(new_n783), .B2(G116), .ZN(new_n1143));
  OAI221_X1 g0943(.A(new_n1143), .B1(new_n780), .B2(new_n223), .C1(new_n852), .C2(new_n786), .ZN(new_n1144));
  AOI211_X1 g0944(.A(new_n799), .B(new_n1144), .C1(G97), .C2(new_n805), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1145), .B1(new_n202), .B2(new_n794), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n820), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n863), .B1(new_n589), .B2(new_n1147), .ZN(new_n1148));
  XOR2_X1   g0948(.A(new_n1148), .B(KEYINPUT116), .Z(new_n1149));
  XNOR2_X1  g0949(.A(KEYINPUT54), .B(G143), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n804), .A2(new_n1150), .B1(new_n780), .B2(new_n1010), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(G159), .B2(new_n795), .ZN(new_n1152));
  XOR2_X1   g0952(.A(new_n1152), .B(KEYINPUT114), .Z(new_n1153));
  NAND2_X1  g0953(.A1(new_n822), .A2(G150), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(new_n1154), .B(KEYINPUT53), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(new_n785), .A2(G128), .B1(G132), .B2(new_n783), .ZN(new_n1156));
  XOR2_X1   g0956(.A(new_n1156), .B(KEYINPUT115), .Z(new_n1157));
  INV_X1    g0957(.A(G125), .ZN(new_n1158));
  OAI221_X1 g0958(.A(new_n299), .B1(new_n787), .B2(new_n811), .C1(new_n1147), .C2(new_n1158), .ZN(new_n1159));
  OR3_X1    g0959(.A1(new_n1155), .A2(new_n1157), .A3(new_n1159), .ZN(new_n1160));
  OAI22_X1  g0960(.A1(new_n1146), .A2(new_n1149), .B1(new_n1153), .B2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1142), .B1(new_n1161), .B2(new_n773), .ZN(new_n1162));
  AND3_X1   g0962(.A1(new_n1141), .A2(KEYINPUT117), .A3(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(KEYINPUT117), .B1(new_n1141), .B2(new_n1162), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1140), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1136), .A2(new_n1166), .ZN(G378));
  NAND2_X1  g0967(.A1(new_n658), .A2(new_n659), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n279), .A2(new_n691), .ZN(new_n1169));
  INV_X1    g0969(.A(KEYINPUT118), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(new_n1169), .B(new_n1170), .ZN(new_n1171));
  AND3_X1   g0971(.A1(new_n1168), .A2(new_n311), .A3(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1171), .B1(new_n1168), .B2(new_n311), .ZN(new_n1173));
  XOR2_X1   g0973(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  NOR3_X1   g0975(.A1(new_n1172), .A2(new_n1173), .A3(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1171), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n331), .A2(new_n1177), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1168), .A2(new_n1171), .A3(new_n311), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1174), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n1176), .A2(new_n1180), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n1181), .A2(new_n771), .ZN(new_n1182));
  INV_X1    g0982(.A(G128), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n786), .A2(new_n1158), .B1(new_n1183), .B2(new_n784), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1184), .B1(G132), .B2(new_n779), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1150), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(new_n805), .A2(G137), .B1(new_n822), .B2(new_n1186), .ZN(new_n1187));
  OAI211_X1 g0987(.A(new_n1185), .B(new_n1187), .C1(new_n270), .C2(new_n794), .ZN(new_n1188));
  OR2_X1    g0988(.A1(new_n1188), .A2(KEYINPUT59), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1188), .A2(KEYINPUT59), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n267), .A2(new_n284), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n811), .A2(new_n808), .ZN(new_n1192));
  AOI211_X1 g0992(.A(new_n1191), .B(new_n1192), .C1(G124), .C2(new_n1059), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1189), .A2(new_n1190), .A3(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n812), .A2(G58), .ZN(new_n1195));
  OAI221_X1 g0995(.A(new_n1195), .B1(new_n443), .B2(new_n804), .C1(new_n852), .C2(new_n1147), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(new_n779), .A2(G97), .B1(G107), .B2(new_n783), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1197), .B1(new_n493), .B2(new_n786), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n475), .B(new_n586), .C1(new_n798), .C2(new_n202), .ZN(new_n1199));
  NOR4_X1   g0999(.A1(new_n1196), .A2(new_n1009), .A3(new_n1198), .A4(new_n1199), .ZN(new_n1200));
  OR2_X1    g1000(.A1(new_n1200), .A2(KEYINPUT58), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1200), .A2(KEYINPUT58), .ZN(new_n1202));
  OAI211_X1 g1002(.A(new_n787), .B(new_n1191), .C1(new_n556), .C2(new_n288), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1194), .A2(new_n1201), .A3(new_n1202), .A4(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1204), .A2(new_n773), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n1205), .B(new_n757), .C1(G50), .C2(new_n849), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n1182), .A2(new_n1206), .ZN(new_n1207));
  AND2_X1   g1007(.A1(new_n954), .A2(G330), .ZN(new_n1208));
  OR2_X1    g1008(.A1(new_n1176), .A2(new_n1180), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n950), .A2(new_n1208), .A3(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n944), .B1(new_n1107), .B2(new_n1112), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n954), .A2(G330), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1181), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  AND3_X1   g1013(.A1(new_n1210), .A2(new_n937), .A3(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n937), .B1(new_n1210), .B2(new_n1213), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1207), .B1(new_n1216), .B2(new_n756), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n1137), .B(new_n1128), .C1(new_n1139), .C2(new_n1118), .ZN(new_n1218));
  AND2_X1   g1018(.A1(new_n1218), .A2(new_n1130), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n915), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1220), .B1(new_n1138), .B2(new_n1100), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1209), .B1(new_n950), .B2(new_n1208), .ZN(new_n1222));
  NOR3_X1   g1022(.A1(new_n1211), .A2(new_n1212), .A3(new_n1181), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1221), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1210), .A2(new_n937), .A3(new_n1213), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1224), .A2(KEYINPUT57), .A3(new_n1225), .ZN(new_n1226));
  OAI21_X1  g1026(.A(KEYINPUT119), .B1(new_n1219), .B2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1218), .A2(new_n1130), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT119), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n1228), .A2(new_n1216), .A3(new_n1229), .A4(KEYINPUT57), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1227), .A2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1232), .B1(new_n1130), .B2(new_n1218), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1066), .B1(new_n1233), .B2(KEYINPUT57), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1217), .B1(new_n1231), .B2(new_n1234), .ZN(G375));
  INV_X1    g1035(.A(new_n1133), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n986), .ZN(new_n1237));
  OR2_X1    g1037(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1236), .A2(new_n1237), .A3(new_n1238), .ZN(new_n1239));
  OAI22_X1  g1039(.A1(new_n780), .A2(new_n1150), .B1(new_n784), .B2(new_n1010), .ZN(new_n1240));
  OAI22_X1  g1040(.A1(new_n1147), .A2(new_n1183), .B1(new_n804), .B2(new_n270), .ZN(new_n1241));
  OAI211_X1 g1041(.A(new_n1195), .B(new_n556), .C1(new_n787), .C2(new_n794), .ZN(new_n1242));
  AOI211_X1 g1042(.A(new_n1241), .B(new_n1242), .C1(G159), .C2(new_n822), .ZN(new_n1243));
  XOR2_X1   g1043(.A(new_n1243), .B(KEYINPUT120), .Z(new_n1244));
  AOI211_X1 g1044(.A(new_n1240), .B(new_n1244), .C1(G132), .C2(new_n785), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n299), .B1(new_n783), .B2(G283), .ZN(new_n1246));
  OAI221_X1 g1046(.A(new_n1246), .B1(new_n780), .B2(new_n493), .C1(new_n589), .C2(new_n786), .ZN(new_n1247));
  OAI22_X1  g1047(.A1(new_n1147), .A2(new_n481), .B1(new_n497), .B2(new_n798), .ZN(new_n1248));
  OAI22_X1  g1048(.A1(new_n804), .A2(new_n223), .B1(new_n811), .B2(new_n202), .ZN(new_n1249));
  NOR4_X1   g1049(.A1(new_n1247), .A2(new_n1248), .A3(new_n1046), .A4(new_n1249), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n773), .B1(new_n1245), .B2(new_n1250), .ZN(new_n1251));
  OAI211_X1 g1051(.A(new_n1251), .B(new_n757), .C1(G68), .C2(new_n849), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1252), .B1(new_n770), .B2(new_n1122), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1253), .B1(new_n1128), .B2(new_n756), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1239), .A2(new_n1254), .ZN(G381));
  INV_X1    g1055(.A(G390), .ZN(new_n1256));
  NOR3_X1   g1056(.A1(G384), .A2(G396), .A3(G393), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1256), .A2(new_n1254), .A3(new_n1239), .A4(new_n1257), .ZN(new_n1258));
  OR4_X1    g1058(.A1(G387), .A2(G375), .A3(new_n1258), .A4(G378), .ZN(G407));
  AOI21_X1  g1059(.A(new_n1165), .B1(new_n1135), .B2(new_n1066), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1260), .A2(G213), .A3(new_n692), .ZN(new_n1261));
  OAI211_X1 g1061(.A(G407), .B(G213), .C1(G375), .C2(new_n1261), .ZN(G409));
  OAI211_X1 g1062(.A(G378), .B(new_n1217), .C1(new_n1231), .C2(new_n1234), .ZN(new_n1263));
  OAI21_X1  g1063(.A(KEYINPUT121), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT121), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1224), .A2(new_n1265), .A3(new_n1225), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1264), .A2(new_n756), .A3(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1228), .A2(new_n1216), .A3(new_n1237), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1207), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1267), .A2(new_n1268), .A3(new_n1269), .ZN(new_n1270));
  AND3_X1   g1070(.A1(new_n1270), .A2(new_n1260), .A3(KEYINPUT122), .ZN(new_n1271));
  AOI21_X1  g1071(.A(KEYINPUT122), .B1(new_n1270), .B2(new_n1260), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1263), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT123), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n692), .A2(G213), .ZN(new_n1276));
  OAI211_X1 g1076(.A(new_n1263), .B(KEYINPUT123), .C1(new_n1271), .C2(new_n1272), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1275), .A2(new_n1276), .A3(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT60), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1238), .A2(new_n1279), .ZN(new_n1280));
  OR3_X1    g1080(.A1(new_n1128), .A2(new_n1130), .A3(new_n1279), .ZN(new_n1281));
  NAND4_X1  g1081(.A1(new_n1280), .A2(new_n1066), .A3(new_n1236), .A4(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(new_n1254), .ZN(new_n1283));
  INV_X1    g1083(.A(G384), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1284), .A2(KEYINPUT124), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT124), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(G384), .A2(new_n1286), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1283), .A2(new_n1285), .A3(new_n1287), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1282), .A2(new_n1284), .A3(KEYINPUT124), .A4(new_n1254), .ZN(new_n1289));
  AND3_X1   g1089(.A1(new_n1288), .A2(KEYINPUT125), .A3(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(KEYINPUT125), .B1(new_n1288), .B2(new_n1289), .ZN(new_n1291));
  INV_X1    g1091(.A(G2897), .ZN(new_n1292));
  OAI22_X1  g1092(.A1(new_n1290), .A2(new_n1291), .B1(new_n1292), .B2(new_n1276), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1294));
  OR3_X1    g1094(.A1(new_n1294), .A2(new_n1292), .A3(new_n1276), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1278), .A2(new_n1293), .A3(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1291), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1288), .A2(KEYINPUT125), .A3(new_n1289), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  NAND4_X1  g1099(.A1(new_n1275), .A2(new_n1276), .A3(new_n1299), .A4(new_n1277), .ZN(new_n1300));
  XOR2_X1   g1100(.A(KEYINPUT126), .B(KEYINPUT63), .Z(new_n1301));
  NAND2_X1  g1101(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1302));
  NOR2_X1   g1102(.A1(new_n1256), .A2(G387), .ZN(new_n1303));
  AOI21_X1  g1103(.A(G390), .B1(new_n1003), .B2(new_n1030), .ZN(new_n1304));
  OAI21_X1  g1104(.A(KEYINPUT127), .B1(new_n1303), .B2(new_n1304), .ZN(new_n1305));
  XNOR2_X1  g1105(.A(G393), .B(new_n829), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT61), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1306), .ZN(new_n1309));
  OAI211_X1 g1109(.A(KEYINPUT127), .B(new_n1309), .C1(new_n1303), .C2(new_n1304), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1307), .A2(new_n1308), .A3(new_n1310), .ZN(new_n1311));
  AND2_X1   g1111(.A1(new_n1299), .A2(KEYINPUT63), .ZN(new_n1312));
  AND2_X1   g1112(.A1(new_n1273), .A2(new_n1276), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1311), .B1(new_n1312), .B2(new_n1313), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1296), .A2(new_n1302), .A3(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1293), .A2(new_n1295), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1308), .B1(new_n1313), .B2(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT62), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1300), .A2(new_n1318), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1313), .A2(KEYINPUT62), .A3(new_n1299), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1317), .B1(new_n1319), .B2(new_n1320), .ZN(new_n1321));
  AND2_X1   g1121(.A1(new_n1307), .A2(new_n1310), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1315), .B1(new_n1321), .B2(new_n1322), .ZN(G405));
  XNOR2_X1  g1123(.A(G375), .B(G378), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1324), .A2(new_n1294), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1325), .B1(new_n1299), .B2(new_n1324), .ZN(new_n1326));
  XNOR2_X1  g1126(.A(new_n1326), .B(new_n1322), .ZN(G402));
endmodule


