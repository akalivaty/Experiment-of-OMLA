//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 0 0 1 0 0 0 0 1 0 0 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 0 0 1 0 1 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 0 1 0 1 1 0 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:38 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n772, new_n773, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n796, new_n797, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1061, new_n1062, new_n1063, new_n1064, new_n1065, new_n1066,
    new_n1067, new_n1068, new_n1069, new_n1070, new_n1071, new_n1072,
    new_n1073, new_n1074, new_n1075, new_n1076, new_n1077, new_n1078,
    new_n1079, new_n1080, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1106, new_n1107, new_n1108, new_n1109,
    new_n1110, new_n1111, new_n1112, new_n1113, new_n1114, new_n1115;
  XNOR2_X1  g000(.A(KEYINPUT66), .B(G146), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  XNOR2_X1  g002(.A(KEYINPUT65), .B(G143), .ZN(new_n189));
  AOI22_X1  g003(.A1(new_n188), .A2(G143), .B1(new_n189), .B2(G146), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT1), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(KEYINPUT70), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT70), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(KEYINPUT1), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G128), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G107), .ZN(new_n198));
  OAI21_X1  g012(.A(KEYINPUT78), .B1(new_n198), .B2(G104), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT78), .ZN(new_n200));
  INV_X1    g014(.A(G104), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n200), .A2(new_n201), .A3(G107), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n198), .A2(G104), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n199), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G101), .ZN(new_n205));
  INV_X1    g019(.A(G101), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n201), .A2(G107), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n198), .A2(KEYINPUT3), .A3(G104), .ZN(new_n208));
  INV_X1    g022(.A(new_n208), .ZN(new_n209));
  AOI21_X1  g023(.A(KEYINPUT3), .B1(new_n198), .B2(G104), .ZN(new_n210));
  OAI211_X1 g024(.A(new_n206), .B(new_n207), .C1(new_n209), .C2(new_n210), .ZN(new_n211));
  AOI22_X1  g025(.A1(new_n190), .A2(new_n197), .B1(new_n205), .B2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G146), .ZN(new_n213));
  INV_X1    g027(.A(G143), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(KEYINPUT65), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT65), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G143), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g032(.A1(new_n213), .A2(new_n218), .B1(new_n187), .B2(new_n214), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT66), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(new_n213), .ZN(new_n221));
  NAND2_X1  g035(.A1(KEYINPUT66), .A2(G146), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n221), .A2(G143), .A3(new_n222), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n196), .B1(new_n223), .B2(new_n195), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT71), .ZN(new_n225));
  NOR3_X1   g039(.A1(new_n219), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  AND2_X1   g040(.A1(KEYINPUT66), .A2(G146), .ZN(new_n227));
  NOR2_X1   g041(.A1(KEYINPUT66), .A2(G146), .ZN(new_n228));
  NOR3_X1   g042(.A1(new_n227), .A2(new_n228), .A3(new_n214), .ZN(new_n229));
  XNOR2_X1  g043(.A(KEYINPUT70), .B(KEYINPUT1), .ZN(new_n230));
  OAI21_X1  g044(.A(G128), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n214), .B1(new_n227), .B2(new_n228), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n232), .B1(new_n189), .B2(G146), .ZN(new_n233));
  AOI21_X1  g047(.A(KEYINPUT71), .B1(new_n231), .B2(new_n233), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n212), .B1(new_n226), .B2(new_n234), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n223), .B1(new_n218), .B2(new_n213), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n191), .B1(new_n218), .B2(new_n213), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n236), .B1(new_n237), .B2(new_n196), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n189), .A2(G146), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n197), .A2(new_n223), .A3(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  AND2_X1   g055(.A1(new_n205), .A2(new_n211), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n235), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(G137), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n245), .A2(KEYINPUT11), .A3(G134), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT11), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(G137), .ZN(new_n248));
  AND2_X1   g062(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(G134), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(KEYINPUT67), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT67), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G134), .ZN(new_n253));
  OAI211_X1 g067(.A(new_n251), .B(new_n253), .C1(new_n247), .C2(G137), .ZN(new_n254));
  NAND2_X1  g068(.A1(KEYINPUT68), .A2(G131), .ZN(new_n255));
  AND3_X1   g069(.A1(new_n249), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n255), .B1(new_n249), .B2(new_n254), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  AOI21_X1  g073(.A(KEYINPUT12), .B1(new_n244), .B2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT12), .ZN(new_n261));
  AOI211_X1 g075(.A(new_n261), .B(new_n258), .C1(new_n235), .C2(new_n243), .ZN(new_n262));
  OAI21_X1  g076(.A(KEYINPUT80), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n225), .B1(new_n219), .B2(new_n224), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n231), .A2(KEYINPUT71), .A3(new_n233), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  AOI22_X1  g080(.A1(new_n266), .A2(new_n212), .B1(new_n241), .B2(new_n242), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n261), .B1(new_n267), .B2(new_n258), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n244), .A2(KEYINPUT12), .A3(new_n259), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT80), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n268), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  XNOR2_X1  g085(.A(G110), .B(G140), .ZN(new_n272));
  INV_X1    g086(.A(G953), .ZN(new_n273));
  AND2_X1   g087(.A1(new_n273), .A2(G227), .ZN(new_n274));
  XNOR2_X1  g088(.A(new_n272), .B(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n205), .A2(new_n211), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n276), .B1(new_n238), .B2(new_n240), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n207), .B1(new_n209), .B2(new_n210), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT4), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n278), .A2(new_n279), .A3(G101), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n211), .A2(KEYINPUT4), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT3), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n282), .B1(new_n201), .B2(G107), .ZN(new_n283));
  AOI22_X1  g097(.A1(new_n283), .A2(new_n208), .B1(new_n201), .B2(G107), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n284), .A2(new_n206), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n280), .B1(new_n281), .B2(new_n285), .ZN(new_n286));
  OR3_X1    g100(.A1(KEYINPUT64), .A2(KEYINPUT0), .A3(G128), .ZN(new_n287));
  OAI21_X1  g101(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n288));
  AOI22_X1  g102(.A1(new_n287), .A2(new_n288), .B1(KEYINPUT0), .B2(G128), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n233), .A2(new_n289), .ZN(new_n290));
  NAND4_X1  g104(.A1(new_n239), .A2(KEYINPUT0), .A3(G128), .A4(new_n223), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  OAI22_X1  g106(.A1(new_n277), .A2(KEYINPUT10), .B1(new_n286), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n242), .A2(KEYINPUT10), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n294), .B1(new_n266), .B2(new_n240), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n275), .B1(new_n296), .B2(new_n258), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n263), .A2(new_n271), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(KEYINPUT81), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT81), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n263), .A2(new_n300), .A3(new_n271), .A4(new_n297), .ZN(new_n301));
  INV_X1    g115(.A(new_n293), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n240), .B1(new_n226), .B2(new_n234), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n303), .A2(KEYINPUT10), .A3(new_n242), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n302), .A2(new_n304), .A3(new_n258), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n259), .B1(new_n293), .B2(new_n295), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(new_n275), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n299), .A2(new_n301), .A3(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(G469), .ZN(new_n310));
  INV_X1    g124(.A(G902), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n309), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT79), .ZN(new_n313));
  INV_X1    g127(.A(new_n275), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n268), .A2(new_n269), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n314), .B1(new_n315), .B2(new_n305), .ZN(new_n316));
  AND3_X1   g130(.A1(new_n305), .A2(new_n314), .A3(new_n306), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n311), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n313), .B1(new_n318), .B2(G469), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n318), .A2(new_n313), .A3(G469), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n312), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  XNOR2_X1  g136(.A(KEYINPUT9), .B(G234), .ZN(new_n323));
  OAI21_X1  g137(.A(G221), .B1(new_n323), .B2(G902), .ZN(new_n324));
  XOR2_X1   g138(.A(new_n324), .B(KEYINPUT77), .Z(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n322), .A2(new_n326), .ZN(new_n327));
  OAI21_X1  g141(.A(G210), .B1(G237), .B2(G902), .ZN(new_n328));
  XNOR2_X1  g142(.A(new_n328), .B(KEYINPUT85), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT84), .ZN(new_n330));
  XOR2_X1   g144(.A(G110), .B(G122), .Z(new_n331));
  XNOR2_X1  g145(.A(KEYINPUT83), .B(KEYINPUT8), .ZN(new_n332));
  XNOR2_X1  g146(.A(new_n331), .B(new_n332), .ZN(new_n333));
  OR2_X1    g147(.A1(KEYINPUT72), .A2(G116), .ZN(new_n334));
  NAND2_X1  g148(.A1(KEYINPUT72), .A2(G116), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n334), .A2(G119), .A3(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(G116), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n337), .A2(G119), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n336), .A2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  XOR2_X1   g155(.A(KEYINPUT2), .B(G113), .Z(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT5), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n338), .A2(new_n344), .ZN(new_n345));
  OAI211_X1 g159(.A(G113), .B(new_n345), .C1(new_n340), .C2(new_n344), .ZN(new_n346));
  AND3_X1   g160(.A1(new_n242), .A2(new_n343), .A3(new_n346), .ZN(new_n347));
  AOI22_X1  g161(.A1(new_n343), .A2(new_n346), .B1(new_n211), .B2(new_n205), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n333), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n242), .A2(new_n346), .A3(new_n343), .ZN(new_n350));
  INV_X1    g164(.A(new_n331), .ZN(new_n351));
  XNOR2_X1  g165(.A(new_n340), .B(new_n342), .ZN(new_n352));
  OAI211_X1 g166(.A(new_n350), .B(new_n351), .C1(new_n352), .C2(new_n286), .ZN(new_n353));
  INV_X1    g167(.A(G125), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n354), .B1(new_n290), .B2(new_n291), .ZN(new_n355));
  AND3_X1   g169(.A1(new_n197), .A2(new_n223), .A3(new_n239), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n356), .B1(new_n264), .B2(new_n265), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n355), .B1(new_n357), .B2(new_n354), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n273), .A2(G224), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(KEYINPUT7), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  OAI211_X1 g175(.A(new_n349), .B(new_n353), .C1(new_n358), .C2(new_n361), .ZN(new_n362));
  AOI211_X1 g176(.A(G125), .B(new_n356), .C1(new_n264), .C2(new_n265), .ZN(new_n363));
  NOR3_X1   g177(.A1(new_n363), .A2(new_n355), .A3(new_n360), .ZN(new_n364));
  OAI211_X1 g178(.A(new_n330), .B(new_n311), .C1(new_n362), .C2(new_n364), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n350), .B1(new_n352), .B2(new_n286), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(new_n331), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n367), .A2(KEYINPUT6), .A3(new_n353), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT6), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n366), .A2(new_n369), .A3(new_n331), .ZN(new_n370));
  XOR2_X1   g184(.A(new_n359), .B(KEYINPUT82), .Z(new_n371));
  AND2_X1   g185(.A1(new_n358), .A2(new_n371), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n358), .A2(new_n371), .ZN(new_n373));
  OAI211_X1 g187(.A(new_n368), .B(new_n370), .C1(new_n372), .C2(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n365), .A2(new_n374), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n360), .B1(new_n363), .B2(new_n355), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n358), .A2(new_n361), .ZN(new_n377));
  NAND4_X1  g191(.A1(new_n376), .A2(new_n377), .A3(new_n353), .A4(new_n349), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n330), .B1(new_n378), .B2(new_n311), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n329), .B1(new_n375), .B2(new_n379), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n311), .B1(new_n362), .B2(new_n364), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(KEYINPUT84), .ZN(new_n382));
  INV_X1    g196(.A(new_n329), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n382), .A2(new_n383), .A3(new_n374), .A4(new_n365), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n380), .A2(KEYINPUT86), .A3(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(new_n375), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT86), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n386), .A2(new_n387), .A3(new_n383), .A4(new_n382), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n385), .A2(new_n388), .ZN(new_n389));
  OAI21_X1  g203(.A(G214), .B1(G237), .B2(G902), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  OAI21_X1  g205(.A(KEYINPUT87), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT87), .ZN(new_n393));
  NAND4_X1  g207(.A1(new_n385), .A2(new_n393), .A3(new_n390), .A4(new_n388), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n327), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(G472), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT73), .ZN(new_n397));
  OAI211_X1 g211(.A(new_n290), .B(new_n291), .C1(new_n256), .C2(new_n257), .ZN(new_n398));
  AOI21_X1  g212(.A(G137), .B1(new_n251), .B2(new_n253), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n245), .A2(G134), .ZN(new_n400));
  OAI21_X1  g214(.A(G131), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(G131), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n249), .A2(new_n254), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  OAI211_X1 g218(.A(new_n352), .B(new_n398), .C1(new_n357), .C2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT30), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n404), .A2(KEYINPUT69), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT69), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n401), .A2(new_n403), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  OAI211_X1 g225(.A(new_n407), .B(new_n398), .C1(new_n411), .C2(new_n357), .ZN(new_n412));
  INV_X1    g226(.A(new_n398), .ZN(new_n413));
  INV_X1    g227(.A(new_n404), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n413), .B1(new_n303), .B2(new_n414), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n412), .B1(new_n415), .B2(new_n407), .ZN(new_n416));
  INV_X1    g230(.A(new_n352), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n406), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(G237), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n419), .A2(new_n273), .A3(G210), .ZN(new_n420));
  XOR2_X1   g234(.A(new_n420), .B(KEYINPUT27), .Z(new_n421));
  XNOR2_X1  g235(.A(KEYINPUT26), .B(G101), .ZN(new_n422));
  XNOR2_X1  g236(.A(new_n421), .B(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n397), .B1(new_n418), .B2(new_n424), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n404), .B1(new_n266), .B2(new_n240), .ZN(new_n426));
  OAI21_X1  g240(.A(KEYINPUT30), .B1(new_n426), .B2(new_n413), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n352), .B1(new_n427), .B2(new_n412), .ZN(new_n428));
  NOR4_X1   g242(.A1(new_n428), .A2(KEYINPUT73), .A3(new_n406), .A4(new_n423), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT31), .ZN(new_n430));
  NOR3_X1   g244(.A1(new_n425), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n418), .A2(new_n430), .A3(new_n424), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n406), .A2(KEYINPUT28), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT28), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n405), .A2(new_n434), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n398), .B1(new_n411), .B2(new_n357), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(new_n417), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n433), .A2(new_n435), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(new_n423), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n432), .A2(new_n439), .ZN(new_n440));
  OAI211_X1 g254(.A(new_n396), .B(new_n311), .C1(new_n431), .C2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT32), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND4_X1  g257(.A1(new_n433), .A2(new_n424), .A3(new_n435), .A4(new_n437), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT29), .ZN(new_n445));
  OAI211_X1 g259(.A(new_n444), .B(new_n445), .C1(new_n418), .C2(new_n424), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n417), .B1(new_n426), .B2(new_n413), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n434), .B1(new_n447), .B2(new_n405), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT74), .ZN(new_n449));
  AOI22_X1  g263(.A1(new_n448), .A2(new_n449), .B1(new_n434), .B2(new_n405), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n447), .A2(new_n405), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(KEYINPUT28), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(KEYINPUT74), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n450), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n424), .A2(KEYINPUT29), .ZN(new_n455));
  OAI211_X1 g269(.A(new_n446), .B(new_n311), .C1(new_n454), .C2(new_n455), .ZN(new_n456));
  AND2_X1   g270(.A1(new_n456), .A2(G472), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n416), .A2(new_n417), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n459), .A2(new_n405), .A3(new_n424), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(KEYINPUT73), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n418), .A2(new_n397), .A3(new_n424), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n461), .A2(KEYINPUT31), .A3(new_n462), .ZN(new_n463));
  AND2_X1   g277(.A1(new_n432), .A2(new_n439), .ZN(new_n464));
  AOI21_X1  g278(.A(G902), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n465), .A2(KEYINPUT32), .A3(new_n396), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n443), .A2(new_n458), .A3(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(G217), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n468), .B1(G234), .B2(new_n311), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(G119), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n471), .A2(G128), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n471), .A2(G128), .ZN(new_n474));
  AND2_X1   g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  XNOR2_X1  g289(.A(KEYINPUT24), .B(G110), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n196), .A2(KEYINPUT23), .A3(G119), .ZN(new_n478));
  OAI211_X1 g292(.A(new_n478), .B(new_n474), .C1(new_n472), .C2(KEYINPUT23), .ZN(new_n479));
  OAI22_X1  g293(.A1(new_n475), .A2(new_n477), .B1(G110), .B2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(G140), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(G125), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n354), .A2(G140), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n482), .A2(new_n483), .A3(KEYINPUT16), .ZN(new_n484));
  NOR3_X1   g298(.A1(new_n354), .A2(KEYINPUT16), .A3(G140), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n484), .A2(G146), .A3(new_n486), .ZN(new_n487));
  XNOR2_X1  g301(.A(G125), .B(G140), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n188), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n480), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n486), .A2(new_n484), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(new_n213), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(new_n487), .ZN(new_n493));
  INV_X1    g307(.A(new_n475), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n493), .B1(new_n494), .B2(new_n476), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n479), .A2(G110), .ZN(new_n496));
  XNOR2_X1  g310(.A(new_n496), .B(KEYINPUT75), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n490), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  XNOR2_X1  g312(.A(KEYINPUT22), .B(G137), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n273), .A2(G221), .A3(G234), .ZN(new_n500));
  XNOR2_X1  g314(.A(new_n499), .B(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  OR2_X1    g316(.A1(new_n498), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n498), .A2(new_n502), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  NOR2_X1   g320(.A1(KEYINPUT76), .A2(KEYINPUT25), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n506), .A2(new_n311), .A3(new_n508), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n507), .B1(new_n505), .B2(G902), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n470), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NOR3_X1   g325(.A1(new_n505), .A2(G902), .A3(new_n469), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n489), .B1(new_n213), .B2(new_n488), .ZN(new_n514));
  NAND4_X1  g328(.A1(new_n419), .A2(new_n273), .A3(G143), .A4(G214), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT18), .ZN(new_n516));
  AND3_X1   g330(.A1(new_n419), .A2(new_n273), .A3(G214), .ZN(new_n517));
  OAI221_X1 g331(.A(new_n515), .B1(new_n516), .B2(new_n402), .C1(new_n218), .C2(new_n517), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n515), .B1(new_n218), .B2(new_n517), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(G131), .ZN(new_n520));
  OAI211_X1 g334(.A(new_n514), .B(new_n518), .C1(new_n516), .C2(new_n520), .ZN(new_n521));
  XNOR2_X1  g335(.A(G113), .B(G122), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n522), .B(new_n201), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT17), .ZN(new_n524));
  OAI211_X1 g338(.A(new_n402), .B(new_n515), .C1(new_n218), .C2(new_n517), .ZN(new_n525));
  AND3_X1   g339(.A1(new_n520), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  OAI211_X1 g340(.A(new_n492), .B(new_n487), .C1(new_n520), .C2(new_n524), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n521), .B(new_n523), .C1(new_n526), .C2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT88), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n482), .A2(new_n483), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT19), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n488), .A2(KEYINPUT19), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n187), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  AND3_X1   g348(.A1(new_n486), .A2(new_n484), .A3(G146), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n529), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n520), .A2(new_n525), .ZN(new_n537));
  AND3_X1   g351(.A1(new_n482), .A2(new_n483), .A3(KEYINPUT19), .ZN(new_n538));
  AOI21_X1  g352(.A(KEYINPUT19), .B1(new_n482), .B2(new_n483), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n188), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n540), .A2(KEYINPUT88), .A3(new_n487), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n536), .A2(new_n537), .A3(new_n541), .ZN(new_n542));
  AND2_X1   g356(.A1(new_n542), .A2(new_n521), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n528), .B1(new_n543), .B2(new_n523), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT89), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT20), .ZN(new_n546));
  NOR2_X1   g360(.A1(G475), .A2(G902), .ZN(new_n547));
  NAND4_X1  g361(.A1(new_n544), .A2(new_n545), .A3(new_n546), .A4(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(new_n528), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n523), .B1(new_n542), .B2(new_n521), .ZN(new_n550));
  OAI211_X1 g364(.A(new_n546), .B(new_n547), .C1(new_n549), .C2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(KEYINPUT89), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n547), .B1(new_n549), .B2(new_n550), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(KEYINPUT20), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n548), .A2(new_n552), .A3(new_n554), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n521), .B1(new_n526), .B2(new_n527), .ZN(new_n556));
  INV_X1    g370(.A(new_n523), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  AND2_X1   g372(.A1(new_n558), .A2(new_n528), .ZN(new_n559));
  OAI21_X1  g373(.A(G475), .B1(new_n559), .B2(G902), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n555), .A2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(G234), .A2(G237), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n563), .A2(G952), .A3(new_n273), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n563), .A2(G902), .A3(G953), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  XNOR2_X1  g381(.A(KEYINPUT21), .B(G898), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n565), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n562), .A2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(G478), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n572), .A2(KEYINPUT15), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n214), .A2(G128), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n574), .B1(new_n189), .B2(G128), .ZN(new_n575));
  AND2_X1   g389(.A1(new_n251), .A2(new_n253), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n575), .B(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n334), .A2(G122), .A3(new_n335), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT90), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n337), .A2(G122), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n578), .A2(new_n579), .A3(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n579), .B1(new_n578), .B2(new_n581), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n198), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  AND2_X1   g399(.A1(KEYINPUT72), .A2(G116), .ZN(new_n586));
  NOR2_X1   g400(.A1(KEYINPUT72), .A2(G116), .ZN(new_n587));
  INV_X1    g401(.A(G122), .ZN(new_n588));
  NOR3_X1   g402(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n198), .B1(new_n589), .B2(KEYINPUT14), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT14), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n578), .A2(new_n591), .A3(new_n581), .ZN(new_n592));
  AND3_X1   g406(.A1(new_n590), .A2(KEYINPUT91), .A3(new_n592), .ZN(new_n593));
  AOI21_X1  g407(.A(KEYINPUT91), .B1(new_n590), .B2(new_n592), .ZN(new_n594));
  OAI211_X1 g408(.A(new_n577), .B(new_n585), .C1(new_n593), .C2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n575), .A2(KEYINPUT13), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT13), .ZN(new_n597));
  NAND4_X1  g411(.A1(new_n215), .A2(new_n217), .A3(new_n597), .A4(G128), .ZN(new_n598));
  AND2_X1   g412(.A1(new_n598), .A2(G134), .ZN(new_n599));
  AOI22_X1  g413(.A1(new_n596), .A2(new_n599), .B1(new_n576), .B2(new_n575), .ZN(new_n600));
  NOR3_X1   g414(.A1(new_n583), .A2(new_n584), .A3(new_n198), .ZN(new_n601));
  OAI21_X1  g415(.A(KEYINPUT90), .B1(new_n589), .B2(new_n580), .ZN(new_n602));
  AOI21_X1  g416(.A(G107), .B1(new_n602), .B2(new_n582), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n600), .B1(new_n601), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n595), .A2(new_n604), .ZN(new_n605));
  NOR3_X1   g419(.A1(new_n323), .A2(new_n468), .A3(G953), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n595), .A2(new_n604), .A3(new_n606), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  AOI21_X1  g424(.A(KEYINPUT92), .B1(new_n610), .B2(new_n311), .ZN(new_n611));
  AND3_X1   g425(.A1(new_n595), .A2(new_n604), .A3(new_n606), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n606), .B1(new_n595), .B2(new_n604), .ZN(new_n613));
  OAI211_X1 g427(.A(KEYINPUT92), .B(new_n311), .C1(new_n612), .C2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n573), .B1(new_n611), .B2(new_n615), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n311), .B1(new_n612), .B2(new_n613), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT92), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n573), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n616), .A2(new_n621), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n571), .A2(new_n622), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n395), .A2(new_n467), .A3(new_n513), .A4(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(G101), .ZN(G3));
  INV_X1    g439(.A(KEYINPUT94), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT93), .ZN(new_n627));
  OAI21_X1  g441(.A(G472), .B1(new_n465), .B2(new_n627), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n425), .A2(new_n429), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n440), .B1(new_n629), .B2(KEYINPUT31), .ZN(new_n630));
  NOR3_X1   g444(.A1(new_n630), .A2(KEYINPUT93), .A3(G902), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n628), .A2(new_n631), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n322), .A2(new_n441), .A3(new_n513), .A4(new_n326), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n626), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  OAI21_X1  g448(.A(KEYINPUT93), .B1(new_n630), .B2(G902), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n465), .A2(new_n627), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n635), .A2(new_n636), .A3(G472), .ZN(new_n637));
  AOI211_X1 g451(.A(G472), .B(G902), .C1(new_n463), .C2(new_n464), .ZN(new_n638));
  INV_X1    g452(.A(new_n513), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n305), .A2(new_n306), .A3(new_n314), .ZN(new_n641));
  AOI22_X1  g455(.A1(new_n269), .A2(new_n268), .B1(new_n296), .B2(new_n258), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n641), .B1(new_n642), .B2(new_n314), .ZN(new_n643));
  AOI211_X1 g457(.A(KEYINPUT79), .B(new_n310), .C1(new_n643), .C2(new_n311), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n644), .A2(new_n319), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n325), .B1(new_n645), .B2(new_n312), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n637), .A2(KEYINPUT94), .A3(new_n640), .A4(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n634), .A2(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT95), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT33), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(KEYINPUT95), .A2(KEYINPUT33), .ZN(new_n653));
  OAI211_X1 g467(.A(new_n652), .B(new_n653), .C1(new_n612), .C2(new_n613), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n608), .A2(new_n650), .A3(new_n651), .A4(new_n609), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n572), .A2(G902), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n617), .A2(new_n572), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n561), .A2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(new_n570), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n391), .B1(new_n380), .B2(new_n384), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n649), .A2(new_n666), .ZN(new_n667));
  XOR2_X1   g481(.A(KEYINPUT34), .B(G104), .Z(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G6));
  INV_X1    g483(.A(new_n622), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n554), .A2(new_n551), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT96), .ZN(new_n672));
  OAI211_X1 g486(.A(new_n672), .B(G475), .C1(new_n559), .C2(G902), .ZN(new_n673));
  AOI21_X1  g487(.A(G902), .B1(new_n558), .B2(new_n528), .ZN(new_n674));
  INV_X1    g488(.A(G475), .ZN(new_n675));
  OAI21_X1  g489(.A(KEYINPUT96), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n671), .A2(new_n673), .A3(new_n676), .ZN(new_n677));
  NOR4_X1   g491(.A1(new_n665), .A2(new_n569), .A3(new_n670), .A4(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n649), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(KEYINPUT97), .ZN(new_n680));
  XOR2_X1   g494(.A(KEYINPUT35), .B(G107), .Z(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(G9));
  NAND2_X1  g496(.A1(new_n463), .A2(new_n464), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(new_n311), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n396), .B1(new_n684), .B2(KEYINPUT93), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n638), .B1(new_n685), .B2(new_n636), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n502), .A2(KEYINPUT36), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n498), .B(new_n687), .ZN(new_n688));
  AND3_X1   g502(.A1(new_n688), .A2(new_n311), .A3(new_n470), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n511), .A2(new_n689), .ZN(new_n690));
  NOR3_X1   g504(.A1(new_n571), .A2(new_n690), .A3(new_n622), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n395), .A2(new_n686), .A3(new_n691), .ZN(new_n692));
  XOR2_X1   g506(.A(KEYINPUT37), .B(G110), .Z(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(G12));
  INV_X1    g508(.A(new_n677), .ZN(new_n695));
  XOR2_X1   g509(.A(new_n564), .B(KEYINPUT98), .Z(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(G900), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n697), .B1(new_n698), .B2(new_n567), .ZN(new_n699));
  INV_X1    g513(.A(new_n699), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n622), .A2(new_n695), .A3(new_n700), .ZN(new_n701));
  AOI211_X1 g515(.A(new_n325), .B(new_n701), .C1(new_n645), .C2(new_n312), .ZN(new_n702));
  INV_X1    g516(.A(new_n690), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(new_n664), .ZN(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n467), .A2(new_n702), .A3(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G128), .ZN(G30));
  NAND2_X1  g521(.A1(new_n461), .A2(new_n462), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n708), .B1(new_n423), .B2(new_n451), .ZN(new_n709));
  OAI21_X1  g523(.A(G472), .B1(new_n709), .B2(G902), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n443), .A2(new_n710), .A3(new_n466), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n389), .A2(KEYINPUT38), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT38), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n713), .B1(new_n385), .B2(new_n388), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  AOI22_X1  g529(.A1(new_n616), .A2(new_n621), .B1(new_n555), .B2(new_n560), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n703), .A2(new_n391), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n711), .A2(new_n715), .A3(new_n716), .A4(new_n717), .ZN(new_n718));
  XOR2_X1   g532(.A(new_n699), .B(KEYINPUT39), .Z(new_n719));
  NAND3_X1  g533(.A1(new_n322), .A2(new_n326), .A3(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT40), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n720), .A2(new_n721), .ZN(new_n723));
  INV_X1    g537(.A(new_n723), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n718), .B1(new_n722), .B2(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(new_n189), .ZN(G45));
  NAND3_X1  g540(.A1(new_n561), .A2(new_n660), .A3(new_n700), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(KEYINPUT99), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT99), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n561), .A2(new_n660), .A3(new_n729), .A4(new_n700), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(new_n731), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n467), .A2(new_n646), .A3(new_n705), .A4(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(KEYINPUT100), .B(G146), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n733), .B(new_n734), .ZN(G48));
  AOI22_X1  g549(.A1(new_n298), .A2(KEYINPUT81), .B1(new_n275), .B2(new_n307), .ZN(new_n736));
  AOI211_X1 g550(.A(G469), .B(G902), .C1(new_n736), .C2(new_n301), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n310), .B1(new_n309), .B2(new_n311), .ZN(new_n738));
  NOR3_X1   g552(.A1(new_n737), .A2(new_n738), .A3(new_n325), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n467), .A2(new_n513), .A3(new_n666), .A4(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(KEYINPUT41), .B(G113), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n740), .B(new_n741), .ZN(G15));
  NAND4_X1  g556(.A1(new_n467), .A2(new_n678), .A3(new_n513), .A4(new_n739), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G116), .ZN(G18));
  NAND2_X1  g558(.A1(new_n309), .A2(new_n311), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n745), .A2(G469), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n746), .A2(new_n326), .A3(new_n312), .A4(new_n664), .ZN(new_n747));
  INV_X1    g561(.A(new_n747), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n748), .A2(new_n467), .A3(new_n691), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G119), .ZN(G21));
  NOR2_X1   g564(.A1(new_n737), .A2(new_n738), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n380), .A2(new_n384), .ZN(new_n752));
  AND4_X1   g566(.A1(new_n570), .A2(new_n752), .A3(new_n390), .A4(new_n716), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n751), .A2(new_n753), .A3(new_n326), .ZN(new_n754));
  NOR3_X1   g568(.A1(new_n428), .A2(new_n406), .A3(new_n423), .ZN(new_n755));
  AOI22_X1  g569(.A1(new_n454), .A2(new_n423), .B1(new_n430), .B2(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(new_n463), .ZN(new_n757));
  NOR2_X1   g571(.A1(G472), .A2(G902), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(KEYINPUT101), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  OAI211_X1 g574(.A(new_n760), .B(new_n513), .C1(new_n396), .C2(new_n465), .ZN(new_n761));
  OAI21_X1  g575(.A(KEYINPUT102), .B1(new_n754), .B2(new_n761), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n396), .B1(new_n683), .B2(new_n311), .ZN(new_n763));
  INV_X1    g577(.A(new_n759), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n764), .B1(new_n756), .B2(new_n463), .ZN(new_n765));
  NOR3_X1   g579(.A1(new_n763), .A2(new_n639), .A3(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT102), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n766), .A2(new_n767), .A3(new_n739), .A4(new_n753), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n762), .A2(new_n768), .ZN(new_n769));
  XOR2_X1   g583(.A(KEYINPUT103), .B(G122), .Z(new_n770));
  XNOR2_X1  g584(.A(new_n769), .B(new_n770), .ZN(G24));
  NOR3_X1   g585(.A1(new_n763), .A2(new_n690), .A3(new_n765), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n748), .A2(new_n772), .A3(new_n732), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G125), .ZN(G27));
  AOI21_X1  g588(.A(new_n391), .B1(new_n385), .B2(new_n388), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n318), .A2(G469), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n312), .A2(new_n776), .ZN(new_n777));
  AND3_X1   g591(.A1(new_n775), .A2(new_n777), .A3(new_n326), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n467), .A2(new_n778), .A3(new_n513), .A4(new_n732), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT42), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT104), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n443), .A2(new_n782), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n457), .B1(new_n638), .B2(KEYINPUT32), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n441), .A2(KEYINPUT104), .A3(new_n442), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n783), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n389), .A2(new_n390), .A3(new_n326), .ZN(new_n787));
  INV_X1    g601(.A(new_n776), .ZN(new_n788));
  AOI21_X1  g602(.A(G902), .B1(new_n736), .B2(new_n301), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n788), .B1(new_n789), .B2(new_n310), .ZN(new_n790));
  NOR3_X1   g604(.A1(new_n787), .A2(new_n731), .A3(new_n790), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n786), .A2(KEYINPUT42), .A3(new_n513), .A4(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n781), .A2(new_n792), .ZN(new_n793));
  XOR2_X1   g607(.A(KEYINPUT105), .B(G131), .Z(new_n794));
  XNOR2_X1  g608(.A(new_n793), .B(new_n794), .ZN(G33));
  INV_X1    g609(.A(new_n701), .ZN(new_n796));
  AND4_X1   g610(.A1(new_n467), .A2(new_n778), .A3(new_n513), .A4(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(new_n250), .ZN(G36));
  INV_X1    g612(.A(new_n719), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n310), .A2(new_n311), .ZN(new_n800));
  INV_X1    g614(.A(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT45), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n310), .B1(new_n643), .B2(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT106), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(new_n805), .ZN(new_n806));
  OAI22_X1  g620(.A1(new_n803), .A2(new_n804), .B1(new_n802), .B2(new_n643), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n801), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT46), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n737), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n316), .A2(new_n317), .ZN(new_n811));
  OAI21_X1  g625(.A(G469), .B1(new_n811), .B2(KEYINPUT45), .ZN(new_n812));
  AOI22_X1  g626(.A1(new_n812), .A2(KEYINPUT106), .B1(KEYINPUT45), .B2(new_n811), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n800), .B1(new_n813), .B2(new_n805), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(KEYINPUT46), .ZN(new_n815));
  AOI211_X1 g629(.A(new_n325), .B(new_n799), .C1(new_n810), .C2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT44), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n562), .A2(new_n660), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(KEYINPUT43), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT43), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n562), .A2(new_n820), .A3(new_n660), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n819), .A2(new_n703), .A3(new_n821), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n817), .B1(new_n686), .B2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(new_n822), .ZN(new_n824));
  OAI211_X1 g638(.A(KEYINPUT44), .B(new_n824), .C1(new_n632), .C2(new_n638), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n816), .A2(new_n823), .A3(new_n775), .A4(new_n825), .ZN(new_n826));
  XNOR2_X1  g640(.A(KEYINPUT107), .B(G137), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n826), .B(new_n827), .ZN(G39));
  INV_X1    g642(.A(new_n775), .ZN(new_n829));
  NOR4_X1   g643(.A1(new_n467), .A2(new_n513), .A3(new_n731), .A4(new_n829), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n325), .B1(new_n810), .B2(new_n815), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n831), .A2(KEYINPUT47), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT47), .ZN(new_n833));
  AOI211_X1 g647(.A(new_n833), .B(new_n325), .C1(new_n810), .C2(new_n815), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n830), .B1(new_n832), .B2(new_n834), .ZN(new_n835));
  XOR2_X1   g649(.A(KEYINPUT108), .B(G140), .Z(new_n836));
  XNOR2_X1  g650(.A(new_n835), .B(new_n836), .ZN(G42));
  INV_X1    g651(.A(KEYINPUT51), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n312), .B1(new_n814), .B2(KEYINPUT46), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n808), .A2(new_n809), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n326), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n841), .A2(new_n833), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n831), .A2(KEYINPUT47), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n751), .A2(new_n325), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n842), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  AND3_X1   g659(.A1(new_n819), .A2(new_n697), .A3(new_n821), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n766), .A2(new_n846), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n847), .A2(new_n829), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n838), .B1(new_n845), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n751), .A2(new_n326), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n513), .A2(new_n565), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n850), .A2(new_n829), .A3(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(new_n711), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n561), .A2(new_n660), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n852), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT114), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NOR4_X1   g671(.A1(new_n711), .A2(new_n850), .A3(new_n829), .A4(new_n851), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n858), .A2(KEYINPUT114), .A3(new_n854), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n846), .A2(new_n739), .A3(new_n775), .ZN(new_n860));
  INV_X1    g674(.A(new_n860), .ZN(new_n861));
  AOI22_X1  g675(.A1(new_n857), .A2(new_n859), .B1(new_n772), .B2(new_n861), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n847), .A2(new_n715), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n746), .A2(new_n391), .A3(new_n326), .A4(new_n312), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT113), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n864), .B(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n863), .A2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT50), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n863), .A2(new_n866), .A3(KEYINPUT50), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n849), .A2(new_n862), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n872), .A2(KEYINPUT115), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT115), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n849), .A2(new_n862), .A3(new_n874), .A4(new_n871), .ZN(new_n875));
  OAI211_X1 g689(.A(G952), .B(new_n273), .C1(new_n847), .C2(new_n747), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n876), .B1(new_n662), .B2(new_n858), .ZN(new_n877));
  AND2_X1   g691(.A1(new_n786), .A2(new_n513), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n878), .A2(KEYINPUT116), .A3(KEYINPUT48), .A4(new_n861), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n861), .A2(new_n513), .A3(new_n786), .ZN(new_n880));
  XOR2_X1   g694(.A(KEYINPUT116), .B(KEYINPUT48), .Z(new_n881));
  NAND2_X1  g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n877), .A2(new_n879), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n883), .A2(KEYINPUT117), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT117), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n877), .A2(new_n879), .A3(new_n885), .A4(new_n882), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n873), .A2(new_n875), .A3(new_n887), .ZN(new_n888));
  OR3_X1    g702(.A1(new_n832), .A2(new_n834), .A3(KEYINPUT112), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n842), .A2(new_n843), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n890), .A2(KEYINPUT112), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n889), .A2(new_n891), .A3(new_n844), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(new_n848), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n862), .A2(new_n871), .ZN(new_n894));
  INV_X1    g708(.A(new_n894), .ZN(new_n895));
  AOI21_X1  g709(.A(KEYINPUT51), .B1(new_n893), .B2(new_n895), .ZN(new_n896));
  OAI21_X1  g710(.A(KEYINPUT118), .B1(new_n888), .B2(new_n896), .ZN(new_n897));
  AOI22_X1  g711(.A1(new_n872), .A2(KEYINPUT115), .B1(new_n884), .B2(new_n886), .ZN(new_n898));
  INV_X1    g712(.A(new_n848), .ZN(new_n899));
  AOI22_X1  g713(.A1(new_n890), .A2(KEYINPUT112), .B1(new_n325), .B2(new_n751), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n899), .B1(new_n900), .B2(new_n889), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n838), .B1(new_n901), .B2(new_n894), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT118), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n898), .A2(new_n902), .A3(new_n903), .A4(new_n875), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n897), .A2(new_n904), .ZN(new_n905));
  XNOR2_X1  g719(.A(KEYINPUT111), .B(KEYINPUT53), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT109), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n663), .B1(new_n392), .B2(new_n394), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n634), .A2(new_n647), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n907), .B1(new_n909), .B2(new_n624), .ZN(new_n910));
  AOI211_X1 g724(.A(new_n571), .B(new_n670), .C1(new_n392), .C2(new_n394), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n634), .A2(new_n911), .A3(new_n647), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(new_n692), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n910), .A2(new_n913), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n769), .A2(new_n740), .A3(new_n743), .A4(new_n749), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n829), .A2(new_n325), .ZN(new_n916));
  NOR4_X1   g730(.A1(new_n690), .A2(new_n622), .A3(new_n677), .A4(new_n699), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n467), .A2(new_n916), .A3(new_n322), .A4(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n791), .A2(new_n772), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n915), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n909), .A2(new_n907), .A3(new_n624), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n797), .B1(new_n781), .B2(new_n792), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n914), .A2(new_n921), .A3(new_n922), .A4(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n704), .B1(new_n784), .B2(new_n443), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n747), .A2(new_n731), .ZN(new_n926));
  AOI22_X1  g740(.A1(new_n925), .A2(new_n702), .B1(new_n926), .B2(new_n772), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT52), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n325), .B1(new_n699), .B2(KEYINPUT110), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n929), .B1(KEYINPUT110), .B2(new_n699), .ZN(new_n930));
  NOR3_X1   g744(.A1(new_n511), .A2(new_n689), .A3(new_n930), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n931), .A2(new_n664), .A3(new_n716), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n932), .A2(new_n790), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n711), .A2(new_n933), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n927), .A2(new_n928), .A3(new_n733), .A4(new_n934), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n733), .A2(new_n773), .A3(new_n706), .A4(new_n934), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(KEYINPUT52), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n906), .B1(new_n924), .B2(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT54), .ZN(new_n940));
  AND3_X1   g754(.A1(new_n769), .A2(new_n740), .A3(new_n749), .ZN(new_n941));
  INV_X1    g755(.A(new_n920), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n941), .A2(new_n923), .A3(new_n743), .A4(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(new_n922), .ZN(new_n945));
  NOR3_X1   g759(.A1(new_n945), .A2(new_n910), .A3(new_n913), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n773), .A2(new_n706), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(KEYINPUT52), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n935), .A2(new_n937), .A3(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(new_n949), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n944), .A2(new_n946), .A3(KEYINPUT53), .A4(new_n950), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n939), .A2(new_n940), .A3(new_n951), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n924), .A2(new_n938), .ZN(new_n953));
  INV_X1    g767(.A(new_n906), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n944), .A2(new_n946), .A3(new_n950), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT53), .ZN(new_n956));
  AOI22_X1  g770(.A1(new_n953), .A2(new_n954), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n952), .B1(new_n957), .B2(new_n940), .ZN(new_n958));
  OAI22_X1  g772(.A1(new_n905), .A2(new_n958), .B1(G952), .B2(G953), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n513), .A2(new_n390), .A3(new_n326), .ZN(new_n960));
  INV_X1    g774(.A(new_n751), .ZN(new_n961));
  AOI211_X1 g775(.A(new_n818), .B(new_n960), .C1(new_n961), .C2(KEYINPUT49), .ZN(new_n962));
  INV_X1    g776(.A(new_n715), .ZN(new_n963));
  OR2_X1    g777(.A1(new_n961), .A2(KEYINPUT49), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n962), .A2(new_n963), .A3(new_n853), .A4(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n959), .A2(new_n965), .ZN(G75));
  NOR2_X1   g780(.A1(new_n372), .A2(new_n373), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n368), .A2(new_n370), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n969), .A2(new_n374), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n970), .B(KEYINPUT55), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n311), .B1(new_n939), .B2(new_n951), .ZN(new_n972));
  AOI211_X1 g786(.A(KEYINPUT56), .B(new_n971), .C1(new_n972), .C2(new_n329), .ZN(new_n973));
  INV_X1    g787(.A(new_n971), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n939), .A2(new_n951), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n975), .A2(G902), .A3(new_n329), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT56), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n974), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n273), .A2(G952), .ZN(new_n979));
  NOR3_X1   g793(.A1(new_n973), .A2(new_n978), .A3(new_n979), .ZN(G51));
  XNOR2_X1  g794(.A(new_n800), .B(KEYINPUT57), .ZN(new_n981));
  AND3_X1   g795(.A1(new_n939), .A2(new_n940), .A3(new_n951), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n940), .B1(new_n939), .B2(new_n951), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n981), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n984), .A2(new_n309), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n972), .A2(new_n805), .A3(new_n813), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n979), .B1(new_n985), .B2(new_n986), .ZN(G54));
  AND2_X1   g801(.A1(KEYINPUT58), .A2(G475), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n972), .A2(new_n988), .ZN(new_n989));
  INV_X1    g803(.A(new_n544), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n979), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  NAND4_X1  g805(.A1(new_n972), .A2(KEYINPUT119), .A3(new_n544), .A4(new_n988), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n972), .A2(new_n544), .A3(new_n988), .ZN(new_n993));
  INV_X1    g807(.A(KEYINPUT119), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  AND3_X1   g809(.A1(new_n991), .A2(new_n992), .A3(new_n995), .ZN(G60));
  NAND2_X1  g810(.A1(G478), .A2(G902), .ZN(new_n997));
  XOR2_X1   g811(.A(new_n997), .B(KEYINPUT59), .Z(new_n998));
  INV_X1    g812(.A(new_n998), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n656), .B1(new_n958), .B2(new_n999), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n998), .B1(new_n654), .B2(new_n655), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n1001), .B1(new_n982), .B2(new_n983), .ZN(new_n1002));
  INV_X1    g816(.A(new_n979), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NOR2_X1   g818(.A1(new_n1000), .A2(new_n1004), .ZN(G63));
  NAND2_X1  g819(.A1(G217), .A2(G902), .ZN(new_n1006));
  XNOR2_X1  g820(.A(new_n1006), .B(KEYINPUT60), .ZN(new_n1007));
  INV_X1    g821(.A(new_n1007), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n975), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1009), .A2(new_n505), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n1007), .B1(new_n939), .B2(new_n951), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n979), .B1(new_n1011), .B2(new_n688), .ZN(new_n1012));
  INV_X1    g826(.A(KEYINPUT120), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n1013), .B1(new_n1011), .B2(new_n688), .ZN(new_n1014));
  OAI211_X1 g828(.A(new_n1010), .B(new_n1012), .C1(new_n1014), .C2(KEYINPUT61), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n909), .A2(new_n624), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1016), .A2(KEYINPUT109), .ZN(new_n1017));
  AND2_X1   g831(.A1(new_n912), .A2(new_n692), .ZN(new_n1018));
  NAND3_X1  g832(.A1(new_n1017), .A2(new_n922), .A3(new_n1018), .ZN(new_n1019));
  NOR2_X1   g833(.A1(new_n1019), .A2(new_n943), .ZN(new_n1020));
  INV_X1    g834(.A(new_n938), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n954), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  NOR4_X1   g836(.A1(new_n1019), .A2(new_n943), .A3(new_n949), .A4(new_n956), .ZN(new_n1023));
  OAI211_X1 g837(.A(new_n688), .B(new_n1008), .C1(new_n1022), .C2(new_n1023), .ZN(new_n1024));
  OAI211_X1 g838(.A(new_n1024), .B(new_n1003), .C1(new_n506), .C2(new_n1011), .ZN(new_n1025));
  AOI21_X1  g839(.A(KEYINPUT61), .B1(new_n1024), .B2(KEYINPUT120), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n1015), .A2(new_n1027), .ZN(G66));
  INV_X1    g842(.A(new_n568), .ZN(new_n1029));
  AOI21_X1  g843(.A(new_n273), .B1(new_n1029), .B2(G224), .ZN(new_n1030));
  NOR2_X1   g844(.A1(new_n1019), .A2(new_n915), .ZN(new_n1031));
  INV_X1    g845(.A(new_n1031), .ZN(new_n1032));
  AOI21_X1  g846(.A(new_n1030), .B1(new_n1032), .B2(new_n273), .ZN(new_n1033));
  OAI21_X1  g847(.A(new_n968), .B1(G898), .B2(new_n273), .ZN(new_n1034));
  XOR2_X1   g848(.A(new_n1033), .B(new_n1034), .Z(G69));
  AOI21_X1  g849(.A(new_n273), .B1(G227), .B2(G900), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n532), .A2(new_n533), .ZN(new_n1037));
  XOR2_X1   g851(.A(new_n416), .B(new_n1037), .Z(new_n1038));
  NAND2_X1  g852(.A1(new_n698), .A2(G953), .ZN(new_n1039));
  XOR2_X1   g853(.A(new_n1039), .B(KEYINPUT125), .Z(new_n1040));
  NAND4_X1  g854(.A1(new_n878), .A2(new_n816), .A3(new_n664), .A4(new_n716), .ZN(new_n1041));
  NAND3_X1  g855(.A1(new_n835), .A2(new_n1041), .A3(new_n923), .ZN(new_n1042));
  INV_X1    g856(.A(KEYINPUT126), .ZN(new_n1043));
  NAND3_X1  g857(.A1(new_n733), .A2(new_n773), .A3(new_n706), .ZN(new_n1044));
  INV_X1    g858(.A(new_n1044), .ZN(new_n1045));
  AOI21_X1  g859(.A(new_n1043), .B1(new_n826), .B2(new_n1045), .ZN(new_n1046));
  INV_X1    g860(.A(new_n1046), .ZN(new_n1047));
  NAND3_X1  g861(.A1(new_n826), .A2(new_n1043), .A3(new_n1045), .ZN(new_n1048));
  AOI21_X1  g862(.A(new_n1042), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g863(.A(new_n1040), .B1(new_n1049), .B2(G953), .ZN(new_n1050));
  NAND2_X1  g864(.A1(new_n1050), .A2(KEYINPUT127), .ZN(new_n1051));
  AND2_X1   g865(.A1(new_n835), .A2(new_n1041), .ZN(new_n1052));
  AND3_X1   g866(.A1(new_n826), .A2(new_n1043), .A3(new_n1045), .ZN(new_n1053));
  OAI211_X1 g867(.A(new_n1052), .B(new_n923), .C1(new_n1053), .C2(new_n1046), .ZN(new_n1054));
  NAND2_X1  g868(.A1(new_n1054), .A2(new_n273), .ZN(new_n1055));
  INV_X1    g869(.A(KEYINPUT127), .ZN(new_n1056));
  NAND3_X1  g870(.A1(new_n1055), .A2(new_n1056), .A3(new_n1040), .ZN(new_n1057));
  AOI21_X1  g871(.A(new_n1038), .B1(new_n1051), .B2(new_n1057), .ZN(new_n1058));
  INV_X1    g872(.A(new_n1038), .ZN(new_n1059));
  INV_X1    g873(.A(new_n835), .ZN(new_n1060));
  INV_X1    g874(.A(KEYINPUT122), .ZN(new_n1061));
  NAND2_X1  g875(.A1(new_n467), .A2(new_n513), .ZN(new_n1062));
  AOI21_X1  g876(.A(new_n620), .B1(new_n619), .B2(new_n614), .ZN(new_n1063));
  NOR2_X1   g877(.A1(new_n611), .A2(new_n573), .ZN(new_n1064));
  OAI211_X1 g878(.A(new_n560), .B(new_n555), .C1(new_n1063), .C2(new_n1064), .ZN(new_n1065));
  AND3_X1   g879(.A1(new_n661), .A2(new_n1065), .A3(KEYINPUT121), .ZN(new_n1066));
  AOI21_X1  g880(.A(KEYINPUT121), .B1(new_n661), .B2(new_n1065), .ZN(new_n1067));
  NOR2_X1   g881(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND4_X1  g882(.A1(new_n1068), .A2(new_n646), .A3(new_n719), .A4(new_n775), .ZN(new_n1069));
  OAI21_X1  g883(.A(new_n1061), .B1(new_n1062), .B2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g884(.A(new_n639), .B1(new_n784), .B2(new_n443), .ZN(new_n1071));
  INV_X1    g885(.A(new_n720), .ZN(new_n1072));
  NOR3_X1   g886(.A1(new_n829), .A2(new_n1066), .A3(new_n1067), .ZN(new_n1073));
  NAND4_X1  g887(.A1(new_n1071), .A2(KEYINPUT122), .A3(new_n1072), .A4(new_n1073), .ZN(new_n1074));
  AND2_X1   g888(.A1(new_n1070), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g889(.A1(new_n1075), .A2(new_n826), .ZN(new_n1076));
  INV_X1    g890(.A(KEYINPUT123), .ZN(new_n1077));
  NAND2_X1  g891(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g892(.A1(new_n1075), .A2(new_n826), .A3(KEYINPUT123), .ZN(new_n1079));
  AOI21_X1  g893(.A(new_n1060), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  AND2_X1   g894(.A1(new_n724), .A2(new_n722), .ZN(new_n1081));
  OAI211_X1 g895(.A(new_n1045), .B(KEYINPUT62), .C1(new_n1081), .C2(new_n718), .ZN(new_n1082));
  INV_X1    g896(.A(KEYINPUT62), .ZN(new_n1083));
  OAI21_X1  g897(.A(new_n1083), .B1(new_n725), .B2(new_n1044), .ZN(new_n1084));
  NAND2_X1  g898(.A1(new_n1082), .A2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g899(.A1(new_n1080), .A2(KEYINPUT124), .A3(new_n1085), .ZN(new_n1086));
  AND3_X1   g900(.A1(new_n1075), .A2(new_n826), .A3(KEYINPUT123), .ZN(new_n1087));
  AOI21_X1  g901(.A(KEYINPUT123), .B1(new_n1075), .B2(new_n826), .ZN(new_n1088));
  OAI211_X1 g902(.A(new_n1085), .B(new_n835), .C1(new_n1087), .C2(new_n1088), .ZN(new_n1089));
  INV_X1    g903(.A(KEYINPUT124), .ZN(new_n1090));
  NAND2_X1  g904(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g905(.A1(new_n1086), .A2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g906(.A(new_n1059), .B1(new_n1092), .B2(new_n273), .ZN(new_n1093));
  OAI21_X1  g907(.A(new_n1036), .B1(new_n1058), .B2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g908(.A(KEYINPUT124), .B1(new_n1080), .B2(new_n1085), .ZN(new_n1095));
  NOR2_X1   g909(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1096));
  OAI21_X1  g910(.A(new_n273), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g911(.A1(new_n1097), .A2(new_n1038), .ZN(new_n1098));
  AOI21_X1  g912(.A(new_n1056), .B1(new_n1055), .B2(new_n1040), .ZN(new_n1099));
  INV_X1    g913(.A(new_n1040), .ZN(new_n1100));
  AOI211_X1 g914(.A(KEYINPUT127), .B(new_n1100), .C1(new_n1054), .C2(new_n273), .ZN(new_n1101));
  OAI21_X1  g915(.A(new_n1059), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g916(.A(new_n1036), .ZN(new_n1103));
  NAND3_X1  g917(.A1(new_n1098), .A2(new_n1102), .A3(new_n1103), .ZN(new_n1104));
  NAND2_X1  g918(.A1(new_n1094), .A2(new_n1104), .ZN(G72));
  NAND3_X1  g919(.A1(new_n1086), .A2(new_n1091), .A3(new_n1031), .ZN(new_n1106));
  NAND2_X1  g920(.A1(G472), .A2(G902), .ZN(new_n1107));
  XOR2_X1   g921(.A(new_n1107), .B(KEYINPUT63), .Z(new_n1108));
  AOI211_X1 g922(.A(new_n418), .B(new_n423), .C1(new_n1106), .C2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g923(.A(new_n1108), .B1(new_n1032), .B2(new_n1054), .ZN(new_n1110));
  NOR3_X1   g924(.A1(new_n428), .A2(new_n406), .A3(new_n424), .ZN(new_n1111));
  AOI21_X1  g925(.A(new_n979), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  NOR2_X1   g926(.A1(new_n418), .A2(new_n424), .ZN(new_n1113));
  OAI21_X1  g927(.A(new_n1108), .B1(new_n708), .B2(new_n1113), .ZN(new_n1114));
  OAI21_X1  g928(.A(new_n1112), .B1(new_n957), .B2(new_n1114), .ZN(new_n1115));
  NOR2_X1   g929(.A1(new_n1109), .A2(new_n1115), .ZN(G57));
endmodule


