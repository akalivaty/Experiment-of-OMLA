//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 1 1 1 1 1 1 1 0 1 1 1 0 1 0 0 1 1 0 0 0 0 1 1 1 1 0 1 0 1 0 0 1 1 1 0 0 0 1 0 1 0 0 1 1 0 1 0 1 1 0 0 0 1 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:09 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1079, new_n1080, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1143, new_n1144, new_n1145,
    new_n1146, new_n1147, new_n1148, new_n1149, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1169, new_n1170, new_n1171,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1242, new_n1243;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G13), .ZN(new_n204));
  OAI211_X1 g0004(.A(new_n204), .B(G250), .C1(G257), .C2(G264), .ZN(new_n205));
  XOR2_X1   g0005(.A(new_n205), .B(KEYINPUT0), .Z(new_n206));
  AOI22_X1  g0006(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  XOR2_X1   g0009(.A(KEYINPUT64), .B(G244), .Z(new_n210));
  AOI21_X1  g0010(.A(new_n209), .B1(G77), .B2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(G58), .ZN(new_n212));
  INV_X1    g0012(.A(G232), .ZN(new_n213));
  INV_X1    g0013(.A(G97), .ZN(new_n214));
  INV_X1    g0014(.A(G257), .ZN(new_n215));
  OAI221_X1 g0015(.A(new_n211), .B1(new_n212), .B2(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(G50), .ZN(new_n217));
  INV_X1    g0017(.A(G226), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n203), .B1(new_n216), .B2(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n220), .B1(KEYINPUT65), .B2(KEYINPUT1), .ZN(new_n221));
  NAND2_X1  g0021(.A1(KEYINPUT65), .A2(KEYINPUT1), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n221), .B(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G13), .ZN(new_n224));
  INV_X1    g0024(.A(G20), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NOR2_X1   g0026(.A1(G58), .A2(G68), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n228), .A2(G50), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  AOI211_X1 g0030(.A(new_n206), .B(new_n223), .C1(new_n226), .C2(new_n230), .ZN(G361));
  XNOR2_X1  g0031(.A(KEYINPUT2), .B(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(new_n213), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT66), .B(G264), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n235), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G68), .B(G77), .Z(new_n241));
  XNOR2_X1  g0041(.A(G50), .B(G58), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G107), .B(G116), .Z(new_n244));
  XNOR2_X1  g0044(.A(G87), .B(G97), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  AOI21_X1  g0047(.A(new_n224), .B1(G33), .B2(G41), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n215), .A2(G1698), .ZN(new_n249));
  AND2_X1   g0049(.A1(KEYINPUT3), .A2(G33), .ZN(new_n250));
  NOR2_X1   g0050(.A1(KEYINPUT3), .A2(G33), .ZN(new_n251));
  OAI221_X1 g0051(.A(new_n249), .B1(G250), .B2(G1698), .C1(new_n250), .C2(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(G33), .A2(G294), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G45), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n255), .A2(G1), .ZN(new_n256));
  AND2_X1   g0056(.A1(KEYINPUT5), .A2(G41), .ZN(new_n257));
  NOR2_X1   g0057(.A1(KEYINPUT5), .A2(G41), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n256), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(G33), .A2(G41), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n260), .A2(G1), .A3(G13), .ZN(new_n261));
  AND2_X1   g0061(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  AOI22_X1  g0062(.A1(new_n248), .A2(new_n254), .B1(new_n262), .B2(G264), .ZN(new_n263));
  OAI211_X1 g0063(.A(new_n256), .B(G274), .C1(new_n258), .C2(new_n257), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G200), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n261), .B1(new_n252), .B2(new_n253), .ZN(new_n268));
  OR2_X1    g0068(.A1(new_n268), .A2(KEYINPUT78), .ZN(new_n269));
  INV_X1    g0069(.A(new_n264), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n270), .B1(new_n268), .B2(KEYINPUT78), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n262), .A2(G264), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n269), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n267), .B1(G190), .B2(new_n273), .ZN(new_n274));
  NAND3_X1  g0074(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n275));
  AND2_X1   g0075(.A1(new_n275), .A2(new_n224), .ZN(new_n276));
  INV_X1    g0076(.A(G1), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G33), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n277), .A2(G13), .A3(G20), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n276), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G107), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  OAI211_X1 g0082(.A(new_n225), .B(G87), .C1(new_n250), .C2(new_n251), .ZN(new_n283));
  NAND2_X1  g0083(.A1(KEYINPUT77), .A2(KEYINPUT22), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT3), .ZN(new_n287));
  INV_X1    g0087(.A(G33), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(KEYINPUT3), .A2(G33), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND4_X1  g0091(.A1(new_n291), .A2(new_n225), .A3(G87), .A4(new_n284), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n286), .A2(new_n292), .ZN(new_n293));
  XNOR2_X1  g0093(.A(KEYINPUT74), .B(G116), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n288), .A2(G20), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n281), .A2(G20), .ZN(new_n297));
  XNOR2_X1  g0097(.A(new_n297), .B(KEYINPUT23), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n293), .A2(new_n296), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(KEYINPUT24), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT24), .ZN(new_n302));
  NAND4_X1  g0102(.A1(new_n293), .A2(new_n302), .A3(new_n296), .A4(new_n299), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n275), .A2(new_n224), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n282), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n279), .A2(G107), .ZN(new_n307));
  XNOR2_X1  g0107(.A(new_n307), .B(KEYINPUT25), .ZN(new_n308));
  AND3_X1   g0108(.A1(new_n274), .A2(new_n306), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n273), .A2(G169), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n263), .A2(G179), .A3(new_n264), .ZN(new_n311));
  AOI22_X1  g0111(.A1(new_n306), .A2(new_n308), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n309), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(G1698), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(G222), .ZN(new_n315));
  NAND2_X1  g0115(.A1(G223), .A2(G1698), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n291), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  OAI211_X1 g0117(.A(new_n317), .B(new_n248), .C1(G77), .C2(new_n291), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n277), .B1(G41), .B2(G45), .ZN(new_n319));
  INV_X1    g0119(.A(G274), .ZN(new_n320));
  OR2_X1    g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n261), .A2(new_n319), .ZN(new_n322));
  OAI211_X1 g0122(.A(new_n318), .B(new_n321), .C1(new_n218), .C2(new_n322), .ZN(new_n323));
  OR2_X1    g0123(.A1(new_n323), .A2(G179), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n276), .A2(KEYINPUT67), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n225), .A2(G1), .ZN(new_n326));
  AND3_X1   g0126(.A1(new_n275), .A2(KEYINPUT67), .A3(new_n224), .ZN(new_n327));
  NOR3_X1   g0127(.A1(new_n325), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(G50), .ZN(new_n329));
  OAI21_X1  g0129(.A(G20), .B1(new_n228), .B2(G50), .ZN(new_n330));
  INV_X1    g0130(.A(G150), .ZN(new_n331));
  NOR2_X1   g0131(.A1(G20), .A2(G33), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(new_n295), .ZN(new_n334));
  XNOR2_X1  g0134(.A(KEYINPUT8), .B(G58), .ZN(new_n335));
  OAI221_X1 g0135(.A(new_n330), .B1(new_n331), .B2(new_n333), .C1(new_n334), .C2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(new_n305), .ZN(new_n337));
  OAI211_X1 g0137(.A(new_n329), .B(new_n337), .C1(G50), .C2(new_n279), .ZN(new_n338));
  INV_X1    g0138(.A(G169), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n323), .A2(new_n339), .ZN(new_n340));
  AND3_X1   g0140(.A1(new_n324), .A2(new_n338), .A3(new_n340), .ZN(new_n341));
  XNOR2_X1  g0141(.A(new_n338), .B(KEYINPUT9), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(G190), .ZN(new_n344));
  OR2_X1    g0144(.A1(new_n323), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n323), .A2(G200), .ZN(new_n346));
  AND2_X1   g0146(.A1(new_n346), .A2(KEYINPUT70), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n346), .A2(KEYINPUT70), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n345), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  OAI21_X1  g0149(.A(KEYINPUT10), .B1(new_n343), .B2(new_n349), .ZN(new_n350));
  OR2_X1    g0150(.A1(new_n347), .A2(new_n348), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT10), .ZN(new_n352));
  NAND4_X1  g0152(.A1(new_n351), .A2(new_n352), .A3(new_n342), .A4(new_n345), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n341), .B1(new_n350), .B2(new_n353), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n319), .A2(new_n320), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n218), .A2(new_n314), .ZN(new_n356));
  OAI211_X1 g0156(.A(new_n291), .B(new_n356), .C1(G232), .C2(new_n314), .ZN(new_n357));
  NAND2_X1  g0157(.A1(G33), .A2(G97), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n355), .B1(new_n359), .B2(new_n248), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT13), .ZN(new_n361));
  INV_X1    g0161(.A(new_n322), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(G238), .ZN(new_n363));
  AND3_X1   g0163(.A1(new_n360), .A2(new_n361), .A3(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n361), .B1(new_n360), .B2(new_n363), .ZN(new_n365));
  OAI21_X1  g0165(.A(G169), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(KEYINPUT14), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n364), .A2(new_n365), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(G179), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT14), .ZN(new_n370));
  OAI211_X1 g0170(.A(new_n370), .B(G169), .C1(new_n364), .C2(new_n365), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n367), .A2(new_n369), .A3(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(G68), .ZN(new_n373));
  AOI22_X1  g0173(.A1(new_n295), .A2(G77), .B1(G20), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n332), .A2(G50), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n276), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  XOR2_X1   g0176(.A(new_n376), .B(KEYINPUT11), .Z(new_n377));
  INV_X1    g0177(.A(KEYINPUT69), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n279), .A2(new_n378), .ZN(new_n379));
  NAND4_X1  g0179(.A1(new_n277), .A2(KEYINPUT69), .A3(G13), .A4(G20), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n381), .A2(KEYINPUT12), .A3(new_n373), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT12), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n279), .A2(new_n383), .ZN(new_n384));
  NOR3_X1   g0184(.A1(new_n381), .A2(new_n305), .A3(new_n326), .ZN(new_n385));
  OAI21_X1  g0185(.A(G68), .B1(new_n385), .B2(new_n383), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n377), .A2(new_n382), .A3(new_n384), .A4(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n372), .A2(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n387), .B1(new_n368), .B2(G190), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n389), .B1(new_n266), .B2(new_n368), .ZN(new_n390));
  XOR2_X1   g0190(.A(KEYINPUT8), .B(G58), .Z(new_n391));
  NAND2_X1  g0191(.A1(new_n333), .A2(KEYINPUT68), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT68), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n332), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n391), .A2(new_n392), .A3(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(G77), .ZN(new_n396));
  XNOR2_X1  g0196(.A(KEYINPUT15), .B(G87), .ZN(new_n397));
  OAI221_X1 g0197(.A(new_n395), .B1(new_n225), .B2(new_n396), .C1(new_n334), .C2(new_n397), .ZN(new_n398));
  AOI22_X1  g0198(.A1(new_n398), .A2(new_n305), .B1(G77), .B2(new_n385), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n381), .A2(new_n396), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(G238), .A2(G1698), .ZN(new_n402));
  OAI211_X1 g0202(.A(new_n291), .B(new_n402), .C1(new_n213), .C2(G1698), .ZN(new_n403));
  OAI211_X1 g0203(.A(new_n403), .B(new_n248), .C1(G107), .C2(new_n291), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n362), .A2(new_n210), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n404), .A2(new_n321), .A3(new_n405), .ZN(new_n406));
  AND2_X1   g0206(.A1(new_n406), .A2(G200), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n406), .A2(new_n344), .ZN(new_n408));
  OR3_X1    g0208(.A1(new_n401), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n354), .A2(new_n388), .A3(new_n390), .A4(new_n409), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n391), .A2(new_n279), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n411), .B1(new_n328), .B2(new_n391), .ZN(new_n412));
  INV_X1    g0212(.A(new_n412), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n212), .A2(new_n373), .ZN(new_n414));
  OAI21_X1  g0214(.A(G20), .B1(new_n414), .B2(new_n227), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n332), .A2(G159), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n250), .A2(new_n251), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n418), .A2(KEYINPUT7), .A3(new_n225), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n289), .A2(new_n225), .A3(new_n290), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT71), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT7), .ZN(new_n422));
  AND3_X1   g0222(.A1(new_n420), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n421), .B1(new_n420), .B2(new_n422), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n419), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n417), .B1(new_n425), .B2(G68), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n276), .B1(new_n426), .B2(KEYINPUT16), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT16), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n420), .A2(new_n422), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n373), .B1(new_n429), .B2(new_n419), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n428), .B1(new_n430), .B2(new_n417), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n413), .B1(new_n427), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n218), .A2(G1698), .ZN(new_n433));
  OAI221_X1 g0233(.A(new_n433), .B1(G223), .B2(G1698), .C1(new_n250), .C2(new_n251), .ZN(new_n434));
  NAND2_X1  g0234(.A1(G33), .A2(G87), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n261), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n321), .B1(new_n322), .B2(new_n213), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(G200), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n438), .A2(G190), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n432), .A2(KEYINPUT17), .A3(new_n440), .A4(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n417), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n420), .A2(new_n422), .ZN(new_n444));
  NOR3_X1   g0244(.A1(new_n250), .A2(new_n251), .A3(G20), .ZN(new_n445));
  OAI21_X1  g0245(.A(KEYINPUT71), .B1(new_n445), .B2(KEYINPUT7), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n420), .A2(new_n421), .A3(new_n422), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n444), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  OAI211_X1 g0248(.A(KEYINPUT16), .B(new_n443), .C1(new_n448), .C2(new_n373), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n449), .A2(new_n305), .A3(new_n431), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n450), .A2(new_n440), .A3(new_n441), .A4(new_n412), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT17), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n442), .A2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n450), .A2(new_n412), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n434), .A2(new_n435), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(new_n248), .ZN(new_n458));
  INV_X1    g0258(.A(new_n437), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n339), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(G179), .ZN(new_n461));
  NOR3_X1   g0261(.A1(new_n436), .A2(new_n437), .A3(new_n461), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(KEYINPUT18), .B1(new_n456), .B2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT18), .ZN(new_n466));
  AOI211_X1 g0266(.A(new_n466), .B(new_n463), .C1(new_n450), .C2(new_n412), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n455), .A2(new_n469), .ZN(new_n470));
  OR2_X1    g0270(.A1(new_n406), .A2(G179), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n406), .A2(new_n339), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n401), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  NOR3_X1   g0274(.A1(new_n410), .A2(new_n470), .A3(new_n474), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n294), .B1(new_n379), .B2(new_n380), .ZN(new_n476));
  INV_X1    g0276(.A(G116), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n477), .B1(new_n277), .B2(G33), .ZN(new_n478));
  AND4_X1   g0278(.A1(new_n276), .A2(new_n379), .A3(new_n380), .A4(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(G33), .A2(G283), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n480), .B(new_n225), .C1(G33), .C2(new_n214), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n305), .B(new_n481), .C1(new_n294), .C2(new_n225), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT20), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n477), .A2(KEYINPUT74), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT74), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(G116), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(G20), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n489), .A2(KEYINPUT20), .A3(new_n305), .A4(new_n481), .ZN(new_n490));
  AOI211_X1 g0290(.A(new_n476), .B(new_n479), .C1(new_n484), .C2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT75), .ZN(new_n492));
  INV_X1    g0292(.A(G303), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n289), .A2(new_n493), .A3(new_n290), .ZN(new_n494));
  NAND2_X1  g0294(.A1(G264), .A2(G1698), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n495), .B1(new_n215), .B2(G1698), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n494), .B(new_n248), .C1(new_n418), .C2(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n259), .A2(G270), .A3(new_n261), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n497), .A2(new_n264), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(G200), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n497), .A2(new_n498), .A3(G190), .A4(new_n264), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n491), .A2(new_n492), .A3(new_n500), .A4(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n484), .A2(new_n490), .ZN(new_n503));
  INV_X1    g0303(.A(new_n476), .ZN(new_n504));
  INV_X1    g0304(.A(new_n479), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n503), .A2(new_n501), .A3(new_n504), .A4(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(new_n500), .ZN(new_n507));
  OAI21_X1  g0307(.A(KEYINPUT75), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  AND2_X1   g0308(.A1(new_n502), .A2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT21), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n499), .A2(G169), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n510), .B1(new_n491), .B2(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n503), .A2(new_n504), .A3(new_n505), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n499), .A2(new_n461), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(new_n511), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n516), .A2(new_n513), .A3(KEYINPUT21), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n512), .A2(new_n515), .A3(new_n517), .ZN(new_n518));
  OAI21_X1  g0318(.A(KEYINPUT76), .B1(new_n509), .B2(new_n518), .ZN(new_n519));
  NOR3_X1   g0319(.A1(new_n491), .A2(new_n510), .A3(new_n511), .ZN(new_n520));
  AOI21_X1  g0320(.A(KEYINPUT21), .B1(new_n516), .B2(new_n513), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n502), .A2(new_n508), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT76), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n522), .A2(new_n523), .A3(new_n524), .A4(new_n515), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n519), .A2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT4), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n527), .A2(G1698), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n528), .B(G244), .C1(new_n251), .C2(new_n250), .ZN(new_n529));
  INV_X1    g0329(.A(G244), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n530), .B1(new_n289), .B2(new_n290), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n529), .B(new_n480), .C1(new_n531), .C2(KEYINPUT4), .ZN(new_n532));
  OAI21_X1  g0332(.A(G250), .B1(new_n250), .B2(new_n251), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n314), .B1(new_n533), .B2(KEYINPUT4), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n248), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT72), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n270), .B1(new_n262), .B2(G257), .ZN(new_n538));
  OAI211_X1 g0338(.A(KEYINPUT72), .B(new_n248), .C1(new_n532), .C2(new_n534), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(G200), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n279), .A2(G97), .ZN(new_n542));
  INV_X1    g0342(.A(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(new_n280), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(G97), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n281), .B1(new_n429), .B2(new_n419), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n333), .A2(new_n396), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT6), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n214), .A2(new_n281), .ZN(new_n549));
  NOR2_X1   g0349(.A1(G97), .A2(G107), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n548), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n281), .A2(KEYINPUT6), .A3(G97), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n225), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NOR3_X1   g0353(.A1(new_n546), .A2(new_n547), .A3(new_n553), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n543), .B(new_n545), .C1(new_n554), .C2(new_n276), .ZN(new_n555));
  INV_X1    g0355(.A(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n535), .A2(G190), .A3(new_n538), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n541), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n530), .A2(G1698), .ZN(new_n559));
  OAI221_X1 g0359(.A(new_n559), .B1(G238), .B2(G1698), .C1(new_n250), .C2(new_n251), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n294), .A2(G33), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n261), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(G250), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n320), .B1(new_n563), .B2(KEYINPUT73), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n256), .ZN(new_n565));
  OAI211_X1 g0365(.A(KEYINPUT73), .B(G250), .C1(new_n255), .C2(G1), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n248), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  OR2_X1    g0367(.A1(new_n562), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(new_n339), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n291), .A2(new_n225), .A3(G68), .ZN(new_n570));
  INV_X1    g0370(.A(G87), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n550), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n358), .A2(new_n225), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n572), .A2(KEYINPUT19), .A3(new_n573), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n358), .A2(G20), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n570), .B(new_n574), .C1(KEYINPUT19), .C2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(new_n305), .ZN(new_n577));
  INV_X1    g0377(.A(new_n397), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n544), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n381), .A2(new_n397), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n577), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n562), .A2(new_n567), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n461), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n569), .A2(new_n581), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n582), .A2(G190), .ZN(new_n585));
  AOI22_X1  g0385(.A1(new_n576), .A2(new_n305), .B1(new_n381), .B2(new_n397), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n544), .A2(G87), .ZN(new_n587));
  OAI21_X1  g0387(.A(G200), .B1(new_n562), .B2(new_n567), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n585), .A2(new_n586), .A3(new_n587), .A4(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n584), .A2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(new_n590), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n537), .A2(new_n461), .A3(new_n538), .A4(new_n539), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n535), .A2(new_n538), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(new_n339), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n592), .A2(new_n555), .A3(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n558), .A2(new_n591), .A3(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  AND4_X1   g0397(.A1(new_n313), .A2(new_n475), .A3(new_n526), .A4(new_n597), .ZN(G372));
  INV_X1    g0398(.A(new_n584), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n304), .A2(new_n305), .ZN(new_n600));
  INV_X1    g0400(.A(new_n282), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n600), .A2(new_n601), .A3(new_n308), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n310), .A2(new_n311), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(new_n518), .ZN(new_n605));
  AND3_X1   g0405(.A1(new_n600), .A2(new_n601), .A3(new_n308), .ZN(new_n606));
  AOI22_X1  g0406(.A1(new_n604), .A2(new_n605), .B1(new_n606), .B2(new_n274), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n599), .B1(new_n607), .B2(new_n597), .ZN(new_n608));
  INV_X1    g0408(.A(new_n595), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n609), .A2(new_n591), .A3(KEYINPUT26), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT79), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n609), .A2(new_n591), .A3(KEYINPUT79), .A4(KEYINPUT26), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT26), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n614), .B1(new_n595), .B2(new_n590), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n612), .A2(new_n613), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n608), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n475), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n388), .A2(new_n473), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n619), .A2(new_n390), .A3(new_n455), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(new_n469), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n350), .A2(new_n353), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n341), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n618), .A2(new_n623), .ZN(G369));
  INV_X1    g0424(.A(G13), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n625), .A2(G20), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(new_n277), .ZN(new_n627));
  OR2_X1    g0427(.A1(new_n627), .A2(KEYINPUT27), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(KEYINPUT27), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n628), .A2(G213), .A3(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(G343), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n513), .A2(new_n632), .ZN(new_n633));
  MUX2_X1   g0433(.A(new_n518), .B(new_n526), .S(new_n633), .Z(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(G330), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n632), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n313), .B1(new_n606), .B2(new_n637), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n638), .B1(new_n604), .B2(new_n637), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n636), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n607), .A2(new_n637), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(new_n641), .ZN(G399));
  INV_X1    g0442(.A(new_n204), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n643), .A2(G41), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n572), .A2(G116), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n645), .A2(G1), .A3(new_n646), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n647), .B1(new_n229), .B2(new_n645), .ZN(new_n648));
  XNOR2_X1  g0448(.A(new_n648), .B(KEYINPUT28), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n610), .A2(new_n615), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n274), .A2(new_n306), .A3(new_n308), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n651), .B1(new_n312), .B2(new_n518), .ZN(new_n652));
  OAI211_X1 g0452(.A(new_n650), .B(new_n584), .C1(new_n652), .C2(new_n596), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT82), .ZN(new_n654));
  AND3_X1   g0454(.A1(new_n653), .A2(new_n654), .A3(new_n637), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n654), .B1(new_n653), .B2(new_n637), .ZN(new_n656));
  OAI21_X1  g0456(.A(KEYINPUT29), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n632), .B1(new_n608), .B2(new_n616), .ZN(new_n658));
  OR2_X1    g0458(.A1(new_n658), .A2(KEYINPUT29), .ZN(new_n659));
  AND3_X1   g0459(.A1(new_n497), .A2(new_n264), .A3(new_n498), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n660), .A2(G179), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n540), .A2(new_n265), .A3(new_n568), .A4(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT30), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n663), .A2(KEYINPUT80), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  AND4_X1   g0465(.A1(new_n263), .A2(new_n535), .A3(new_n582), .A4(new_n538), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n663), .A2(KEYINPUT80), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n660), .A2(G179), .A3(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n665), .B1(new_n666), .B2(new_n669), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n263), .A2(new_n535), .A3(new_n582), .A4(new_n538), .ZN(new_n671));
  NOR3_X1   g0471(.A1(new_n671), .A2(new_n664), .A3(new_n668), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n662), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT81), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  OAI211_X1 g0475(.A(KEYINPUT81), .B(new_n662), .C1(new_n670), .C2(new_n672), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n675), .A2(new_n632), .A3(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT31), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n526), .A2(new_n313), .A3(new_n597), .A4(new_n637), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n673), .A2(KEYINPUT31), .A3(new_n632), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n679), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  AOI22_X1  g0482(.A1(new_n657), .A2(new_n659), .B1(G330), .B2(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n649), .B1(new_n683), .B2(G1), .ZN(G364));
  NAND2_X1  g0484(.A1(new_n626), .A2(G45), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n645), .A2(G1), .A3(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n634), .A2(G330), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n686), .B1(new_n636), .B2(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n344), .A2(G200), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(new_n461), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(G20), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(G294), .ZN(new_n692));
  NAND2_X1  g0492(.A1(G20), .A2(G179), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT85), .ZN(new_n694));
  XNOR2_X1  g0494(.A(new_n693), .B(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n266), .A2(G190), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  XOR2_X1   g0497(.A(KEYINPUT33), .B(G317), .Z(new_n698));
  NOR2_X1   g0498(.A1(new_n344), .A2(new_n266), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n225), .A2(G179), .ZN(new_n700));
  AND2_X1   g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  OR2_X1    g0501(.A1(new_n701), .A2(KEYINPUT88), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(KEYINPUT88), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  OAI221_X1 g0504(.A(new_n692), .B1(new_n697), .B2(new_n698), .C1(new_n704), .C2(new_n493), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n695), .A2(new_n689), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n705), .B1(G322), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n695), .A2(new_n699), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  XOR2_X1   g0510(.A(KEYINPUT89), .B(G326), .Z(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(G190), .A2(G200), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n695), .A2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n291), .B1(new_n715), .B2(G311), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n700), .A2(new_n696), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n700), .A2(new_n713), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  AOI22_X1  g0520(.A1(G283), .A2(new_n718), .B1(new_n720), .B2(G329), .ZN(new_n721));
  XNOR2_X1  g0521(.A(new_n721), .B(KEYINPUT90), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n708), .A2(new_n712), .A3(new_n716), .A4(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n704), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(G87), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n691), .A2(G97), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n710), .A2(G50), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n718), .A2(G107), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n725), .A2(new_n726), .A3(new_n727), .A4(new_n728), .ZN(new_n729));
  XNOR2_X1  g0529(.A(new_n706), .B(KEYINPUT86), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n729), .B1(G58), .B2(new_n730), .ZN(new_n731));
  XOR2_X1   g0531(.A(KEYINPUT87), .B(G159), .Z(new_n732));
  NAND2_X1  g0532(.A1(new_n720), .A2(new_n732), .ZN(new_n733));
  AND2_X1   g0533(.A1(new_n733), .A2(KEYINPUT32), .ZN(new_n734));
  INV_X1    g0534(.A(new_n697), .ZN(new_n735));
  AOI211_X1 g0535(.A(new_n418), .B(new_n734), .C1(G68), .C2(new_n735), .ZN(new_n736));
  OAI211_X1 g0536(.A(new_n731), .B(new_n736), .C1(new_n396), .C2(new_n714), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n733), .A2(KEYINPUT32), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n723), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n224), .B1(G20), .B2(new_n339), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(G13), .A2(G33), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(G20), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n741), .B1(new_n634), .B2(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n744), .A2(new_n740), .ZN(new_n747));
  XOR2_X1   g0547(.A(new_n747), .B(KEYINPUT84), .Z(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n291), .A2(G355), .A3(new_n204), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n418), .A2(new_n204), .ZN(new_n751));
  XNOR2_X1  g0551(.A(new_n751), .B(KEYINPUT83), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n752), .B1(G45), .B2(new_n229), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n243), .A2(new_n255), .ZN(new_n754));
  OAI221_X1 g0554(.A(new_n750), .B1(G116), .B2(new_n204), .C1(new_n753), .C2(new_n754), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n746), .B1(new_n749), .B2(new_n755), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n688), .B1(new_n756), .B2(new_n686), .ZN(new_n757));
  XOR2_X1   g0557(.A(new_n757), .B(KEYINPUT91), .Z(G396));
  NOR2_X1   g0558(.A1(new_n740), .A2(new_n742), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n686), .B1(new_n396), .B2(new_n759), .ZN(new_n760));
  XNOR2_X1  g0560(.A(new_n760), .B(KEYINPUT92), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n473), .A2(new_n632), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n401), .A2(new_n632), .ZN(new_n764));
  AND2_X1   g0564(.A1(new_n409), .A2(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n763), .B1(new_n765), .B2(new_n474), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(G132), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n291), .B1(new_n719), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n730), .A2(G143), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n715), .A2(new_n732), .ZN(new_n771));
  AOI22_X1  g0571(.A1(G137), .A2(new_n710), .B1(new_n735), .B2(G150), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n770), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  XOR2_X1   g0573(.A(new_n773), .B(KEYINPUT34), .Z(new_n774));
  AOI211_X1 g0574(.A(new_n769), .B(new_n774), .C1(G68), .C2(new_n718), .ZN(new_n775));
  INV_X1    g0575(.A(new_n691), .ZN(new_n776));
  OAI221_X1 g0576(.A(new_n775), .B1(new_n217), .B2(new_n704), .C1(new_n212), .C2(new_n776), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n418), .B1(new_n704), .B2(new_n281), .ZN(new_n778));
  OAI22_X1  g0578(.A1(new_n493), .A2(new_n709), .B1(new_n714), .B2(new_n488), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n717), .A2(new_n571), .ZN(new_n780));
  INV_X1    g0580(.A(G311), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n726), .B1(new_n781), .B2(new_n719), .ZN(new_n782));
  NOR4_X1   g0582(.A1(new_n778), .A2(new_n779), .A3(new_n780), .A4(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(G294), .ZN(new_n784));
  OR2_X1    g0584(.A1(new_n697), .A2(KEYINPUT93), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n697), .A2(KEYINPUT93), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  XOR2_X1   g0587(.A(KEYINPUT94), .B(G283), .Z(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  OAI221_X1 g0589(.A(new_n783), .B1(new_n784), .B2(new_n706), .C1(new_n787), .C2(new_n789), .ZN(new_n790));
  AND2_X1   g0590(.A1(new_n777), .A2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n740), .ZN(new_n792));
  OAI221_X1 g0592(.A(new_n761), .B1(new_n743), .B2(new_n767), .C1(new_n791), .C2(new_n792), .ZN(new_n793));
  XNOR2_X1  g0593(.A(new_n658), .B(new_n766), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n682), .A2(G330), .ZN(new_n795));
  XOR2_X1   g0595(.A(new_n794), .B(new_n795), .Z(new_n796));
  INV_X1    g0596(.A(new_n686), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n793), .B1(new_n796), .B2(new_n797), .ZN(G384));
  INV_X1    g0598(.A(G330), .ZN(new_n799));
  NAND4_X1  g0599(.A1(new_n675), .A2(KEYINPUT31), .A3(new_n632), .A4(new_n676), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n679), .A2(new_n680), .A3(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n475), .A2(new_n801), .ZN(new_n802));
  XOR2_X1   g0602(.A(new_n802), .B(KEYINPUT98), .Z(new_n803));
  INV_X1    g0603(.A(new_n630), .ZN(new_n804));
  OAI211_X1 g0604(.A(new_n456), .B(new_n804), .C1(new_n454), .C2(new_n468), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n463), .A2(new_n630), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n456), .A2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(KEYINPUT37), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n807), .A2(new_n808), .A3(new_n451), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n808), .B1(new_n807), .B2(new_n451), .ZN(new_n811));
  OR2_X1    g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(KEYINPUT38), .B1(new_n805), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n449), .A2(new_n305), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n425), .A2(G68), .ZN(new_n815));
  AOI21_X1  g0615(.A(KEYINPUT16), .B1(new_n815), .B2(new_n443), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n412), .B1(new_n814), .B2(new_n816), .ZN(new_n817));
  OAI211_X1 g0617(.A(new_n804), .B(new_n817), .C1(new_n454), .C2(new_n468), .ZN(new_n818));
  INV_X1    g0618(.A(KEYINPUT95), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n817), .A2(new_n806), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n808), .B1(new_n820), .B2(new_n451), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n819), .B1(new_n810), .B2(new_n821), .ZN(new_n822));
  AND2_X1   g0622(.A1(new_n820), .A2(new_n451), .ZN(new_n823));
  OAI211_X1 g0623(.A(KEYINPUT95), .B(new_n809), .C1(new_n823), .C2(new_n808), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n818), .A2(new_n822), .A3(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n813), .B1(new_n826), .B2(KEYINPUT38), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n387), .A2(new_n632), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n388), .A2(new_n390), .A3(new_n828), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n372), .A2(new_n387), .A3(new_n632), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n766), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n801), .A2(new_n831), .ZN(new_n832));
  OAI21_X1  g0632(.A(KEYINPUT40), .B1(new_n827), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n832), .A2(KEYINPUT97), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT38), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n825), .A2(new_n835), .ZN(new_n836));
  NAND4_X1  g0636(.A1(new_n818), .A2(new_n824), .A3(new_n822), .A4(KEYINPUT38), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT40), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n839), .A2(KEYINPUT97), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n801), .A2(new_n831), .A3(new_n840), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n834), .A2(new_n838), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n833), .A2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n799), .B1(new_n803), .B2(new_n844), .ZN(new_n845));
  XOR2_X1   g0645(.A(new_n845), .B(KEYINPUT99), .Z(new_n846));
  OAI21_X1  g0646(.A(new_n846), .B1(new_n844), .B2(new_n803), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n762), .B1(new_n658), .B2(new_n767), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n829), .A2(new_n830), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  AOI22_X1  g0651(.A1(new_n851), .A2(new_n838), .B1(new_n468), .B2(new_n630), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n836), .A2(KEYINPUT39), .A3(new_n837), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n372), .A2(new_n387), .A3(new_n637), .ZN(new_n854));
  XOR2_X1   g0654(.A(new_n854), .B(KEYINPUT96), .Z(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  OAI211_X1 g0656(.A(new_n853), .B(new_n856), .C1(new_n827), .C2(KEYINPUT39), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n852), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n657), .A2(new_n475), .A3(new_n659), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n859), .A2(new_n623), .ZN(new_n860));
  XOR2_X1   g0660(.A(new_n858), .B(new_n860), .Z(new_n861));
  XNOR2_X1  g0661(.A(new_n847), .B(new_n861), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n862), .B1(new_n277), .B2(new_n626), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n551), .A2(new_n552), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n477), .B1(new_n864), .B2(KEYINPUT35), .ZN(new_n865));
  OAI211_X1 g0665(.A(new_n865), .B(new_n226), .C1(KEYINPUT35), .C2(new_n864), .ZN(new_n866));
  XNOR2_X1  g0666(.A(new_n866), .B(KEYINPUT36), .ZN(new_n867));
  OAI21_X1  g0667(.A(G77), .B1(new_n212), .B2(new_n373), .ZN(new_n868));
  OAI22_X1  g0668(.A1(new_n229), .A2(new_n868), .B1(G50), .B2(new_n373), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n869), .A2(G1), .A3(new_n625), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n863), .A2(new_n867), .A3(new_n870), .ZN(G367));
  OAI211_X1 g0671(.A(new_n558), .B(new_n595), .C1(new_n556), .C2(new_n637), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n872), .B1(new_n595), .B2(new_n637), .ZN(new_n873));
  XOR2_X1   g0673(.A(new_n873), .B(KEYINPUT100), .Z(new_n874));
  OR2_X1    g0674(.A1(new_n874), .A2(new_n604), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n632), .B1(new_n875), .B2(new_n595), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n605), .A2(new_n632), .ZN(new_n877));
  AND2_X1   g0677(.A1(new_n313), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(new_n873), .ZN(new_n879));
  XNOR2_X1  g0679(.A(new_n879), .B(KEYINPUT42), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT43), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n637), .B1(new_n586), .B2(new_n587), .ZN(new_n882));
  MUX2_X1   g0682(.A(new_n590), .B(new_n584), .S(new_n882), .Z(new_n883));
  OAI22_X1  g0683(.A1(new_n876), .A2(new_n880), .B1(new_n881), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n881), .ZN(new_n885));
  XOR2_X1   g0685(.A(new_n884), .B(new_n885), .Z(new_n886));
  NOR2_X1   g0686(.A1(new_n640), .A2(new_n874), .ZN(new_n887));
  XNOR2_X1  g0687(.A(new_n886), .B(new_n887), .ZN(new_n888));
  XNOR2_X1  g0688(.A(new_n644), .B(KEYINPUT41), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n878), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n891), .B1(new_n639), .B2(new_n877), .ZN(new_n892));
  XNOR2_X1  g0692(.A(new_n636), .B(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(new_n683), .ZN(new_n894));
  INV_X1    g0694(.A(new_n640), .ZN(new_n895));
  AND2_X1   g0695(.A1(new_n895), .A2(KEYINPUT102), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n641), .A2(new_n873), .ZN(new_n897));
  XOR2_X1   g0697(.A(new_n897), .B(KEYINPUT45), .Z(new_n898));
  NAND3_X1  g0698(.A1(new_n607), .A2(new_n637), .A3(new_n872), .ZN(new_n899));
  XOR2_X1   g0699(.A(KEYINPUT101), .B(KEYINPUT44), .Z(new_n900));
  XNOR2_X1  g0700(.A(new_n899), .B(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n898), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n894), .B1(new_n896), .B2(new_n902), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n903), .B1(new_n896), .B2(new_n902), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n890), .B1(new_n904), .B2(new_n683), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n685), .A2(G1), .ZN(new_n906));
  XOR2_X1   g0706(.A(new_n906), .B(KEYINPUT103), .Z(new_n907));
  OAI21_X1  g0707(.A(new_n888), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n748), .B1(new_n239), .B2(new_n752), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n578), .A2(new_n643), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n686), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  XOR2_X1   g0711(.A(new_n911), .B(KEYINPUT104), .Z(new_n912));
  INV_X1    g0712(.A(new_n787), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n732), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n707), .A2(G150), .ZN(new_n915));
  AOI22_X1  g0715(.A1(new_n724), .A2(G58), .B1(G50), .B2(new_n715), .ZN(new_n916));
  XNOR2_X1  g0716(.A(KEYINPUT106), .B(G137), .ZN(new_n917));
  AOI22_X1  g0717(.A1(G68), .A2(new_n691), .B1(new_n720), .B2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(G143), .ZN(new_n919));
  OAI211_X1 g0719(.A(new_n918), .B(new_n291), .C1(new_n919), .C2(new_n709), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n717), .A2(new_n396), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND4_X1  g0722(.A1(new_n914), .A2(new_n915), .A3(new_n916), .A4(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(KEYINPUT46), .B1(new_n724), .B2(new_n294), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n720), .A2(G317), .ZN(new_n925));
  AOI22_X1  g0725(.A1(new_n715), .A2(new_n788), .B1(G107), .B2(new_n691), .ZN(new_n926));
  OAI221_X1 g0726(.A(new_n925), .B1(new_n781), .B2(new_n709), .C1(new_n926), .C2(KEYINPUT105), .ZN(new_n927));
  AOI211_X1 g0727(.A(new_n924), .B(new_n927), .C1(G294), .C2(new_n913), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n730), .A2(G303), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n291), .B1(new_n926), .B2(KEYINPUT105), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n724), .A2(KEYINPUT46), .A3(G116), .ZN(new_n931));
  NAND4_X1  g0731(.A1(new_n928), .A2(new_n929), .A3(new_n930), .A4(new_n931), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n717), .A2(new_n214), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n923), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  XOR2_X1   g0734(.A(new_n934), .B(KEYINPUT47), .Z(new_n935));
  OAI21_X1  g0735(.A(new_n912), .B1(new_n935), .B2(new_n792), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n936), .B1(new_n744), .B2(new_n883), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n937), .B(KEYINPUT107), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n908), .A2(new_n938), .ZN(G387));
  NOR2_X1   g0739(.A1(new_n335), .A2(G50), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n940), .B(KEYINPUT50), .ZN(new_n941));
  NAND2_X1  g0741(.A1(G68), .A2(G77), .ZN(new_n942));
  NAND4_X1  g0742(.A1(new_n941), .A2(new_n255), .A3(new_n942), .A4(new_n646), .ZN(new_n943));
  INV_X1    g0743(.A(new_n752), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n944), .B1(new_n235), .B2(G45), .ZN(new_n945));
  NOR3_X1   g0745(.A1(new_n646), .A2(new_n418), .A3(new_n643), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n943), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n643), .A2(new_n281), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n748), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n776), .A2(new_n397), .ZN(new_n950));
  OAI221_X1 g0750(.A(new_n291), .B1(new_n714), .B2(new_n373), .C1(new_n217), .C2(new_n706), .ZN(new_n951));
  AOI211_X1 g0751(.A(new_n950), .B(new_n951), .C1(G150), .C2(new_n720), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n724), .A2(G77), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n710), .A2(G159), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n933), .B1(new_n735), .B2(new_n391), .ZN(new_n955));
  NAND4_X1  g0755(.A1(new_n952), .A2(new_n953), .A3(new_n954), .A4(new_n955), .ZN(new_n956));
  AOI22_X1  g0756(.A1(new_n730), .A2(G317), .B1(G322), .B2(new_n710), .ZN(new_n957));
  OAI221_X1 g0757(.A(new_n957), .B1(new_n493), .B2(new_n714), .C1(new_n781), .C2(new_n787), .ZN(new_n958));
  XOR2_X1   g0758(.A(new_n958), .B(KEYINPUT108), .Z(new_n959));
  AND2_X1   g0759(.A1(new_n959), .A2(KEYINPUT48), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n959), .A2(KEYINPUT48), .ZN(new_n961));
  OAI22_X1  g0761(.A1(new_n704), .A2(new_n784), .B1(new_n776), .B2(new_n789), .ZN(new_n962));
  NOR3_X1   g0762(.A1(new_n960), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(KEYINPUT49), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n718), .A2(new_n294), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n720), .A2(new_n711), .ZN(new_n966));
  NAND4_X1  g0766(.A1(new_n964), .A2(new_n418), .A3(new_n965), .A4(new_n966), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n963), .A2(KEYINPUT49), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n956), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  AOI211_X1 g0769(.A(new_n686), .B(new_n949), .C1(new_n969), .C2(new_n740), .ZN(new_n970));
  OR2_X1    g0770(.A1(new_n639), .A2(new_n745), .ZN(new_n971));
  AOI22_X1  g0771(.A1(new_n970), .A2(new_n971), .B1(new_n893), .B2(new_n907), .ZN(new_n972));
  INV_X1    g0772(.A(new_n894), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n644), .B1(new_n893), .B2(new_n683), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n972), .B1(new_n973), .B2(new_n974), .ZN(G393));
  AOI22_X1  g0775(.A1(G311), .A2(new_n707), .B1(new_n710), .B2(G317), .ZN(new_n976));
  XOR2_X1   g0776(.A(new_n976), .B(KEYINPUT52), .Z(new_n977));
  OAI211_X1 g0777(.A(new_n977), .B(new_n418), .C1(new_n493), .C2(new_n787), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n704), .A2(new_n789), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n776), .A2(new_n488), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n720), .A2(G322), .ZN(new_n981));
  OAI211_X1 g0781(.A(new_n728), .B(new_n981), .C1(new_n714), .C2(new_n784), .ZN(new_n982));
  NOR4_X1   g0782(.A1(new_n978), .A2(new_n979), .A3(new_n980), .A4(new_n982), .ZN(new_n983));
  AOI22_X1  g0783(.A1(new_n691), .A2(G77), .B1(new_n720), .B2(G143), .ZN(new_n984));
  OAI211_X1 g0784(.A(new_n291), .B(new_n984), .C1(new_n704), .C2(new_n373), .ZN(new_n985));
  INV_X1    g0785(.A(G159), .ZN(new_n986));
  OAI22_X1  g0786(.A1(new_n331), .A2(new_n709), .B1(new_n706), .B2(new_n986), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT51), .ZN(new_n988));
  OAI221_X1 g0788(.A(new_n988), .B1(new_n571), .B2(new_n717), .C1(new_n335), .C2(new_n714), .ZN(new_n989));
  AOI211_X1 g0789(.A(new_n985), .B(new_n989), .C1(G50), .C2(new_n913), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n740), .B1(new_n983), .B2(new_n990), .ZN(new_n991));
  OAI221_X1 g0791(.A(new_n749), .B1(new_n214), .B2(new_n204), .C1(new_n246), .C2(new_n944), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n991), .A2(new_n797), .A3(new_n992), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n993), .B1(new_n874), .B2(new_n744), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n902), .B1(new_n895), .B2(KEYINPUT109), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n895), .A2(KEYINPUT109), .ZN(new_n996));
  XOR2_X1   g0796(.A(new_n995), .B(new_n996), .Z(new_n997));
  AOI21_X1  g0797(.A(new_n994), .B1(new_n997), .B2(new_n907), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n904), .B1(new_n997), .B2(new_n973), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n998), .B1(new_n999), .B2(new_n645), .ZN(G390));
  AND3_X1   g0800(.A1(new_n836), .A2(KEYINPUT39), .A3(new_n837), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n813), .ZN(new_n1002));
  AOI21_X1  g0802(.A(KEYINPUT39), .B1(new_n1002), .B2(new_n837), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n742), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n759), .A2(new_n335), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n418), .B1(new_n719), .B2(new_n784), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n710), .A2(G283), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n725), .A2(new_n1007), .ZN(new_n1008));
  AOI211_X1 g0808(.A(new_n1006), .B(new_n1008), .C1(G68), .C2(new_n718), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n715), .A2(G97), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(new_n913), .A2(G107), .B1(G77), .B2(new_n691), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1009), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1012), .B1(G116), .B2(new_n707), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n776), .A2(new_n986), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n724), .A2(G150), .ZN(new_n1015));
  OR2_X1    g0815(.A1(new_n1015), .A2(KEYINPUT53), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n1015), .A2(KEYINPUT53), .B1(G132), .B2(new_n707), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n913), .A2(new_n917), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n291), .B1(new_n717), .B2(new_n217), .ZN(new_n1019));
  INV_X1    g0819(.A(G128), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n709), .A2(new_n1020), .ZN(new_n1021));
  AOI211_X1 g0821(.A(new_n1019), .B(new_n1021), .C1(G125), .C2(new_n720), .ZN(new_n1022));
  NAND4_X1  g0822(.A1(new_n1016), .A2(new_n1017), .A3(new_n1018), .A4(new_n1022), .ZN(new_n1023));
  XOR2_X1   g0823(.A(KEYINPUT54), .B(G143), .Z(new_n1024));
  AOI211_X1 g0824(.A(new_n1014), .B(new_n1023), .C1(new_n715), .C2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n740), .B1(new_n1013), .B2(new_n1025), .ZN(new_n1026));
  NAND4_X1  g0826(.A1(new_n1004), .A2(new_n797), .A3(new_n1005), .A4(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT112), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n653), .A2(new_n637), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1029), .A2(KEYINPUT82), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n653), .A2(new_n654), .A3(new_n637), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1030), .A2(new_n1031), .A3(new_n763), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT110), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n849), .B(new_n1033), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n765), .A2(new_n474), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n1035), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1032), .A2(new_n1034), .A3(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1002), .A2(new_n837), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1037), .A2(new_n1038), .A3(new_n855), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n855), .B1(new_n848), .B2(new_n850), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1040), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1041));
  NAND4_X1  g0841(.A1(new_n682), .A2(G330), .A3(new_n767), .A4(new_n849), .ZN(new_n1042));
  AND3_X1   g0842(.A1(new_n1039), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n832), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1044), .A2(G330), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1045), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n1043), .A2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1028), .B1(new_n1047), .B2(new_n907), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n1045), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1039), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1052));
  AND4_X1   g0852(.A1(new_n1028), .A2(new_n1051), .A3(new_n907), .A4(new_n1052), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1027), .B1(new_n1048), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT113), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n850), .B1(new_n795), .B2(new_n766), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1045), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n848), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1032), .A2(new_n1036), .ZN(new_n1061));
  AND3_X1   g0861(.A1(new_n801), .A2(G330), .A3(new_n767), .ZN(new_n1062));
  OAI211_X1 g0862(.A(new_n1061), .B(new_n1042), .C1(new_n1034), .C2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1060), .A2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n475), .A2(G330), .A3(new_n801), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n859), .A2(new_n623), .A3(new_n1065), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1064), .A2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1068), .B1(new_n1043), .B2(new_n1046), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1066), .B1(new_n1060), .B2(new_n1063), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1051), .A2(new_n1070), .A3(new_n1052), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1069), .A2(new_n644), .A3(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(KEYINPUT111), .ZN(new_n1073));
  INV_X1    g0873(.A(KEYINPUT111), .ZN(new_n1074));
  NAND4_X1  g0874(.A1(new_n1069), .A2(new_n1071), .A3(new_n1074), .A4(new_n644), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1076));
  OAI211_X1 g0876(.A(KEYINPUT113), .B(new_n1027), .C1(new_n1048), .C2(new_n1053), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1056), .A2(new_n1076), .A3(new_n1077), .ZN(G378));
  OAI21_X1  g0878(.A(new_n217), .B1(new_n250), .B2(G41), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(G132), .A2(new_n735), .B1(new_n715), .B2(G137), .ZN(new_n1080));
  XOR2_X1   g0880(.A(new_n1080), .B(KEYINPUT115), .Z(new_n1081));
  NAND2_X1  g0881(.A1(new_n724), .A2(new_n1024), .ZN(new_n1082));
  OAI211_X1 g0882(.A(new_n1081), .B(new_n1082), .C1(new_n331), .C2(new_n776), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(G125), .B2(new_n710), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1084), .B1(new_n1020), .B2(new_n706), .ZN(new_n1085));
  AOI21_X1  g0885(.A(G41), .B1(new_n1085), .B2(KEYINPUT59), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n718), .A2(new_n732), .ZN(new_n1087));
  AOI21_X1  g0887(.A(G33), .B1(new_n720), .B2(G124), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1086), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n1085), .A2(KEYINPUT59), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1079), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n707), .A2(G107), .ZN(new_n1092));
  XOR2_X1   g0892(.A(new_n1092), .B(KEYINPUT114), .Z(new_n1093));
  OAI22_X1  g0893(.A1(new_n697), .A2(new_n214), .B1(new_n212), .B2(new_n717), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n715), .A2(new_n578), .B1(G68), .B2(new_n691), .ZN(new_n1096));
  INV_X1    g0896(.A(G283), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n418), .B1(new_n719), .B2(new_n1097), .ZN(new_n1098));
  AOI211_X1 g0898(.A(G41), .B(new_n1098), .C1(new_n710), .C2(G116), .ZN(new_n1099));
  NAND4_X1  g0899(.A1(new_n1095), .A2(new_n953), .A3(new_n1096), .A4(new_n1099), .ZN(new_n1100));
  XOR2_X1   g0900(.A(new_n1100), .B(KEYINPUT58), .Z(new_n1101));
  OAI21_X1  g0901(.A(new_n740), .B1(new_n1091), .B2(new_n1101), .ZN(new_n1102));
  XOR2_X1   g0902(.A(new_n1102), .B(KEYINPUT116), .Z(new_n1103));
  INV_X1    g0903(.A(new_n759), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n1104), .A2(G50), .ZN(new_n1105));
  XOR2_X1   g0905(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1106));
  AND2_X1   g0906(.A1(new_n350), .A2(new_n353), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1106), .B1(new_n1107), .B2(new_n341), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n338), .A2(new_n804), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1106), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n354), .A2(new_n1111), .ZN(new_n1112));
  AND3_X1   g0912(.A1(new_n1108), .A2(new_n1110), .A3(new_n1112), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1110), .B1(new_n1108), .B2(new_n1112), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n797), .B1(new_n1115), .B2(new_n743), .ZN(new_n1116));
  OR3_X1    g0916(.A1(new_n1103), .A2(new_n1105), .A3(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1071), .A2(new_n1067), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n858), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1115), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1121), .B1(new_n843), .B2(G330), .ZN(new_n1122));
  AOI211_X1 g0922(.A(new_n799), .B(new_n1115), .C1(new_n833), .C2(new_n842), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1120), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  AND3_X1   g0924(.A1(new_n834), .A2(new_n838), .A3(new_n841), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n839), .B1(new_n1038), .B2(new_n1044), .ZN(new_n1126));
  OAI21_X1  g0926(.A(G330), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1127), .A2(new_n1115), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n843), .A2(G330), .A3(new_n1121), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1128), .A2(new_n858), .A3(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1124), .A2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1119), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT57), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n645), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1124), .A2(new_n1130), .A3(KEYINPUT117), .ZN(new_n1135));
  INV_X1    g0935(.A(KEYINPUT117), .ZN(new_n1136));
  NAND4_X1  g0936(.A1(new_n1128), .A2(new_n1136), .A3(new_n858), .A4(new_n1129), .ZN(new_n1137));
  NAND4_X1  g0937(.A1(new_n1135), .A2(new_n1119), .A3(KEYINPUT57), .A4(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1118), .B1(new_n1134), .B2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1131), .A2(new_n907), .ZN(new_n1140));
  AND2_X1   g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(G375));
  NOR2_X1   g0942(.A1(new_n1034), .A2(new_n743), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n1104), .A2(G68), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n709), .A2(new_n784), .ZN(new_n1145));
  AOI211_X1 g0945(.A(new_n1145), .B(new_n950), .C1(G283), .C2(new_n707), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n291), .B1(new_n720), .B2(G303), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n921), .B1(new_n724), .B2(G97), .ZN(new_n1148));
  AND3_X1   g0948(.A1(new_n1146), .A2(new_n1147), .A3(new_n1148), .ZN(new_n1149));
  OAI221_X1 g0949(.A(new_n1149), .B1(new_n281), .B2(new_n714), .C1(new_n488), .C2(new_n787), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n291), .B1(new_n776), .B2(new_n217), .ZN(new_n1151));
  OAI22_X1  g0951(.A1(new_n704), .A2(new_n986), .B1(new_n212), .B2(new_n717), .ZN(new_n1152));
  AOI211_X1 g0952(.A(new_n1151), .B(new_n1152), .C1(G132), .C2(new_n710), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n730), .A2(new_n917), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n720), .A2(G128), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(new_n913), .A2(new_n1024), .B1(G150), .B2(new_n715), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n1153), .A2(new_n1154), .A3(new_n1155), .A4(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n792), .B1(new_n1150), .B2(new_n1157), .ZN(new_n1158));
  NOR4_X1   g0958(.A1(new_n1143), .A2(new_n686), .A3(new_n1144), .A4(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1159), .B1(new_n1064), .B2(new_n907), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1060), .A2(new_n1063), .A3(new_n1066), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1161), .A2(new_n889), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1160), .B1(new_n1162), .B2(new_n1070), .ZN(G381));
  NAND3_X1  g0963(.A1(new_n1056), .A2(new_n1077), .A3(new_n1072), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(G375), .A2(new_n1164), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(G387), .A2(G381), .ZN(new_n1166));
  NOR4_X1   g0966(.A1(G390), .A2(G396), .A3(G393), .A4(G384), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1165), .A2(new_n1166), .A3(new_n1167), .ZN(G407));
  NAND2_X1  g0968(.A1(new_n631), .A2(G213), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(new_n1169), .B(KEYINPUT118), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1165), .A2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(G407), .A2(G213), .A3(new_n1171), .ZN(G409));
  INV_X1    g0972(.A(KEYINPUT125), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT120), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1161), .A2(new_n1174), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n644), .B(new_n1068), .C1(new_n1175), .C2(KEYINPUT60), .ZN(new_n1176));
  AND2_X1   g0976(.A1(new_n1175), .A2(KEYINPUT60), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1160), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(new_n1178), .B(G384), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1135), .A2(new_n907), .A3(new_n1137), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1181), .A2(new_n1117), .ZN(new_n1182));
  INV_X1    g0982(.A(KEYINPUT119), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1119), .A2(new_n1131), .A3(new_n889), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1181), .A2(KEYINPUT119), .A3(new_n1117), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1184), .A2(new_n1185), .A3(new_n1186), .ZN(new_n1187));
  AND3_X1   g0987(.A1(new_n1056), .A2(new_n1077), .A3(new_n1072), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1139), .A2(G378), .A3(new_n1140), .ZN(new_n1190));
  AOI211_X1 g0990(.A(new_n1170), .B(new_n1180), .C1(new_n1189), .C2(new_n1190), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1173), .B1(new_n1191), .B2(KEYINPUT62), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1170), .ZN(new_n1194));
  NAND4_X1  g0994(.A1(new_n1193), .A2(KEYINPUT62), .A3(new_n1194), .A4(new_n1179), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT126), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1170), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1198));
  NAND4_X1  g0998(.A1(new_n1198), .A2(KEYINPUT126), .A3(KEYINPUT62), .A4(new_n1179), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1186), .ZN(new_n1200));
  AOI21_X1  g1000(.A(KEYINPUT119), .B1(new_n1181), .B2(new_n1117), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1164), .B1(new_n1202), .B2(new_n1185), .ZN(new_n1203));
  AND3_X1   g1003(.A1(new_n1139), .A2(G378), .A3(new_n1140), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n1194), .B(new_n1179), .C1(new_n1203), .C2(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(KEYINPUT62), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1205), .A2(KEYINPUT125), .A3(new_n1206), .ZN(new_n1207));
  NAND4_X1  g1007(.A1(new_n1192), .A2(new_n1197), .A3(new_n1199), .A4(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1198), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1170), .A2(G2897), .ZN(new_n1210));
  XOR2_X1   g1010(.A(new_n1179), .B(new_n1210), .Z(new_n1211));
  AOI21_X1  g1011(.A(KEYINPUT61), .B1(new_n1209), .B2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1208), .A2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1213), .A2(KEYINPUT127), .ZN(new_n1214));
  XOR2_X1   g1014(.A(G393), .B(G396), .Z(new_n1215));
  NAND3_X1  g1015(.A1(new_n908), .A2(new_n938), .A3(G390), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(G390), .B1(new_n908), .B2(new_n938), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1215), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1219), .A2(KEYINPUT122), .ZN(new_n1220));
  INV_X1    g1020(.A(KEYINPUT122), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n1221), .B(new_n1215), .C1(new_n1217), .C2(new_n1218), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT123), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1218), .B1(new_n1217), .B2(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1215), .B1(new_n1216), .B2(KEYINPUT123), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(new_n1220), .A2(new_n1222), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT127), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1208), .A2(new_n1227), .A3(new_n1212), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1214), .A2(new_n1226), .A3(new_n1228), .ZN(new_n1229));
  XNOR2_X1  g1029(.A(new_n1205), .B(KEYINPUT63), .ZN(new_n1230));
  XNOR2_X1  g1030(.A(new_n1211), .B(KEYINPUT121), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1231), .A2(new_n1209), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1220), .A2(new_n1222), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT61), .ZN(new_n1236));
  AOI21_X1  g1036(.A(KEYINPUT124), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT124), .ZN(new_n1238));
  NOR3_X1   g1038(.A1(new_n1226), .A2(new_n1238), .A3(KEYINPUT61), .ZN(new_n1239));
  OAI211_X1 g1039(.A(new_n1230), .B(new_n1232), .C1(new_n1237), .C2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1229), .A2(new_n1240), .ZN(G405));
  OAI21_X1  g1041(.A(new_n1190), .B1(new_n1141), .B2(new_n1164), .ZN(new_n1242));
  XNOR2_X1  g1042(.A(new_n1242), .B(new_n1179), .ZN(new_n1243));
  XNOR2_X1  g1043(.A(new_n1226), .B(new_n1243), .ZN(G402));
endmodule


