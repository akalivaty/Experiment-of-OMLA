

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785;

  XNOR2_X2 U374 ( .A(n569), .B(n568), .ZN(n732) );
  BUF_X4 U375 ( .A(n606), .Z(n353) );
  XNOR2_X1 U376 ( .A(n538), .B(n537), .ZN(n541) );
  INV_X1 U377 ( .A(G953), .ZN(n778) );
  NOR2_X1 U378 ( .A1(n714), .A2(n648), .ZN(n649) );
  XNOR2_X1 U379 ( .A(n420), .B(KEYINPUT66), .ZN(n597) );
  NAND2_X1 U380 ( .A1(n541), .A2(n735), .ZN(n373) );
  INV_X1 U381 ( .A(G143), .ZN(n447) );
  XNOR2_X1 U382 ( .A(n656), .B(KEYINPUT85), .ZN(n408) );
  AND2_X1 U383 ( .A1(n388), .A2(n387), .ZN(n386) );
  AND2_X1 U384 ( .A1(n406), .A2(KEYINPUT45), .ZN(n355) );
  AND2_X1 U385 ( .A1(n413), .A2(n411), .ZN(n410) );
  XNOR2_X1 U386 ( .A(n580), .B(KEYINPUT32), .ZN(n602) );
  INV_X1 U387 ( .A(n734), .ZN(n404) );
  XNOR2_X1 U388 ( .A(n458), .B(n435), .ZN(n621) );
  XNOR2_X1 U389 ( .A(n494), .B(n493), .ZN(n722) );
  XNOR2_X1 U390 ( .A(n474), .B(n455), .ZN(n659) );
  XNOR2_X1 U391 ( .A(n524), .B(n441), .ZN(n497) );
  XNOR2_X1 U392 ( .A(n447), .B(G128), .ZN(n524) );
  XNOR2_X1 U393 ( .A(KEYINPUT18), .B(KEYINPUT81), .ZN(n522) );
  INV_X1 U394 ( .A(n757), .ZN(n354) );
  NAND2_X1 U395 ( .A1(n386), .A2(n383), .ZN(n756) );
  XNOR2_X2 U396 ( .A(n353), .B(n555), .ZN(n590) );
  XNOR2_X2 U397 ( .A(n373), .B(KEYINPUT89), .ZN(n626) );
  XNOR2_X2 U398 ( .A(n497), .B(n437), .ZN(n772) );
  XNOR2_X1 U399 ( .A(n614), .B(n613), .ZN(n736) );
  AND2_X1 U400 ( .A1(n620), .A2(n736), .ZN(n436) );
  NAND2_X1 U401 ( .A1(n416), .A2(n722), .ZN(n607) );
  NOR2_X1 U402 ( .A1(n556), .A2(n723), .ZN(n416) );
  NAND2_X1 U403 ( .A1(n535), .A2(G214), .ZN(n735) );
  XNOR2_X1 U404 ( .A(KEYINPUT15), .B(G902), .ZN(n651) );
  XNOR2_X1 U405 ( .A(G116), .B(G113), .ZN(n449) );
  XNOR2_X1 U406 ( .A(n391), .B(n365), .ZN(n643) );
  NOR2_X1 U407 ( .A1(G953), .A2(G237), .ZN(n514) );
  XNOR2_X1 U408 ( .A(n418), .B(n417), .ZN(n499) );
  INV_X1 U409 ( .A(KEYINPUT8), .ZN(n417) );
  NAND2_X1 U410 ( .A1(n778), .A2(G234), .ZN(n418) );
  XNOR2_X1 U411 ( .A(G113), .B(G143), .ZN(n510) );
  INV_X1 U412 ( .A(n654), .ZN(n423) );
  INV_X1 U413 ( .A(n425), .ZN(n377) );
  NAND2_X1 U414 ( .A1(n643), .A2(n645), .ZN(n381) );
  INV_X1 U415 ( .A(G237), .ZN(n457) );
  XNOR2_X1 U416 ( .A(KEYINPUT10), .B(G140), .ZN(n479) );
  INV_X1 U417 ( .A(G134), .ZN(n441) );
  XNOR2_X1 U418 ( .A(n498), .B(n356), .ZN(n445) );
  NAND2_X1 U419 ( .A1(n362), .A2(n392), .ZN(n747) );
  NOR2_X1 U420 ( .A1(n738), .A2(n394), .ZN(n393) );
  AND2_X1 U421 ( .A1(n621), .A2(n622), .ZN(n429) );
  XNOR2_X1 U422 ( .A(n415), .B(n610), .ZN(n612) );
  XNOR2_X1 U423 ( .A(n609), .B(KEYINPUT111), .ZN(n610) );
  NOR2_X1 U424 ( .A1(n608), .A2(n607), .ZN(n415) );
  XNOR2_X1 U425 ( .A(n505), .B(n504), .ZN(n589) );
  XNOR2_X1 U426 ( .A(n587), .B(n366), .ZN(n402) );
  XNOR2_X1 U427 ( .A(n584), .B(KEYINPUT98), .ZN(n401) );
  NOR2_X1 U428 ( .A1(n639), .A2(n412), .ZN(n411) );
  INV_X1 U429 ( .A(n640), .ZN(n412) );
  AND2_X1 U430 ( .A1(n635), .A2(n704), .ZN(n636) );
  XNOR2_X1 U431 ( .A(n440), .B(G131), .ZN(n509) );
  INV_X1 U432 ( .A(KEYINPUT67), .ZN(n440) );
  INV_X1 U433 ( .A(KEYINPUT41), .ZN(n398) );
  XNOR2_X1 U434 ( .A(G101), .B(KEYINPUT69), .ZN(n448) );
  XNOR2_X1 U435 ( .A(n509), .B(n438), .ZN(n437) );
  XNOR2_X1 U436 ( .A(n439), .B(G137), .ZN(n438) );
  INV_X1 U437 ( .A(KEYINPUT4), .ZN(n439) );
  NOR2_X1 U438 ( .A1(n422), .A2(n368), .ZN(n421) );
  XNOR2_X1 U439 ( .A(KEYINPUT4), .B(KEYINPUT17), .ZN(n527) );
  NAND2_X1 U440 ( .A1(G234), .A2(G237), .ZN(n459) );
  NAND2_X1 U441 ( .A1(n735), .A2(n398), .ZN(n394) );
  OR2_X1 U442 ( .A1(n736), .A2(n398), .ZN(n397) );
  NAND2_X1 U443 ( .A1(n396), .A2(KEYINPUT41), .ZN(n395) );
  NAND2_X1 U444 ( .A1(n615), .A2(n735), .ZN(n396) );
  INV_X1 U445 ( .A(G902), .ZN(n519) );
  XNOR2_X1 U446 ( .A(G107), .B(G104), .ZN(n468) );
  XNOR2_X1 U447 ( .A(G119), .B(G128), .ZN(n481) );
  XNOR2_X1 U448 ( .A(n518), .B(n517), .ZN(n666) );
  XNOR2_X1 U449 ( .A(n516), .B(n515), .ZN(n517) );
  NOR2_X1 U450 ( .A1(n378), .A2(n377), .ZN(n376) );
  NAND2_X1 U451 ( .A1(n381), .A2(n358), .ZN(n378) );
  NAND2_X1 U452 ( .A1(n385), .A2(n384), .ZN(n383) );
  XNOR2_X1 U453 ( .A(n560), .B(KEYINPUT110), .ZN(n625) );
  NOR2_X1 U454 ( .A1(n623), .A2(n607), .ZN(n559) );
  AND2_X1 U455 ( .A1(n433), .A2(n431), .ZN(n430) );
  OR2_X1 U456 ( .A1(n436), .A2(n622), .ZN(n433) );
  XOR2_X1 U457 ( .A(n570), .B(KEYINPUT34), .Z(n571) );
  INV_X1 U458 ( .A(KEYINPUT30), .ZN(n435) );
  XNOR2_X1 U459 ( .A(n626), .B(n443), .ZN(n547) );
  INV_X1 U460 ( .A(KEYINPUT19), .ZN(n443) );
  XNOR2_X1 U461 ( .A(n659), .B(KEYINPUT62), .ZN(n660) );
  XNOR2_X1 U462 ( .A(n503), .B(n444), .ZN(n687) );
  XNOR2_X1 U463 ( .A(n497), .B(n445), .ZN(n444) );
  XOR2_X1 U464 ( .A(n666), .B(KEYINPUT59), .Z(n667) );
  XNOR2_X1 U465 ( .A(n673), .B(n675), .ZN(n676) );
  XNOR2_X1 U466 ( .A(n619), .B(n618), .ZN(n784) );
  OR2_X1 U467 ( .A1(n402), .A2(n623), .ZN(n709) );
  OR2_X1 U468 ( .A1(n401), .A2(n623), .ZN(n697) );
  NAND2_X1 U469 ( .A1(n589), .A2(n588), .ZN(n623) );
  XOR2_X1 U470 ( .A(KEYINPUT104), .B(KEYINPUT9), .Z(n356) );
  XNOR2_X1 U471 ( .A(n521), .B(n520), .ZN(n557) );
  XNOR2_X1 U472 ( .A(n552), .B(n551), .ZN(n593) );
  XOR2_X1 U473 ( .A(n369), .B(KEYINPUT78), .Z(n357) );
  AND2_X1 U474 ( .A1(n649), .A2(KEYINPUT2), .ZN(n358) );
  AND2_X1 U475 ( .A1(n605), .A2(KEYINPUT45), .ZN(n359) );
  AND2_X1 U476 ( .A1(n407), .A2(n421), .ZN(n360) );
  AND2_X1 U477 ( .A1(n428), .A2(n708), .ZN(n361) );
  AND2_X1 U478 ( .A1(n397), .A2(n395), .ZN(n362) );
  AND2_X1 U479 ( .A1(n602), .A2(n600), .ZN(n363) );
  AND2_X1 U480 ( .A1(n615), .A2(n550), .ZN(n364) );
  XOR2_X1 U481 ( .A(KEYINPUT46), .B(KEYINPUT87), .Z(n365) );
  NOR2_X1 U482 ( .A1(n634), .A2(n382), .ZN(n704) );
  XNOR2_X1 U483 ( .A(KEYINPUT99), .B(KEYINPUT31), .ZN(n366) );
  XOR2_X1 U484 ( .A(n548), .B(KEYINPUT0), .Z(n367) );
  INV_X1 U485 ( .A(n622), .ZN(n434) );
  INV_X1 U486 ( .A(KEYINPUT45), .ZN(n389) );
  NOR2_X1 U487 ( .A1(n655), .A2(KEYINPUT65), .ZN(n368) );
  INV_X1 U488 ( .A(n623), .ZN(n708) );
  NAND2_X1 U489 ( .A1(n354), .A2(n408), .ZN(n369) );
  NAND2_X1 U490 ( .A1(n756), .A2(n408), .ZN(n374) );
  XNOR2_X1 U491 ( .A(n374), .B(KEYINPUT78), .ZN(n715) );
  NAND2_X1 U492 ( .A1(n405), .A2(n406), .ZN(n370) );
  NAND2_X1 U493 ( .A1(n355), .A2(n405), .ZN(n388) );
  AND2_X1 U494 ( .A1(n370), .A2(n389), .ZN(n385) );
  XNOR2_X2 U495 ( .A(n371), .B(n575), .ZN(n420) );
  NAND2_X1 U496 ( .A1(n372), .A2(n574), .ZN(n371) );
  XNOR2_X1 U497 ( .A(n572), .B(n571), .ZN(n372) );
  NAND2_X1 U498 ( .A1(n547), .A2(n446), .ZN(n549) );
  INV_X1 U499 ( .A(n696), .ZN(n442) );
  NAND2_X1 U500 ( .A1(n375), .A2(n363), .ZN(n399) );
  INV_X1 U501 ( .A(n597), .ZN(n375) );
  NAND2_X1 U502 ( .A1(n390), .A2(n359), .ZN(n387) );
  OR2_X1 U503 ( .A1(n402), .A2(n646), .ZN(n711) );
  OR2_X1 U504 ( .A1(n401), .A2(n646), .ZN(n700) );
  NAND2_X1 U505 ( .A1(n381), .A2(n649), .ZN(n380) );
  NAND2_X1 U506 ( .A1(n376), .A2(n409), .ZN(n656) );
  NOR2_X1 U507 ( .A1(n380), .A2(n379), .ZN(n775) );
  NAND2_X1 U508 ( .A1(n409), .A2(n425), .ZN(n379) );
  INV_X1 U509 ( .A(n547), .ZN(n382) );
  NAND2_X1 U510 ( .A1(n390), .A2(n605), .ZN(n384) );
  NAND2_X1 U511 ( .A1(n399), .A2(n598), .ZN(n390) );
  NAND2_X1 U512 ( .A1(n581), .A2(n732), .ZN(n572) );
  XNOR2_X2 U513 ( .A(n549), .B(n367), .ZN(n581) );
  BUF_X2 U514 ( .A(n689), .Z(n685) );
  NAND2_X1 U515 ( .A1(n782), .A2(n784), .ZN(n391) );
  NAND2_X1 U516 ( .A1(n736), .A2(n735), .ZN(n733) );
  NAND2_X1 U517 ( .A1(n736), .A2(n393), .ZN(n392) );
  NAND2_X1 U518 ( .A1(n400), .A2(n404), .ZN(n403) );
  NAND2_X1 U519 ( .A1(n402), .A2(n401), .ZN(n400) );
  NAND2_X1 U520 ( .A1(n403), .A2(n442), .ZN(n596) );
  OR2_X1 U521 ( .A1(n596), .A2(n595), .ZN(n405) );
  NAND2_X1 U522 ( .A1(n594), .A2(n597), .ZN(n406) );
  NAND2_X1 U523 ( .A1(n360), .A2(n715), .ZN(n658) );
  NAND2_X1 U524 ( .A1(n424), .A2(n423), .ZN(n407) );
  NAND2_X1 U525 ( .A1(n426), .A2(n427), .ZN(n409) );
  NAND2_X1 U526 ( .A1(n641), .A2(n410), .ZN(n642) );
  XNOR2_X1 U527 ( .A(n636), .B(n414), .ZN(n413) );
  INV_X1 U528 ( .A(KEYINPUT74), .ZN(n414) );
  NAND2_X1 U529 ( .A1(n420), .A2(KEYINPUT88), .ZN(n604) );
  XNOR2_X1 U530 ( .A(n420), .B(n419), .ZN(G24) );
  INV_X1 U531 ( .A(G122), .ZN(n419) );
  AND2_X1 U532 ( .A1(n354), .A2(n775), .ZN(n716) );
  NOR2_X1 U533 ( .A1(n775), .A2(n654), .ZN(n422) );
  INV_X1 U534 ( .A(n756), .ZN(n424) );
  NAND2_X1 U535 ( .A1(n642), .A2(n645), .ZN(n425) );
  NOR2_X1 U536 ( .A1(n642), .A2(n645), .ZN(n426) );
  INV_X1 U537 ( .A(n643), .ZN(n427) );
  NAND2_X1 U538 ( .A1(n430), .A2(n428), .ZN(n647) );
  NAND2_X1 U539 ( .A1(n361), .A2(n430), .ZN(n624) );
  NAND2_X1 U540 ( .A1(n436), .A2(n429), .ZN(n428) );
  NAND2_X1 U541 ( .A1(n432), .A2(n434), .ZN(n431) );
  INV_X1 U542 ( .A(n621), .ZN(n432) );
  NAND2_X1 U543 ( .A1(n581), .A2(n364), .ZN(n552) );
  NOR2_X1 U544 ( .A1(n596), .A2(n598), .ZN(n594) );
  INV_X1 U545 ( .A(n589), .ZN(n558) );
  BUF_X1 U546 ( .A(n581), .Z(n586) );
  XOR2_X1 U547 ( .A(n546), .B(n545), .Z(n446) );
  XNOR2_X1 U548 ( .A(n611), .B(KEYINPUT1), .ZN(n566) );
  BUF_X1 U549 ( .A(n566), .Z(n718) );
  XNOR2_X2 U550 ( .A(n772), .B(G146), .ZN(n474) );
  XNOR2_X1 U551 ( .A(n449), .B(n448), .ZN(n451) );
  XNOR2_X1 U552 ( .A(KEYINPUT3), .B(G119), .ZN(n450) );
  XNOR2_X1 U553 ( .A(n451), .B(n450), .ZN(n533) );
  XOR2_X1 U554 ( .A(KEYINPUT5), .B(KEYINPUT76), .Z(n453) );
  NAND2_X1 U555 ( .A1(n514), .A2(G210), .ZN(n452) );
  XNOR2_X1 U556 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U557 ( .A(n533), .B(n454), .ZN(n455) );
  NAND2_X1 U558 ( .A1(n659), .A2(n519), .ZN(n456) );
  XNOR2_X2 U559 ( .A(n456), .B(G472), .ZN(n606) );
  NAND2_X1 U560 ( .A1(n519), .A2(n457), .ZN(n535) );
  NAND2_X1 U561 ( .A1(n353), .A2(n735), .ZN(n458) );
  XNOR2_X1 U562 ( .A(n459), .B(KEYINPUT94), .ZN(n460) );
  XNOR2_X1 U563 ( .A(KEYINPUT14), .B(n460), .ZN(n462) );
  NAND2_X1 U564 ( .A1(n462), .A2(G952), .ZN(n461) );
  XOR2_X1 U565 ( .A(KEYINPUT95), .B(n461), .Z(n746) );
  NOR2_X1 U566 ( .A1(G953), .A2(n746), .ZN(n544) );
  AND2_X1 U567 ( .A1(n462), .A2(G953), .ZN(n463) );
  NAND2_X1 U568 ( .A1(G902), .A2(n463), .ZN(n542) );
  XNOR2_X1 U569 ( .A(n542), .B(KEYINPUT108), .ZN(n464) );
  NOR2_X1 U570 ( .A1(G900), .A2(n464), .ZN(n465) );
  XOR2_X1 U571 ( .A(KEYINPUT109), .B(n465), .Z(n466) );
  NOR2_X1 U572 ( .A1(n544), .A2(n466), .ZN(n556) );
  XNOR2_X1 U573 ( .A(KEYINPUT77), .B(G110), .ZN(n467) );
  XNOR2_X1 U574 ( .A(n468), .B(n467), .ZN(n764) );
  XNOR2_X1 U575 ( .A(n764), .B(KEYINPUT70), .ZN(n530) );
  NAND2_X1 U576 ( .A1(G227), .A2(n778), .ZN(n469) );
  XNOR2_X1 U577 ( .A(n469), .B(G140), .ZN(n471) );
  XNOR2_X1 U578 ( .A(G101), .B(KEYINPUT80), .ZN(n470) );
  XNOR2_X1 U579 ( .A(n471), .B(n470), .ZN(n472) );
  XNOR2_X1 U580 ( .A(n530), .B(n472), .ZN(n473) );
  XNOR2_X1 U581 ( .A(n474), .B(n473), .ZN(n691) );
  NAND2_X1 U582 ( .A1(n691), .A2(n519), .ZN(n475) );
  XNOR2_X2 U583 ( .A(n475), .B(G469), .ZN(n611) );
  NAND2_X1 U584 ( .A1(n651), .A2(G234), .ZN(n476) );
  XNOR2_X1 U585 ( .A(n476), .B(KEYINPUT20), .ZN(n488) );
  AND2_X1 U586 ( .A1(n488), .A2(G221), .ZN(n478) );
  INV_X1 U587 ( .A(KEYINPUT21), .ZN(n477) );
  XNOR2_X1 U588 ( .A(n478), .B(n477), .ZN(n723) );
  XNOR2_X2 U589 ( .A(G146), .B(G125), .ZN(n523) );
  BUF_X1 U590 ( .A(n523), .Z(n480) );
  XNOR2_X1 U591 ( .A(n480), .B(n479), .ZN(n771) );
  XOR2_X1 U592 ( .A(G110), .B(G137), .Z(n482) );
  XNOR2_X1 U593 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U594 ( .A(n771), .B(n483), .ZN(n487) );
  NAND2_X1 U595 ( .A1(G221), .A2(n499), .ZN(n485) );
  XNOR2_X1 U596 ( .A(KEYINPUT23), .B(KEYINPUT24), .ZN(n484) );
  XNOR2_X1 U597 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U598 ( .A(n487), .B(n486), .ZN(n682) );
  NAND2_X1 U599 ( .A1(n682), .A2(n519), .ZN(n494) );
  XOR2_X1 U600 ( .A(KEYINPUT97), .B(KEYINPUT79), .Z(n490) );
  NAND2_X1 U601 ( .A1(n488), .A2(G217), .ZN(n489) );
  XNOR2_X1 U602 ( .A(n490), .B(n489), .ZN(n492) );
  INV_X1 U603 ( .A(KEYINPUT25), .ZN(n491) );
  XNOR2_X1 U604 ( .A(n492), .B(n491), .ZN(n493) );
  NOR2_X1 U605 ( .A1(n723), .A2(n722), .ZN(n719) );
  NAND2_X1 U606 ( .A1(n611), .A2(n719), .ZN(n582) );
  NOR2_X1 U607 ( .A1(n556), .A2(n582), .ZN(n620) );
  AND2_X1 U608 ( .A1(n621), .A2(n620), .ZN(n540) );
  XOR2_X1 U609 ( .A(KEYINPUT106), .B(KEYINPUT103), .Z(n496) );
  XNOR2_X1 U610 ( .A(G107), .B(KEYINPUT7), .ZN(n495) );
  XNOR2_X1 U611 ( .A(n496), .B(n495), .ZN(n498) );
  NAND2_X1 U612 ( .A1(G217), .A2(n499), .ZN(n502) );
  XOR2_X1 U613 ( .A(G116), .B(G122), .Z(n500) );
  XNOR2_X1 U614 ( .A(KEYINPUT105), .B(n500), .ZN(n501) );
  XNOR2_X1 U615 ( .A(n502), .B(n501), .ZN(n503) );
  NAND2_X1 U616 ( .A1(n687), .A2(n519), .ZN(n505) );
  XNOR2_X1 U617 ( .A(KEYINPUT107), .B(G478), .ZN(n504) );
  XOR2_X1 U618 ( .A(KEYINPUT12), .B(KEYINPUT100), .Z(n507) );
  XNOR2_X1 U619 ( .A(KEYINPUT102), .B(KEYINPUT101), .ZN(n506) );
  XNOR2_X1 U620 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U621 ( .A(n771), .B(n508), .ZN(n518) );
  XNOR2_X1 U622 ( .A(n509), .B(KEYINPUT11), .ZN(n513) );
  XNOR2_X1 U623 ( .A(G104), .B(G122), .ZN(n511) );
  XNOR2_X1 U624 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U625 ( .A(n513), .B(n512), .ZN(n516) );
  NAND2_X1 U626 ( .A1(G214), .A2(n514), .ZN(n515) );
  NAND2_X1 U627 ( .A1(n666), .A2(n519), .ZN(n521) );
  XNOR2_X1 U628 ( .A(KEYINPUT13), .B(G475), .ZN(n520) );
  INV_X1 U629 ( .A(n557), .ZN(n588) );
  NAND2_X1 U630 ( .A1(n558), .A2(n588), .ZN(n573) );
  XNOR2_X1 U631 ( .A(n523), .B(n522), .ZN(n525) );
  XNOR2_X1 U632 ( .A(n525), .B(n524), .ZN(n529) );
  NAND2_X1 U633 ( .A1(n778), .A2(G224), .ZN(n526) );
  XNOR2_X1 U634 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U635 ( .A(n529), .B(n528), .ZN(n531) );
  XNOR2_X1 U636 ( .A(n531), .B(n530), .ZN(n534) );
  XNOR2_X1 U637 ( .A(KEYINPUT16), .B(G122), .ZN(n532) );
  XNOR2_X1 U638 ( .A(n533), .B(n532), .ZN(n766) );
  XNOR2_X1 U639 ( .A(n534), .B(n766), .ZN(n672) );
  INV_X1 U640 ( .A(n651), .ZN(n655) );
  OR2_X2 U641 ( .A1(n672), .A2(n655), .ZN(n538) );
  NAND2_X1 U642 ( .A1(n535), .A2(G210), .ZN(n536) );
  XNOR2_X1 U643 ( .A(n536), .B(KEYINPUT93), .ZN(n537) );
  BUF_X1 U644 ( .A(n541), .Z(n614) );
  INV_X1 U645 ( .A(n614), .ZN(n563) );
  NOR2_X1 U646 ( .A1(n573), .A2(n563), .ZN(n539) );
  NAND2_X1 U647 ( .A1(n540), .A2(n539), .ZN(n640) );
  XNOR2_X1 U648 ( .A(n640), .B(G143), .ZN(G45) );
  NOR2_X1 U649 ( .A1(G898), .A2(n542), .ZN(n543) );
  OR2_X1 U650 ( .A1(n544), .A2(n543), .ZN(n546) );
  INV_X1 U651 ( .A(KEYINPUT96), .ZN(n545) );
  INV_X1 U652 ( .A(KEYINPUT91), .ZN(n548) );
  AND2_X1 U653 ( .A1(n589), .A2(n557), .ZN(n615) );
  INV_X1 U654 ( .A(n723), .ZN(n550) );
  XNOR2_X1 U655 ( .A(KEYINPUT73), .B(KEYINPUT22), .ZN(n551) );
  INV_X1 U656 ( .A(n722), .ZN(n577) );
  OR2_X1 U657 ( .A1(n353), .A2(n577), .ZN(n553) );
  NOR2_X1 U658 ( .A1(n718), .A2(n553), .ZN(n554) );
  NAND2_X1 U659 ( .A1(n593), .A2(n554), .ZN(n600) );
  XNOR2_X1 U660 ( .A(n600), .B(G110), .ZN(G12) );
  INV_X1 U661 ( .A(KEYINPUT6), .ZN(n555) );
  NAND2_X1 U662 ( .A1(n590), .A2(n559), .ZN(n560) );
  NOR2_X1 U663 ( .A1(n625), .A2(n718), .ZN(n561) );
  NAND2_X1 U664 ( .A1(n561), .A2(n735), .ZN(n562) );
  XNOR2_X1 U665 ( .A(n562), .B(KEYINPUT43), .ZN(n564) );
  AND2_X1 U666 ( .A1(n564), .A2(n563), .ZN(n648) );
  XNOR2_X1 U667 ( .A(G140), .B(KEYINPUT118), .ZN(n565) );
  XOR2_X1 U668 ( .A(n648), .B(n565), .Z(G42) );
  AND2_X1 U669 ( .A1(n566), .A2(n719), .ZN(n585) );
  NAND2_X1 U670 ( .A1(n585), .A2(n590), .ZN(n569) );
  INV_X1 U671 ( .A(KEYINPUT71), .ZN(n567) );
  XNOR2_X1 U672 ( .A(n567), .B(KEYINPUT33), .ZN(n568) );
  INV_X1 U673 ( .A(KEYINPUT83), .ZN(n570) );
  INV_X1 U674 ( .A(n573), .ZN(n574) );
  XNOR2_X1 U675 ( .A(KEYINPUT82), .B(KEYINPUT35), .ZN(n575) );
  INV_X1 U676 ( .A(KEYINPUT92), .ZN(n576) );
  XNOR2_X1 U677 ( .A(n718), .B(n576), .ZN(n631) );
  OR2_X1 U678 ( .A1(n590), .A2(n577), .ZN(n578) );
  NOR2_X1 U679 ( .A1(n631), .A2(n578), .ZN(n579) );
  NAND2_X1 U680 ( .A1(n593), .A2(n579), .ZN(n580) );
  XNOR2_X1 U681 ( .A(n602), .B(G119), .ZN(G21) );
  NOR2_X1 U682 ( .A1(n582), .A2(n353), .ZN(n583) );
  NAND2_X1 U683 ( .A1(n586), .A2(n583), .ZN(n584) );
  AND2_X1 U684 ( .A1(n585), .A2(n353), .ZN(n729) );
  NAND2_X1 U685 ( .A1(n586), .A2(n729), .ZN(n587) );
  OR2_X1 U686 ( .A1(n589), .A2(n588), .ZN(n646) );
  INV_X1 U687 ( .A(n646), .ZN(n710) );
  NOR2_X1 U688 ( .A1(n708), .A2(n710), .ZN(n734) );
  OR2_X1 U689 ( .A1(n718), .A2(n722), .ZN(n591) );
  NOR2_X1 U690 ( .A1(n591), .A2(n590), .ZN(n592) );
  AND2_X1 U691 ( .A1(n593), .A2(n592), .ZN(n696) );
  INV_X1 U692 ( .A(KEYINPUT88), .ZN(n595) );
  INV_X1 U693 ( .A(KEYINPUT44), .ZN(n598) );
  AND2_X1 U694 ( .A1(KEYINPUT66), .A2(KEYINPUT44), .ZN(n599) );
  AND2_X1 U695 ( .A1(n600), .A2(n599), .ZN(n601) );
  AND2_X1 U696 ( .A1(n602), .A2(n601), .ZN(n603) );
  NAND2_X1 U697 ( .A1(n604), .A2(n603), .ZN(n605) );
  INV_X1 U698 ( .A(n353), .ZN(n608) );
  INV_X1 U699 ( .A(KEYINPUT28), .ZN(n609) );
  NAND2_X1 U700 ( .A1(n612), .A2(n611), .ZN(n634) );
  INV_X1 U701 ( .A(n634), .ZN(n616) );
  XNOR2_X1 U702 ( .A(KEYINPUT75), .B(KEYINPUT38), .ZN(n613) );
  INV_X1 U703 ( .A(n615), .ZN(n738) );
  NAND2_X1 U704 ( .A1(n616), .A2(n747), .ZN(n619) );
  XOR2_X1 U705 ( .A(KEYINPUT113), .B(KEYINPUT42), .Z(n617) );
  XNOR2_X1 U706 ( .A(KEYINPUT112), .B(n617), .ZN(n618) );
  XNOR2_X1 U707 ( .A(KEYINPUT39), .B(KEYINPUT72), .ZN(n622) );
  XNOR2_X1 U708 ( .A(n624), .B(KEYINPUT40), .ZN(n782) );
  INV_X1 U709 ( .A(n625), .ZN(n628) );
  BUF_X1 U710 ( .A(n626), .Z(n627) );
  NAND2_X1 U711 ( .A1(n628), .A2(n627), .ZN(n629) );
  XNOR2_X1 U712 ( .A(n629), .B(KEYINPUT36), .ZN(n630) );
  NOR2_X1 U713 ( .A1(n631), .A2(n630), .ZN(n712) );
  AND2_X1 U714 ( .A1(n734), .A2(KEYINPUT47), .ZN(n632) );
  NOR2_X1 U715 ( .A1(KEYINPUT84), .A2(n632), .ZN(n633) );
  NOR2_X1 U716 ( .A1(n712), .A2(n633), .ZN(n641) );
  NOR2_X1 U717 ( .A1(n734), .A2(KEYINPUT47), .ZN(n635) );
  NAND2_X1 U718 ( .A1(KEYINPUT84), .A2(n734), .ZN(n637) );
  NAND2_X1 U719 ( .A1(n704), .A2(n637), .ZN(n638) );
  AND2_X1 U720 ( .A1(n638), .A2(KEYINPUT47), .ZN(n639) );
  XNOR2_X1 U721 ( .A(KEYINPUT48), .B(KEYINPUT68), .ZN(n644) );
  XNOR2_X1 U722 ( .A(n644), .B(KEYINPUT86), .ZN(n645) );
  NOR2_X1 U723 ( .A1(n647), .A2(n646), .ZN(n714) );
  NAND2_X1 U724 ( .A1(KEYINPUT2), .A2(KEYINPUT65), .ZN(n650) );
  NOR2_X1 U725 ( .A1(n651), .A2(n650), .ZN(n653) );
  NOR2_X1 U726 ( .A1(KEYINPUT2), .A2(KEYINPUT65), .ZN(n652) );
  NOR2_X1 U727 ( .A1(n653), .A2(n652), .ZN(n654) );
  INV_X1 U728 ( .A(KEYINPUT64), .ZN(n657) );
  XNOR2_X2 U729 ( .A(n658), .B(n657), .ZN(n689) );
  NAND2_X1 U730 ( .A1(n689), .A2(G472), .ZN(n661) );
  XNOR2_X1 U731 ( .A(n661), .B(n660), .ZN(n663) );
  INV_X1 U732 ( .A(G952), .ZN(n662) );
  NAND2_X1 U733 ( .A1(n662), .A2(G953), .ZN(n683) );
  NAND2_X1 U734 ( .A1(n663), .A2(n683), .ZN(n665) );
  XNOR2_X1 U735 ( .A(KEYINPUT114), .B(KEYINPUT63), .ZN(n664) );
  XNOR2_X1 U736 ( .A(n665), .B(n664), .ZN(G57) );
  NAND2_X1 U737 ( .A1(n689), .A2(G475), .ZN(n668) );
  XNOR2_X1 U738 ( .A(n668), .B(n667), .ZN(n669) );
  NAND2_X1 U739 ( .A1(n669), .A2(n683), .ZN(n671) );
  INV_X1 U740 ( .A(KEYINPUT60), .ZN(n670) );
  XNOR2_X1 U741 ( .A(n671), .B(n670), .ZN(G60) );
  NAND2_X1 U742 ( .A1(n689), .A2(G210), .ZN(n677) );
  BUF_X1 U743 ( .A(n672), .Z(n673) );
  XNOR2_X1 U744 ( .A(KEYINPUT90), .B(KEYINPUT54), .ZN(n674) );
  XNOR2_X1 U745 ( .A(n674), .B(KEYINPUT55), .ZN(n675) );
  XNOR2_X1 U746 ( .A(n677), .B(n676), .ZN(n678) );
  NAND2_X1 U747 ( .A1(n678), .A2(n683), .ZN(n680) );
  INV_X1 U748 ( .A(KEYINPUT56), .ZN(n679) );
  XNOR2_X1 U749 ( .A(n680), .B(n679), .ZN(G51) );
  AND2_X1 U750 ( .A1(n685), .A2(G217), .ZN(n681) );
  XNOR2_X1 U751 ( .A(n682), .B(n681), .ZN(n684) );
  INV_X1 U752 ( .A(n683), .ZN(n694) );
  NOR2_X1 U753 ( .A1(n684), .A2(n694), .ZN(G66) );
  AND2_X1 U754 ( .A1(n685), .A2(G478), .ZN(n686) );
  XNOR2_X1 U755 ( .A(n687), .B(n686), .ZN(n688) );
  NOR2_X1 U756 ( .A1(n688), .A2(n694), .ZN(G63) );
  NAND2_X1 U757 ( .A1(n685), .A2(G469), .ZN(n693) );
  XNOR2_X1 U758 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n690) );
  XNOR2_X1 U759 ( .A(n691), .B(n690), .ZN(n692) );
  XNOR2_X1 U760 ( .A(n693), .B(n692), .ZN(n695) );
  NOR2_X1 U761 ( .A1(n695), .A2(n694), .ZN(G54) );
  XOR2_X1 U762 ( .A(G101), .B(n696), .Z(G3) );
  XOR2_X1 U763 ( .A(KEYINPUT115), .B(KEYINPUT116), .Z(n698) );
  XNOR2_X1 U764 ( .A(n698), .B(n697), .ZN(n699) );
  XNOR2_X1 U765 ( .A(G104), .B(n699), .ZN(G6) );
  XOR2_X1 U766 ( .A(KEYINPUT117), .B(KEYINPUT26), .Z(n701) );
  XNOR2_X1 U767 ( .A(n701), .B(n700), .ZN(n703) );
  XOR2_X1 U768 ( .A(G107), .B(KEYINPUT27), .Z(n702) );
  XNOR2_X1 U769 ( .A(n703), .B(n702), .ZN(G9) );
  XOR2_X1 U770 ( .A(G128), .B(KEYINPUT29), .Z(n706) );
  NAND2_X1 U771 ( .A1(n704), .A2(n710), .ZN(n705) );
  XNOR2_X1 U772 ( .A(n706), .B(n705), .ZN(G30) );
  NAND2_X1 U773 ( .A1(n704), .A2(n708), .ZN(n707) );
  XNOR2_X1 U774 ( .A(n707), .B(G146), .ZN(G48) );
  XNOR2_X1 U775 ( .A(n709), .B(G113), .ZN(G15) );
  XNOR2_X1 U776 ( .A(n711), .B(G116), .ZN(G18) );
  XNOR2_X1 U777 ( .A(G125), .B(n712), .ZN(n713) );
  XNOR2_X1 U778 ( .A(n713), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U779 ( .A(G134), .B(n714), .Z(G36) );
  NOR2_X1 U780 ( .A1(n716), .A2(KEYINPUT2), .ZN(n717) );
  NOR2_X1 U781 ( .A1(n357), .A2(n717), .ZN(n754) );
  NOR2_X1 U782 ( .A1(n719), .A2(n718), .ZN(n721) );
  XNOR2_X1 U783 ( .A(KEYINPUT50), .B(KEYINPUT119), .ZN(n720) );
  XNOR2_X1 U784 ( .A(n721), .B(n720), .ZN(n726) );
  NAND2_X1 U785 ( .A1(n723), .A2(n722), .ZN(n724) );
  XOR2_X1 U786 ( .A(KEYINPUT49), .B(n724), .Z(n725) );
  NAND2_X1 U787 ( .A1(n726), .A2(n725), .ZN(n727) );
  NOR2_X1 U788 ( .A1(n353), .A2(n727), .ZN(n728) );
  NOR2_X1 U789 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U790 ( .A(KEYINPUT51), .B(n730), .ZN(n731) );
  NAND2_X1 U791 ( .A1(n747), .A2(n731), .ZN(n743) );
  NOR2_X1 U792 ( .A1(n734), .A2(n733), .ZN(n740) );
  NOR2_X1 U793 ( .A1(n736), .A2(n735), .ZN(n737) );
  NOR2_X1 U794 ( .A1(n738), .A2(n737), .ZN(n739) );
  OR2_X1 U795 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U796 ( .A1(n732), .A2(n741), .ZN(n742) );
  NAND2_X1 U797 ( .A1(n743), .A2(n742), .ZN(n744) );
  XOR2_X1 U798 ( .A(KEYINPUT52), .B(n744), .Z(n745) );
  NOR2_X1 U799 ( .A1(n746), .A2(n745), .ZN(n750) );
  NAND2_X1 U800 ( .A1(n747), .A2(n732), .ZN(n748) );
  XOR2_X1 U801 ( .A(KEYINPUT120), .B(n748), .Z(n749) );
  NOR2_X1 U802 ( .A1(n750), .A2(n749), .ZN(n751) );
  XOR2_X1 U803 ( .A(KEYINPUT121), .B(n751), .Z(n752) );
  NAND2_X1 U804 ( .A1(n752), .A2(n778), .ZN(n753) );
  NOR2_X1 U805 ( .A1(n754), .A2(n753), .ZN(n755) );
  XNOR2_X1 U806 ( .A(KEYINPUT53), .B(n755), .ZN(G75) );
  INV_X1 U807 ( .A(n756), .ZN(n757) );
  NOR2_X1 U808 ( .A1(n757), .A2(G953), .ZN(n763) );
  NAND2_X1 U809 ( .A1(G224), .A2(G953), .ZN(n758) );
  XNOR2_X1 U810 ( .A(n758), .B(KEYINPUT122), .ZN(n759) );
  XNOR2_X1 U811 ( .A(KEYINPUT61), .B(n759), .ZN(n760) );
  NAND2_X1 U812 ( .A1(n760), .A2(G898), .ZN(n761) );
  XNOR2_X1 U813 ( .A(n761), .B(KEYINPUT123), .ZN(n762) );
  NOR2_X1 U814 ( .A1(n763), .A2(n762), .ZN(n770) );
  NOR2_X1 U815 ( .A1(G898), .A2(n778), .ZN(n768) );
  XNOR2_X1 U816 ( .A(n764), .B(KEYINPUT124), .ZN(n765) );
  XNOR2_X1 U817 ( .A(n766), .B(n765), .ZN(n767) );
  NOR2_X1 U818 ( .A1(n768), .A2(n767), .ZN(n769) );
  XOR2_X1 U819 ( .A(n770), .B(n769), .Z(G69) );
  XNOR2_X1 U820 ( .A(n772), .B(n771), .ZN(n776) );
  XNOR2_X1 U821 ( .A(G227), .B(n776), .ZN(n773) );
  NAND2_X1 U822 ( .A1(n773), .A2(G900), .ZN(n774) );
  NAND2_X1 U823 ( .A1(n774), .A2(G953), .ZN(n781) );
  XNOR2_X1 U824 ( .A(n776), .B(n775), .ZN(n777) );
  XNOR2_X1 U825 ( .A(n777), .B(KEYINPUT125), .ZN(n779) );
  NAND2_X1 U826 ( .A1(n779), .A2(n778), .ZN(n780) );
  NAND2_X1 U827 ( .A1(n781), .A2(n780), .ZN(G72) );
  XOR2_X1 U828 ( .A(n782), .B(G131), .Z(n783) );
  XNOR2_X1 U829 ( .A(KEYINPUT127), .B(n783), .ZN(G33) );
  XNOR2_X1 U830 ( .A(G137), .B(KEYINPUT126), .ZN(n785) );
  XNOR2_X1 U831 ( .A(n785), .B(n784), .ZN(G39) );
endmodule

