

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586;

  XNOR2_X1 U326 ( .A(n359), .B(n358), .ZN(n442) );
  XNOR2_X2 U327 ( .A(n477), .B(n476), .ZN(n534) );
  NOR2_X2 U328 ( .A1(n536), .A2(n485), .ZN(n564) );
  XNOR2_X1 U329 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U330 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n476) );
  XNOR2_X1 U331 ( .A(KEYINPUT54), .B(KEYINPUT122), .ZN(n479) );
  XNOR2_X1 U332 ( .A(n456), .B(n455), .ZN(n462) );
  XNOR2_X1 U333 ( .A(n454), .B(n453), .ZN(n455) );
  XOR2_X1 U334 ( .A(KEYINPUT28), .B(n482), .Z(n539) );
  XOR2_X2 U335 ( .A(KEYINPUT124), .B(n572), .Z(n579) );
  XOR2_X2 U336 ( .A(KEYINPUT41), .B(n462), .Z(n551) );
  NOR2_X1 U337 ( .A1(n374), .A2(n373), .ZN(n375) );
  XNOR2_X1 U338 ( .A(n467), .B(KEYINPUT47), .ZN(n468) );
  XNOR2_X1 U339 ( .A(n469), .B(n468), .ZN(n475) );
  XNOR2_X1 U340 ( .A(n446), .B(n445), .ZN(n449) );
  XNOR2_X1 U341 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U342 ( .A(KEYINPUT55), .B(KEYINPUT123), .ZN(n483) );
  XNOR2_X1 U343 ( .A(KEYINPUT101), .B(KEYINPUT26), .ZN(n370) );
  XNOR2_X1 U344 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U345 ( .A(n371), .B(n370), .ZN(n549) );
  XOR2_X1 U346 ( .A(n334), .B(n333), .Z(n527) );
  XNOR2_X1 U347 ( .A(n458), .B(n457), .ZN(n507) );
  XNOR2_X1 U348 ( .A(n486), .B(G176GAT), .ZN(n487) );
  XNOR2_X1 U349 ( .A(n459), .B(G29GAT), .ZN(n460) );
  XNOR2_X1 U350 ( .A(n488), .B(n487), .ZN(G1349GAT) );
  XNOR2_X1 U351 ( .A(n461), .B(n460), .ZN(G1328GAT) );
  NAND2_X1 U352 ( .A1(G225GAT), .A2(G233GAT), .ZN(n299) );
  XOR2_X1 U353 ( .A(G85GAT), .B(G155GAT), .Z(n295) );
  XNOR2_X1 U354 ( .A(G127GAT), .B(G120GAT), .ZN(n294) );
  XNOR2_X1 U355 ( .A(n295), .B(n294), .ZN(n297) );
  XOR2_X1 U356 ( .A(G29GAT), .B(G162GAT), .Z(n296) );
  XNOR2_X1 U357 ( .A(n297), .B(n296), .ZN(n298) );
  XNOR2_X1 U358 ( .A(n299), .B(n298), .ZN(n316) );
  XOR2_X1 U359 ( .A(KEYINPUT96), .B(KEYINPUT97), .Z(n301) );
  XNOR2_X1 U360 ( .A(G1GAT), .B(KEYINPUT1), .ZN(n300) );
  XNOR2_X1 U361 ( .A(n301), .B(n300), .ZN(n314) );
  XOR2_X1 U362 ( .A(KEYINPUT94), .B(KEYINPUT95), .Z(n303) );
  XNOR2_X1 U363 ( .A(G148GAT), .B(G57GAT), .ZN(n302) );
  XNOR2_X1 U364 ( .A(n303), .B(n302), .ZN(n307) );
  XOR2_X1 U365 ( .A(KEYINPUT6), .B(KEYINPUT4), .Z(n305) );
  XNOR2_X1 U366 ( .A(KEYINPUT98), .B(KEYINPUT5), .ZN(n304) );
  XNOR2_X1 U367 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U368 ( .A(n307), .B(n306), .Z(n312) );
  XNOR2_X1 U369 ( .A(G113GAT), .B(G134GAT), .ZN(n308) );
  XNOR2_X1 U370 ( .A(n308), .B(KEYINPUT0), .ZN(n322) );
  XOR2_X1 U371 ( .A(KEYINPUT2), .B(KEYINPUT3), .Z(n310) );
  XNOR2_X1 U372 ( .A(G141GAT), .B(KEYINPUT92), .ZN(n309) );
  XNOR2_X1 U373 ( .A(n310), .B(n309), .ZN(n361) );
  XNOR2_X1 U374 ( .A(n322), .B(n361), .ZN(n311) );
  XNOR2_X1 U375 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U376 ( .A(n314), .B(n313), .Z(n315) );
  XNOR2_X1 U377 ( .A(n316), .B(n315), .ZN(n522) );
  XNOR2_X1 U378 ( .A(KEYINPUT107), .B(KEYINPUT38), .ZN(n458) );
  XOR2_X1 U379 ( .A(KEYINPUT20), .B(KEYINPUT84), .Z(n318) );
  XNOR2_X1 U380 ( .A(G190GAT), .B(KEYINPUT86), .ZN(n317) );
  XNOR2_X1 U381 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U382 ( .A(n319), .B(G99GAT), .Z(n321) );
  XOR2_X1 U383 ( .A(G120GAT), .B(G71GAT), .Z(n441) );
  XNOR2_X1 U384 ( .A(G43GAT), .B(n441), .ZN(n320) );
  XNOR2_X1 U385 ( .A(n321), .B(n320), .ZN(n326) );
  XOR2_X1 U386 ( .A(G15GAT), .B(G127GAT), .Z(n412) );
  XOR2_X1 U387 ( .A(n322), .B(n412), .Z(n324) );
  NAND2_X1 U388 ( .A1(G227GAT), .A2(G233GAT), .ZN(n323) );
  XNOR2_X1 U389 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U390 ( .A(n326), .B(n325), .Z(n334) );
  XOR2_X1 U391 ( .A(KEYINPUT17), .B(KEYINPUT19), .Z(n328) );
  XNOR2_X1 U392 ( .A(KEYINPUT18), .B(KEYINPUT85), .ZN(n327) );
  XNOR2_X1 U393 ( .A(n328), .B(n327), .ZN(n329) );
  XOR2_X1 U394 ( .A(G169GAT), .B(n329), .Z(n348) );
  XOR2_X1 U395 ( .A(G176GAT), .B(G183GAT), .Z(n331) );
  XNOR2_X1 U396 ( .A(KEYINPUT83), .B(KEYINPUT87), .ZN(n330) );
  XNOR2_X1 U397 ( .A(n331), .B(n330), .ZN(n332) );
  XNOR2_X1 U398 ( .A(n348), .B(n332), .ZN(n333) );
  XNOR2_X1 U399 ( .A(G8GAT), .B(G183GAT), .ZN(n335) );
  XNOR2_X1 U400 ( .A(n335), .B(KEYINPUT77), .ZN(n409) );
  XOR2_X1 U401 ( .A(KEYINPUT99), .B(n409), .Z(n337) );
  NAND2_X1 U402 ( .A1(G226GAT), .A2(G233GAT), .ZN(n336) );
  XNOR2_X1 U403 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U404 ( .A(G36GAT), .B(G190GAT), .Z(n385) );
  XOR2_X1 U405 ( .A(n338), .B(n385), .Z(n347) );
  XNOR2_X1 U406 ( .A(G211GAT), .B(KEYINPUT90), .ZN(n339) );
  XNOR2_X1 U407 ( .A(n339), .B(KEYINPUT21), .ZN(n340) );
  XOR2_X1 U408 ( .A(n340), .B(KEYINPUT91), .Z(n342) );
  XNOR2_X1 U409 ( .A(G197GAT), .B(G218GAT), .ZN(n341) );
  XNOR2_X1 U410 ( .A(n342), .B(n341), .ZN(n362) );
  XOR2_X1 U411 ( .A(G92GAT), .B(KEYINPUT74), .Z(n344) );
  XNOR2_X1 U412 ( .A(G176GAT), .B(G64GAT), .ZN(n343) );
  XNOR2_X1 U413 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U414 ( .A(G204GAT), .B(n345), .Z(n454) );
  XNOR2_X1 U415 ( .A(n362), .B(n454), .ZN(n346) );
  XNOR2_X1 U416 ( .A(n347), .B(n346), .ZN(n349) );
  XNOR2_X1 U417 ( .A(n349), .B(n348), .ZN(n524) );
  NAND2_X1 U418 ( .A1(n527), .A2(n524), .ZN(n367) );
  XOR2_X1 U419 ( .A(G50GAT), .B(KEYINPUT75), .Z(n350) );
  XOR2_X1 U420 ( .A(G162GAT), .B(n350), .Z(n399) );
  XOR2_X1 U421 ( .A(n399), .B(KEYINPUT23), .Z(n352) );
  NAND2_X1 U422 ( .A1(G228GAT), .A2(G233GAT), .ZN(n351) );
  XNOR2_X1 U423 ( .A(n352), .B(n351), .ZN(n366) );
  XOR2_X1 U424 ( .A(KEYINPUT89), .B(KEYINPUT93), .Z(n354) );
  XNOR2_X1 U425 ( .A(KEYINPUT24), .B(KEYINPUT88), .ZN(n353) );
  XNOR2_X1 U426 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U427 ( .A(n355), .B(KEYINPUT22), .Z(n357) );
  XOR2_X1 U428 ( .A(G22GAT), .B(G155GAT), .Z(n411) );
  XNOR2_X1 U429 ( .A(n411), .B(G204GAT), .ZN(n356) );
  XNOR2_X1 U430 ( .A(n357), .B(n356), .ZN(n360) );
  XOR2_X1 U431 ( .A(G78GAT), .B(G148GAT), .Z(n359) );
  XNOR2_X1 U432 ( .A(G106GAT), .B(KEYINPUT71), .ZN(n358) );
  XOR2_X1 U433 ( .A(n360), .B(n442), .Z(n364) );
  XNOR2_X1 U434 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U435 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U436 ( .A(n366), .B(n365), .ZN(n482) );
  NAND2_X1 U437 ( .A1(n367), .A2(n482), .ZN(n368) );
  XNOR2_X1 U438 ( .A(n368), .B(KEYINPUT103), .ZN(n369) );
  XOR2_X1 U439 ( .A(KEYINPUT25), .B(n369), .Z(n374) );
  XNOR2_X1 U440 ( .A(n524), .B(KEYINPUT27), .ZN(n378) );
  NOR2_X1 U441 ( .A1(n527), .A2(n482), .ZN(n371) );
  INV_X1 U442 ( .A(n549), .ZN(n570) );
  NAND2_X1 U443 ( .A1(n378), .A2(n570), .ZN(n372) );
  XOR2_X1 U444 ( .A(KEYINPUT102), .B(n372), .Z(n373) );
  XNOR2_X1 U445 ( .A(n375), .B(KEYINPUT104), .ZN(n376) );
  NOR2_X1 U446 ( .A1(n522), .A2(n376), .ZN(n377) );
  XNOR2_X1 U447 ( .A(n377), .B(KEYINPUT105), .ZN(n382) );
  NAND2_X1 U448 ( .A1(n522), .A2(n378), .ZN(n533) );
  NOR2_X1 U449 ( .A1(n533), .A2(n539), .ZN(n379) );
  XNOR2_X1 U450 ( .A(KEYINPUT100), .B(n379), .ZN(n380) );
  INV_X1 U451 ( .A(n527), .ZN(n536) );
  NAND2_X1 U452 ( .A1(n380), .A2(n536), .ZN(n381) );
  NAND2_X1 U453 ( .A1(n382), .A2(n381), .ZN(n492) );
  XOR2_X1 U454 ( .A(G29GAT), .B(G43GAT), .Z(n384) );
  XNOR2_X1 U455 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n383) );
  XNOR2_X1 U456 ( .A(n384), .B(n383), .ZN(n428) );
  XOR2_X1 U457 ( .A(n385), .B(KEYINPUT11), .Z(n388) );
  XNOR2_X1 U458 ( .A(G99GAT), .B(G85GAT), .ZN(n386) );
  XNOR2_X1 U459 ( .A(n386), .B(KEYINPUT72), .ZN(n447) );
  XNOR2_X1 U460 ( .A(G218GAT), .B(n447), .ZN(n387) );
  XNOR2_X1 U461 ( .A(n388), .B(n387), .ZN(n392) );
  XOR2_X1 U462 ( .A(G106GAT), .B(KEYINPUT10), .Z(n390) );
  NAND2_X1 U463 ( .A1(G232GAT), .A2(G233GAT), .ZN(n389) );
  XNOR2_X1 U464 ( .A(n390), .B(n389), .ZN(n391) );
  XOR2_X1 U465 ( .A(n392), .B(n391), .Z(n397) );
  XOR2_X1 U466 ( .A(KEYINPUT76), .B(KEYINPUT65), .Z(n394) );
  XNOR2_X1 U467 ( .A(G92GAT), .B(KEYINPUT9), .ZN(n393) );
  XNOR2_X1 U468 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U469 ( .A(G134GAT), .B(n395), .ZN(n396) );
  XNOR2_X1 U470 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U471 ( .A(n428), .B(n398), .ZN(n400) );
  XOR2_X1 U472 ( .A(n400), .B(n399), .Z(n489) );
  INV_X1 U473 ( .A(n489), .ZN(n563) );
  XOR2_X1 U474 ( .A(KEYINPUT36), .B(n563), .Z(n584) );
  XOR2_X1 U475 ( .A(KEYINPUT79), .B(G78GAT), .Z(n402) );
  XNOR2_X1 U476 ( .A(G71GAT), .B(G211GAT), .ZN(n401) );
  XNOR2_X1 U477 ( .A(n402), .B(n401), .ZN(n406) );
  XOR2_X1 U478 ( .A(KEYINPUT81), .B(KEYINPUT80), .Z(n404) );
  XNOR2_X1 U479 ( .A(G64GAT), .B(KEYINPUT78), .ZN(n403) );
  XNOR2_X1 U480 ( .A(n404), .B(n403), .ZN(n405) );
  XOR2_X1 U481 ( .A(n406), .B(n405), .Z(n408) );
  XOR2_X1 U482 ( .A(G1GAT), .B(KEYINPUT69), .Z(n425) );
  XOR2_X1 U483 ( .A(G57GAT), .B(KEYINPUT13), .Z(n452) );
  XNOR2_X1 U484 ( .A(n425), .B(n452), .ZN(n407) );
  XNOR2_X1 U485 ( .A(n408), .B(n407), .ZN(n410) );
  XOR2_X1 U486 ( .A(n410), .B(n409), .Z(n414) );
  XNOR2_X1 U487 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U488 ( .A(n414), .B(n413), .ZN(n419) );
  XOR2_X1 U489 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n416) );
  NAND2_X1 U490 ( .A1(G231GAT), .A2(G233GAT), .ZN(n415) );
  XNOR2_X1 U491 ( .A(n416), .B(n415), .ZN(n417) );
  XOR2_X1 U492 ( .A(KEYINPUT15), .B(n417), .Z(n418) );
  XOR2_X1 U493 ( .A(n419), .B(n418), .Z(n580) );
  NOR2_X1 U494 ( .A1(n584), .A2(n580), .ZN(n420) );
  NAND2_X1 U495 ( .A1(n492), .A2(n420), .ZN(n421) );
  XOR2_X1 U496 ( .A(KEYINPUT37), .B(n421), .Z(n521) );
  XOR2_X1 U497 ( .A(G15GAT), .B(G113GAT), .Z(n423) );
  XNOR2_X1 U498 ( .A(G50GAT), .B(G36GAT), .ZN(n422) );
  XNOR2_X1 U499 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U500 ( .A(n424), .B(G22GAT), .Z(n427) );
  XNOR2_X1 U501 ( .A(G169GAT), .B(n425), .ZN(n426) );
  XNOR2_X1 U502 ( .A(n427), .B(n426), .ZN(n432) );
  XOR2_X1 U503 ( .A(n428), .B(KEYINPUT66), .Z(n430) );
  NAND2_X1 U504 ( .A1(G229GAT), .A2(G233GAT), .ZN(n429) );
  XNOR2_X1 U505 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U506 ( .A(n432), .B(n431), .Z(n440) );
  XOR2_X1 U507 ( .A(KEYINPUT70), .B(G8GAT), .Z(n434) );
  XNOR2_X1 U508 ( .A(G141GAT), .B(G197GAT), .ZN(n433) );
  XNOR2_X1 U509 ( .A(n434), .B(n433), .ZN(n438) );
  XOR2_X1 U510 ( .A(KEYINPUT68), .B(KEYINPUT67), .Z(n436) );
  XNOR2_X1 U511 ( .A(KEYINPUT30), .B(KEYINPUT29), .ZN(n435) );
  XNOR2_X1 U512 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U513 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U514 ( .A(n440), .B(n439), .Z(n560) );
  INV_X1 U515 ( .A(n560), .ZN(n573) );
  XNOR2_X1 U516 ( .A(n442), .B(n441), .ZN(n446) );
  AND2_X1 U517 ( .A1(G230GAT), .A2(G233GAT), .ZN(n444) );
  INV_X1 U518 ( .A(KEYINPUT33), .ZN(n443) );
  XNOR2_X1 U519 ( .A(n447), .B(KEYINPUT73), .ZN(n448) );
  XNOR2_X1 U520 ( .A(n449), .B(n448), .ZN(n451) );
  INV_X1 U521 ( .A(KEYINPUT32), .ZN(n450) );
  XNOR2_X1 U522 ( .A(n451), .B(n450), .ZN(n456) );
  XNOR2_X1 U523 ( .A(n452), .B(KEYINPUT31), .ZN(n453) );
  BUF_X1 U524 ( .A(n462), .Z(n576) );
  OR2_X1 U525 ( .A1(n573), .A2(n576), .ZN(n494) );
  OR2_X1 U526 ( .A1(n521), .A2(n494), .ZN(n457) );
  NAND2_X1 U527 ( .A1(n522), .A2(n507), .ZN(n461) );
  XOR2_X1 U528 ( .A(KEYINPUT39), .B(KEYINPUT108), .Z(n459) );
  XOR2_X1 U529 ( .A(KEYINPUT121), .B(n524), .Z(n478) );
  AND2_X1 U530 ( .A1(n560), .A2(n551), .ZN(n463) );
  XNOR2_X1 U531 ( .A(n463), .B(KEYINPUT46), .ZN(n464) );
  NOR2_X1 U532 ( .A1(n580), .A2(n464), .ZN(n465) );
  XNOR2_X1 U533 ( .A(n465), .B(KEYINPUT115), .ZN(n466) );
  NOR2_X1 U534 ( .A1(n563), .A2(n466), .ZN(n469) );
  XOR2_X1 U535 ( .A(KEYINPUT116), .B(KEYINPUT117), .Z(n467) );
  INV_X1 U536 ( .A(n580), .ZN(n470) );
  NOR2_X1 U537 ( .A1(n584), .A2(n470), .ZN(n471) );
  XOR2_X1 U538 ( .A(KEYINPUT45), .B(n471), .Z(n472) );
  NOR2_X1 U539 ( .A1(n576), .A2(n472), .ZN(n473) );
  NAND2_X1 U540 ( .A1(n473), .A2(n573), .ZN(n474) );
  NAND2_X1 U541 ( .A1(n475), .A2(n474), .ZN(n477) );
  NAND2_X1 U542 ( .A1(n478), .A2(n534), .ZN(n480) );
  NOR2_X1 U543 ( .A1(n522), .A2(n481), .ZN(n571) );
  NAND2_X1 U544 ( .A1(n482), .A2(n571), .ZN(n484) );
  NAND2_X1 U545 ( .A1(n564), .A2(n551), .ZN(n488) );
  XOR2_X1 U546 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n486) );
  XOR2_X1 U547 ( .A(KEYINPUT16), .B(KEYINPUT82), .Z(n491) );
  NAND2_X1 U548 ( .A1(n580), .A2(n489), .ZN(n490) );
  XNOR2_X1 U549 ( .A(n491), .B(n490), .ZN(n493) );
  NAND2_X1 U550 ( .A1(n493), .A2(n492), .ZN(n509) );
  NOR2_X1 U551 ( .A1(n494), .A2(n509), .ZN(n501) );
  NAND2_X1 U552 ( .A1(n501), .A2(n522), .ZN(n495) );
  XNOR2_X1 U553 ( .A(n495), .B(KEYINPUT34), .ZN(n496) );
  XNOR2_X1 U554 ( .A(G1GAT), .B(n496), .ZN(G1324GAT) );
  NAND2_X1 U555 ( .A1(n524), .A2(n501), .ZN(n497) );
  XNOR2_X1 U556 ( .A(n497), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U557 ( .A(KEYINPUT35), .B(KEYINPUT106), .Z(n499) );
  NAND2_X1 U558 ( .A1(n501), .A2(n527), .ZN(n498) );
  XNOR2_X1 U559 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U560 ( .A(G15GAT), .B(n500), .ZN(G1326GAT) );
  NAND2_X1 U561 ( .A1(n539), .A2(n501), .ZN(n502) );
  XNOR2_X1 U562 ( .A(n502), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U563 ( .A(G36GAT), .B(KEYINPUT109), .Z(n504) );
  NAND2_X1 U564 ( .A1(n507), .A2(n524), .ZN(n503) );
  XNOR2_X1 U565 ( .A(n504), .B(n503), .ZN(G1329GAT) );
  NAND2_X1 U566 ( .A1(n507), .A2(n527), .ZN(n505) );
  XNOR2_X1 U567 ( .A(n505), .B(KEYINPUT40), .ZN(n506) );
  XNOR2_X1 U568 ( .A(G43GAT), .B(n506), .ZN(G1330GAT) );
  NAND2_X1 U569 ( .A1(n507), .A2(n539), .ZN(n508) );
  XNOR2_X1 U570 ( .A(n508), .B(G50GAT), .ZN(G1331GAT) );
  NAND2_X1 U571 ( .A1(n551), .A2(n573), .ZN(n520) );
  NOR2_X1 U572 ( .A1(n520), .A2(n509), .ZN(n515) );
  NAND2_X1 U573 ( .A1(n522), .A2(n515), .ZN(n510) );
  XNOR2_X1 U574 ( .A(KEYINPUT42), .B(n510), .ZN(n511) );
  XNOR2_X1 U575 ( .A(G57GAT), .B(n511), .ZN(G1332GAT) );
  NAND2_X1 U576 ( .A1(n524), .A2(n515), .ZN(n512) );
  XNOR2_X1 U577 ( .A(n512), .B(KEYINPUT110), .ZN(n513) );
  XNOR2_X1 U578 ( .A(G64GAT), .B(n513), .ZN(G1333GAT) );
  NAND2_X1 U579 ( .A1(n527), .A2(n515), .ZN(n514) );
  XNOR2_X1 U580 ( .A(n514), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U581 ( .A(KEYINPUT112), .B(KEYINPUT43), .Z(n517) );
  NAND2_X1 U582 ( .A1(n515), .A2(n539), .ZN(n516) );
  XNOR2_X1 U583 ( .A(n517), .B(n516), .ZN(n519) );
  XOR2_X1 U584 ( .A(G78GAT), .B(KEYINPUT111), .Z(n518) );
  XNOR2_X1 U585 ( .A(n519), .B(n518), .ZN(G1335GAT) );
  NOR2_X1 U586 ( .A1(n521), .A2(n520), .ZN(n529) );
  NAND2_X1 U587 ( .A1(n522), .A2(n529), .ZN(n523) );
  XNOR2_X1 U588 ( .A(G85GAT), .B(n523), .ZN(G1336GAT) );
  XOR2_X1 U589 ( .A(G92GAT), .B(KEYINPUT113), .Z(n526) );
  NAND2_X1 U590 ( .A1(n529), .A2(n524), .ZN(n525) );
  XNOR2_X1 U591 ( .A(n526), .B(n525), .ZN(G1337GAT) );
  NAND2_X1 U592 ( .A1(n527), .A2(n529), .ZN(n528) );
  XNOR2_X1 U593 ( .A(n528), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U594 ( .A(KEYINPUT44), .B(KEYINPUT114), .Z(n531) );
  NAND2_X1 U595 ( .A1(n529), .A2(n539), .ZN(n530) );
  XNOR2_X1 U596 ( .A(n531), .B(n530), .ZN(n532) );
  XOR2_X1 U597 ( .A(G106GAT), .B(n532), .Z(G1339GAT) );
  INV_X1 U598 ( .A(n533), .ZN(n535) );
  NAND2_X1 U599 ( .A1(n535), .A2(n534), .ZN(n548) );
  NOR2_X1 U600 ( .A1(n536), .A2(n548), .ZN(n537) );
  XOR2_X1 U601 ( .A(KEYINPUT118), .B(n537), .Z(n538) );
  NOR2_X1 U602 ( .A1(n539), .A2(n538), .ZN(n545) );
  NAND2_X1 U603 ( .A1(n560), .A2(n545), .ZN(n540) );
  XNOR2_X1 U604 ( .A(n540), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U605 ( .A(G120GAT), .B(KEYINPUT49), .Z(n542) );
  NAND2_X1 U606 ( .A1(n545), .A2(n551), .ZN(n541) );
  XNOR2_X1 U607 ( .A(n542), .B(n541), .ZN(G1341GAT) );
  NAND2_X1 U608 ( .A1(n545), .A2(n580), .ZN(n543) );
  XNOR2_X1 U609 ( .A(n543), .B(KEYINPUT50), .ZN(n544) );
  XNOR2_X1 U610 ( .A(G127GAT), .B(n544), .ZN(G1342GAT) );
  XOR2_X1 U611 ( .A(G134GAT), .B(KEYINPUT51), .Z(n547) );
  NAND2_X1 U612 ( .A1(n545), .A2(n563), .ZN(n546) );
  XNOR2_X1 U613 ( .A(n547), .B(n546), .ZN(G1343GAT) );
  NOR2_X1 U614 ( .A1(n549), .A2(n548), .ZN(n557) );
  NAND2_X1 U615 ( .A1(n557), .A2(n560), .ZN(n550) );
  XNOR2_X1 U616 ( .A(G141GAT), .B(n550), .ZN(G1344GAT) );
  XOR2_X1 U617 ( .A(KEYINPUT119), .B(KEYINPUT53), .Z(n553) );
  NAND2_X1 U618 ( .A1(n557), .A2(n551), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n553), .B(n552), .ZN(n555) );
  XOR2_X1 U620 ( .A(G148GAT), .B(KEYINPUT52), .Z(n554) );
  XNOR2_X1 U621 ( .A(n555), .B(n554), .ZN(G1345GAT) );
  NAND2_X1 U622 ( .A1(n557), .A2(n580), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n556), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U624 ( .A1(n557), .A2(n563), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n558), .B(KEYINPUT120), .ZN(n559) );
  XNOR2_X1 U626 ( .A(G162GAT), .B(n559), .ZN(G1347GAT) );
  NAND2_X1 U627 ( .A1(n560), .A2(n564), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n561), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U629 ( .A1(n564), .A2(n580), .ZN(n562) );
  XNOR2_X1 U630 ( .A(n562), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U631 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n565), .B(KEYINPUT58), .ZN(n566) );
  XNOR2_X1 U633 ( .A(G190GAT), .B(n566), .ZN(G1351GAT) );
  XOR2_X1 U634 ( .A(KEYINPUT126), .B(KEYINPUT60), .Z(n568) );
  XNOR2_X1 U635 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n567) );
  XNOR2_X1 U636 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U637 ( .A(KEYINPUT125), .B(n569), .ZN(n575) );
  NAND2_X1 U638 ( .A1(n571), .A2(n570), .ZN(n572) );
  INV_X1 U639 ( .A(n579), .ZN(n583) );
  NOR2_X1 U640 ( .A1(n573), .A2(n583), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(G1352GAT) );
  XOR2_X1 U642 ( .A(G204GAT), .B(KEYINPUT61), .Z(n578) );
  NAND2_X1 U643 ( .A1(n579), .A2(n576), .ZN(n577) );
  XNOR2_X1 U644 ( .A(n578), .B(n577), .ZN(G1353GAT) );
  XOR2_X1 U645 ( .A(G211GAT), .B(KEYINPUT127), .Z(n582) );
  NAND2_X1 U646 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(G1354GAT) );
  NOR2_X1 U648 ( .A1(n584), .A2(n583), .ZN(n585) );
  XOR2_X1 U649 ( .A(KEYINPUT62), .B(n585), .Z(n586) );
  XNOR2_X1 U650 ( .A(G218GAT), .B(n586), .ZN(G1355GAT) );
endmodule

