//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 0 1 1 1 0 0 1 0 0 0 0 1 1 0 1 0 0 1 1 1 0 0 0 1 0 0 1 1 1 0 0 1 0 0 1 1 1 1 1 0 0 1 0 1 1 1 1 0 0 1 0 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:21 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n447, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n544, new_n545, new_n546, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n604, new_n605, new_n608, new_n609, new_n611, new_n612,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1159, new_n1160,
    new_n1161;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT64), .B(G2066), .ZN(G411));
  XNOR2_X1  g006(.A(KEYINPUT65), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT66), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT67), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  XNOR2_X1  g017(.A(KEYINPUT68), .B(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  NAND2_X1  g021(.A1(G94), .A2(G452), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n447), .B(KEYINPUT69), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  OR4_X1    g027(.A1(G221), .A2(G220), .A3(G219), .A4(G218), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n455), .A2(new_n456), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  INV_X1    g034(.A(G567), .ZN(new_n460));
  OAI21_X1  g035(.A(new_n459), .B1(new_n460), .B2(new_n456), .ZN(new_n461));
  XNOR2_X1  g036(.A(new_n461), .B(KEYINPUT70), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  XNOR2_X1  g038(.A(KEYINPUT3), .B(G2104), .ZN(new_n464));
  AND2_X1   g039(.A1(new_n464), .A2(G125), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  XOR2_X1   g041(.A(new_n466), .B(KEYINPUT71), .Z(new_n467));
  OAI21_X1  g042(.A(G2105), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  AND2_X1   g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  NOR2_X1   g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n471), .A2(G2105), .ZN(new_n472));
  INV_X1    g047(.A(G2105), .ZN(new_n473));
  AND2_X1   g048(.A1(new_n473), .A2(G2104), .ZN(new_n474));
  AOI22_X1  g049(.A1(new_n472), .A2(G137), .B1(G101), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n468), .A2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(G160));
  NAND2_X1  g052(.A1(new_n472), .A2(G136), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n471), .A2(new_n473), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  OR2_X1    g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n481), .B(G2104), .C1(G112), .C2(new_n473), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n478), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G162));
  AND2_X1   g059(.A1(G126), .A2(G2105), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n485), .B1(new_n469), .B2(new_n470), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(KEYINPUT72), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT72), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n488), .B(new_n485), .C1(new_n469), .C2(new_n470), .ZN(new_n489));
  AND2_X1   g064(.A1(KEYINPUT73), .A2(G114), .ZN(new_n490));
  NOR2_X1   g065(.A1(KEYINPUT73), .A2(G114), .ZN(new_n491));
  OAI21_X1  g066(.A(G2105), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  OAI21_X1  g067(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  AOI22_X1  g069(.A1(new_n487), .A2(new_n489), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  OAI211_X1 g070(.A(G138), .B(new_n473), .C1(new_n469), .C2(new_n470), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n464), .A2(new_n498), .A3(G138), .A4(new_n473), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n495), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(G164));
  INV_X1    g077(.A(G50), .ZN(new_n503));
  AND2_X1   g078(.A1(KEYINPUT6), .A2(G651), .ZN(new_n504));
  NOR2_X1   g079(.A1(KEYINPUT6), .A2(G651), .ZN(new_n505));
  OR2_X1    g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(G543), .ZN(new_n507));
  NOR2_X1   g082(.A1(KEYINPUT5), .A2(G543), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n506), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G88), .ZN(new_n513));
  OAI22_X1  g088(.A1(new_n503), .A2(new_n507), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n511), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n514), .A2(new_n517), .ZN(G166));
  NAND3_X1  g093(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n519));
  XNOR2_X1  g094(.A(new_n519), .B(KEYINPUT7), .ZN(new_n520));
  INV_X1    g095(.A(G51), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n520), .B1(new_n507), .B2(new_n521), .ZN(new_n522));
  AND2_X1   g097(.A1(KEYINPUT5), .A2(G543), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n523), .A2(new_n508), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n506), .A2(G89), .ZN(new_n525));
  NAND2_X1  g100(.A1(G63), .A2(G651), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n522), .A2(new_n527), .ZN(G168));
  INV_X1    g103(.A(G52), .ZN(new_n529));
  INV_X1    g104(.A(G90), .ZN(new_n530));
  OAI22_X1  g105(.A1(new_n529), .A2(new_n507), .B1(new_n512), .B2(new_n530), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n511), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n532), .A2(new_n516), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n531), .A2(new_n533), .ZN(G171));
  INV_X1    g109(.A(G43), .ZN(new_n535));
  INV_X1    g110(.A(G81), .ZN(new_n536));
  OAI22_X1  g111(.A1(new_n535), .A2(new_n507), .B1(new_n512), .B2(new_n536), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n511), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n538), .A2(new_n516), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G860), .ZN(new_n541));
  XOR2_X1   g116(.A(new_n541), .B(KEYINPUT74), .Z(G153));
  NAND4_X1  g117(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g118(.A1(G1), .A2(G3), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n544), .B(KEYINPUT75), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT8), .ZN(new_n546));
  NAND4_X1  g121(.A1(G319), .A2(G483), .A3(G661), .A4(new_n546), .ZN(G188));
  XNOR2_X1  g122(.A(new_n524), .B(KEYINPUT76), .ZN(new_n548));
  AND2_X1   g123(.A1(new_n548), .A2(G65), .ZN(new_n549));
  AND2_X1   g124(.A1(G78), .A2(G543), .ZN(new_n550));
  OAI21_X1  g125(.A(G651), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(G53), .ZN(new_n552));
  OR3_X1    g127(.A1(new_n507), .A2(KEYINPUT9), .A3(new_n552), .ZN(new_n553));
  OAI21_X1  g128(.A(KEYINPUT9), .B1(new_n507), .B2(new_n552), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n504), .A2(new_n505), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n555), .A2(new_n524), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n553), .A2(new_n554), .B1(G91), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n551), .A2(new_n557), .ZN(G299));
  INV_X1    g133(.A(G171), .ZN(G301));
  INV_X1    g134(.A(G168), .ZN(G286));
  INV_X1    g135(.A(G166), .ZN(G303));
  NAND2_X1  g136(.A1(new_n556), .A2(G87), .ZN(new_n562));
  INV_X1    g137(.A(G543), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n555), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G49), .ZN(new_n565));
  OAI21_X1  g140(.A(G651), .B1(new_n511), .B2(G74), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n562), .A2(new_n565), .A3(new_n566), .ZN(G288));
  OAI21_X1  g142(.A(G61), .B1(new_n523), .B2(new_n508), .ZN(new_n568));
  OR2_X1    g143(.A1(new_n568), .A2(KEYINPUT77), .ZN(new_n569));
  AOI22_X1  g144(.A1(new_n568), .A2(KEYINPUT77), .B1(G73), .B2(G543), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(G651), .ZN(new_n572));
  AOI22_X1  g147(.A1(G86), .A2(new_n556), .B1(new_n564), .B2(G48), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n572), .A2(new_n573), .ZN(G305));
  INV_X1    g149(.A(G85), .ZN(new_n575));
  XNOR2_X1  g150(.A(KEYINPUT78), .B(G47), .ZN(new_n576));
  OAI22_X1  g151(.A1(new_n575), .A2(new_n512), .B1(new_n507), .B2(new_n576), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n511), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n578));
  NOR2_X1   g153(.A1(new_n578), .A2(new_n516), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(G290));
  INV_X1    g156(.A(G868), .ZN(new_n582));
  NOR2_X1   g157(.A1(G171), .A2(new_n582), .ZN(new_n583));
  XNOR2_X1  g158(.A(new_n583), .B(KEYINPUT79), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT10), .ZN(new_n585));
  INV_X1    g160(.A(G92), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n512), .B2(new_n586), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n556), .A2(KEYINPUT10), .A3(G92), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n587), .A2(new_n588), .B1(G54), .B2(new_n564), .ZN(new_n589));
  NAND2_X1  g164(.A1(G79), .A2(G543), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n511), .B(KEYINPUT76), .ZN(new_n591));
  INV_X1    g166(.A(G66), .ZN(new_n592));
  OAI211_X1 g167(.A(KEYINPUT80), .B(new_n590), .C1(new_n591), .C2(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n593), .A2(G651), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n548), .A2(G66), .ZN(new_n595));
  AOI21_X1  g170(.A(KEYINPUT80), .B1(new_n595), .B2(new_n590), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n589), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT81), .ZN(new_n598));
  AND2_X1   g173(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n597), .A2(new_n598), .ZN(new_n600));
  OR2_X1    g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n584), .B1(new_n601), .B2(G868), .ZN(G284));
  OAI21_X1  g177(.A(new_n584), .B1(new_n601), .B2(G868), .ZN(G321));
  NAND2_X1  g178(.A1(G286), .A2(G868), .ZN(new_n604));
  INV_X1    g179(.A(G299), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n605), .B2(G868), .ZN(G280));
  XOR2_X1   g181(.A(G280), .B(KEYINPUT82), .Z(G297));
  NOR2_X1   g182(.A1(new_n599), .A2(new_n600), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n608), .A2(G559), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n609), .B1(G860), .B2(new_n601), .ZN(G148));
  OR2_X1    g185(.A1(new_n537), .A2(new_n539), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n611), .A2(new_n582), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n612), .B1(new_n609), .B2(new_n582), .ZN(G323));
  XNOR2_X1  g188(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g189(.A1(new_n472), .A2(G135), .ZN(new_n615));
  XOR2_X1   g190(.A(new_n615), .B(KEYINPUT84), .Z(new_n616));
  OAI21_X1  g191(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n617));
  INV_X1    g192(.A(G111), .ZN(new_n618));
  AOI21_X1  g193(.A(new_n617), .B1(new_n618), .B2(G2105), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n619), .B1(new_n479), .B2(G123), .ZN(new_n620));
  AND2_X1   g195(.A1(new_n616), .A2(new_n620), .ZN(new_n621));
  INV_X1    g196(.A(new_n621), .ZN(new_n622));
  OR2_X1    g197(.A1(new_n622), .A2(G2096), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n464), .A2(new_n474), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT12), .ZN(new_n625));
  XNOR2_X1  g200(.A(KEYINPUT83), .B(KEYINPUT13), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  INV_X1    g202(.A(new_n627), .ZN(new_n628));
  OR2_X1    g203(.A1(new_n628), .A2(G2100), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n628), .A2(G2100), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n622), .A2(G2096), .ZN(new_n631));
  NAND4_X1  g206(.A1(new_n623), .A2(new_n629), .A3(new_n630), .A4(new_n631), .ZN(G156));
  XNOR2_X1  g207(.A(G2427), .B(G2438), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2430), .ZN(new_n634));
  XNOR2_X1  g209(.A(KEYINPUT15), .B(G2435), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n634), .A2(new_n635), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n636), .A2(KEYINPUT14), .A3(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2443), .B(G2446), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(G1341), .B(G1348), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(G2451), .B(G2454), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT16), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT85), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n643), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n643), .A2(new_n646), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n647), .A2(G14), .A3(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n649), .B(KEYINPUT86), .Z(G401));
  XOR2_X1   g225(.A(G2072), .B(G2078), .Z(new_n651));
  XOR2_X1   g226(.A(new_n651), .B(KEYINPUT87), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT17), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2067), .B(G2678), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2084), .B(G2090), .ZN(new_n655));
  NOR3_X1   g230(.A1(new_n653), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  OAI21_X1  g231(.A(new_n655), .B1(new_n652), .B2(new_n654), .ZN(new_n657));
  AOI21_X1  g232(.A(new_n657), .B1(new_n653), .B2(new_n654), .ZN(new_n658));
  INV_X1    g233(.A(new_n654), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n659), .A2(new_n655), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n652), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT18), .ZN(new_n662));
  NOR3_X1   g237(.A1(new_n656), .A2(new_n658), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2096), .B(G2100), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(G227));
  XOR2_X1   g240(.A(G1971), .B(G1976), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT19), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1956), .B(G2474), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1961), .B(G1966), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  AND2_X1   g245(.A1(new_n668), .A2(new_n669), .ZN(new_n671));
  NOR3_X1   g246(.A1(new_n667), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n667), .A2(new_n670), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n673), .B(KEYINPUT20), .Z(new_n674));
  AOI211_X1 g249(.A(new_n672), .B(new_n674), .C1(new_n667), .C2(new_n671), .ZN(new_n675));
  XOR2_X1   g250(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1991), .B(G1996), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1981), .B(G1986), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(G229));
  NAND2_X1  g256(.A1(new_n472), .A2(G139), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n473), .A2(G103), .A3(G2104), .ZN(new_n683));
  INV_X1    g258(.A(KEYINPUT25), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n464), .A2(G127), .ZN(new_n687));
  NAND2_X1  g262(.A1(G115), .A2(G2104), .ZN(new_n688));
  AOI21_X1  g263(.A(new_n473), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT93), .ZN(new_n691));
  MUX2_X1   g266(.A(G33), .B(new_n691), .S(G29), .Z(new_n692));
  NOR2_X1   g267(.A1(new_n692), .A2(G2072), .ZN(new_n693));
  XOR2_X1   g268(.A(new_n693), .B(KEYINPUT94), .Z(new_n694));
  INV_X1    g269(.A(G16), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n695), .A2(G20), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT23), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n697), .B1(new_n605), .B2(new_n695), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT98), .B(G1956), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  AND2_X1   g276(.A1(new_n692), .A2(G2072), .ZN(new_n702));
  AND2_X1   g277(.A1(new_n699), .A2(new_n700), .ZN(new_n703));
  NOR4_X1   g278(.A1(new_n694), .A2(new_n701), .A3(new_n702), .A4(new_n703), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n601), .A2(new_n695), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n705), .B1(G4), .B2(new_n695), .ZN(new_n706));
  INV_X1    g281(.A(G1348), .ZN(new_n707));
  OR2_X1    g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n706), .A2(new_n707), .ZN(new_n709));
  NOR2_X1   g284(.A1(G171), .A2(new_n695), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n710), .B1(G5), .B2(new_n695), .ZN(new_n711));
  INV_X1    g286(.A(G1961), .ZN(new_n712));
  NOR2_X1   g287(.A1(G16), .A2(G19), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n713), .B1(new_n540), .B2(G16), .ZN(new_n714));
  OAI22_X1  g289(.A1(new_n711), .A2(new_n712), .B1(new_n714), .B2(G1341), .ZN(new_n715));
  XOR2_X1   g290(.A(KEYINPUT88), .B(G29), .Z(new_n716));
  INV_X1    g291(.A(KEYINPUT24), .ZN(new_n717));
  OR2_X1    g292(.A1(new_n717), .A2(G34), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n717), .A2(G34), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n716), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(G29), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n720), .B1(new_n476), .B2(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(G2084), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n715), .A2(new_n724), .ZN(new_n725));
  AOI22_X1  g300(.A1(new_n711), .A2(new_n712), .B1(G1341), .B2(new_n714), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n721), .A2(G32), .ZN(new_n727));
  AOI22_X1  g302(.A1(new_n472), .A2(G141), .B1(G105), .B2(new_n474), .ZN(new_n728));
  NAND3_X1  g303(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n729), .B(KEYINPUT26), .Z(new_n730));
  INV_X1    g305(.A(G129), .ZN(new_n731));
  INV_X1    g306(.A(new_n479), .ZN(new_n732));
  OAI211_X1 g307(.A(new_n728), .B(new_n730), .C1(new_n731), .C2(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(new_n733), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n727), .B1(new_n734), .B2(new_n721), .ZN(new_n735));
  XNOR2_X1  g310(.A(KEYINPUT27), .B(G1996), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT95), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n735), .B(new_n737), .ZN(new_n738));
  NAND3_X1  g313(.A1(new_n725), .A2(new_n726), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n716), .A2(G26), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT28), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n472), .A2(G140), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n479), .A2(G128), .ZN(new_n743));
  OR2_X1    g318(.A1(G104), .A2(G2105), .ZN(new_n744));
  OAI211_X1 g319(.A(new_n744), .B(G2104), .C1(G116), .C2(new_n473), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n742), .A2(new_n743), .A3(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(new_n746), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n741), .B1(new_n747), .B2(new_n721), .ZN(new_n748));
  INV_X1    g323(.A(G2067), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(new_n716), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n751), .A2(G35), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(G162), .B2(new_n751), .ZN(new_n753));
  XNOR2_X1  g328(.A(KEYINPUT97), .B(KEYINPUT29), .ZN(new_n754));
  INV_X1    g329(.A(G2090), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n753), .B(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT31), .ZN(new_n758));
  OR2_X1    g333(.A1(new_n758), .A2(G11), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n758), .A2(G11), .ZN(new_n760));
  INV_X1    g335(.A(KEYINPUT30), .ZN(new_n761));
  AND2_X1   g336(.A1(new_n761), .A2(G28), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n721), .B1(new_n761), .B2(G28), .ZN(new_n763));
  OAI211_X1 g338(.A(new_n759), .B(new_n760), .C1(new_n762), .C2(new_n763), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(new_n621), .B2(new_n751), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n695), .A2(G21), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(G168), .B2(new_n695), .ZN(new_n767));
  OR2_X1    g342(.A1(new_n767), .A2(G1966), .ZN(new_n768));
  NAND4_X1  g343(.A1(new_n750), .A2(new_n757), .A3(new_n765), .A4(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n767), .A2(G1966), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(KEYINPUT96), .Z(new_n771));
  NOR2_X1   g346(.A1(new_n751), .A2(G27), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(G164), .B2(new_n751), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(G2078), .ZN(new_n774));
  NOR4_X1   g349(.A1(new_n739), .A2(new_n769), .A3(new_n771), .A4(new_n774), .ZN(new_n775));
  NAND4_X1  g350(.A1(new_n704), .A2(new_n708), .A3(new_n709), .A4(new_n775), .ZN(new_n776));
  NOR2_X1   g351(.A1(G16), .A2(G23), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT91), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G288), .B2(new_n695), .ZN(new_n779));
  XOR2_X1   g354(.A(KEYINPUT33), .B(G1976), .Z(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(KEYINPUT92), .ZN(new_n782));
  OR2_X1    g357(.A1(G6), .A2(G16), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G305), .B2(new_n695), .ZN(new_n784));
  XNOR2_X1  g359(.A(KEYINPUT32), .B(G1981), .ZN(new_n785));
  INV_X1    g360(.A(new_n785), .ZN(new_n786));
  AOI22_X1  g361(.A1(new_n781), .A2(new_n782), .B1(new_n784), .B2(new_n786), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(new_n782), .B2(new_n781), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n695), .A2(G22), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(G166), .B2(new_n695), .ZN(new_n790));
  OR2_X1    g365(.A1(new_n790), .A2(G1971), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n790), .A2(G1971), .ZN(new_n792));
  OAI211_X1 g367(.A(new_n791), .B(new_n792), .C1(new_n784), .C2(new_n786), .ZN(new_n793));
  OR3_X1    g368(.A1(new_n788), .A2(KEYINPUT34), .A3(new_n793), .ZN(new_n794));
  OAI21_X1  g369(.A(KEYINPUT34), .B1(new_n788), .B2(new_n793), .ZN(new_n795));
  AND2_X1   g370(.A1(new_n716), .A2(G25), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n479), .A2(G119), .ZN(new_n797));
  XOR2_X1   g372(.A(new_n797), .B(KEYINPUT89), .Z(new_n798));
  OAI21_X1  g373(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n799));
  INV_X1    g374(.A(G107), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n799), .B1(new_n800), .B2(G2105), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(new_n472), .B2(G131), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n798), .A2(new_n802), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n796), .B1(new_n803), .B2(new_n751), .ZN(new_n804));
  XOR2_X1   g379(.A(KEYINPUT35), .B(G1991), .Z(new_n805));
  AND2_X1   g380(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n804), .A2(new_n805), .ZN(new_n807));
  INV_X1    g382(.A(G24), .ZN(new_n808));
  OR3_X1    g383(.A1(new_n808), .A2(KEYINPUT90), .A3(G16), .ZN(new_n809));
  OAI21_X1  g384(.A(KEYINPUT90), .B1(new_n808), .B2(G16), .ZN(new_n810));
  OAI211_X1 g385(.A(new_n809), .B(new_n810), .C1(new_n580), .C2(new_n695), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(G1986), .ZN(new_n812));
  NOR3_X1   g387(.A1(new_n806), .A2(new_n807), .A3(new_n812), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n794), .A2(new_n795), .A3(new_n813), .ZN(new_n814));
  XOR2_X1   g389(.A(new_n814), .B(KEYINPUT36), .Z(new_n815));
  NOR2_X1   g390(.A1(new_n776), .A2(new_n815), .ZN(G311));
  INV_X1    g391(.A(G311), .ZN(G150));
  NAND2_X1  g392(.A1(new_n601), .A2(G559), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT38), .ZN(new_n819));
  INV_X1    g394(.A(G93), .ZN(new_n820));
  XNOR2_X1  g395(.A(KEYINPUT99), .B(G55), .ZN(new_n821));
  OAI22_X1  g396(.A1(new_n820), .A2(new_n512), .B1(new_n507), .B2(new_n821), .ZN(new_n822));
  AOI22_X1  g397(.A1(new_n511), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n823), .A2(new_n516), .ZN(new_n824));
  OR2_X1    g399(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n825), .A2(new_n611), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n822), .A2(new_n824), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n540), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n819), .B(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT39), .ZN(new_n831));
  AOI21_X1  g406(.A(G860), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n832), .B1(new_n831), .B2(new_n830), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n825), .A2(G860), .ZN(new_n834));
  XOR2_X1   g409(.A(KEYINPUT100), .B(KEYINPUT37), .Z(new_n835));
  XNOR2_X1  g410(.A(new_n834), .B(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n833), .A2(new_n836), .ZN(G145));
  INV_X1    g412(.A(G37), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n733), .B(new_n747), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT102), .ZN(new_n840));
  AND3_X1   g415(.A1(new_n495), .A2(new_n840), .A3(new_n500), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n840), .B1(new_n495), .B2(new_n500), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n839), .B(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(new_n690), .ZN(new_n845));
  OR2_X1    g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n844), .A2(new_n691), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n803), .B(new_n625), .ZN(new_n849));
  OAI21_X1  g424(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n850));
  INV_X1    g425(.A(G118), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n850), .B1(new_n851), .B2(G2105), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n479), .A2(G130), .ZN(new_n853));
  XOR2_X1   g428(.A(new_n853), .B(KEYINPUT103), .Z(new_n854));
  AOI211_X1 g429(.A(new_n852), .B(new_n854), .C1(G142), .C2(new_n472), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n849), .B(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n848), .A2(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(G162), .B(new_n476), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(KEYINPUT101), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(new_n622), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n856), .A2(new_n846), .A3(new_n847), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n858), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n861), .B1(new_n858), .B2(new_n862), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT104), .ZN(new_n865));
  AND2_X1   g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n864), .A2(new_n865), .ZN(new_n867));
  OAI211_X1 g442(.A(new_n838), .B(new_n863), .C1(new_n866), .C2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g444(.A(new_n829), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n609), .B(new_n870), .ZN(new_n871));
  XOR2_X1   g446(.A(KEYINPUT105), .B(KEYINPUT41), .Z(new_n872));
  OR2_X1    g447(.A1(new_n597), .A2(G299), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n597), .A2(G299), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n872), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n873), .A2(new_n874), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n876), .A2(KEYINPUT41), .ZN(new_n877));
  OR3_X1    g452(.A1(new_n871), .A2(new_n875), .A3(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n871), .A2(new_n876), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n580), .B(G288), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT106), .ZN(new_n881));
  AND2_X1   g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n880), .A2(new_n881), .ZN(new_n883));
  XNOR2_X1  g458(.A(G305), .B(G166), .ZN(new_n884));
  OR3_X1    g459(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n883), .A2(new_n884), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(KEYINPUT42), .ZN(new_n888));
  AND3_X1   g463(.A1(new_n878), .A2(new_n879), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n888), .B1(new_n878), .B2(new_n879), .ZN(new_n890));
  OAI21_X1  g465(.A(G868), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n891), .B1(G868), .B2(new_n827), .ZN(G295));
  OAI21_X1  g467(.A(new_n891), .B1(G868), .B2(new_n827), .ZN(G331));
  NOR2_X1   g468(.A1(new_n829), .A2(G171), .ZN(new_n894));
  AOI21_X1  g469(.A(G301), .B1(new_n826), .B2(new_n828), .ZN(new_n895));
  OR3_X1    g470(.A1(new_n894), .A2(G286), .A3(new_n895), .ZN(new_n896));
  OAI21_X1  g471(.A(G286), .B1(new_n894), .B2(new_n895), .ZN(new_n897));
  OAI211_X1 g472(.A(new_n896), .B(new_n897), .C1(new_n877), .C2(new_n875), .ZN(new_n898));
  INV_X1    g473(.A(new_n887), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n896), .A2(new_n897), .ZN(new_n900));
  INV_X1    g475(.A(new_n876), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n898), .A2(new_n899), .A3(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT107), .ZN(new_n904));
  AOI21_X1  g479(.A(G37), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n898), .A2(new_n902), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n906), .A2(new_n887), .ZN(new_n907));
  NAND4_X1  g482(.A1(new_n898), .A2(new_n899), .A3(new_n902), .A4(KEYINPUT107), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n905), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT43), .ZN(new_n910));
  AND2_X1   g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  OAI211_X1 g486(.A(new_n896), .B(new_n897), .C1(new_n901), .C2(KEYINPUT41), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n876), .A2(new_n872), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n902), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(new_n887), .ZN(new_n915));
  AND4_X1   g490(.A1(KEYINPUT43), .A2(new_n905), .A3(new_n908), .A4(new_n915), .ZN(new_n916));
  OAI21_X1  g491(.A(KEYINPUT44), .B1(new_n911), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n909), .A2(KEYINPUT43), .ZN(new_n918));
  NAND4_X1  g493(.A1(new_n905), .A2(new_n910), .A3(new_n908), .A4(new_n915), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT44), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n917), .A2(new_n922), .ZN(G397));
  INV_X1    g498(.A(G1384), .ZN(new_n924));
  AOI21_X1  g499(.A(KEYINPUT45), .B1(new_n843), .B2(new_n924), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n468), .A2(new_n475), .A3(G40), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(new_n928), .ZN(new_n929));
  XOR2_X1   g504(.A(new_n733), .B(G1996), .Z(new_n930));
  XNOR2_X1  g505(.A(new_n746), .B(new_n749), .ZN(new_n931));
  INV_X1    g506(.A(new_n805), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n803), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n798), .A2(new_n805), .A3(new_n802), .ZN(new_n934));
  NAND4_X1  g509(.A1(new_n930), .A2(new_n931), .A3(new_n933), .A4(new_n934), .ZN(new_n935));
  XOR2_X1   g510(.A(new_n580), .B(G1986), .Z(new_n936));
  OAI21_X1  g511(.A(new_n929), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(G303), .A2(G8), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n938), .B(KEYINPUT55), .ZN(new_n939));
  AOI21_X1  g514(.A(KEYINPUT109), .B1(new_n501), .B2(new_n924), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT109), .ZN(new_n941));
  AOI211_X1 g516(.A(new_n941), .B(G1384), .C1(new_n495), .C2(new_n500), .ZN(new_n942));
  OAI21_X1  g517(.A(KEYINPUT50), .B1(new_n940), .B2(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(G1384), .B1(new_n495), .B2(new_n500), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT50), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n926), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n943), .A2(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(G2090), .B1(new_n947), .B2(KEYINPUT114), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT114), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n943), .A2(new_n949), .A3(new_n946), .ZN(new_n950));
  AND2_X1   g525(.A1(new_n497), .A2(new_n499), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n492), .A2(new_n494), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n488), .B1(new_n464), .B2(new_n485), .ZN(new_n953));
  INV_X1    g528(.A(new_n489), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n952), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(KEYINPUT102), .B1(new_n951), .B2(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n495), .A2(new_n840), .A3(new_n500), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT45), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n958), .A2(G1384), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n956), .A2(new_n957), .A3(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT108), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n956), .A2(KEYINPUT108), .A3(new_n957), .A4(new_n959), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n927), .B1(new_n944), .B2(KEYINPUT45), .ZN(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(G1971), .ZN(new_n968));
  AOI22_X1  g543(.A1(new_n948), .A2(new_n950), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(G8), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n939), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n924), .B1(new_n951), .B2(new_n955), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT110), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n972), .A2(new_n973), .A3(KEYINPUT50), .ZN(new_n974));
  OAI21_X1  g549(.A(KEYINPUT110), .B1(new_n944), .B2(new_n945), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n972), .A2(new_n941), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n944), .A2(KEYINPUT109), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n977), .A2(new_n945), .A3(new_n978), .ZN(new_n979));
  NAND4_X1  g554(.A1(new_n976), .A2(new_n979), .A3(new_n755), .A4(new_n927), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n965), .B1(new_n962), .B2(new_n963), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n980), .B1(new_n981), .B2(G1971), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(KEYINPUT111), .ZN(new_n983));
  INV_X1    g558(.A(new_n939), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT111), .ZN(new_n985));
  OAI211_X1 g560(.A(new_n980), .B(new_n985), .C1(new_n981), .C2(G1971), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n983), .A2(G8), .A3(new_n984), .A4(new_n986), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n977), .A2(new_n927), .A3(new_n978), .ZN(new_n988));
  INV_X1    g563(.A(G288), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(G1976), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n988), .A2(G8), .A3(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(KEYINPUT52), .ZN(new_n992));
  INV_X1    g567(.A(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(G305), .A2(G1981), .ZN(new_n994));
  INV_X1    g569(.A(G1981), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n572), .A2(new_n995), .A3(new_n573), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n994), .A2(KEYINPUT49), .A3(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT49), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n995), .B1(new_n572), .B2(new_n573), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n516), .B1(new_n569), .B2(new_n570), .ZN(new_n1000));
  INV_X1    g575(.A(G48), .ZN(new_n1001));
  INV_X1    g576(.A(G86), .ZN(new_n1002));
  OAI22_X1  g577(.A1(new_n1001), .A2(new_n507), .B1(new_n512), .B2(new_n1002), .ZN(new_n1003));
  NOR3_X1   g578(.A1(new_n1000), .A2(new_n1003), .A3(G1981), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n998), .B1(new_n999), .B2(new_n1004), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n997), .A2(new_n1005), .A3(new_n988), .A4(G8), .ZN(new_n1006));
  INV_X1    g581(.A(G1976), .ZN(new_n1007));
  AOI21_X1  g582(.A(KEYINPUT52), .B1(G288), .B2(new_n1007), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n988), .A2(G8), .A3(new_n990), .A4(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1006), .A2(new_n1009), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n993), .A2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n971), .A2(new_n987), .A3(new_n1011), .ZN(new_n1012));
  NOR2_X1   g587(.A1(G168), .A2(new_n970), .ZN(new_n1013));
  INV_X1    g588(.A(G1966), .ZN(new_n1014));
  AOI21_X1  g589(.A(KEYINPUT45), .B1(new_n977), .B2(new_n978), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n927), .B1(new_n972), .B2(new_n958), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1014), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n976), .A2(new_n979), .A3(new_n723), .A4(new_n927), .ZN(new_n1018));
  AND3_X1   g593(.A1(new_n1017), .A2(new_n1018), .A3(KEYINPUT121), .ZN(new_n1019));
  AOI21_X1  g594(.A(KEYINPUT121), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1013), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(G8), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1013), .A2(KEYINPUT51), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NOR3_X1   g600(.A1(new_n1019), .A2(new_n1020), .A3(G286), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT51), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1027), .A2(new_n970), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1028), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1025), .B1(new_n1026), .B2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1012), .B1(new_n1021), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT53), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1032), .B1(new_n967), .B2(G2078), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n976), .A2(new_n979), .A3(new_n927), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(KEYINPUT117), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT117), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n976), .A2(new_n979), .A3(new_n1036), .A4(new_n927), .ZN(new_n1037));
  XOR2_X1   g612(.A(KEYINPUT122), .B(G1961), .Z(new_n1038));
  NAND3_X1  g613(.A1(new_n1035), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1039));
  OR4_X1    g614(.A1(new_n1032), .A2(new_n1015), .A3(G2078), .A4(new_n1016), .ZN(new_n1040));
  AND3_X1   g615(.A1(new_n1039), .A2(KEYINPUT123), .A3(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(KEYINPUT123), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1042));
  OAI211_X1 g617(.A(G301), .B(new_n1033), .C1(new_n1041), .C2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT124), .ZN(new_n1044));
  AND3_X1   g619(.A1(new_n1035), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1045));
  OR3_X1    g620(.A1(new_n926), .A2(new_n1032), .A3(G2078), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n925), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(new_n964), .ZN(new_n1048));
  AOI211_X1 g623(.A(G2078), .B(new_n965), .C1(new_n962), .C2(new_n963), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1048), .B1(new_n1049), .B2(KEYINPUT53), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1044), .B1(new_n1045), .B2(new_n1050), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1039), .A2(new_n1033), .A3(KEYINPUT124), .A4(new_n1048), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1051), .A2(G171), .A3(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1043), .A2(KEYINPUT54), .A3(new_n1053), .ZN(new_n1054));
  NOR3_X1   g629(.A1(new_n1045), .A2(new_n1050), .A3(G171), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1033), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1055), .B1(new_n1056), .B2(G171), .ZN(new_n1057));
  OAI211_X1 g632(.A(new_n1031), .B(new_n1054), .C1(new_n1057), .C2(KEYINPUT54), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1035), .A2(new_n707), .A3(new_n1037), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n977), .A2(new_n749), .A3(new_n927), .A4(new_n978), .ZN(new_n1060));
  XOR2_X1   g635(.A(new_n1060), .B(KEYINPUT116), .Z(new_n1061));
  NAND2_X1  g636(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1062));
  XOR2_X1   g637(.A(G299), .B(KEYINPUT57), .Z(new_n1063));
  INV_X1    g638(.A(G1956), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n947), .A2(new_n1064), .ZN(new_n1065));
  XNOR2_X1  g640(.A(KEYINPUT56), .B(G2072), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n981), .A2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1063), .A2(new_n1065), .A3(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1062), .A2(new_n601), .A3(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1063), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1067), .A2(new_n1065), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1069), .A2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1059), .A2(new_n1061), .A3(KEYINPUT60), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(KEYINPUT120), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT120), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1059), .A2(new_n1061), .A3(new_n1076), .A4(KEYINPUT60), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1075), .A2(new_n601), .A3(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1074), .A2(KEYINPUT120), .A3(new_n608), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT60), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1062), .A2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1078), .A2(new_n1079), .A3(new_n1081), .ZN(new_n1082));
  XNOR2_X1  g657(.A(KEYINPUT118), .B(G1996), .ZN(new_n1083));
  AOI211_X1 g658(.A(new_n1083), .B(new_n965), .C1(new_n962), .C2(new_n963), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT119), .ZN(new_n1085));
  INV_X1    g660(.A(new_n988), .ZN(new_n1086));
  XNOR2_X1  g661(.A(KEYINPUT58), .B(G1341), .ZN(new_n1087));
  OAI22_X1  g662(.A1(new_n1084), .A2(new_n1085), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  NOR3_X1   g663(.A1(new_n967), .A2(KEYINPUT119), .A3(new_n1083), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n540), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(KEYINPUT59), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT59), .ZN(new_n1092));
  OAI211_X1 g667(.A(new_n1092), .B(new_n540), .C1(new_n1088), .C2(new_n1089), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1068), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1063), .B1(new_n1067), .B2(new_n1065), .ZN(new_n1095));
  OAI21_X1  g670(.A(KEYINPUT61), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT61), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1072), .A2(new_n1097), .A3(new_n1068), .ZN(new_n1098));
  AOI22_X1  g673(.A1(new_n1091), .A2(new_n1093), .B1(new_n1096), .B2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1073), .B1(new_n1082), .B2(new_n1099), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1058), .A2(new_n1100), .ZN(new_n1101));
  AND2_X1   g676(.A1(new_n1056), .A2(G171), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1012), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT62), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1030), .A2(new_n1104), .A3(new_n1021), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT121), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1022), .A2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1017), .A2(new_n1018), .A3(KEYINPUT121), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1107), .A2(G168), .A3(new_n1108), .ZN(new_n1109));
  AOI22_X1  g684(.A1(new_n1109), .A2(new_n1028), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1021), .ZN(new_n1111));
  OAI21_X1  g686(.A(KEYINPUT62), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1102), .A2(new_n1103), .A3(new_n1105), .A4(new_n1112), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n983), .A2(G8), .A3(new_n986), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(new_n939), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1022), .A2(KEYINPUT63), .A3(G8), .A4(G168), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT112), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1117), .B1(new_n993), .B2(new_n1010), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n992), .A2(KEYINPUT112), .A3(new_n1009), .A4(new_n1006), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1116), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1115), .A2(new_n987), .A3(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT115), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT63), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1022), .A2(G8), .A3(G168), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1124), .B1(new_n1012), .B2(new_n1125), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1115), .A2(new_n1120), .A3(KEYINPUT115), .A4(new_n987), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1123), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n987), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n988), .A2(G8), .ZN(new_n1130));
  XNOR2_X1  g705(.A(new_n1130), .B(KEYINPUT113), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1006), .A2(new_n1007), .A3(new_n989), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1131), .B1(new_n1132), .B2(new_n996), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1129), .A2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1113), .A2(new_n1128), .A3(new_n1134), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n937), .B1(new_n1101), .B2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n928), .B1(new_n734), .B2(new_n931), .ZN(new_n1137));
  OR3_X1    g712(.A1(new_n928), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1138));
  OAI21_X1  g713(.A(KEYINPUT46), .B1(new_n928), .B2(G1996), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1137), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  XOR2_X1   g715(.A(new_n1140), .B(KEYINPUT47), .Z(new_n1141));
  NAND2_X1  g716(.A1(new_n930), .A2(new_n931), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n929), .A2(new_n1142), .ZN(new_n1143));
  XOR2_X1   g718(.A(new_n934), .B(KEYINPUT125), .Z(new_n1144));
  AOI22_X1  g719(.A1(new_n1143), .A2(new_n1144), .B1(new_n749), .B2(new_n747), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT126), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n928), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1147), .B1(new_n1146), .B2(new_n1145), .ZN(new_n1148));
  OR3_X1    g723(.A1(new_n928), .A2(G1986), .A3(G290), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1149), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1150), .A2(KEYINPUT48), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n929), .A2(new_n935), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT48), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1152), .B1(new_n1149), .B2(new_n1153), .ZN(new_n1154));
  OAI211_X1 g729(.A(new_n1141), .B(new_n1148), .C1(new_n1151), .C2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1136), .A2(new_n1156), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g732(.A1(new_n462), .A2(G227), .ZN(new_n1159));
  NAND2_X1  g733(.A1(new_n649), .A2(new_n1159), .ZN(new_n1160));
  NOR2_X1   g734(.A1(G229), .A2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g735(.A1(new_n1161), .A2(new_n920), .A3(new_n868), .ZN(G225));
  INV_X1    g736(.A(G225), .ZN(G308));
endmodule


