//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 1 0 1 0 0 0 1 0 1 1 1 1 1 0 1 1 0 1 0 1 0 0 0 0 0 0 1 1 1 0 0 0 0 1 0 1 0 0 1 0 1 0 1 1 0 1 1 1 0 1 1 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:37 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1341,
    new_n1342, new_n1343;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G50), .ZN(new_n204));
  INV_X1    g0004(.A(G77), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n206), .B(KEYINPUT64), .ZN(G353));
  OAI21_X1  g0007(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n210));
  INV_X1    g0010(.A(G232), .ZN(new_n211));
  INV_X1    g0011(.A(G238), .ZN(new_n212));
  OAI221_X1 g0012(.A(new_n210), .B1(new_n201), .B2(new_n211), .C1(new_n202), .C2(new_n212), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G50), .A2(G226), .B1(G87), .B2(G250), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  OAI21_X1  g0016(.A(new_n209), .B1(new_n213), .B2(new_n216), .ZN(new_n217));
  XNOR2_X1  g0017(.A(new_n217), .B(KEYINPUT1), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n209), .A2(G13), .ZN(new_n219));
  OAI211_X1 g0019(.A(new_n219), .B(G250), .C1(G257), .C2(G264), .ZN(new_n220));
  INV_X1    g0020(.A(KEYINPUT0), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n203), .A2(G50), .ZN(new_n222));
  INV_X1    g0022(.A(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G13), .ZN(new_n224));
  INV_X1    g0024(.A(G20), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  AOI22_X1  g0026(.A1(new_n220), .A2(new_n221), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n227), .B1(new_n221), .B2(new_n220), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n218), .A2(new_n228), .ZN(G361));
  XOR2_X1   g0029(.A(G226), .B(G232), .Z(new_n230));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(KEYINPUT65), .B(KEYINPUT2), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G250), .B(G257), .Z(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XOR2_X1   g0038(.A(G107), .B(G116), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT66), .ZN(new_n240));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n242), .B(new_n245), .Z(G351));
  INV_X1    g0046(.A(G1), .ZN(new_n247));
  NAND3_X1  g0047(.A1(new_n247), .A2(G13), .A3(G20), .ZN(new_n248));
  INV_X1    g0048(.A(KEYINPUT71), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND4_X1  g0050(.A1(new_n247), .A2(KEYINPUT71), .A3(G13), .A4(G20), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(new_n202), .ZN(new_n254));
  OR2_X1    g0054(.A1(new_n254), .A2(KEYINPUT12), .ZN(new_n255));
  AND2_X1   g0055(.A1(new_n255), .A2(KEYINPUT73), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n254), .A2(KEYINPUT12), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n257), .B1(new_n255), .B2(KEYINPUT73), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g0059(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(new_n224), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n225), .A2(G33), .ZN(new_n262));
  OAI22_X1  g0062(.A1(new_n262), .A2(new_n205), .B1(new_n225), .B2(G68), .ZN(new_n263));
  INV_X1    g0063(.A(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n225), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G50), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n261), .B1(new_n263), .B2(new_n267), .ZN(new_n268));
  XNOR2_X1  g0068(.A(new_n268), .B(KEYINPUT11), .ZN(new_n269));
  INV_X1    g0069(.A(new_n261), .ZN(new_n270));
  OAI211_X1 g0070(.A(new_n252), .B(new_n270), .C1(G1), .C2(new_n225), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n269), .B1(new_n202), .B2(new_n271), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n259), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G169), .ZN(new_n275));
  NAND2_X1  g0075(.A1(G33), .A2(G41), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n276), .A2(G1), .A3(G13), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(KEYINPUT68), .ZN(new_n278));
  AND2_X1   g0078(.A1(G1), .A2(G13), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT68), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n279), .A2(new_n280), .A3(new_n276), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n278), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(G33), .A2(G97), .ZN(new_n283));
  XNOR2_X1  g0083(.A(KEYINPUT3), .B(G33), .ZN(new_n284));
  INV_X1    g0084(.A(G1698), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G226), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n283), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n284), .A2(G1698), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n289), .A2(new_n211), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n282), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G41), .ZN(new_n292));
  INV_X1    g0092(.A(G45), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  AOI22_X1  g0094(.A1(new_n247), .A2(new_n294), .B1(new_n279), .B2(new_n276), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(G238), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n247), .B1(G41), .B2(G45), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT67), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n247), .B(KEYINPUT67), .C1(G41), .C2(G45), .ZN(new_n300));
  NAND4_X1  g0100(.A1(new_n299), .A2(G274), .A3(new_n277), .A4(new_n300), .ZN(new_n301));
  AND3_X1   g0101(.A1(new_n296), .A2(new_n301), .A3(KEYINPUT72), .ZN(new_n302));
  AOI21_X1  g0102(.A(KEYINPUT72), .B1(new_n296), .B2(new_n301), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n291), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(KEYINPUT13), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT13), .ZN(new_n306));
  OAI211_X1 g0106(.A(new_n291), .B(new_n306), .C1(new_n302), .C2(new_n303), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n275), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT14), .ZN(new_n309));
  AND2_X1   g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n305), .A2(G179), .A3(new_n307), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n311), .B1(new_n308), .B2(new_n309), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n274), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  AND2_X1   g0113(.A1(new_n305), .A2(new_n307), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(G190), .ZN(new_n315));
  INV_X1    g0115(.A(G200), .ZN(new_n316));
  OAI211_X1 g0116(.A(new_n315), .B(new_n273), .C1(new_n316), .C2(new_n314), .ZN(new_n317));
  AND3_X1   g0117(.A1(new_n313), .A2(KEYINPUT74), .A3(new_n317), .ZN(new_n318));
  XNOR2_X1  g0118(.A(KEYINPUT8), .B(G58), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT69), .ZN(new_n320));
  XNOR2_X1  g0120(.A(new_n319), .B(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n271), .A2(new_n321), .ZN(new_n322));
  XNOR2_X1  g0122(.A(new_n319), .B(KEYINPUT69), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(new_n252), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT7), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n327), .B1(new_n284), .B2(G20), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n264), .A2(KEYINPUT3), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT3), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(G33), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n332), .A2(KEYINPUT7), .A3(new_n225), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n328), .A2(new_n333), .A3(KEYINPUT76), .ZN(new_n334));
  AOI21_X1  g0134(.A(KEYINPUT7), .B1(new_n332), .B2(new_n225), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT76), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n334), .A2(new_n337), .A3(G68), .ZN(new_n338));
  AND2_X1   g0138(.A1(G58), .A2(G68), .ZN(new_n339));
  NOR2_X1   g0139(.A1(G58), .A2(G68), .ZN(new_n340));
  OAI21_X1  g0140(.A(G20), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NOR2_X1   g0141(.A1(G20), .A2(G33), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(G159), .ZN(new_n343));
  AND3_X1   g0143(.A1(new_n341), .A2(KEYINPUT75), .A3(new_n343), .ZN(new_n344));
  AOI21_X1  g0144(.A(KEYINPUT75), .B1(new_n341), .B2(new_n343), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n338), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT16), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT75), .ZN(new_n350));
  NAND2_X1  g0150(.A1(G58), .A2(G68), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n225), .B1(new_n203), .B2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(new_n343), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n350), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n341), .A2(KEYINPUT75), .A3(new_n343), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n202), .B1(new_n328), .B2(new_n333), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n270), .B1(new_n358), .B2(KEYINPUT16), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n326), .B1(new_n349), .B2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT77), .ZN(new_n361));
  AND3_X1   g0161(.A1(new_n300), .A2(new_n277), .A3(G274), .ZN(new_n362));
  AOI22_X1  g0162(.A1(new_n362), .A2(new_n299), .B1(G232), .B2(new_n295), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n329), .A2(new_n331), .A3(G226), .A4(G1698), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n329), .A2(new_n331), .A3(G223), .A4(new_n285), .ZN(new_n365));
  NAND2_X1  g0165(.A1(G33), .A2(G87), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n364), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(new_n282), .ZN(new_n368));
  INV_X1    g0168(.A(G190), .ZN(new_n369));
  AND3_X1   g0169(.A1(new_n363), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  AOI21_X1  g0170(.A(G200), .B1(new_n363), .B2(new_n368), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n361), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n363), .A2(new_n368), .A3(new_n369), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n277), .A2(G232), .A3(new_n297), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n301), .A2(new_n374), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n375), .B1(new_n282), .B2(new_n367), .ZN(new_n376));
  OAI211_X1 g0176(.A(KEYINPUT77), .B(new_n373), .C1(new_n376), .C2(G200), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n372), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n360), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(KEYINPUT17), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT17), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n360), .A2(new_n378), .A3(new_n381), .ZN(new_n382));
  NOR3_X1   g0182(.A1(new_n284), .A2(new_n327), .A3(G20), .ZN(new_n383));
  OAI21_X1  g0183(.A(G68), .B1(new_n383), .B2(new_n335), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n346), .A2(new_n384), .A3(KEYINPUT16), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(new_n261), .ZN(new_n386));
  AOI21_X1  g0186(.A(KEYINPUT16), .B1(new_n338), .B2(new_n346), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n325), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n376), .A2(G179), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n389), .B1(new_n376), .B2(new_n275), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT18), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n388), .A2(KEYINPUT18), .A3(new_n390), .ZN(new_n394));
  AOI22_X1  g0194(.A1(new_n380), .A2(new_n382), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT9), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT70), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n397), .B1(new_n204), .B2(new_n225), .ZN(new_n398));
  OAI211_X1 g0198(.A(KEYINPUT70), .B(G20), .C1(new_n203), .C2(G50), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n342), .A2(G150), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n398), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n264), .A2(G20), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n321), .A2(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n270), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n253), .A2(new_n266), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n406), .B1(new_n271), .B2(new_n266), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n396), .B1(new_n405), .B2(new_n407), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n323), .A2(new_n262), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n261), .B1(new_n409), .B2(new_n401), .ZN(new_n410));
  OR2_X1    g0210(.A1(new_n271), .A2(new_n266), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n410), .A2(KEYINPUT9), .A3(new_n406), .A4(new_n411), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n284), .A2(G222), .A3(new_n285), .ZN(new_n413));
  INV_X1    g0213(.A(G223), .ZN(new_n414));
  OAI221_X1 g0214(.A(new_n413), .B1(new_n205), .B2(new_n284), .C1(new_n289), .C2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(new_n282), .ZN(new_n416));
  AOI22_X1  g0216(.A1(new_n362), .A2(new_n299), .B1(G226), .B2(new_n295), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(G200), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n416), .A2(G190), .A3(new_n417), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n408), .A2(new_n412), .A3(new_n419), .A4(new_n420), .ZN(new_n421));
  XNOR2_X1  g0221(.A(new_n421), .B(KEYINPUT10), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n418), .A2(new_n275), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n410), .A2(new_n406), .A3(new_n411), .ZN(new_n424));
  OAI211_X1 g0224(.A(new_n423), .B(new_n424), .C1(G179), .C2(new_n418), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n295), .A2(G244), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(new_n301), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n332), .A2(G107), .ZN(new_n428));
  OAI221_X1 g0228(.A(new_n428), .B1(new_n286), .B2(new_n211), .C1(new_n212), .C2(new_n289), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n427), .B1(new_n429), .B2(new_n282), .ZN(new_n430));
  INV_X1    g0230(.A(G179), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  OR2_X1    g0232(.A1(new_n271), .A2(new_n205), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n253), .A2(new_n205), .ZN(new_n434));
  XOR2_X1   g0234(.A(KEYINPUT15), .B(G87), .Z(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n436), .A2(new_n262), .ZN(new_n437));
  OAI22_X1  g0237(.A1(new_n319), .A2(new_n265), .B1(new_n225), .B2(new_n205), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n261), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n433), .A2(new_n434), .A3(new_n439), .ZN(new_n440));
  OAI211_X1 g0240(.A(new_n432), .B(new_n440), .C1(G169), .C2(new_n430), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  AND2_X1   g0242(.A1(new_n430), .A2(G190), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n430), .A2(new_n316), .ZN(new_n444));
  NOR3_X1   g0244(.A1(new_n443), .A2(new_n444), .A3(new_n440), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n442), .A2(new_n445), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n395), .A2(new_n422), .A3(new_n425), .A4(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(KEYINPUT74), .B1(new_n313), .B2(new_n317), .ZN(new_n448));
  NOR3_X1   g0248(.A1(new_n318), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n329), .A2(new_n331), .A3(G250), .A4(new_n285), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n329), .A2(new_n331), .A3(G257), .A4(G1698), .ZN(new_n451));
  NAND2_X1  g0251(.A1(G33), .A2(G294), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n450), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(new_n282), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n247), .B(G45), .C1(new_n292), .C2(KEYINPUT5), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT5), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n456), .A2(G41), .ZN(new_n457));
  OAI211_X1 g0257(.A(G264), .B(new_n277), .C1(new_n455), .C2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n454), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n247), .A2(G45), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n292), .A2(KEYINPUT5), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n456), .A2(G41), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n462), .A2(new_n463), .A3(new_n464), .A4(G274), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n275), .B1(new_n460), .B2(new_n465), .ZN(new_n466));
  AND3_X1   g0266(.A1(new_n454), .A2(KEYINPUT85), .A3(new_n458), .ZN(new_n467));
  AOI21_X1  g0267(.A(KEYINPUT85), .B1(new_n454), .B2(new_n458), .ZN(new_n468));
  OAI211_X1 g0268(.A(G179), .B(new_n465), .C1(new_n467), .C2(new_n468), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n466), .B1(new_n469), .B2(KEYINPUT86), .ZN(new_n470));
  INV_X1    g0270(.A(new_n465), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT85), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n459), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n454), .A2(KEYINPUT85), .A3(new_n458), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n471), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT86), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n475), .A2(new_n476), .A3(G179), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n470), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n247), .A2(G33), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n252), .A2(new_n270), .A3(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(G107), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n252), .A2(G107), .ZN(new_n483));
  XNOR2_X1  g0283(.A(new_n483), .B(KEYINPUT25), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT23), .ZN(new_n485));
  NOR3_X1   g0285(.A1(new_n485), .A2(new_n225), .A3(G107), .ZN(new_n486));
  INV_X1    g0286(.A(G107), .ZN(new_n487));
  AOI21_X1  g0287(.A(KEYINPUT23), .B1(new_n487), .B2(G20), .ZN(new_n488));
  NAND2_X1  g0288(.A1(G33), .A2(G116), .ZN(new_n489));
  OAI22_X1  g0289(.A1(new_n486), .A2(new_n488), .B1(G20), .B2(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n284), .A2(new_n225), .A3(G87), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(KEYINPUT22), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT22), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n284), .A2(new_n493), .A3(new_n225), .A4(G87), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n490), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  AND2_X1   g0295(.A1(new_n495), .A2(KEYINPUT24), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n261), .B1(new_n495), .B2(KEYINPUT24), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n482), .B(new_n484), .C1(new_n496), .C2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n478), .A2(new_n498), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n329), .A2(new_n331), .A3(G257), .A4(new_n285), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n329), .A2(new_n331), .A3(G264), .A4(G1698), .ZN(new_n501));
  INV_X1    g0301(.A(G303), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n500), .B(new_n501), .C1(new_n502), .C2(new_n284), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(new_n282), .ZN(new_n504));
  OAI211_X1 g0304(.A(G270), .B(new_n277), .C1(new_n455), .C2(new_n457), .ZN(new_n505));
  AND2_X1   g0305(.A1(new_n505), .A2(new_n465), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n316), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(new_n507), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n252), .A2(G116), .A3(new_n270), .A4(new_n479), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n509), .B1(G116), .B2(new_n252), .ZN(new_n510));
  INV_X1    g0310(.A(G116), .ZN(new_n511));
  AOI22_X1  g0311(.A1(new_n260), .A2(new_n224), .B1(G20), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(G33), .A2(G283), .ZN(new_n513));
  INV_X1    g0313(.A(G97), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n513), .B(new_n225), .C1(G33), .C2(new_n514), .ZN(new_n515));
  AND3_X1   g0315(.A1(new_n512), .A2(KEYINPUT20), .A3(new_n515), .ZN(new_n516));
  AOI21_X1  g0316(.A(KEYINPUT20), .B1(new_n512), .B2(new_n515), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n510), .A2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT84), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n508), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  OAI221_X1 g0321(.A(new_n509), .B1(G116), .B2(new_n252), .C1(new_n517), .C2(new_n516), .ZN(new_n522));
  OAI21_X1  g0322(.A(KEYINPUT84), .B1(new_n522), .B2(new_n507), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n504), .A2(new_n506), .ZN(new_n524));
  INV_X1    g0324(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(G190), .ZN(new_n526));
  AND3_X1   g0326(.A1(new_n521), .A2(new_n523), .A3(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT21), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n524), .A2(G169), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n528), .B1(new_n529), .B2(new_n519), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n522), .A2(KEYINPUT21), .A3(G169), .A4(new_n524), .ZN(new_n531));
  AND3_X1   g0331(.A1(new_n504), .A2(G179), .A3(new_n506), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(new_n522), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n530), .A2(new_n531), .A3(new_n533), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n527), .A2(new_n534), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n465), .B1(new_n467), .B2(new_n468), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(new_n316), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n460), .A2(new_n369), .A3(new_n465), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n498), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(new_n539), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n499), .A2(new_n535), .A3(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT6), .ZN(new_n542));
  AND2_X1   g0342(.A1(G97), .A2(G107), .ZN(new_n543));
  NOR2_X1   g0343(.A1(G97), .A2(G107), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n542), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n487), .A2(KEYINPUT78), .A3(KEYINPUT6), .A4(G97), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT78), .ZN(new_n547));
  NAND2_X1  g0347(.A1(KEYINPUT6), .A2(G97), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n547), .B1(new_n548), .B2(G107), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n545), .A2(new_n546), .A3(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT79), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n545), .A2(KEYINPUT79), .A3(new_n546), .A4(new_n549), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n552), .A2(G20), .A3(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT80), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n342), .A2(G77), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n334), .A2(new_n337), .A3(G107), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n555), .B1(new_n554), .B2(new_n556), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n261), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n252), .A2(G97), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n562), .B1(new_n481), .B2(G97), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n329), .A2(new_n331), .A3(G244), .A4(new_n285), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT4), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n284), .A2(KEYINPUT4), .A3(G244), .A4(new_n285), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n284), .A2(G250), .A3(G1698), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n567), .A2(new_n568), .A3(new_n513), .A4(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(new_n282), .ZN(new_n571));
  OAI211_X1 g0371(.A(G257), .B(new_n277), .C1(new_n455), .C2(new_n457), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n465), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n575), .A2(G179), .ZN(new_n576));
  AOI21_X1  g0376(.A(KEYINPUT81), .B1(new_n571), .B2(new_n574), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT81), .ZN(new_n578));
  AOI211_X1 g0378(.A(new_n578), .B(new_n573), .C1(new_n570), .C2(new_n282), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n576), .B1(new_n580), .B2(new_n275), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n564), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n481), .A2(new_n435), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT19), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n225), .B1(new_n283), .B2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(G87), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n544), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  AOI21_X1  g0388(.A(KEYINPUT19), .B1(new_n403), .B2(G97), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n588), .B1(new_n589), .B2(KEYINPUT82), .ZN(new_n590));
  OAI211_X1 g0390(.A(KEYINPUT82), .B(new_n584), .C1(new_n262), .C2(new_n514), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n329), .A2(new_n331), .A3(new_n225), .A4(G68), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n261), .B1(new_n590), .B2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT83), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n252), .A2(new_n435), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n594), .A2(new_n595), .A3(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(new_n598), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n595), .B1(new_n594), .B2(new_n597), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n583), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n224), .B1(G33), .B2(G41), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n461), .A2(G250), .ZN(new_n603));
  INV_X1    g0403(.A(G274), .ZN(new_n604));
  OAI22_X1  g0404(.A1(new_n602), .A2(new_n603), .B1(new_n604), .B2(new_n461), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n329), .A2(new_n331), .A3(G238), .A4(new_n285), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n329), .A2(new_n331), .A3(G244), .A4(G1698), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n606), .A2(new_n607), .A3(new_n489), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n605), .B1(new_n608), .B2(new_n282), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n609), .A2(G169), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n610), .B1(new_n431), .B2(new_n609), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n480), .A2(new_n586), .ZN(new_n612));
  AND2_X1   g0412(.A1(new_n591), .A2(new_n592), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n584), .B1(new_n262), .B2(new_n514), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT82), .ZN(new_n615));
  AOI22_X1  g0415(.A1(new_n614), .A2(new_n615), .B1(new_n585), .B2(new_n587), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n270), .B1(new_n613), .B2(new_n616), .ZN(new_n617));
  OAI21_X1  g0417(.A(KEYINPUT83), .B1(new_n617), .B2(new_n596), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n612), .B1(new_n618), .B2(new_n598), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n609), .A2(new_n316), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n620), .B1(G190), .B2(new_n609), .ZN(new_n621));
  AOI22_X1  g0421(.A1(new_n601), .A2(new_n611), .B1(new_n619), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n575), .A2(G200), .ZN(new_n623));
  OAI21_X1  g0423(.A(G190), .B1(new_n577), .B2(new_n579), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n561), .A2(new_n563), .A3(new_n623), .A4(new_n624), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n582), .A2(new_n622), .A3(new_n625), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n541), .A2(new_n626), .ZN(new_n627));
  AND2_X1   g0427(.A1(new_n449), .A2(new_n627), .ZN(G372));
  NOR2_X1   g0428(.A1(new_n496), .A2(new_n497), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n484), .A2(new_n482), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n631), .B1(new_n470), .B2(new_n477), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n540), .B1(new_n632), .B2(new_n534), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n633), .A2(new_n626), .ZN(new_n634));
  AND2_X1   g0434(.A1(new_n601), .A2(new_n611), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n622), .A2(new_n564), .A3(new_n581), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n635), .B1(new_n636), .B2(KEYINPUT26), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n575), .A2(new_n578), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n573), .B1(new_n570), .B2(new_n282), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(KEYINPUT81), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n638), .A2(new_n275), .A3(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n576), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  AOI22_X1  g0443(.A1(new_n643), .A2(KEYINPUT87), .B1(new_n561), .B2(new_n563), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT26), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT87), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n641), .A2(new_n646), .A3(new_n642), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n644), .A2(new_n645), .A3(new_n622), .A4(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n637), .A2(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n449), .B1(new_n634), .B2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n425), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n393), .A2(new_n394), .ZN(new_n652));
  AND2_X1   g0452(.A1(new_n313), .A2(new_n441), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n380), .A2(new_n382), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(new_n317), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n652), .B1(new_n653), .B2(new_n655), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n651), .B1(new_n656), .B2(new_n422), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n650), .A2(new_n657), .ZN(new_n658));
  XOR2_X1   g0458(.A(new_n658), .B(KEYINPUT88), .Z(G369));
  INV_X1    g0459(.A(KEYINPUT27), .ZN(new_n660));
  AND2_X1   g0460(.A1(new_n225), .A2(G13), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT89), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n661), .A2(new_n662), .A3(new_n247), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n247), .A2(new_n225), .A3(G13), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(KEYINPUT89), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n660), .B1(new_n663), .B2(new_n665), .ZN(new_n666));
  XNOR2_X1  g0466(.A(new_n666), .B(KEYINPUT91), .ZN(new_n667));
  INV_X1    g0467(.A(G213), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n663), .A2(new_n665), .A3(new_n660), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT90), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n663), .A2(new_n665), .A3(KEYINPUT90), .A4(new_n660), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n668), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n667), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(G343), .ZN(new_n675));
  OR3_X1    g0475(.A1(new_n674), .A2(KEYINPUT92), .A3(new_n675), .ZN(new_n676));
  OAI21_X1  g0476(.A(KEYINPUT92), .B1(new_n674), .B2(new_n675), .ZN(new_n677));
  AND2_X1   g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n678), .A2(new_n519), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(new_n534), .ZN(new_n680));
  INV_X1    g0480(.A(new_n535), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n680), .B1(new_n681), .B2(new_n679), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(G330), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n632), .A2(new_n539), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n676), .A2(new_n677), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(new_n498), .ZN(new_n686));
  AOI22_X1  g0486(.A1(new_n684), .A2(new_n686), .B1(new_n632), .B2(new_n685), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n683), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n684), .A2(new_n534), .A3(new_n678), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n690), .B1(new_n499), .B2(new_n685), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n689), .A2(new_n692), .ZN(G399));
  INV_X1    g0493(.A(new_n219), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n694), .A2(G41), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n587), .A2(G116), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n696), .A2(G1), .A3(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n698), .B1(new_n222), .B2(new_n696), .ZN(new_n699));
  XNOR2_X1  g0499(.A(new_n699), .B(KEYINPUT28), .ZN(new_n700));
  NOR3_X1   g0500(.A1(new_n577), .A2(new_n579), .A3(G169), .ZN(new_n701));
  OAI21_X1  g0501(.A(KEYINPUT87), .B1(new_n701), .B2(new_n576), .ZN(new_n702));
  AND3_X1   g0502(.A1(new_n702), .A2(new_n564), .A3(new_n647), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT95), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n703), .A2(new_n704), .A3(KEYINPUT26), .A4(new_n622), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n702), .A2(new_n622), .A3(new_n564), .A4(new_n647), .ZN(new_n706));
  OAI21_X1  g0506(.A(KEYINPUT95), .B1(new_n706), .B2(new_n645), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n636), .A2(new_n645), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT96), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n636), .A2(KEYINPUT96), .A3(new_n645), .ZN(new_n711));
  AND4_X1   g0511(.A1(new_n705), .A2(new_n707), .A3(new_n710), .A4(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n635), .ZN(new_n713));
  AND3_X1   g0513(.A1(new_n582), .A2(KEYINPUT97), .A3(new_n625), .ZN(new_n714));
  AOI21_X1  g0514(.A(KEYINPUT97), .B1(new_n582), .B2(new_n625), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  OAI211_X1 g0516(.A(new_n540), .B(new_n622), .C1(new_n632), .C2(new_n534), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n713), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  OAI211_X1 g0518(.A(KEYINPUT29), .B(new_n678), .C1(new_n712), .C2(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n678), .B1(new_n649), .B2(new_n634), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT29), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n719), .A2(new_n722), .ZN(new_n723));
  AND3_X1   g0523(.A1(new_n582), .A2(new_n622), .A3(new_n625), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n724), .A2(new_n535), .A3(new_n684), .A4(new_n678), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT30), .ZN(new_n726));
  OAI211_X1 g0526(.A(new_n532), .B(new_n609), .C1(new_n467), .C2(new_n468), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n726), .B1(new_n580), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n638), .A2(new_n640), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n609), .A2(new_n504), .A3(G179), .A4(new_n506), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n730), .B1(new_n473), .B2(new_n474), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n729), .A2(KEYINPUT30), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n728), .A2(new_n732), .ZN(new_n733));
  NOR3_X1   g0533(.A1(new_n525), .A2(G179), .A3(new_n609), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(KEYINPUT93), .B1(new_n475), .B2(new_n639), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT93), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n536), .A2(new_n737), .A3(new_n575), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n735), .B1(new_n736), .B2(new_n738), .ZN(new_n739));
  OAI211_X1 g0539(.A(KEYINPUT31), .B(new_n685), .C1(new_n733), .C2(new_n739), .ZN(new_n740));
  NOR3_X1   g0540(.A1(new_n475), .A2(KEYINPUT93), .A3(new_n639), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n737), .B1(new_n536), .B2(new_n575), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n734), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n733), .B1(new_n743), .B2(KEYINPUT94), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT94), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n739), .A2(new_n745), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n678), .B1(new_n744), .B2(new_n746), .ZN(new_n747));
  OAI211_X1 g0547(.A(new_n725), .B(new_n740), .C1(new_n747), .C2(KEYINPUT31), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(G330), .ZN(new_n749));
  AND2_X1   g0549(.A1(new_n723), .A2(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n700), .B1(new_n750), .B2(G1), .ZN(G364));
  AOI21_X1  g0551(.A(new_n247), .B1(new_n661), .B2(G45), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n753), .A2(new_n695), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n754), .B1(new_n682), .B2(G330), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n755), .B1(G330), .B2(new_n682), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n694), .A2(new_n332), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(G355), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n758), .B1(G116), .B2(new_n219), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n694), .A2(new_n284), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n761), .B1(new_n293), .B2(new_n223), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n245), .A2(G45), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n759), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(G13), .A2(G33), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(G20), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n224), .B1(G20), .B2(new_n275), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n754), .B1(new_n764), .B2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n225), .A2(new_n369), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n431), .A2(G200), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n316), .A2(G179), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n772), .A2(new_n775), .ZN(new_n776));
  OAI22_X1  g0576(.A1(new_n201), .A2(new_n774), .B1(new_n776), .B2(new_n586), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n225), .A2(G190), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n778), .A2(G179), .A3(G200), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  AOI211_X1 g0580(.A(new_n332), .B(new_n777), .C1(G68), .C2(new_n780), .ZN(new_n781));
  NOR4_X1   g0581(.A1(new_n225), .A2(new_n431), .A3(new_n369), .A4(new_n316), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n775), .A2(new_n778), .ZN(new_n784));
  OAI22_X1  g0584(.A1(new_n783), .A2(new_n266), .B1(new_n784), .B2(new_n487), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n778), .A2(new_n773), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n785), .B1(G77), .B2(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(G179), .A2(G200), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n225), .B1(new_n789), .B2(G190), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(G97), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n778), .A2(new_n789), .ZN(new_n793));
  INV_X1    g0593(.A(G159), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  XNOR2_X1  g0595(.A(KEYINPUT98), .B(KEYINPUT32), .ZN(new_n796));
  XNOR2_X1  g0596(.A(new_n795), .B(new_n796), .ZN(new_n797));
  NAND4_X1  g0597(.A1(new_n781), .A2(new_n788), .A3(new_n792), .A4(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(G283), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n332), .B1(new_n784), .B2(new_n799), .ZN(new_n800));
  XOR2_X1   g0600(.A(KEYINPUT33), .B(G317), .Z(new_n801));
  NOR2_X1   g0601(.A1(new_n801), .A2(new_n779), .ZN(new_n802));
  AOI211_X1 g0602(.A(new_n800), .B(new_n802), .C1(G311), .C2(new_n787), .ZN(new_n803));
  XOR2_X1   g0603(.A(KEYINPUT99), .B(G326), .Z(new_n804));
  AOI22_X1  g0604(.A1(new_n782), .A2(new_n804), .B1(new_n791), .B2(G294), .ZN(new_n805));
  OR2_X1    g0605(.A1(new_n805), .A2(KEYINPUT100), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n805), .A2(KEYINPUT100), .ZN(new_n807));
  INV_X1    g0607(.A(G322), .ZN(new_n808));
  INV_X1    g0608(.A(G329), .ZN(new_n809));
  OAI22_X1  g0609(.A1(new_n774), .A2(new_n808), .B1(new_n793), .B2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n776), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n810), .B1(G303), .B2(new_n811), .ZN(new_n812));
  NAND4_X1  g0612(.A1(new_n803), .A2(new_n806), .A3(new_n807), .A4(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n798), .A2(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n771), .B1(new_n814), .B2(new_n768), .ZN(new_n815));
  INV_X1    g0615(.A(new_n767), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n815), .B1(new_n682), .B2(new_n816), .ZN(new_n817));
  AND2_X1   g0617(.A1(new_n756), .A2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(G396));
  INV_X1    g0619(.A(new_n440), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n820), .B1(new_n676), .B2(new_n677), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n441), .B1(new_n821), .B2(new_n445), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n678), .A2(new_n442), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n720), .A2(new_n824), .ZN(new_n825));
  AND2_X1   g0625(.A1(new_n822), .A2(new_n823), .ZN(new_n826));
  OAI211_X1 g0626(.A(new_n678), .B(new_n826), .C1(new_n649), .C2(new_n634), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n754), .B1(new_n828), .B2(new_n749), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n829), .B1(new_n749), .B2(new_n828), .ZN(new_n830));
  INV_X1    g0630(.A(new_n754), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n768), .A2(new_n765), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n831), .B1(new_n205), .B2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n768), .ZN(new_n834));
  AOI22_X1  g0634(.A1(G137), .A2(new_n782), .B1(new_n787), .B2(G159), .ZN(new_n835));
  INV_X1    g0635(.A(G143), .ZN(new_n836));
  INV_X1    g0636(.A(G150), .ZN(new_n837));
  OAI221_X1 g0637(.A(new_n835), .B1(new_n836), .B2(new_n774), .C1(new_n837), .C2(new_n779), .ZN(new_n838));
  XNOR2_X1  g0638(.A(new_n838), .B(KEYINPUT34), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n284), .B1(new_n776), .B2(new_n266), .ZN(new_n840));
  INV_X1    g0640(.A(new_n784), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(G68), .ZN(new_n842));
  INV_X1    g0642(.A(G132), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n842), .B1(new_n843), .B2(new_n793), .ZN(new_n844));
  AOI211_X1 g0644(.A(new_n840), .B(new_n844), .C1(G58), .C2(new_n791), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n784), .A2(new_n586), .ZN(new_n846));
  INV_X1    g0646(.A(new_n793), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n846), .B1(G311), .B2(new_n847), .ZN(new_n848));
  XNOR2_X1  g0648(.A(new_n848), .B(KEYINPUT101), .ZN(new_n849));
  AOI22_X1  g0649(.A1(G283), .A2(new_n780), .B1(new_n811), .B2(G107), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n850), .B1(new_n502), .B2(new_n783), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n332), .B1(new_n786), .B2(new_n511), .ZN(new_n852));
  NOR3_X1   g0652(.A1(new_n849), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(G294), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n792), .B1(new_n854), .B2(new_n774), .ZN(new_n855));
  XNOR2_X1  g0655(.A(new_n855), .B(KEYINPUT102), .ZN(new_n856));
  AOI22_X1  g0656(.A1(new_n839), .A2(new_n845), .B1(new_n853), .B2(new_n856), .ZN(new_n857));
  OAI221_X1 g0657(.A(new_n833), .B1(new_n834), .B2(new_n857), .C1(new_n826), .C2(new_n766), .ZN(new_n858));
  AND2_X1   g0658(.A1(new_n830), .A2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(G384));
  INV_X1    g0660(.A(G330), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT31), .ZN(new_n862));
  OAI211_X1 g0662(.A(new_n728), .B(new_n732), .C1(new_n739), .C2(new_n745), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n743), .A2(KEYINPUT94), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n685), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  AOI22_X1  g0665(.A1(new_n862), .A2(new_n865), .B1(new_n627), .B2(new_n678), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n747), .A2(KEYINPUT31), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n861), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(new_n449), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n865), .A2(new_n862), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n867), .A2(new_n870), .A3(new_n725), .ZN(new_n871));
  AND3_X1   g0671(.A1(new_n360), .A2(new_n378), .A3(new_n381), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n381), .B1(new_n360), .B2(new_n378), .ZN(new_n873));
  AND3_X1   g0673(.A1(new_n388), .A2(KEYINPUT18), .A3(new_n390), .ZN(new_n874));
  AOI21_X1  g0674(.A(KEYINPUT18), .B1(new_n388), .B2(new_n390), .ZN(new_n875));
  OAI22_X1  g0675(.A1(new_n872), .A2(new_n873), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n674), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n348), .B1(new_n356), .B2(new_n357), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n878), .A2(new_n385), .A3(new_n261), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(new_n325), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n876), .A2(new_n877), .A3(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT103), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT37), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n880), .B1(new_n390), .B2(new_n877), .ZN(new_n884));
  AOI211_X1 g0684(.A(new_n882), .B(new_n883), .C1(new_n379), .C2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n388), .A2(new_n877), .ZN(new_n886));
  NAND4_X1  g0686(.A1(new_n379), .A2(new_n391), .A3(new_n886), .A4(new_n883), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n883), .B1(new_n379), .B2(new_n884), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n887), .B1(new_n888), .B2(KEYINPUT103), .ZN(new_n889));
  OAI211_X1 g0689(.A(new_n881), .B(KEYINPUT38), .C1(new_n885), .C2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT38), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n379), .A2(new_n391), .A3(new_n886), .ZN(new_n892));
  XNOR2_X1  g0692(.A(new_n892), .B(new_n883), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n886), .B1(new_n654), .B2(new_n652), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n891), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n890), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n274), .A2(new_n685), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n313), .A2(new_n317), .A3(new_n897), .ZN(new_n898));
  OAI211_X1 g0698(.A(new_n274), .B(new_n685), .C1(new_n310), .C2(new_n312), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n824), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n871), .A2(new_n896), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n898), .A2(new_n899), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(new_n826), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n903), .B1(new_n866), .B2(new_n867), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n880), .A2(new_n877), .ZN(new_n905));
  OAI22_X1  g0705(.A1(new_n889), .A2(new_n885), .B1(new_n395), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(new_n891), .ZN(new_n907));
  AOI21_X1  g0707(.A(KEYINPUT40), .B1(new_n907), .B2(new_n890), .ZN(new_n908));
  AOI22_X1  g0708(.A1(new_n901), .A2(KEYINPUT40), .B1(new_n904), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n869), .B1(new_n909), .B2(new_n861), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n725), .B1(new_n747), .B2(KEYINPUT31), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n865), .A2(new_n862), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n900), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  AND2_X1   g0713(.A1(new_n890), .A2(new_n895), .ZN(new_n914));
  OAI21_X1  g0714(.A(KEYINPUT40), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n904), .A2(new_n908), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n917), .A2(new_n449), .A3(new_n871), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n910), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n719), .A2(new_n449), .A3(new_n722), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(new_n657), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n919), .B(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n827), .A2(new_n823), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n902), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n906), .A2(new_n891), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n379), .A2(new_n884), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(KEYINPUT37), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(new_n882), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n888), .A2(KEYINPUT103), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n928), .A2(new_n929), .A3(new_n887), .ZN(new_n930));
  AOI21_X1  g0730(.A(KEYINPUT38), .B1(new_n930), .B2(new_n881), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n925), .A2(new_n931), .ZN(new_n932));
  OAI22_X1  g0732(.A1(new_n924), .A2(new_n932), .B1(new_n652), .B2(new_n877), .ZN(new_n933));
  INV_X1    g0733(.A(new_n933), .ZN(new_n934));
  OR2_X1    g0734(.A1(new_n313), .A2(new_n685), .ZN(new_n935));
  INV_X1    g0735(.A(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT39), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n890), .A2(new_n895), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n937), .B1(new_n907), .B2(new_n890), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT104), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n938), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  AOI211_X1 g0741(.A(KEYINPUT104), .B(new_n937), .C1(new_n907), .C2(new_n890), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n936), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n934), .A2(new_n943), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n944), .B(KEYINPUT105), .ZN(new_n945));
  OAI22_X1  g0745(.A1(new_n922), .A2(new_n945), .B1(new_n247), .B2(new_n661), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n946), .B1(new_n922), .B2(new_n945), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n552), .A2(new_n553), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT35), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n552), .A2(KEYINPUT35), .A3(new_n553), .ZN(new_n951));
  NAND4_X1  g0751(.A1(new_n950), .A2(G116), .A3(new_n226), .A4(new_n951), .ZN(new_n952));
  XOR2_X1   g0752(.A(new_n952), .B(KEYINPUT36), .Z(new_n953));
  NAND3_X1  g0753(.A1(new_n223), .A2(G77), .A3(new_n351), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n266), .A2(G68), .ZN(new_n955));
  AOI211_X1 g0755(.A(new_n247), .B(G13), .C1(new_n954), .C2(new_n955), .ZN(new_n956));
  OR3_X1    g0756(.A1(new_n947), .A2(new_n953), .A3(new_n956), .ZN(G367));
  OR2_X1    g0757(.A1(new_n678), .A2(new_n619), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n958), .B(new_n622), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(KEYINPUT106), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT43), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT106), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n959), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n961), .A2(new_n962), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n582), .A2(new_n625), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT97), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n582), .A2(KEYINPUT97), .A3(new_n625), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n685), .A2(new_n564), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n703), .A2(new_n685), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n974), .A2(new_n632), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n685), .B1(new_n975), .B2(new_n582), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n716), .A2(new_n690), .ZN(new_n977));
  XOR2_X1   g0777(.A(new_n977), .B(KEYINPUT42), .Z(new_n978));
  OAI221_X1 g0778(.A(new_n965), .B1(new_n962), .B2(new_n960), .C1(new_n976), .C2(new_n978), .ZN(new_n979));
  OR3_X1    g0779(.A1(new_n976), .A2(new_n978), .A3(new_n965), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(new_n974), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n689), .A2(new_n982), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n981), .B(new_n983), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n695), .B(KEYINPUT41), .ZN(new_n985));
  INV_X1    g0785(.A(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n974), .A2(new_n692), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n987), .A2(KEYINPUT45), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n972), .A2(new_n691), .A3(new_n973), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT44), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n990), .A2(KEYINPUT107), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n988), .A2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT45), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n974), .A2(new_n994), .A3(new_n692), .ZN(new_n995));
  XNOR2_X1  g0795(.A(KEYINPUT107), .B(KEYINPUT44), .ZN(new_n996));
  NAND4_X1  g0796(.A1(new_n972), .A2(new_n691), .A3(new_n973), .A4(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  NOR3_X1   g0798(.A1(new_n993), .A2(new_n688), .A3(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(new_n998), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(new_n987), .A2(KEYINPUT45), .B1(new_n989), .B2(new_n991), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n689), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n999), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n678), .A2(new_n534), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n687), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1005), .A2(new_n690), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n688), .B1(new_n1006), .B2(new_n683), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n723), .A2(new_n1007), .A3(new_n749), .ZN(new_n1008));
  OR2_X1    g0808(.A1(new_n1008), .A2(KEYINPUT108), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(KEYINPUT108), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1003), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n986), .B1(new_n1011), .B2(new_n750), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n984), .B1(new_n1012), .B2(new_n753), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n237), .A2(new_n761), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n769), .B1(new_n219), .B2(new_n436), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n754), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n332), .B1(new_n774), .B2(new_n502), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(KEYINPUT109), .B(G317), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n786), .A2(new_n799), .B1(new_n793), .B2(new_n1018), .ZN(new_n1019));
  AOI211_X1 g0819(.A(new_n1017), .B(new_n1019), .C1(G107), .C2(new_n791), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n811), .A2(G116), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT46), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n782), .A2(G311), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(G294), .A2(new_n780), .B1(new_n841), .B2(G97), .ZN(new_n1024));
  NAND4_X1  g0824(.A1(new_n1020), .A2(new_n1022), .A3(new_n1023), .A4(new_n1024), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1025), .B(KEYINPUT110), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n774), .A2(new_n837), .B1(new_n786), .B2(new_n266), .ZN(new_n1027));
  AOI211_X1 g0827(.A(new_n332), .B(new_n1027), .C1(G58), .C2(new_n811), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(G159), .A2(new_n780), .B1(new_n841), .B2(G77), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(new_n782), .A2(G143), .B1(new_n847), .B2(G137), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n791), .A2(G68), .ZN(new_n1031));
  NAND4_X1  g0831(.A1(new_n1028), .A2(new_n1029), .A3(new_n1030), .A4(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1026), .A2(new_n1032), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(KEYINPUT111), .B(KEYINPUT47), .ZN(new_n1034));
  OR2_X1    g0834(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n834), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1016), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1037), .B1(new_n959), .B2(new_n816), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1013), .A2(new_n1038), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n1039), .A2(KEYINPUT112), .ZN(new_n1040));
  INV_X1    g0840(.A(KEYINPUT112), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1041), .B1(new_n1013), .B2(new_n1038), .ZN(new_n1042));
  OR2_X1    g0842(.A1(new_n1040), .A2(new_n1042), .ZN(G387));
  OAI22_X1  g0843(.A1(new_n776), .A2(new_n205), .B1(new_n786), .B2(new_n202), .ZN(new_n1044));
  AOI211_X1 g0844(.A(new_n332), .B(new_n1044), .C1(G97), .C2(new_n841), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n791), .A2(new_n435), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n321), .A2(new_n780), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n774), .A2(new_n266), .B1(new_n793), .B2(new_n837), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1048), .B1(G159), .B2(new_n782), .ZN(new_n1049));
  NAND4_X1  g0849(.A1(new_n1045), .A2(new_n1046), .A3(new_n1047), .A4(new_n1049), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n847), .A2(new_n804), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n284), .B1(new_n841), .B2(G116), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(G311), .A2(new_n780), .B1(new_n782), .B2(G322), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n1053), .B1(new_n502), .B2(new_n786), .C1(new_n774), .C2(new_n1018), .ZN(new_n1054));
  XOR2_X1   g0854(.A(new_n1054), .B(KEYINPUT48), .Z(new_n1055));
  OAI22_X1  g0855(.A1(new_n776), .A2(new_n854), .B1(new_n790), .B2(new_n799), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n1051), .B(new_n1052), .C1(new_n1057), .C2(KEYINPUT49), .ZN(new_n1058));
  AND2_X1   g0858(.A1(new_n1057), .A2(KEYINPUT49), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1050), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1060), .A2(new_n768), .ZN(new_n1061));
  OR2_X1    g0861(.A1(new_n234), .A2(new_n293), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n697), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n1062), .A2(new_n760), .B1(new_n1063), .B2(new_n757), .ZN(new_n1064));
  AOI21_X1  g0864(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1065));
  OR2_X1    g0865(.A1(new_n319), .A2(G50), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n697), .B(new_n1065), .C1(new_n1066), .C2(KEYINPUT50), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1067), .B1(KEYINPUT50), .B2(new_n1066), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n1064), .A2(new_n1068), .B1(G107), .B2(new_n219), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n831), .B1(new_n1069), .B2(new_n769), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1061), .A2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1071), .B1(new_n687), .B2(new_n767), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1072), .B1(new_n1007), .B2(new_n753), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n750), .A2(new_n1007), .ZN(new_n1074));
  XOR2_X1   g0874(.A(new_n695), .B(KEYINPUT113), .Z(new_n1075));
  INV_X1    g0875(.A(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1008), .A2(new_n1076), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1073), .B1(new_n1074), .B2(new_n1077), .ZN(G393));
  NOR2_X1   g0878(.A1(new_n242), .A2(new_n761), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n769), .B1(new_n514), .B2(new_n219), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(G50), .A2(new_n780), .B1(new_n811), .B2(G68), .ZN(new_n1081));
  OAI221_X1 g0881(.A(new_n1081), .B1(new_n836), .B2(new_n793), .C1(new_n319), .C2(new_n786), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n790), .A2(new_n205), .ZN(new_n1083));
  NOR4_X1   g0883(.A1(new_n1082), .A2(new_n332), .A3(new_n846), .A4(new_n1083), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n783), .A2(new_n837), .B1(new_n774), .B2(new_n794), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n1085), .B(KEYINPUT51), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n332), .B1(new_n790), .B2(new_n511), .C1(new_n487), .C2(new_n784), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n502), .A2(new_n779), .B1(new_n776), .B2(new_n799), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n786), .A2(new_n854), .B1(new_n793), .B2(new_n808), .ZN(new_n1089));
  NOR3_X1   g0889(.A1(new_n1087), .A2(new_n1088), .A3(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n774), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n1091), .A2(G311), .B1(new_n782), .B2(G317), .ZN(new_n1092));
  XOR2_X1   g0892(.A(KEYINPUT115), .B(KEYINPUT52), .Z(new_n1093));
  XNOR2_X1  g0893(.A(new_n1092), .B(new_n1093), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n1084), .A2(new_n1086), .B1(new_n1090), .B2(new_n1094), .ZN(new_n1095));
  OAI221_X1 g0895(.A(new_n754), .B1(new_n1079), .B2(new_n1080), .C1(new_n1095), .C2(new_n834), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1096), .B1(new_n982), .B2(new_n767), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n688), .B1(new_n993), .B2(new_n998), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1000), .A2(new_n1001), .A3(new_n689), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(KEYINPUT114), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n752), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1003), .A2(KEYINPUT114), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1097), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1075), .B1(new_n1100), .B2(new_n1008), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1011), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1104), .A2(new_n1106), .ZN(G390));
  NAND3_X1  g0907(.A1(new_n748), .A2(G330), .A3(new_n826), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n902), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n868), .A2(new_n900), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n923), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n902), .B1(new_n868), .B2(new_n826), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n678), .B(new_n822), .C1(new_n712), .C2(new_n718), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n748), .A2(G330), .A3(new_n900), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1113), .A2(new_n823), .A3(new_n1114), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n1110), .A2(new_n1111), .B1(new_n1112), .B2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n920), .A2(new_n657), .A3(new_n869), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n924), .A2(new_n935), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n939), .A2(new_n940), .ZN(new_n1121));
  OAI21_X1  g0921(.A(KEYINPUT39), .B1(new_n925), .B2(new_n931), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(KEYINPUT104), .ZN(new_n1123));
  NAND4_X1  g0923(.A1(new_n1120), .A2(new_n1121), .A3(new_n1123), .A4(new_n938), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(new_n935), .B(KEYINPUT116), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1125), .A2(new_n896), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n717), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n635), .B1(new_n970), .B2(new_n1128), .ZN(new_n1129));
  NAND4_X1  g0929(.A1(new_n705), .A2(new_n710), .A3(new_n707), .A4(new_n711), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n685), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n1131), .A2(new_n822), .B1(new_n442), .B2(new_n678), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1127), .B1(new_n1132), .B2(new_n1109), .ZN(new_n1133));
  AND3_X1   g0933(.A1(new_n1124), .A2(new_n1133), .A3(new_n1114), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n871), .A2(G330), .A3(new_n900), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1135), .B1(new_n1124), .B2(new_n1133), .ZN(new_n1136));
  OAI211_X1 g0936(.A(KEYINPUT117), .B(new_n1119), .C1(new_n1134), .C2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1124), .A2(new_n1133), .A3(new_n1114), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1135), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n936), .B1(new_n923), .B2(new_n902), .ZN(new_n1140));
  NOR3_X1   g0940(.A1(new_n941), .A2(new_n1140), .A3(new_n942), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1113), .A2(new_n823), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1126), .B1(new_n1142), .B2(new_n902), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1139), .B1(new_n1141), .B2(new_n1143), .ZN(new_n1144));
  AND2_X1   g0944(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n923), .B1(new_n1145), .B2(new_n1139), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n871), .A2(G330), .A3(new_n826), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1147), .A2(new_n1109), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1148), .A2(new_n1132), .A3(new_n1114), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1117), .B1(new_n1146), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(KEYINPUT117), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n1138), .B(new_n1144), .C1(new_n1150), .C2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1137), .A2(new_n1076), .A3(new_n1152), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1144), .A2(new_n753), .A3(new_n1138), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n832), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n754), .B1(new_n321), .B2(new_n1155), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n776), .A2(new_n837), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(new_n1157), .B(KEYINPUT53), .ZN(new_n1158));
  XOR2_X1   g0958(.A(KEYINPUT54), .B(G143), .Z(new_n1159));
  AOI22_X1  g0959(.A1(new_n787), .A2(new_n1159), .B1(new_n841), .B2(G50), .ZN(new_n1160));
  INV_X1    g0960(.A(G128), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n1158), .B(new_n1160), .C1(new_n1161), .C2(new_n783), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(G137), .A2(new_n780), .B1(new_n1091), .B2(G132), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n332), .B1(new_n847), .B2(G125), .ZN(new_n1164));
  OAI211_X1 g0964(.A(new_n1163), .B(new_n1164), .C1(new_n794), .C2(new_n790), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(G283), .A2(new_n782), .B1(new_n787), .B2(G97), .ZN(new_n1166));
  OAI221_X1 g0966(.A(new_n1166), .B1(new_n487), .B2(new_n779), .C1(new_n511), .C2(new_n774), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n284), .B1(new_n811), .B2(G87), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1083), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n847), .A2(G294), .ZN(new_n1170));
  NAND4_X1  g0970(.A1(new_n1168), .A2(new_n842), .A3(new_n1169), .A4(new_n1170), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n1162), .A2(new_n1165), .B1(new_n1167), .B2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1156), .B1(new_n1172), .B2(new_n768), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1123), .A2(new_n1121), .A3(new_n938), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1173), .B1(new_n1174), .B2(new_n766), .ZN(new_n1175));
  AND2_X1   g0975(.A1(new_n1154), .A2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1153), .A2(new_n1176), .ZN(G378));
  NAND3_X1  g0977(.A1(new_n1144), .A2(new_n1138), .A3(new_n1116), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n877), .A2(new_n424), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n422), .A2(new_n425), .A3(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1181), .B1(new_n422), .B2(new_n425), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1180), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1184), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1186), .A2(new_n1182), .A3(new_n1179), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1185), .A2(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1188), .B1(new_n917), .B2(G330), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1188), .ZN(new_n1190));
  AOI211_X1 g0990(.A(new_n861), .B(new_n1190), .C1(new_n915), .C2(new_n916), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n944), .B1(new_n1189), .B2(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n933), .B1(new_n1174), .B2(new_n936), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1190), .B1(new_n909), .B2(new_n861), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n917), .A2(G330), .A3(new_n1188), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1193), .A2(new_n1194), .A3(new_n1195), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(new_n1178), .A2(new_n1118), .B1(new_n1192), .B2(new_n1196), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1076), .B1(new_n1197), .B2(KEYINPUT57), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1178), .A2(new_n1118), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1192), .A2(new_n1196), .ZN(new_n1200));
  AND3_X1   g1000(.A1(new_n1199), .A2(KEYINPUT57), .A3(new_n1200), .ZN(new_n1201));
  OR2_X1    g1001(.A1(new_n1198), .A2(new_n1201), .ZN(new_n1202));
  AND3_X1   g1002(.A1(new_n1193), .A2(new_n1195), .A3(new_n1194), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n1194), .A2(new_n1195), .B1(new_n943), .B2(new_n934), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n753), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n831), .B1(new_n266), .B2(new_n832), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(G97), .A2(new_n780), .B1(new_n1091), .B2(G107), .ZN(new_n1207));
  OAI221_X1 g1007(.A(new_n1207), .B1(new_n799), .B2(new_n793), .C1(new_n436), .C2(new_n786), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n790), .A2(new_n202), .ZN(new_n1209));
  OAI211_X1 g1009(.A(new_n292), .B(new_n332), .C1(new_n776), .C2(new_n205), .ZN(new_n1210));
  OAI22_X1  g1010(.A1(new_n783), .A2(new_n511), .B1(new_n784), .B2(new_n201), .ZN(new_n1211));
  NOR4_X1   g1011(.A1(new_n1208), .A2(new_n1209), .A3(new_n1210), .A4(new_n1211), .ZN(new_n1212));
  XOR2_X1   g1012(.A(new_n1212), .B(KEYINPUT58), .Z(new_n1213));
  AOI21_X1  g1013(.A(G50), .B1(new_n264), .B2(new_n292), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1214), .B1(new_n284), .B2(G41), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(G128), .A2(new_n1091), .B1(new_n811), .B2(new_n1159), .ZN(new_n1216));
  INV_X1    g1016(.A(G125), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1216), .B1(new_n1217), .B2(new_n783), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(G132), .A2(new_n780), .B1(new_n787), .B2(G137), .ZN(new_n1219));
  XNOR2_X1  g1019(.A(new_n1219), .B(KEYINPUT118), .ZN(new_n1220));
  AOI211_X1 g1020(.A(new_n1218), .B(new_n1220), .C1(G150), .C2(new_n791), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1222), .A2(KEYINPUT59), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n264), .B(new_n292), .C1(new_n784), .C2(new_n794), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1224), .B1(G124), .B2(new_n847), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT59), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1225), .B1(new_n1221), .B2(new_n1226), .ZN(new_n1227));
  OAI211_X1 g1027(.A(new_n1213), .B(new_n1215), .C1(new_n1223), .C2(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT119), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1231), .A2(new_n768), .ZN(new_n1232));
  OAI221_X1 g1032(.A(new_n1206), .B1(new_n1230), .B2(new_n1232), .C1(new_n1188), .C2(new_n766), .ZN(new_n1233));
  AND2_X1   g1033(.A1(new_n1205), .A2(new_n1233), .ZN(new_n1234));
  AND2_X1   g1034(.A1(new_n1202), .A2(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1235), .ZN(G375));
  AOI21_X1  g1036(.A(new_n752), .B1(new_n1146), .B2(new_n1149), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n831), .B1(new_n202), .B2(new_n832), .ZN(new_n1238));
  OAI22_X1  g1038(.A1(new_n514), .A2(new_n776), .B1(new_n774), .B2(new_n799), .ZN(new_n1239));
  AOI211_X1 g1039(.A(new_n284), .B(new_n1239), .C1(G77), .C2(new_n841), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(G107), .A2(new_n787), .B1(new_n847), .B2(G303), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(G116), .A2(new_n780), .B1(new_n782), .B2(G294), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1240), .A2(new_n1046), .A3(new_n1241), .A4(new_n1242), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n284), .B1(new_n784), .B2(new_n201), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1244), .B1(G50), .B2(new_n791), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(G132), .A2(new_n782), .B1(new_n787), .B2(G150), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(new_n780), .A2(new_n1159), .B1(new_n1091), .B2(G137), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1245), .A2(new_n1246), .A3(new_n1247), .ZN(new_n1248));
  OAI22_X1  g1048(.A1(new_n776), .A2(new_n794), .B1(new_n793), .B2(new_n1161), .ZN(new_n1249));
  XNOR2_X1  g1049(.A(new_n1249), .B(KEYINPUT120), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1243), .B1(new_n1248), .B2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1251), .ZN(new_n1252));
  AND2_X1   g1052(.A1(new_n1252), .A2(KEYINPUT121), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n768), .B1(new_n1252), .B2(KEYINPUT121), .ZN(new_n1254));
  OAI221_X1 g1054(.A(new_n1238), .B1(new_n1253), .B2(new_n1254), .C1(new_n902), .C2(new_n766), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1255), .ZN(new_n1256));
  OR3_X1    g1056(.A1(new_n1237), .A2(KEYINPUT122), .A3(new_n1256), .ZN(new_n1257));
  OAI21_X1  g1057(.A(KEYINPUT122), .B1(new_n1237), .B2(new_n1256), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1116), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1260), .A2(new_n1117), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1261), .A2(new_n985), .A3(new_n1119), .ZN(new_n1262));
  AND2_X1   g1062(.A1(new_n1259), .A2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1263), .ZN(G381));
  AOI21_X1  g1064(.A(KEYINPUT123), .B1(new_n1153), .B2(new_n1176), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1153), .A2(KEYINPUT123), .A3(new_n1176), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1235), .B1(new_n1265), .B2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(G390), .ZN(new_n1269));
  NOR3_X1   g1069(.A1(G393), .A2(G384), .A3(G396), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1263), .A2(new_n1269), .A3(new_n1270), .ZN(new_n1271));
  OR3_X1    g1071(.A1(new_n1268), .A2(G387), .A3(new_n1271), .ZN(G407));
  OAI211_X1 g1072(.A(G407), .B(G213), .C1(G343), .C2(new_n1268), .ZN(G409));
  OAI21_X1  g1073(.A(new_n1269), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1274));
  AND3_X1   g1074(.A1(new_n1013), .A2(new_n1038), .A3(G390), .ZN(new_n1275));
  XNOR2_X1  g1075(.A(G393), .B(new_n818), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1274), .A2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT125), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1039), .A2(new_n1269), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1013), .A2(new_n1038), .A3(G390), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1279), .B1(new_n1282), .B2(new_n1276), .ZN(new_n1283));
  AOI21_X1  g1083(.A(G390), .B1(new_n1013), .B2(new_n1038), .ZN(new_n1284));
  OAI211_X1 g1084(.A(new_n1279), .B(new_n1276), .C1(new_n1275), .C2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1285), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1278), .B1(new_n1283), .B2(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT127), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  OAI211_X1 g1089(.A(new_n1278), .B(KEYINPUT127), .C1(new_n1283), .C2(new_n1286), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT62), .ZN(new_n1292));
  NOR2_X1   g1092(.A1(new_n668), .A2(G343), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT124), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1197), .A2(new_n1295), .A3(new_n985), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1205), .A2(new_n1233), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1199), .A2(new_n985), .A3(new_n1200), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1297), .B1(KEYINPUT124), .B2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT123), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(G378), .A2(new_n1300), .ZN(new_n1301));
  AOI22_X1  g1101(.A1(new_n1296), .A2(new_n1299), .B1(new_n1301), .B2(new_n1266), .ZN(new_n1302));
  OAI211_X1 g1102(.A(G378), .B(new_n1234), .C1(new_n1198), .C2(new_n1201), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1303), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1294), .B1(new_n1302), .B2(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1305), .A2(KEYINPUT126), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1298), .A2(KEYINPUT124), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1307), .A2(new_n1234), .A3(new_n1296), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1308), .B1(new_n1265), .B2(new_n1267), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1309), .A2(new_n1303), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT126), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1310), .A2(new_n1311), .A3(new_n1294), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1306), .A2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT60), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1261), .A2(new_n1314), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1260), .A2(KEYINPUT60), .A3(new_n1117), .ZN(new_n1316));
  NOR2_X1   g1116(.A1(new_n1150), .A2(new_n1075), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1315), .A2(new_n1316), .A3(new_n1317), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1259), .A2(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1319), .A2(new_n859), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1259), .A2(new_n1318), .A3(G384), .ZN(new_n1321));
  AND2_X1   g1121(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1292), .B1(new_n1313), .B2(new_n1322), .ZN(new_n1323));
  AND2_X1   g1123(.A1(new_n1293), .A2(G2897), .ZN(new_n1324));
  XNOR2_X1  g1124(.A(new_n1322), .B(new_n1324), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1306), .A2(new_n1312), .A3(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1327));
  AOI211_X1 g1127(.A(new_n1327), .B(new_n1293), .C1(new_n1309), .C2(new_n1303), .ZN(new_n1328));
  AOI21_X1  g1128(.A(KEYINPUT61), .B1(new_n1328), .B2(new_n1292), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1326), .A2(new_n1329), .ZN(new_n1330));
  OAI21_X1  g1130(.A(new_n1291), .B1(new_n1323), .B2(new_n1330), .ZN(new_n1331));
  XNOR2_X1  g1131(.A(new_n1327), .B(new_n1324), .ZN(new_n1332));
  AOI21_X1  g1132(.A(new_n1332), .B1(new_n1294), .B2(new_n1310), .ZN(new_n1333));
  INV_X1    g1133(.A(KEYINPUT63), .ZN(new_n1334));
  OAI22_X1  g1134(.A1(new_n1333), .A2(new_n1334), .B1(new_n1327), .B2(new_n1305), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1313), .A2(KEYINPUT63), .A3(new_n1322), .ZN(new_n1336));
  INV_X1    g1136(.A(KEYINPUT61), .ZN(new_n1337));
  AND2_X1   g1137(.A1(new_n1287), .A2(new_n1337), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1335), .A2(new_n1336), .A3(new_n1338), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1331), .A2(new_n1339), .ZN(G405));
  NOR2_X1   g1140(.A1(new_n1267), .A2(new_n1265), .ZN(new_n1341));
  OAI21_X1  g1141(.A(new_n1303), .B1(new_n1235), .B2(new_n1341), .ZN(new_n1342));
  XNOR2_X1  g1142(.A(new_n1342), .B(new_n1327), .ZN(new_n1343));
  XNOR2_X1  g1143(.A(new_n1343), .B(new_n1287), .ZN(G402));
endmodule


