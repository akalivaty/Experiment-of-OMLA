

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X2 U555 ( .A1(n551), .A2(n550), .ZN(G164) );
  NOR2_X1 U556 ( .A1(G164), .A2(G1384), .ZN(n697) );
  BUF_X2 U557 ( .A(n619), .Z(n522) );
  NOR2_X1 U558 ( .A1(n715), .A2(n934), .ZN(n717) );
  NAND2_X1 U559 ( .A1(n698), .A2(n815), .ZN(n715) );
  NAND2_X1 U560 ( .A1(n526), .A2(n525), .ZN(n527) );
  INV_X1 U561 ( .A(G2104), .ZN(n526) );
  XOR2_X1 U562 ( .A(KEYINPUT71), .B(n583), .Z(n523) );
  XNOR2_X1 U563 ( .A(KEYINPUT14), .B(n589), .ZN(n524) );
  INV_X1 U564 ( .A(KEYINPUT103), .ZN(n705) );
  INV_X1 U565 ( .A(KEYINPUT29), .ZN(n743) );
  BUF_X1 U566 ( .A(n715), .Z(n748) );
  INV_X1 U567 ( .A(KEYINPUT31), .ZN(n712) );
  XNOR2_X1 U568 ( .A(n713), .B(n712), .ZN(n767) );
  INV_X1 U569 ( .A(KEYINPUT32), .ZN(n763) );
  NOR2_X1 U570 ( .A1(n792), .A2(n791), .ZN(n793) );
  INV_X1 U571 ( .A(G2105), .ZN(n525) );
  AND2_X1 U572 ( .A1(n590), .A2(n524), .ZN(n591) );
  NAND2_X1 U573 ( .A1(n523), .A2(n591), .ZN(n982) );
  XNOR2_X2 U574 ( .A(n527), .B(KEYINPUT17), .ZN(n902) );
  NAND2_X1 U575 ( .A1(n902), .A2(G137), .ZN(n535) );
  INV_X1 U576 ( .A(G2105), .ZN(n529) );
  AND2_X4 U577 ( .A1(n529), .A2(G2104), .ZN(n900) );
  NAND2_X1 U578 ( .A1(G101), .A2(n900), .ZN(n528) );
  XNOR2_X1 U579 ( .A(KEYINPUT23), .B(n528), .ZN(n533) );
  NOR2_X1 U580 ( .A1(G2104), .A2(n529), .ZN(n619) );
  NAND2_X1 U581 ( .A1(G125), .A2(n522), .ZN(n531) );
  AND2_X2 U582 ( .A1(G2105), .A2(G2104), .ZN(n897) );
  NAND2_X1 U583 ( .A1(G113), .A2(n897), .ZN(n530) );
  NAND2_X1 U584 ( .A1(n531), .A2(n530), .ZN(n532) );
  NOR2_X1 U585 ( .A1(n533), .A2(n532), .ZN(n534) );
  AND2_X2 U586 ( .A1(n535), .A2(n534), .ZN(G160) );
  XOR2_X1 U587 ( .A(G2443), .B(G2446), .Z(n537) );
  XNOR2_X1 U588 ( .A(G2427), .B(G2451), .ZN(n536) );
  XNOR2_X1 U589 ( .A(n537), .B(n536), .ZN(n543) );
  XOR2_X1 U590 ( .A(G2430), .B(G2454), .Z(n539) );
  XNOR2_X1 U591 ( .A(G1348), .B(G1341), .ZN(n538) );
  XNOR2_X1 U592 ( .A(n539), .B(n538), .ZN(n541) );
  XOR2_X1 U593 ( .A(G2435), .B(G2438), .Z(n540) );
  XNOR2_X1 U594 ( .A(n541), .B(n540), .ZN(n542) );
  XOR2_X1 U595 ( .A(n543), .B(n542), .Z(n544) );
  AND2_X1 U596 ( .A1(G14), .A2(n544), .ZN(G401) );
  AND2_X1 U597 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U598 ( .A(G57), .ZN(G237) );
  INV_X1 U599 ( .A(G82), .ZN(G220) );
  NAND2_X1 U600 ( .A1(G102), .A2(n900), .ZN(n546) );
  NAND2_X1 U601 ( .A1(G114), .A2(n897), .ZN(n545) );
  AND2_X1 U602 ( .A1(n546), .A2(n545), .ZN(n549) );
  NAND2_X1 U603 ( .A1(n619), .A2(G126), .ZN(n547) );
  XNOR2_X1 U604 ( .A(n547), .B(KEYINPUT90), .ZN(n548) );
  AND2_X1 U605 ( .A1(n549), .A2(n548), .ZN(n551) );
  NAND2_X1 U606 ( .A1(n902), .A2(G138), .ZN(n550) );
  NOR2_X2 U607 ( .A1(G651), .A2(G543), .ZN(n659) );
  NAND2_X1 U608 ( .A1(G88), .A2(n659), .ZN(n552) );
  XNOR2_X1 U609 ( .A(n552), .B(KEYINPUT86), .ZN(n554) );
  XOR2_X1 U610 ( .A(KEYINPUT0), .B(G543), .Z(n647) );
  INV_X1 U611 ( .A(G651), .ZN(n555) );
  NOR2_X2 U612 ( .A1(n647), .A2(n555), .ZN(n658) );
  NAND2_X1 U613 ( .A1(n658), .A2(G75), .ZN(n553) );
  NAND2_X1 U614 ( .A1(n554), .A2(n553), .ZN(n560) );
  NOR2_X1 U615 ( .A1(G543), .A2(n555), .ZN(n556) );
  XOR2_X1 U616 ( .A(KEYINPUT1), .B(n556), .Z(n588) );
  BUF_X1 U617 ( .A(n588), .Z(n662) );
  NAND2_X1 U618 ( .A1(G62), .A2(n662), .ZN(n558) );
  NOR2_X2 U619 ( .A1(G651), .A2(n647), .ZN(n663) );
  NAND2_X1 U620 ( .A1(G50), .A2(n663), .ZN(n557) );
  NAND2_X1 U621 ( .A1(n558), .A2(n557), .ZN(n559) );
  NOR2_X1 U622 ( .A1(n560), .A2(n559), .ZN(G166) );
  NAND2_X1 U623 ( .A1(G64), .A2(n662), .ZN(n561) );
  XNOR2_X1 U624 ( .A(n561), .B(KEYINPUT67), .ZN(n568) );
  NAND2_X1 U625 ( .A1(G77), .A2(n658), .ZN(n563) );
  NAND2_X1 U626 ( .A1(G90), .A2(n659), .ZN(n562) );
  NAND2_X1 U627 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U628 ( .A(n564), .B(KEYINPUT9), .ZN(n566) );
  NAND2_X1 U629 ( .A1(G52), .A2(n663), .ZN(n565) );
  NAND2_X1 U630 ( .A1(n566), .A2(n565), .ZN(n567) );
  NOR2_X1 U631 ( .A1(n568), .A2(n567), .ZN(G171) );
  NAND2_X1 U632 ( .A1(n662), .A2(G63), .ZN(n569) );
  XNOR2_X1 U633 ( .A(n569), .B(KEYINPUT72), .ZN(n571) );
  NAND2_X1 U634 ( .A1(G51), .A2(n663), .ZN(n570) );
  NAND2_X1 U635 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U636 ( .A(KEYINPUT6), .B(n572), .ZN(n578) );
  NAND2_X1 U637 ( .A1(n659), .A2(G89), .ZN(n573) );
  XNOR2_X1 U638 ( .A(n573), .B(KEYINPUT4), .ZN(n575) );
  NAND2_X1 U639 ( .A1(G76), .A2(n658), .ZN(n574) );
  NAND2_X1 U640 ( .A1(n575), .A2(n574), .ZN(n576) );
  XOR2_X1 U641 ( .A(n576), .B(KEYINPUT5), .Z(n577) );
  NOR2_X1 U642 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U643 ( .A(KEYINPUT73), .B(n579), .Z(n580) );
  XOR2_X1 U644 ( .A(KEYINPUT7), .B(n580), .Z(G168) );
  XOR2_X1 U645 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U646 ( .A1(G7), .A2(G661), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n581), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U648 ( .A(G223), .ZN(n852) );
  NAND2_X1 U649 ( .A1(n852), .A2(G567), .ZN(n582) );
  XOR2_X1 U650 ( .A(KEYINPUT11), .B(n582), .Z(G234) );
  NAND2_X1 U651 ( .A1(G43), .A2(n663), .ZN(n583) );
  NAND2_X1 U652 ( .A1(G68), .A2(n658), .ZN(n586) );
  NAND2_X1 U653 ( .A1(n659), .A2(G81), .ZN(n584) );
  XNOR2_X1 U654 ( .A(n584), .B(KEYINPUT12), .ZN(n585) );
  NAND2_X1 U655 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U656 ( .A(n587), .B(KEYINPUT13), .ZN(n590) );
  NAND2_X1 U657 ( .A1(G56), .A2(n588), .ZN(n589) );
  INV_X1 U658 ( .A(G860), .ZN(n611) );
  OR2_X1 U659 ( .A1(n982), .A2(n611), .ZN(G153) );
  INV_X1 U660 ( .A(G171), .ZN(G301) );
  NAND2_X1 U661 ( .A1(G868), .A2(G301), .ZN(n600) );
  NAND2_X1 U662 ( .A1(G79), .A2(n658), .ZN(n593) );
  NAND2_X1 U663 ( .A1(G92), .A2(n659), .ZN(n592) );
  NAND2_X1 U664 ( .A1(n593), .A2(n592), .ZN(n597) );
  NAND2_X1 U665 ( .A1(G66), .A2(n662), .ZN(n595) );
  NAND2_X1 U666 ( .A1(G54), .A2(n663), .ZN(n594) );
  NAND2_X1 U667 ( .A1(n595), .A2(n594), .ZN(n596) );
  NOR2_X1 U668 ( .A1(n597), .A2(n596), .ZN(n598) );
  XOR2_X1 U669 ( .A(KEYINPUT15), .B(n598), .Z(n994) );
  OR2_X1 U670 ( .A1(n994), .A2(G868), .ZN(n599) );
  NAND2_X1 U671 ( .A1(n600), .A2(n599), .ZN(G284) );
  NAND2_X1 U672 ( .A1(G91), .A2(n659), .ZN(n601) );
  XNOR2_X1 U673 ( .A(n601), .B(KEYINPUT68), .ZN(n608) );
  NAND2_X1 U674 ( .A1(G65), .A2(n662), .ZN(n603) );
  NAND2_X1 U675 ( .A1(G53), .A2(n663), .ZN(n602) );
  NAND2_X1 U676 ( .A1(n603), .A2(n602), .ZN(n606) );
  NAND2_X1 U677 ( .A1(G78), .A2(n658), .ZN(n604) );
  XNOR2_X1 U678 ( .A(KEYINPUT69), .B(n604), .ZN(n605) );
  NOR2_X1 U679 ( .A1(n606), .A2(n605), .ZN(n607) );
  NAND2_X1 U680 ( .A1(n608), .A2(n607), .ZN(G299) );
  INV_X1 U681 ( .A(G868), .ZN(n677) );
  NOR2_X1 U682 ( .A1(G286), .A2(n677), .ZN(n610) );
  NOR2_X1 U683 ( .A1(G868), .A2(G299), .ZN(n609) );
  NOR2_X1 U684 ( .A1(n610), .A2(n609), .ZN(G297) );
  NAND2_X1 U685 ( .A1(G559), .A2(n611), .ZN(n612) );
  XNOR2_X1 U686 ( .A(KEYINPUT74), .B(n612), .ZN(n613) );
  NAND2_X1 U687 ( .A1(n613), .A2(n994), .ZN(n615) );
  XOR2_X1 U688 ( .A(KEYINPUT75), .B(KEYINPUT16), .Z(n614) );
  XNOR2_X1 U689 ( .A(n615), .B(n614), .ZN(G148) );
  NOR2_X1 U690 ( .A1(G868), .A2(n982), .ZN(n618) );
  NAND2_X1 U691 ( .A1(G868), .A2(n994), .ZN(n616) );
  NOR2_X1 U692 ( .A1(G559), .A2(n616), .ZN(n617) );
  NOR2_X1 U693 ( .A1(n618), .A2(n617), .ZN(G282) );
  NAND2_X1 U694 ( .A1(G123), .A2(n522), .ZN(n620) );
  XNOR2_X1 U695 ( .A(n620), .B(KEYINPUT76), .ZN(n621) );
  XNOR2_X1 U696 ( .A(n621), .B(KEYINPUT18), .ZN(n623) );
  NAND2_X1 U697 ( .A1(G135), .A2(n902), .ZN(n622) );
  NAND2_X1 U698 ( .A1(n623), .A2(n622), .ZN(n624) );
  XOR2_X1 U699 ( .A(KEYINPUT77), .B(n624), .Z(n631) );
  NAND2_X1 U700 ( .A1(n900), .A2(G99), .ZN(n625) );
  XNOR2_X1 U701 ( .A(KEYINPUT79), .B(n625), .ZN(n628) );
  NAND2_X1 U702 ( .A1(n897), .A2(G111), .ZN(n626) );
  XOR2_X1 U703 ( .A(KEYINPUT78), .B(n626), .Z(n627) );
  NOR2_X1 U704 ( .A1(n628), .A2(n627), .ZN(n629) );
  XOR2_X1 U705 ( .A(KEYINPUT80), .B(n629), .Z(n630) );
  NOR2_X1 U706 ( .A1(n631), .A2(n630), .ZN(n1016) );
  XNOR2_X1 U707 ( .A(n1016), .B(G2096), .ZN(n633) );
  INV_X1 U708 ( .A(G2100), .ZN(n632) );
  NAND2_X1 U709 ( .A1(n633), .A2(n632), .ZN(G156) );
  NAND2_X1 U710 ( .A1(G60), .A2(n662), .ZN(n635) );
  NAND2_X1 U711 ( .A1(G47), .A2(n663), .ZN(n634) );
  NAND2_X1 U712 ( .A1(n635), .A2(n634), .ZN(n640) );
  NAND2_X1 U713 ( .A1(G72), .A2(n658), .ZN(n637) );
  NAND2_X1 U714 ( .A1(G85), .A2(n659), .ZN(n636) );
  NAND2_X1 U715 ( .A1(n637), .A2(n636), .ZN(n638) );
  XOR2_X1 U716 ( .A(KEYINPUT65), .B(n638), .Z(n639) );
  NOR2_X1 U717 ( .A1(n640), .A2(n639), .ZN(n641) );
  XOR2_X1 U718 ( .A(KEYINPUT66), .B(n641), .Z(G290) );
  NAND2_X1 U719 ( .A1(G49), .A2(n663), .ZN(n642) );
  XNOR2_X1 U720 ( .A(n642), .B(KEYINPUT84), .ZN(n645) );
  NAND2_X1 U721 ( .A1(G74), .A2(G651), .ZN(n643) );
  XOR2_X1 U722 ( .A(KEYINPUT85), .B(n643), .Z(n644) );
  NAND2_X1 U723 ( .A1(n645), .A2(n644), .ZN(n646) );
  NOR2_X1 U724 ( .A1(n662), .A2(n646), .ZN(n649) );
  NAND2_X1 U725 ( .A1(n647), .A2(G87), .ZN(n648) );
  NAND2_X1 U726 ( .A1(n649), .A2(n648), .ZN(G288) );
  NAND2_X1 U727 ( .A1(G61), .A2(n662), .ZN(n651) );
  NAND2_X1 U728 ( .A1(G48), .A2(n663), .ZN(n650) );
  NAND2_X1 U729 ( .A1(n651), .A2(n650), .ZN(n654) );
  NAND2_X1 U730 ( .A1(G73), .A2(n658), .ZN(n652) );
  XOR2_X1 U731 ( .A(KEYINPUT2), .B(n652), .Z(n653) );
  NOR2_X1 U732 ( .A1(n654), .A2(n653), .ZN(n656) );
  NAND2_X1 U733 ( .A1(n659), .A2(G86), .ZN(n655) );
  NAND2_X1 U734 ( .A1(n656), .A2(n655), .ZN(G305) );
  NAND2_X1 U735 ( .A1(G559), .A2(n994), .ZN(n657) );
  XNOR2_X1 U736 ( .A(n657), .B(n982), .ZN(n859) );
  NAND2_X1 U737 ( .A1(G80), .A2(n658), .ZN(n661) );
  NAND2_X1 U738 ( .A1(G93), .A2(n659), .ZN(n660) );
  NAND2_X1 U739 ( .A1(n661), .A2(n660), .ZN(n668) );
  NAND2_X1 U740 ( .A1(G67), .A2(n662), .ZN(n665) );
  NAND2_X1 U741 ( .A1(G55), .A2(n663), .ZN(n664) );
  NAND2_X1 U742 ( .A1(n665), .A2(n664), .ZN(n666) );
  XNOR2_X1 U743 ( .A(KEYINPUT82), .B(n666), .ZN(n667) );
  NOR2_X1 U744 ( .A1(n668), .A2(n667), .ZN(n669) );
  XNOR2_X1 U745 ( .A(n669), .B(KEYINPUT83), .ZN(n861) );
  XNOR2_X1 U746 ( .A(G290), .B(n861), .ZN(n675) );
  XOR2_X1 U747 ( .A(KEYINPUT19), .B(KEYINPUT87), .Z(n671) );
  INV_X1 U748 ( .A(G299), .ZN(n999) );
  XNOR2_X1 U749 ( .A(G166), .B(n999), .ZN(n670) );
  XNOR2_X1 U750 ( .A(n671), .B(n670), .ZN(n672) );
  XOR2_X1 U751 ( .A(n672), .B(G305), .Z(n673) );
  XNOR2_X1 U752 ( .A(G288), .B(n673), .ZN(n674) );
  XNOR2_X1 U753 ( .A(n675), .B(n674), .ZN(n920) );
  XNOR2_X1 U754 ( .A(n859), .B(n920), .ZN(n676) );
  NAND2_X1 U755 ( .A1(n676), .A2(G868), .ZN(n679) );
  NAND2_X1 U756 ( .A1(n677), .A2(n861), .ZN(n678) );
  NAND2_X1 U757 ( .A1(n679), .A2(n678), .ZN(G295) );
  NAND2_X1 U758 ( .A1(G2078), .A2(G2084), .ZN(n680) );
  XOR2_X1 U759 ( .A(KEYINPUT20), .B(n680), .Z(n681) );
  NAND2_X1 U760 ( .A1(G2090), .A2(n681), .ZN(n682) );
  XNOR2_X1 U761 ( .A(KEYINPUT21), .B(n682), .ZN(n683) );
  NAND2_X1 U762 ( .A1(n683), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U763 ( .A(KEYINPUT88), .B(G44), .ZN(n684) );
  XNOR2_X1 U764 ( .A(n684), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U765 ( .A(KEYINPUT70), .B(G132), .Z(G219) );
  NOR2_X1 U766 ( .A1(G219), .A2(G220), .ZN(n685) );
  XOR2_X1 U767 ( .A(KEYINPUT22), .B(n685), .Z(n686) );
  NOR2_X1 U768 ( .A1(G218), .A2(n686), .ZN(n687) );
  NAND2_X1 U769 ( .A1(G96), .A2(n687), .ZN(n857) );
  NAND2_X1 U770 ( .A1(G2106), .A2(n857), .ZN(n691) );
  NAND2_X1 U771 ( .A1(G69), .A2(G120), .ZN(n688) );
  NOR2_X1 U772 ( .A1(G237), .A2(n688), .ZN(n689) );
  NAND2_X1 U773 ( .A1(G108), .A2(n689), .ZN(n858) );
  NAND2_X1 U774 ( .A1(G567), .A2(n858), .ZN(n690) );
  NAND2_X1 U775 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U776 ( .A(KEYINPUT89), .B(n692), .ZN(G319) );
  INV_X1 U777 ( .A(G319), .ZN(n694) );
  NAND2_X1 U778 ( .A1(G661), .A2(G483), .ZN(n693) );
  NOR2_X1 U779 ( .A1(n694), .A2(n693), .ZN(n856) );
  NAND2_X1 U780 ( .A1(n856), .A2(G36), .ZN(G176) );
  INV_X1 U781 ( .A(G166), .ZN(G303) );
  NAND2_X1 U782 ( .A1(G40), .A2(G160), .ZN(n695) );
  XNOR2_X1 U783 ( .A(n695), .B(KEYINPUT92), .ZN(n816) );
  INV_X1 U784 ( .A(n816), .ZN(n698) );
  XNOR2_X1 U785 ( .A(n697), .B(KEYINPUT64), .ZN(n815) );
  NAND2_X1 U786 ( .A1(n748), .A2(G1961), .ZN(n701) );
  INV_X1 U787 ( .A(n748), .ZN(n733) );
  XOR2_X1 U788 ( .A(G2078), .B(KEYINPUT98), .Z(n699) );
  XNOR2_X1 U789 ( .A(KEYINPUT25), .B(n699), .ZN(n939) );
  NAND2_X1 U790 ( .A1(n733), .A2(n939), .ZN(n700) );
  NAND2_X1 U791 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U792 ( .A(n702), .B(KEYINPUT99), .ZN(n745) );
  NOR2_X1 U793 ( .A1(G171), .A2(n745), .ZN(n711) );
  INV_X1 U794 ( .A(G1966), .ZN(n704) );
  NAND2_X1 U795 ( .A1(G8), .A2(n715), .ZN(n703) );
  XNOR2_X1 U796 ( .A(KEYINPUT97), .B(n703), .ZN(n750) );
  AND2_X1 U797 ( .A1(n704), .A2(n750), .ZN(n765) );
  NOR2_X1 U798 ( .A1(G2084), .A2(n748), .ZN(n768) );
  NOR2_X1 U799 ( .A1(n765), .A2(n768), .ZN(n706) );
  XNOR2_X1 U800 ( .A(n706), .B(n705), .ZN(n707) );
  NAND2_X1 U801 ( .A1(n707), .A2(G8), .ZN(n708) );
  XNOR2_X1 U802 ( .A(KEYINPUT30), .B(n708), .ZN(n709) );
  NOR2_X1 U803 ( .A1(n709), .A2(G168), .ZN(n710) );
  NOR2_X1 U804 ( .A1(n711), .A2(n710), .ZN(n713) );
  NAND2_X1 U805 ( .A1(n715), .A2(G1341), .ZN(n721) );
  INV_X1 U806 ( .A(n982), .ZN(n714) );
  AND2_X1 U807 ( .A1(n721), .A2(n714), .ZN(n718) );
  INV_X1 U808 ( .A(G1996), .ZN(n934) );
  INV_X1 U809 ( .A(KEYINPUT26), .ZN(n716) );
  XNOR2_X1 U810 ( .A(n717), .B(n716), .ZN(n722) );
  AND2_X1 U811 ( .A1(n718), .A2(n722), .ZN(n719) );
  NOR2_X1 U812 ( .A1(n719), .A2(n994), .ZN(n720) );
  XNOR2_X1 U813 ( .A(n720), .B(KEYINPUT101), .ZN(n730) );
  NAND2_X1 U814 ( .A1(n722), .A2(n721), .ZN(n723) );
  NOR2_X1 U815 ( .A1(n982), .A2(n723), .ZN(n724) );
  NAND2_X1 U816 ( .A1(n724), .A2(n994), .ZN(n728) );
  NOR2_X1 U817 ( .A1(n733), .A2(G1348), .ZN(n726) );
  NOR2_X1 U818 ( .A1(G2067), .A2(n748), .ZN(n725) );
  NOR2_X1 U819 ( .A1(n726), .A2(n725), .ZN(n727) );
  NAND2_X1 U820 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U821 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U822 ( .A(n731), .B(KEYINPUT102), .ZN(n737) );
  NAND2_X1 U823 ( .A1(n733), .A2(G2072), .ZN(n732) );
  XNOR2_X1 U824 ( .A(n732), .B(KEYINPUT27), .ZN(n735) );
  INV_X1 U825 ( .A(G1956), .ZN(n1000) );
  NOR2_X1 U826 ( .A1(n1000), .A2(n733), .ZN(n734) );
  NOR2_X1 U827 ( .A1(n735), .A2(n734), .ZN(n738) );
  NAND2_X1 U828 ( .A1(n738), .A2(n999), .ZN(n736) );
  NAND2_X1 U829 ( .A1(n737), .A2(n736), .ZN(n742) );
  NOR2_X1 U830 ( .A1(n738), .A2(n999), .ZN(n740) );
  XOR2_X1 U831 ( .A(KEYINPUT28), .B(KEYINPUT100), .Z(n739) );
  XNOR2_X1 U832 ( .A(n740), .B(n739), .ZN(n741) );
  NAND2_X1 U833 ( .A1(n742), .A2(n741), .ZN(n744) );
  XNOR2_X1 U834 ( .A(n744), .B(n743), .ZN(n747) );
  NAND2_X1 U835 ( .A1(G171), .A2(n745), .ZN(n746) );
  NAND2_X1 U836 ( .A1(n747), .A2(n746), .ZN(n766) );
  INV_X1 U837 ( .A(G8), .ZN(n756) );
  NOR2_X1 U838 ( .A1(G2090), .A2(n748), .ZN(n749) );
  XNOR2_X1 U839 ( .A(n749), .B(KEYINPUT104), .ZN(n753) );
  BUF_X1 U840 ( .A(n750), .Z(n795) );
  INV_X1 U841 ( .A(n795), .ZN(n751) );
  NOR2_X1 U842 ( .A1(n751), .A2(G1971), .ZN(n752) );
  NOR2_X1 U843 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U844 ( .A1(n754), .A2(G303), .ZN(n755) );
  OR2_X1 U845 ( .A1(n756), .A2(n755), .ZN(n758) );
  AND2_X1 U846 ( .A1(n766), .A2(n758), .ZN(n757) );
  NAND2_X1 U847 ( .A1(n767), .A2(n757), .ZN(n762) );
  INV_X1 U848 ( .A(n758), .ZN(n760) );
  AND2_X1 U849 ( .A1(G286), .A2(G8), .ZN(n759) );
  OR2_X1 U850 ( .A1(n760), .A2(n759), .ZN(n761) );
  NAND2_X1 U851 ( .A1(n762), .A2(n761), .ZN(n764) );
  XNOR2_X1 U852 ( .A(n764), .B(n763), .ZN(n773) );
  NAND2_X1 U853 ( .A1(n766), .A2(n767), .ZN(n770) );
  NAND2_X1 U854 ( .A1(G8), .A2(n768), .ZN(n769) );
  NAND2_X1 U855 ( .A1(n770), .A2(n769), .ZN(n771) );
  NOR2_X1 U856 ( .A1(n765), .A2(n771), .ZN(n772) );
  NOR2_X2 U857 ( .A1(n773), .A2(n772), .ZN(n785) );
  INV_X1 U858 ( .A(n785), .ZN(n776) );
  NOR2_X1 U859 ( .A1(G1971), .A2(G303), .ZN(n774) );
  NOR2_X1 U860 ( .A1(G1976), .A2(G288), .ZN(n998) );
  NOR2_X1 U861 ( .A1(n774), .A2(n998), .ZN(n775) );
  NAND2_X1 U862 ( .A1(n776), .A2(n775), .ZN(n777) );
  NAND2_X1 U863 ( .A1(G1976), .A2(G288), .ZN(n992) );
  NAND2_X1 U864 ( .A1(n777), .A2(n992), .ZN(n778) );
  NOR2_X1 U865 ( .A1(KEYINPUT33), .A2(n778), .ZN(n779) );
  NAND2_X1 U866 ( .A1(n779), .A2(n795), .ZN(n782) );
  NAND2_X1 U867 ( .A1(n998), .A2(n795), .ZN(n780) );
  NAND2_X1 U868 ( .A1(n780), .A2(KEYINPUT33), .ZN(n781) );
  NAND2_X1 U869 ( .A1(n782), .A2(n781), .ZN(n783) );
  XNOR2_X1 U870 ( .A(n783), .B(KEYINPUT105), .ZN(n784) );
  XNOR2_X1 U871 ( .A(G1981), .B(G305), .ZN(n986) );
  NOR2_X1 U872 ( .A1(n784), .A2(n986), .ZN(n792) );
  NAND2_X1 U873 ( .A1(G8), .A2(G166), .ZN(n786) );
  NOR2_X1 U874 ( .A1(G2090), .A2(n786), .ZN(n787) );
  XNOR2_X1 U875 ( .A(n787), .B(KEYINPUT106), .ZN(n788) );
  NOR2_X1 U876 ( .A1(n785), .A2(n788), .ZN(n789) );
  XOR2_X1 U877 ( .A(KEYINPUT107), .B(n789), .Z(n790) );
  NOR2_X1 U878 ( .A1(n795), .A2(n790), .ZN(n791) );
  XNOR2_X1 U879 ( .A(n793), .B(KEYINPUT108), .ZN(n838) );
  NOR2_X1 U880 ( .A1(G1981), .A2(G305), .ZN(n794) );
  XNOR2_X1 U881 ( .A(n794), .B(KEYINPUT24), .ZN(n796) );
  NAND2_X1 U882 ( .A1(n796), .A2(n795), .ZN(n836) );
  NAND2_X1 U883 ( .A1(G105), .A2(n900), .ZN(n797) );
  XNOR2_X1 U884 ( .A(n797), .B(KEYINPUT38), .ZN(n804) );
  NAND2_X1 U885 ( .A1(G129), .A2(n522), .ZN(n799) );
  NAND2_X1 U886 ( .A1(G141), .A2(n902), .ZN(n798) );
  NAND2_X1 U887 ( .A1(n799), .A2(n798), .ZN(n802) );
  NAND2_X1 U888 ( .A1(n897), .A2(G117), .ZN(n800) );
  XOR2_X1 U889 ( .A(KEYINPUT96), .B(n800), .Z(n801) );
  NOR2_X1 U890 ( .A1(n802), .A2(n801), .ZN(n803) );
  NAND2_X1 U891 ( .A1(n804), .A2(n803), .ZN(n914) );
  NOR2_X1 U892 ( .A1(G1996), .A2(n914), .ZN(n1024) );
  NAND2_X1 U893 ( .A1(n900), .A2(G95), .ZN(n805) );
  XNOR2_X1 U894 ( .A(n805), .B(KEYINPUT94), .ZN(n807) );
  NAND2_X1 U895 ( .A1(G131), .A2(n902), .ZN(n806) );
  NAND2_X1 U896 ( .A1(n807), .A2(n806), .ZN(n808) );
  XNOR2_X1 U897 ( .A(KEYINPUT95), .B(n808), .ZN(n812) );
  NAND2_X1 U898 ( .A1(G119), .A2(n522), .ZN(n810) );
  NAND2_X1 U899 ( .A1(G107), .A2(n897), .ZN(n809) );
  AND2_X1 U900 ( .A1(n810), .A2(n809), .ZN(n811) );
  NAND2_X1 U901 ( .A1(n812), .A2(n811), .ZN(n910) );
  AND2_X1 U902 ( .A1(n910), .A2(G1991), .ZN(n814) );
  AND2_X1 U903 ( .A1(n914), .A2(G1996), .ZN(n813) );
  NOR2_X1 U904 ( .A1(n814), .A2(n813), .ZN(n1022) );
  NOR2_X1 U905 ( .A1(n816), .A2(n815), .ZN(n844) );
  INV_X1 U906 ( .A(n844), .ZN(n817) );
  NOR2_X1 U907 ( .A1(n1022), .A2(n817), .ZN(n840) );
  NOR2_X1 U908 ( .A1(G1986), .A2(G290), .ZN(n818) );
  NOR2_X1 U909 ( .A1(G1991), .A2(n910), .ZN(n1015) );
  NOR2_X1 U910 ( .A1(n818), .A2(n1015), .ZN(n819) );
  NOR2_X1 U911 ( .A1(n840), .A2(n819), .ZN(n820) );
  NOR2_X1 U912 ( .A1(n1024), .A2(n820), .ZN(n821) );
  XNOR2_X1 U913 ( .A(n821), .B(KEYINPUT39), .ZN(n832) );
  XNOR2_X1 U914 ( .A(G2067), .B(KEYINPUT37), .ZN(n833) );
  NAND2_X1 U915 ( .A1(G104), .A2(n900), .ZN(n823) );
  NAND2_X1 U916 ( .A1(G140), .A2(n902), .ZN(n822) );
  NAND2_X1 U917 ( .A1(n823), .A2(n822), .ZN(n824) );
  XNOR2_X1 U918 ( .A(KEYINPUT34), .B(n824), .ZN(n829) );
  NAND2_X1 U919 ( .A1(G128), .A2(n522), .ZN(n826) );
  NAND2_X1 U920 ( .A1(G116), .A2(n897), .ZN(n825) );
  NAND2_X1 U921 ( .A1(n826), .A2(n825), .ZN(n827) );
  XOR2_X1 U922 ( .A(n827), .B(KEYINPUT35), .Z(n828) );
  NOR2_X1 U923 ( .A1(n829), .A2(n828), .ZN(n830) );
  XOR2_X1 U924 ( .A(KEYINPUT36), .B(n830), .Z(n831) );
  XNOR2_X1 U925 ( .A(KEYINPUT93), .B(n831), .ZN(n917) );
  NOR2_X1 U926 ( .A1(n833), .A2(n917), .ZN(n1017) );
  NAND2_X1 U927 ( .A1(n844), .A2(n1017), .ZN(n841) );
  NAND2_X1 U928 ( .A1(n832), .A2(n841), .ZN(n834) );
  NAND2_X1 U929 ( .A1(n833), .A2(n917), .ZN(n1021) );
  NAND2_X1 U930 ( .A1(n834), .A2(n1021), .ZN(n835) );
  NAND2_X1 U931 ( .A1(n835), .A2(n844), .ZN(n839) );
  AND2_X1 U932 ( .A1(n836), .A2(n839), .ZN(n837) );
  NAND2_X1 U933 ( .A1(n838), .A2(n837), .ZN(n850) );
  INV_X1 U934 ( .A(n839), .ZN(n848) );
  INV_X1 U935 ( .A(n840), .ZN(n842) );
  NAND2_X1 U936 ( .A1(n842), .A2(n841), .ZN(n846) );
  XOR2_X1 U937 ( .A(KEYINPUT91), .B(G1986), .Z(n843) );
  XNOR2_X1 U938 ( .A(G290), .B(n843), .ZN(n989) );
  AND2_X1 U939 ( .A1(n989), .A2(n844), .ZN(n845) );
  NOR2_X1 U940 ( .A1(n846), .A2(n845), .ZN(n847) );
  OR2_X1 U941 ( .A1(n848), .A2(n847), .ZN(n849) );
  AND2_X1 U942 ( .A1(n850), .A2(n849), .ZN(n851) );
  XNOR2_X1 U943 ( .A(n851), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U944 ( .A1(G2106), .A2(n852), .ZN(G217) );
  NAND2_X1 U945 ( .A1(G15), .A2(G2), .ZN(n853) );
  XNOR2_X1 U946 ( .A(KEYINPUT109), .B(n853), .ZN(n854) );
  NAND2_X1 U947 ( .A1(n854), .A2(G661), .ZN(G259) );
  NAND2_X1 U948 ( .A1(G3), .A2(G1), .ZN(n855) );
  NAND2_X1 U949 ( .A1(n856), .A2(n855), .ZN(G188) );
  INV_X1 U951 ( .A(G120), .ZN(G236) );
  INV_X1 U952 ( .A(G96), .ZN(G221) );
  INV_X1 U953 ( .A(G69), .ZN(G235) );
  NOR2_X1 U954 ( .A1(n858), .A2(n857), .ZN(G325) );
  INV_X1 U955 ( .A(G325), .ZN(G261) );
  XOR2_X1 U956 ( .A(KEYINPUT81), .B(n859), .Z(n860) );
  NOR2_X1 U957 ( .A1(G860), .A2(n860), .ZN(n862) );
  XOR2_X1 U958 ( .A(n862), .B(n861), .Z(G145) );
  XOR2_X1 U959 ( .A(G2100), .B(G2096), .Z(n864) );
  XNOR2_X1 U960 ( .A(KEYINPUT42), .B(G2678), .ZN(n863) );
  XNOR2_X1 U961 ( .A(n864), .B(n863), .ZN(n868) );
  XOR2_X1 U962 ( .A(KEYINPUT43), .B(G2090), .Z(n866) );
  XNOR2_X1 U963 ( .A(G2072), .B(G2067), .ZN(n865) );
  XNOR2_X1 U964 ( .A(n866), .B(n865), .ZN(n867) );
  XOR2_X1 U965 ( .A(n868), .B(n867), .Z(n870) );
  XNOR2_X1 U966 ( .A(G2078), .B(G2084), .ZN(n869) );
  XNOR2_X1 U967 ( .A(n870), .B(n869), .ZN(G227) );
  XOR2_X1 U968 ( .A(G1986), .B(G1956), .Z(n872) );
  XNOR2_X1 U969 ( .A(G1971), .B(G1966), .ZN(n871) );
  XNOR2_X1 U970 ( .A(n872), .B(n871), .ZN(n873) );
  XOR2_X1 U971 ( .A(n873), .B(G2474), .Z(n875) );
  XNOR2_X1 U972 ( .A(G1981), .B(G1961), .ZN(n874) );
  XNOR2_X1 U973 ( .A(n875), .B(n874), .ZN(n879) );
  XOR2_X1 U974 ( .A(KEYINPUT41), .B(G1991), .Z(n877) );
  XNOR2_X1 U975 ( .A(G1976), .B(G1996), .ZN(n876) );
  XNOR2_X1 U976 ( .A(n877), .B(n876), .ZN(n878) );
  XNOR2_X1 U977 ( .A(n879), .B(n878), .ZN(G229) );
  NAND2_X1 U978 ( .A1(G124), .A2(n522), .ZN(n880) );
  XNOR2_X1 U979 ( .A(n880), .B(KEYINPUT44), .ZN(n882) );
  NAND2_X1 U980 ( .A1(n900), .A2(G100), .ZN(n881) );
  NAND2_X1 U981 ( .A1(n882), .A2(n881), .ZN(n886) );
  NAND2_X1 U982 ( .A1(G136), .A2(n902), .ZN(n884) );
  NAND2_X1 U983 ( .A1(G112), .A2(n897), .ZN(n883) );
  NAND2_X1 U984 ( .A1(n884), .A2(n883), .ZN(n885) );
  NOR2_X1 U985 ( .A1(n886), .A2(n885), .ZN(G162) );
  XOR2_X1 U986 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n896) );
  NAND2_X1 U987 ( .A1(G103), .A2(n900), .ZN(n888) );
  NAND2_X1 U988 ( .A1(G139), .A2(n902), .ZN(n887) );
  NAND2_X1 U989 ( .A1(n888), .A2(n887), .ZN(n894) );
  NAND2_X1 U990 ( .A1(G127), .A2(n522), .ZN(n890) );
  NAND2_X1 U991 ( .A1(G115), .A2(n897), .ZN(n889) );
  NAND2_X1 U992 ( .A1(n890), .A2(n889), .ZN(n891) );
  XNOR2_X1 U993 ( .A(KEYINPUT111), .B(n891), .ZN(n892) );
  XNOR2_X1 U994 ( .A(KEYINPUT47), .B(n892), .ZN(n893) );
  NOR2_X1 U995 ( .A1(n894), .A2(n893), .ZN(n1030) );
  XNOR2_X1 U996 ( .A(G164), .B(n1030), .ZN(n895) );
  XNOR2_X1 U997 ( .A(n896), .B(n895), .ZN(n909) );
  NAND2_X1 U998 ( .A1(G130), .A2(n522), .ZN(n899) );
  NAND2_X1 U999 ( .A1(G118), .A2(n897), .ZN(n898) );
  NAND2_X1 U1000 ( .A1(n899), .A2(n898), .ZN(n907) );
  NAND2_X1 U1001 ( .A1(n900), .A2(G106), .ZN(n901) );
  XNOR2_X1 U1002 ( .A(n901), .B(KEYINPUT110), .ZN(n904) );
  NAND2_X1 U1003 ( .A1(G142), .A2(n902), .ZN(n903) );
  NAND2_X1 U1004 ( .A1(n904), .A2(n903), .ZN(n905) );
  XOR2_X1 U1005 ( .A(KEYINPUT45), .B(n905), .Z(n906) );
  NOR2_X1 U1006 ( .A1(n907), .A2(n906), .ZN(n908) );
  XOR2_X1 U1007 ( .A(n909), .B(n908), .Z(n912) );
  XOR2_X1 U1008 ( .A(G160), .B(n910), .Z(n911) );
  XNOR2_X1 U1009 ( .A(n912), .B(n911), .ZN(n913) );
  XOR2_X1 U1010 ( .A(n913), .B(G162), .Z(n916) );
  XOR2_X1 U1011 ( .A(n914), .B(n1016), .Z(n915) );
  XNOR2_X1 U1012 ( .A(n916), .B(n915), .ZN(n918) );
  XOR2_X1 U1013 ( .A(n918), .B(n917), .Z(n919) );
  NOR2_X1 U1014 ( .A1(G37), .A2(n919), .ZN(G395) );
  XOR2_X1 U1015 ( .A(KEYINPUT112), .B(n920), .Z(n922) );
  XNOR2_X1 U1016 ( .A(n994), .B(G286), .ZN(n921) );
  XNOR2_X1 U1017 ( .A(n922), .B(n921), .ZN(n924) );
  XNOR2_X1 U1018 ( .A(n982), .B(G171), .ZN(n923) );
  XNOR2_X1 U1019 ( .A(n924), .B(n923), .ZN(n925) );
  NOR2_X1 U1020 ( .A1(G37), .A2(n925), .ZN(G397) );
  NOR2_X1 U1021 ( .A1(G227), .A2(G229), .ZN(n927) );
  XNOR2_X1 U1022 ( .A(KEYINPUT49), .B(KEYINPUT113), .ZN(n926) );
  XNOR2_X1 U1023 ( .A(n927), .B(n926), .ZN(n930) );
  NOR2_X1 U1024 ( .A1(G395), .A2(G397), .ZN(n928) );
  XNOR2_X1 U1025 ( .A(n928), .B(KEYINPUT114), .ZN(n929) );
  NAND2_X1 U1026 ( .A1(n930), .A2(n929), .ZN(n931) );
  NOR2_X1 U1027 ( .A1(G401), .A2(n931), .ZN(n932) );
  NAND2_X1 U1028 ( .A1(G319), .A2(n932), .ZN(G225) );
  INV_X1 U1029 ( .A(G225), .ZN(G308) );
  INV_X1 U1030 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1031 ( .A(G29), .B(KEYINPUT119), .ZN(n955) );
  XOR2_X1 U1032 ( .A(KEYINPUT55), .B(KEYINPUT118), .Z(n953) );
  XNOR2_X1 U1033 ( .A(G2090), .B(G35), .ZN(n948) );
  XOR2_X1 U1034 ( .A(G25), .B(G1991), .Z(n933) );
  NAND2_X1 U1035 ( .A1(n933), .A2(G28), .ZN(n945) );
  XNOR2_X1 U1036 ( .A(G32), .B(n934), .ZN(n938) );
  XNOR2_X1 U1037 ( .A(G2072), .B(G33), .ZN(n936) );
  XNOR2_X1 U1038 ( .A(G26), .B(G2067), .ZN(n935) );
  NOR2_X1 U1039 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1040 ( .A1(n938), .A2(n937), .ZN(n942) );
  XNOR2_X1 U1041 ( .A(G27), .B(n939), .ZN(n940) );
  XNOR2_X1 U1042 ( .A(KEYINPUT116), .B(n940), .ZN(n941) );
  NOR2_X1 U1043 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1044 ( .A(n943), .B(KEYINPUT117), .ZN(n944) );
  NOR2_X1 U1045 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1046 ( .A(KEYINPUT53), .B(n946), .ZN(n947) );
  NOR2_X1 U1047 ( .A1(n948), .A2(n947), .ZN(n951) );
  XOR2_X1 U1048 ( .A(G2084), .B(G34), .Z(n949) );
  XNOR2_X1 U1049 ( .A(KEYINPUT54), .B(n949), .ZN(n950) );
  NAND2_X1 U1050 ( .A1(n951), .A2(n950), .ZN(n952) );
  XNOR2_X1 U1051 ( .A(n953), .B(n952), .ZN(n954) );
  NAND2_X1 U1052 ( .A1(n955), .A2(n954), .ZN(n1013) );
  XNOR2_X1 U1053 ( .A(G1976), .B(G23), .ZN(n957) );
  XNOR2_X1 U1054 ( .A(G1971), .B(G22), .ZN(n956) );
  NOR2_X1 U1055 ( .A1(n957), .A2(n956), .ZN(n959) );
  XOR2_X1 U1056 ( .A(G1986), .B(G24), .Z(n958) );
  NAND2_X1 U1057 ( .A1(n959), .A2(n958), .ZN(n961) );
  XOR2_X1 U1058 ( .A(KEYINPUT58), .B(KEYINPUT126), .Z(n960) );
  XNOR2_X1 U1059 ( .A(n961), .B(n960), .ZN(n965) );
  XNOR2_X1 U1060 ( .A(G1966), .B(G21), .ZN(n963) );
  XNOR2_X1 U1061 ( .A(G5), .B(G1961), .ZN(n962) );
  NOR2_X1 U1062 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1063 ( .A1(n965), .A2(n964), .ZN(n979) );
  XNOR2_X1 U1064 ( .A(KEYINPUT123), .B(G1981), .ZN(n966) );
  XNOR2_X1 U1065 ( .A(n966), .B(G6), .ZN(n975) );
  XOR2_X1 U1066 ( .A(G1341), .B(G19), .Z(n970) );
  XNOR2_X1 U1067 ( .A(KEYINPUT59), .B(G4), .ZN(n967) );
  XNOR2_X1 U1068 ( .A(n967), .B(KEYINPUT124), .ZN(n968) );
  XNOR2_X1 U1069 ( .A(G1348), .B(n968), .ZN(n969) );
  NAND2_X1 U1070 ( .A1(n970), .A2(n969), .ZN(n973) );
  XOR2_X1 U1071 ( .A(KEYINPUT122), .B(n1000), .Z(n971) );
  XNOR2_X1 U1072 ( .A(G20), .B(n971), .ZN(n972) );
  NOR2_X1 U1073 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1074 ( .A1(n975), .A2(n974), .ZN(n976) );
  XOR2_X1 U1075 ( .A(KEYINPUT60), .B(n976), .Z(n977) );
  XNOR2_X1 U1076 ( .A(KEYINPUT125), .B(n977), .ZN(n978) );
  NOR2_X1 U1077 ( .A1(n979), .A2(n978), .ZN(n980) );
  XOR2_X1 U1078 ( .A(KEYINPUT61), .B(n980), .Z(n981) );
  NOR2_X1 U1079 ( .A1(G16), .A2(n981), .ZN(n1010) );
  XOR2_X1 U1080 ( .A(G16), .B(KEYINPUT56), .Z(n1008) );
  XNOR2_X1 U1081 ( .A(G301), .B(G1961), .ZN(n984) );
  XNOR2_X1 U1082 ( .A(n982), .B(G1341), .ZN(n983) );
  NOR2_X1 U1083 ( .A1(n984), .A2(n983), .ZN(n991) );
  XOR2_X1 U1084 ( .A(G1966), .B(G168), .Z(n985) );
  NOR2_X1 U1085 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1086 ( .A(n987), .B(KEYINPUT57), .ZN(n988) );
  NOR2_X1 U1087 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1088 ( .A1(n991), .A2(n990), .ZN(n1006) );
  XNOR2_X1 U1089 ( .A(G166), .B(G1971), .ZN(n993) );
  NAND2_X1 U1090 ( .A1(n993), .A2(n992), .ZN(n997) );
  XOR2_X1 U1091 ( .A(n994), .B(G1348), .Z(n995) );
  XNOR2_X1 U1092 ( .A(KEYINPUT120), .B(n995), .ZN(n996) );
  NOR2_X1 U1093 ( .A1(n997), .A2(n996), .ZN(n1004) );
  XOR2_X1 U1094 ( .A(n998), .B(KEYINPUT121), .Z(n1002) );
  XNOR2_X1 U1095 ( .A(n1000), .B(n999), .ZN(n1001) );
  NOR2_X1 U1096 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1097 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NOR2_X1 U1098 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NOR2_X1 U1099 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NOR2_X1 U1100 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XOR2_X1 U1101 ( .A(KEYINPUT127), .B(n1011), .Z(n1012) );
  NAND2_X1 U1102 ( .A1(n1013), .A2(n1012), .ZN(n1041) );
  XOR2_X1 U1103 ( .A(G2084), .B(G160), .Z(n1014) );
  NOR2_X1 U1104 ( .A1(n1015), .A2(n1014), .ZN(n1019) );
  NOR2_X1 U1105 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1106 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1107 ( .A(KEYINPUT115), .B(n1020), .ZN(n1029) );
  NAND2_X1 U1108 ( .A1(n1022), .A2(n1021), .ZN(n1027) );
  XOR2_X1 U1109 ( .A(G2090), .B(G162), .Z(n1023) );
  NOR2_X1 U1110 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XNOR2_X1 U1111 ( .A(n1025), .B(KEYINPUT51), .ZN(n1026) );
  NOR2_X1 U1112 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NAND2_X1 U1113 ( .A1(n1029), .A2(n1028), .ZN(n1035) );
  XOR2_X1 U1114 ( .A(G2072), .B(n1030), .Z(n1032) );
  XOR2_X1 U1115 ( .A(G164), .B(G2078), .Z(n1031) );
  NOR2_X1 U1116 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  XOR2_X1 U1117 ( .A(KEYINPUT50), .B(n1033), .Z(n1034) );
  NOR2_X1 U1118 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  XOR2_X1 U1119 ( .A(KEYINPUT52), .B(n1036), .Z(n1037) );
  NOR2_X1 U1120 ( .A1(KEYINPUT55), .A2(n1037), .ZN(n1039) );
  INV_X1 U1121 ( .A(G29), .ZN(n1038) );
  NOR2_X1 U1122 ( .A1(n1039), .A2(n1038), .ZN(n1040) );
  NOR2_X1 U1123 ( .A1(n1041), .A2(n1040), .ZN(n1042) );
  NAND2_X1 U1124 ( .A1(n1042), .A2(G11), .ZN(n1043) );
  XOR2_X1 U1125 ( .A(KEYINPUT62), .B(n1043), .Z(G311) );
  INV_X1 U1126 ( .A(G311), .ZN(G150) );
endmodule

