//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 1 1 0 0 1 0 0 1 0 0 0 0 0 0 0 0 0 1 1 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 1 1 0 1 0 1 1 1 0 0 1 0 1 0 1 0 1 0 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:58 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n669, new_n670, new_n671, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n682, new_n683, new_n684,
    new_n686, new_n687, new_n688, new_n689, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n743, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974;
  INV_X1    g000(.A(G146), .ZN(new_n187));
  NOR2_X1   g001(.A1(new_n187), .A2(G143), .ZN(new_n188));
  XNOR2_X1  g002(.A(KEYINPUT65), .B(G143), .ZN(new_n189));
  AOI21_X1  g003(.A(new_n188), .B1(new_n189), .B2(new_n187), .ZN(new_n190));
  INV_X1    g004(.A(G128), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n187), .A2(G143), .ZN(new_n192));
  AOI21_X1  g006(.A(new_n191), .B1(new_n192), .B2(KEYINPUT1), .ZN(new_n193));
  OAI21_X1  g007(.A(KEYINPUT67), .B1(new_n190), .B2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G143), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(KEYINPUT65), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT65), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G143), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n196), .A2(new_n198), .A3(new_n187), .ZN(new_n199));
  INV_X1    g013(.A(new_n188), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(new_n193), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT67), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g018(.A(KEYINPUT66), .B1(new_n195), .B2(G146), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT66), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n206), .A2(new_n187), .A3(G143), .ZN(new_n207));
  AND2_X1   g021(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n197), .A2(G143), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n195), .A2(KEYINPUT65), .ZN(new_n210));
  OAI21_X1  g024(.A(G146), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n191), .A2(KEYINPUT1), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n208), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n194), .A2(new_n204), .A3(new_n213), .ZN(new_n214));
  OR3_X1    g028(.A1(new_n214), .A2(KEYINPUT81), .A3(G125), .ZN(new_n215));
  NAND2_X1  g029(.A1(KEYINPUT0), .A2(G128), .ZN(new_n216));
  XNOR2_X1  g030(.A(new_n216), .B(KEYINPUT64), .ZN(new_n217));
  OAI211_X1 g031(.A(new_n201), .B(new_n217), .C1(KEYINPUT0), .C2(G128), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n208), .A2(new_n211), .A3(KEYINPUT0), .A4(G128), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G125), .ZN(new_n221));
  OAI21_X1  g035(.A(KEYINPUT81), .B1(new_n214), .B2(G125), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n215), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  XOR2_X1   g037(.A(KEYINPUT82), .B(G224), .Z(new_n224));
  INV_X1    g038(.A(new_n224), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n225), .A2(G953), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n223), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(new_n226), .ZN(new_n228));
  NAND4_X1  g042(.A1(new_n215), .A2(new_n228), .A3(new_n221), .A4(new_n222), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(KEYINPUT7), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT7), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n223), .A2(new_n232), .ZN(new_n233));
  NOR2_X1   g047(.A1(KEYINPUT2), .A2(G113), .ZN(new_n234));
  NAND2_X1  g048(.A1(KEYINPUT2), .A2(G113), .ZN(new_n235));
  OR2_X1    g049(.A1(new_n235), .A2(KEYINPUT69), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(KEYINPUT69), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n234), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  XNOR2_X1  g052(.A(G116), .B(G119), .ZN(new_n239));
  XNOR2_X1  g053(.A(new_n238), .B(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(G104), .ZN(new_n241));
  OAI21_X1  g055(.A(KEYINPUT3), .B1(new_n241), .B2(G107), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT3), .ZN(new_n243));
  INV_X1    g057(.A(G107), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n243), .A2(new_n244), .A3(G104), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n241), .A2(G107), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n242), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT4), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n247), .A2(new_n248), .A3(G101), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n247), .A2(G101), .ZN(new_n250));
  INV_X1    g064(.A(G101), .ZN(new_n251));
  NAND4_X1  g065(.A1(new_n242), .A2(new_n245), .A3(new_n251), .A4(new_n246), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n250), .A2(KEYINPUT4), .A3(new_n252), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n240), .A2(new_n249), .A3(new_n253), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n241), .A2(G107), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n244), .A2(G104), .ZN(new_n256));
  OAI21_X1  g070(.A(G101), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n252), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(KEYINPUT78), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT78), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n252), .A2(new_n257), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n238), .A2(new_n239), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n239), .A2(KEYINPUT5), .ZN(new_n264));
  INV_X1    g078(.A(G119), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(G116), .ZN(new_n266));
  OAI211_X1 g080(.A(new_n264), .B(G113), .C1(KEYINPUT5), .C2(new_n266), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n262), .A2(new_n263), .A3(new_n267), .ZN(new_n268));
  XNOR2_X1  g082(.A(G110), .B(G122), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n254), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(new_n258), .ZN(new_n271));
  AND2_X1   g085(.A1(new_n267), .A2(new_n263), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n268), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  XNOR2_X1  g087(.A(KEYINPUT83), .B(KEYINPUT8), .ZN(new_n274));
  OR2_X1    g088(.A1(new_n269), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n269), .A2(new_n274), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n273), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  AND3_X1   g091(.A1(new_n233), .A2(new_n270), .A3(new_n277), .ZN(new_n278));
  AOI21_X1  g092(.A(G902), .B1(new_n231), .B2(new_n278), .ZN(new_n279));
  OAI21_X1  g093(.A(G210), .B1(G237), .B2(G902), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n254), .A2(new_n268), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT6), .ZN(new_n282));
  INV_X1    g096(.A(new_n269), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n281), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n281), .A2(new_n283), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n285), .A2(KEYINPUT6), .A3(new_n270), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n230), .A2(new_n284), .A3(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n279), .A2(new_n280), .A3(new_n287), .ZN(new_n288));
  XOR2_X1   g102(.A(new_n280), .B(KEYINPUT84), .Z(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(G902), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n232), .B1(new_n227), .B2(new_n229), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n233), .A2(new_n270), .A3(new_n277), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n291), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(new_n230), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n286), .A2(new_n284), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n290), .B1(new_n294), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n288), .A2(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(G214), .B1(G237), .B2(G902), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  XNOR2_X1  g115(.A(G113), .B(G122), .ZN(new_n302));
  XNOR2_X1  g116(.A(new_n302), .B(new_n241), .ZN(new_n303));
  INV_X1    g117(.A(G131), .ZN(new_n304));
  INV_X1    g118(.A(G237), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(KEYINPUT70), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT70), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(G237), .ZN(new_n308));
  AOI21_X1  g122(.A(G953), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n196), .A2(new_n198), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT85), .ZN(new_n311));
  AOI22_X1  g125(.A1(new_n309), .A2(G214), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  XNOR2_X1  g126(.A(KEYINPUT70), .B(G237), .ZN(new_n313));
  NAND2_X1  g127(.A1(KEYINPUT65), .A2(KEYINPUT85), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(new_n195), .ZN(new_n315));
  INV_X1    g129(.A(G214), .ZN(new_n316));
  NOR4_X1   g130(.A1(new_n313), .A2(new_n315), .A3(new_n316), .A4(G953), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n304), .B1(new_n312), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n306), .A2(new_n308), .ZN(new_n319));
  INV_X1    g133(.A(G953), .ZN(new_n320));
  AOI21_X1  g134(.A(G143), .B1(KEYINPUT65), .B2(KEYINPUT85), .ZN(new_n321));
  NAND4_X1  g135(.A1(new_n319), .A2(G214), .A3(new_n320), .A4(new_n321), .ZN(new_n322));
  NOR3_X1   g136(.A1(new_n313), .A2(new_n316), .A3(G953), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n189), .A2(KEYINPUT85), .ZN(new_n324));
  OAI211_X1 g138(.A(G131), .B(new_n322), .C1(new_n323), .C2(new_n324), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n318), .A2(KEYINPUT86), .A3(new_n325), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n322), .B1(new_n323), .B2(new_n324), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT86), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n327), .A2(new_n328), .A3(new_n304), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n326), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(KEYINPUT87), .ZN(new_n331));
  XNOR2_X1  g145(.A(G125), .B(G140), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(KEYINPUT16), .ZN(new_n333));
  INV_X1    g147(.A(G125), .ZN(new_n334));
  OR3_X1    g148(.A1(new_n334), .A2(KEYINPUT16), .A3(G140), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n336), .A2(new_n187), .ZN(new_n337));
  XNOR2_X1  g151(.A(new_n337), .B(KEYINPUT75), .ZN(new_n338));
  XOR2_X1   g152(.A(new_n332), .B(KEYINPUT19), .Z(new_n339));
  OR2_X1    g153(.A1(new_n339), .A2(G146), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT87), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n326), .A2(new_n329), .A3(new_n341), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n331), .A2(new_n338), .A3(new_n340), .A4(new_n342), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n312), .A2(new_n317), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n344), .A2(KEYINPUT18), .A3(G131), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT18), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n327), .A2(new_n346), .ZN(new_n347));
  XNOR2_X1  g161(.A(new_n332), .B(new_n187), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n345), .A2(new_n347), .A3(new_n318), .A4(new_n348), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n303), .B1(new_n343), .B2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT17), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n330), .A2(new_n351), .ZN(new_n352));
  XNOR2_X1  g166(.A(new_n336), .B(G146), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n344), .A2(KEYINPUT88), .A3(KEYINPUT17), .A4(G131), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT88), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n355), .B1(new_n325), .B2(new_n351), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n352), .A2(new_n353), .A3(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n359), .A2(new_n303), .A3(new_n349), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT89), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(new_n349), .ZN(new_n363));
  INV_X1    g177(.A(new_n353), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n364), .B1(new_n330), .B2(new_n351), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n363), .B1(new_n365), .B2(new_n358), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n366), .A2(KEYINPUT89), .A3(new_n303), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n350), .B1(new_n362), .B2(new_n367), .ZN(new_n368));
  NOR2_X1   g182(.A1(G475), .A2(G902), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  OAI21_X1  g184(.A(KEYINPUT20), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n343), .A2(new_n349), .ZN(new_n372));
  INV_X1    g186(.A(new_n303), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g188(.A(KEYINPUT89), .B1(new_n366), .B2(new_n303), .ZN(new_n375));
  AOI21_X1  g189(.A(KEYINPUT17), .B1(new_n326), .B2(new_n329), .ZN(new_n376));
  NOR3_X1   g190(.A1(new_n376), .A2(new_n364), .A3(new_n357), .ZN(new_n377));
  NOR4_X1   g191(.A1(new_n377), .A2(new_n361), .A3(new_n373), .A4(new_n363), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n374), .B1(new_n375), .B2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT20), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n379), .A2(new_n380), .A3(new_n369), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n371), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(G234), .A2(G237), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n383), .A2(G952), .A3(new_n320), .ZN(new_n384));
  XOR2_X1   g198(.A(new_n384), .B(KEYINPUT93), .Z(new_n385));
  XOR2_X1   g199(.A(KEYINPUT21), .B(G898), .Z(new_n386));
  XNOR2_X1  g200(.A(KEYINPUT73), .B(G902), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n387), .A2(G953), .A3(new_n383), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n385), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n195), .A2(G128), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  OAI211_X1 g205(.A(KEYINPUT13), .B(new_n391), .C1(new_n189), .C2(new_n191), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n191), .B1(new_n196), .B2(new_n198), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT13), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n392), .A2(new_n395), .A3(G134), .ZN(new_n396));
  INV_X1    g210(.A(G134), .ZN(new_n397));
  OAI211_X1 g211(.A(new_n397), .B(new_n391), .C1(new_n189), .C2(new_n191), .ZN(new_n398));
  INV_X1    g212(.A(G122), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(G116), .ZN(new_n400));
  INV_X1    g214(.A(G116), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(G122), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n244), .B1(new_n400), .B2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n400), .A2(new_n402), .A3(new_n244), .ZN(new_n405));
  AOI21_X1  g219(.A(KEYINPUT90), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  AND3_X1   g220(.A1(new_n400), .A2(new_n402), .A3(new_n244), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT90), .ZN(new_n408));
  NOR3_X1   g222(.A1(new_n407), .A2(new_n403), .A3(new_n408), .ZN(new_n409));
  OAI211_X1 g223(.A(new_n396), .B(new_n398), .C1(new_n406), .C2(new_n409), .ZN(new_n410));
  OAI21_X1  g224(.A(G134), .B1(new_n393), .B2(new_n390), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(new_n398), .ZN(new_n412));
  XNOR2_X1  g226(.A(new_n405), .B(KEYINPUT91), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n401), .A2(KEYINPUT14), .A3(G122), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n400), .A2(new_n402), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n414), .B(G107), .C1(new_n415), .C2(KEYINPUT14), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n412), .A2(new_n413), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n410), .A2(new_n417), .ZN(new_n418));
  XNOR2_X1  g232(.A(KEYINPUT9), .B(G234), .ZN(new_n419));
  INV_X1    g233(.A(G217), .ZN(new_n420));
  NOR3_X1   g234(.A1(new_n419), .A2(new_n420), .A3(G953), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n418), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n410), .A2(new_n417), .A3(new_n421), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n423), .A2(KEYINPUT92), .A3(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(new_n387), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT92), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n418), .A2(new_n427), .A3(new_n422), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n425), .A2(new_n426), .A3(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(G478), .ZN(new_n430));
  OR2_X1    g244(.A1(new_n430), .A2(KEYINPUT15), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n429), .B(new_n431), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n366), .A2(new_n303), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n433), .B1(new_n362), .B2(new_n367), .ZN(new_n434));
  OAI21_X1  g248(.A(G475), .B1(new_n434), .B2(G902), .ZN(new_n435));
  NAND4_X1  g249(.A1(new_n382), .A2(new_n389), .A3(new_n432), .A4(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT94), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  OAI22_X1  g252(.A1(new_n375), .A2(new_n378), .B1(new_n303), .B2(new_n366), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(new_n291), .ZN(new_n440));
  AOI22_X1  g254(.A1(new_n371), .A2(new_n381), .B1(new_n440), .B2(G475), .ZN(new_n441));
  NAND4_X1  g255(.A1(new_n441), .A2(KEYINPUT94), .A3(new_n389), .A4(new_n432), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n301), .B1(new_n438), .B2(new_n442), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n265), .A2(G128), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n265), .A2(G128), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n444), .B1(KEYINPUT23), .B2(new_n445), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n446), .B1(KEYINPUT23), .B2(new_n444), .ZN(new_n447));
  INV_X1    g261(.A(G110), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(new_n444), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(new_n445), .ZN(new_n451));
  XNOR2_X1  g265(.A(KEYINPUT24), .B(G110), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  AOI22_X1  g267(.A1(new_n449), .A2(new_n453), .B1(new_n187), .B2(new_n332), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n338), .A2(new_n454), .ZN(new_n455));
  OAI22_X1  g269(.A1(new_n447), .A2(new_n448), .B1(new_n451), .B2(new_n452), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n455), .B1(new_n353), .B2(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n320), .A2(G221), .A3(G234), .ZN(new_n458));
  XNOR2_X1  g272(.A(new_n458), .B(KEYINPUT76), .ZN(new_n459));
  XOR2_X1   g273(.A(KEYINPUT22), .B(G137), .Z(new_n460));
  XNOR2_X1  g274(.A(new_n459), .B(new_n460), .ZN(new_n461));
  XNOR2_X1  g275(.A(new_n457), .B(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  NOR2_X1   g277(.A1(KEYINPUT77), .A2(KEYINPUT25), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n463), .A2(new_n426), .A3(new_n464), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n420), .B1(new_n426), .B2(G234), .ZN(new_n466));
  OAI22_X1  g280(.A1(new_n462), .A2(new_n387), .B1(KEYINPUT77), .B2(KEYINPUT25), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n466), .A2(G902), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n463), .A2(new_n469), .ZN(new_n470));
  AND2_X1   g284(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT30), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n472), .A2(KEYINPUT68), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(KEYINPUT68), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  XNOR2_X1  g289(.A(G134), .B(G137), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT11), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n477), .B1(new_n397), .B2(G137), .ZN(new_n478));
  INV_X1    g292(.A(G137), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n479), .A2(KEYINPUT11), .A3(G134), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n397), .A2(G137), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n478), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  MUX2_X1   g296(.A(new_n476), .B(new_n482), .S(new_n304), .Z(new_n483));
  NAND2_X1  g297(.A1(new_n214), .A2(new_n483), .ZN(new_n484));
  XNOR2_X1  g298(.A(new_n482), .B(G131), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n485), .A2(new_n218), .A3(new_n219), .ZN(new_n486));
  AOI211_X1 g300(.A(new_n473), .B(new_n475), .C1(new_n484), .C2(new_n486), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n484), .A2(new_n486), .A3(KEYINPUT68), .A4(new_n472), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n240), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT31), .ZN(new_n491));
  INV_X1    g305(.A(new_n240), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n484), .A2(new_n492), .A3(new_n486), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n309), .A2(G210), .ZN(new_n494));
  XNOR2_X1  g308(.A(new_n494), .B(G101), .ZN(new_n495));
  XNOR2_X1  g309(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n496));
  XNOR2_X1  g310(.A(new_n495), .B(new_n496), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n490), .A2(new_n491), .A3(new_n493), .A4(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(KEYINPUT72), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT28), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n493), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n484), .A2(new_n486), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(new_n240), .ZN(new_n503));
  AND2_X1   g317(.A1(new_n503), .A2(new_n493), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n501), .B1(new_n504), .B2(new_n500), .ZN(new_n505));
  INV_X1    g319(.A(new_n497), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n493), .ZN(new_n508));
  INV_X1    g322(.A(new_n473), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n502), .A2(new_n509), .A3(new_n474), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(new_n488), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n508), .B1(new_n511), .B2(new_n240), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT72), .ZN(new_n513));
  NAND4_X1  g327(.A1(new_n512), .A2(new_n513), .A3(new_n491), .A4(new_n497), .ZN(new_n514));
  AND3_X1   g328(.A1(new_n499), .A2(new_n507), .A3(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT71), .ZN(new_n516));
  AOI211_X1 g330(.A(new_n508), .B(new_n506), .C1(new_n511), .C2(new_n240), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n516), .B1(new_n517), .B2(new_n491), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n512), .A2(new_n497), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n519), .A2(KEYINPUT71), .A3(KEYINPUT31), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n515), .A2(new_n521), .ZN(new_n522));
  NOR2_X1   g336(.A1(G472), .A2(G902), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT32), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT74), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n501), .B(new_n497), .C1(new_n504), .C2(new_n500), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT29), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n426), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n512), .A2(new_n497), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n531), .A2(KEYINPUT29), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n530), .B1(new_n532), .B2(new_n528), .ZN(new_n533));
  INV_X1    g347(.A(G472), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n527), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  OAI211_X1 g349(.A(new_n528), .B(new_n529), .C1(new_n497), .C2(new_n512), .ZN(new_n536));
  OAI211_X1 g350(.A(new_n536), .B(new_n426), .C1(new_n529), .C2(new_n528), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n537), .A2(KEYINPUT74), .A3(G472), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n535), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n522), .A2(KEYINPUT32), .A3(new_n523), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n526), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n205), .A2(new_n207), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n542), .B1(G146), .B2(new_n310), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n191), .B1(new_n199), .B2(KEYINPUT1), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n213), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(new_n271), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT10), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n214), .A2(new_n262), .A3(KEYINPUT10), .ZN(new_n549));
  INV_X1    g363(.A(new_n485), .ZN(new_n550));
  NAND4_X1  g364(.A1(new_n253), .A2(new_n218), .A3(new_n219), .A4(new_n249), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n548), .A2(new_n549), .A3(new_n550), .A4(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT79), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(new_n551), .ZN(new_n555));
  AOI21_X1  g369(.A(KEYINPUT10), .B1(new_n545), .B2(new_n271), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND4_X1  g371(.A1(new_n557), .A2(KEYINPUT79), .A3(new_n550), .A4(new_n549), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n554), .A2(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n546), .B1(new_n214), .B2(new_n262), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT12), .ZN(new_n561));
  AND3_X1   g375(.A1(new_n560), .A2(new_n561), .A3(new_n485), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n561), .B1(new_n560), .B2(new_n485), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  XNOR2_X1  g378(.A(G110), .B(G140), .ZN(new_n565));
  INV_X1    g379(.A(G227), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n566), .A2(G953), .ZN(new_n567));
  XOR2_X1   g381(.A(new_n565), .B(new_n567), .Z(new_n568));
  NAND3_X1  g382(.A1(new_n559), .A2(new_n564), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(KEYINPUT80), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n557), .A2(new_n549), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(new_n485), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n559), .A2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(new_n568), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT80), .ZN(new_n576));
  NAND4_X1  g390(.A1(new_n559), .A2(new_n564), .A3(new_n576), .A4(new_n568), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n570), .A2(new_n575), .A3(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(G469), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n578), .A2(new_n579), .A3(new_n426), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n559), .A2(new_n564), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(new_n574), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n559), .A2(new_n572), .A3(new_n568), .ZN(new_n583));
  AND2_X1   g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(G469), .ZN(new_n585));
  NAND2_X1  g399(.A1(G469), .A2(G902), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n580), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  OAI21_X1  g401(.A(G221), .B1(new_n419), .B2(G902), .ZN(new_n588));
  AND2_X1   g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND4_X1  g403(.A1(new_n443), .A2(new_n471), .A3(new_n541), .A4(new_n589), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n590), .B(G101), .ZN(G3));
  AOI21_X1  g405(.A(new_n387), .B1(new_n515), .B2(new_n521), .ZN(new_n592));
  OR3_X1    g406(.A1(new_n592), .A2(KEYINPUT95), .A3(new_n534), .ZN(new_n593));
  OAI21_X1  g407(.A(KEYINPUT95), .B1(new_n592), .B2(new_n534), .ZN(new_n594));
  AND3_X1   g408(.A1(new_n593), .A2(new_n524), .A3(new_n594), .ZN(new_n595));
  AND3_X1   g409(.A1(new_n595), .A2(new_n471), .A3(new_n589), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT33), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n425), .A2(new_n597), .A3(new_n428), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n423), .A2(KEYINPUT33), .A3(new_n424), .ZN(new_n599));
  AND2_X1   g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n600), .A2(KEYINPUT96), .A3(G478), .A4(new_n426), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n429), .A2(new_n430), .ZN(new_n602));
  NAND4_X1  g416(.A1(new_n598), .A2(G478), .A3(new_n426), .A4(new_n599), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT96), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n601), .A2(new_n602), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n606), .A2(KEYINPUT97), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT97), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n601), .A2(new_n608), .A3(new_n602), .A4(new_n605), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  NOR3_X1   g424(.A1(new_n368), .A2(KEYINPUT20), .A3(new_n370), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n380), .B1(new_n379), .B2(new_n369), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n435), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n610), .A2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n300), .ZN(new_n615));
  INV_X1    g429(.A(new_n280), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n616), .B1(new_n294), .B2(new_n297), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n615), .B1(new_n288), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(new_n389), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n614), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n596), .A2(new_n620), .ZN(new_n621));
  XOR2_X1   g435(.A(KEYINPUT34), .B(G104), .Z(new_n622));
  XNOR2_X1  g436(.A(new_n621), .B(new_n622), .ZN(G6));
  INV_X1    g437(.A(KEYINPUT98), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n381), .A2(new_n624), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n379), .A2(KEYINPUT98), .A3(new_n380), .A4(new_n369), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n625), .A2(new_n371), .A3(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n435), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n628), .A2(new_n432), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n630), .A2(new_n619), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n596), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(KEYINPUT99), .ZN(new_n633));
  XNOR2_X1  g447(.A(KEYINPUT35), .B(G107), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G9));
  NOR2_X1   g449(.A1(new_n461), .A2(KEYINPUT36), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n457), .B(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(new_n469), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n468), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n587), .A2(new_n588), .A3(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n595), .A2(new_n443), .A3(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT37), .B(G110), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G12));
  AND2_X1   g458(.A1(new_n541), .A2(new_n618), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n388), .A2(G900), .ZN(new_n646));
  XOR2_X1   g460(.A(new_n646), .B(KEYINPUT100), .Z(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n385), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n627), .A2(new_n629), .A3(new_n648), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n649), .A2(new_n640), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n645), .A2(new_n650), .ZN(new_n651));
  XOR2_X1   g465(.A(KEYINPUT101), .B(G128), .Z(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G30));
  XNOR2_X1  g467(.A(KEYINPUT102), .B(KEYINPUT39), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n648), .B(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n589), .A2(new_n655), .ZN(new_n656));
  AND2_X1   g470(.A1(new_n656), .A2(KEYINPUT40), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n656), .A2(KEYINPUT40), .ZN(new_n658));
  NOR4_X1   g472(.A1(new_n657), .A2(new_n658), .A3(new_n432), .A4(new_n441), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n512), .A2(new_n506), .ZN(new_n660));
  INV_X1    g474(.A(new_n504), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n291), .B1(new_n661), .B2(new_n497), .ZN(new_n662));
  OAI21_X1  g476(.A(G472), .B1(new_n660), .B2(new_n662), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n526), .A2(new_n540), .A3(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n299), .B(KEYINPUT38), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n639), .A2(new_n615), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n659), .A2(new_n664), .A3(new_n665), .A4(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(new_n189), .ZN(G45));
  NAND3_X1  g482(.A1(new_n610), .A2(new_n613), .A3(new_n648), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n669), .A2(new_n640), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n645), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G146), .ZN(G48));
  NAND2_X1  g486(.A1(new_n578), .A2(new_n426), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT103), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n674), .A2(new_n579), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  OAI211_X1 g490(.A(new_n578), .B(new_n426), .C1(new_n674), .C2(new_n579), .ZN(new_n677));
  AND3_X1   g491(.A1(new_n676), .A2(new_n588), .A3(new_n677), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n541), .A2(new_n620), .A3(new_n471), .A4(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(KEYINPUT41), .B(G113), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(G15));
  NAND4_X1  g495(.A1(new_n676), .A2(new_n588), .A3(new_n677), .A4(new_n389), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n630), .A2(new_n682), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n683), .A2(new_n541), .A3(new_n471), .A4(new_n618), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G116), .ZN(G18));
  NAND3_X1  g499(.A1(new_n541), .A2(new_n618), .A3(new_n639), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n438), .A2(new_n442), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(new_n678), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(new_n265), .ZN(G21));
  NAND2_X1  g504(.A1(new_n522), .A2(new_n426), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n499), .A2(new_n514), .A3(new_n507), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n517), .A2(new_n491), .ZN(new_n693));
  OR2_X1    g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  AOI22_X1  g508(.A1(new_n691), .A2(G472), .B1(new_n523), .B2(new_n694), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n695), .A2(new_n678), .A3(new_n471), .A4(new_n389), .ZN(new_n696));
  OAI21_X1  g510(.A(KEYINPUT104), .B1(new_n441), .B2(new_n432), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT104), .ZN(new_n698));
  INV_X1    g512(.A(new_n432), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n613), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n697), .A2(new_n700), .A3(new_n618), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(KEYINPUT105), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT105), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n697), .A2(new_n700), .A3(new_n703), .A4(new_n618), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n696), .B1(new_n702), .B2(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(new_n399), .ZN(G24));
  AOI21_X1  g520(.A(new_n441), .B1(new_n609), .B2(new_n607), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n695), .A2(new_n707), .A3(new_n648), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n678), .A2(new_n618), .A3(new_n639), .ZN(new_n709));
  OAI21_X1  g523(.A(KEYINPUT106), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n523), .B1(new_n692), .B2(new_n693), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n711), .B1(new_n592), .B2(new_n534), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n669), .A2(new_n712), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n618), .A2(new_n676), .A3(new_n588), .A4(new_n677), .ZN(new_n714));
  INV_X1    g528(.A(new_n639), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT106), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n713), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n710), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G125), .ZN(G27));
  INV_X1    g534(.A(KEYINPUT42), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n288), .A2(new_n298), .A3(new_n300), .ZN(new_n722));
  INV_X1    g536(.A(new_n588), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  OR2_X1    g538(.A1(new_n583), .A2(KEYINPUT107), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n583), .A2(KEYINPUT107), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n725), .A2(G469), .A3(new_n582), .A4(new_n726), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n580), .A2(new_n586), .A3(new_n727), .ZN(new_n728));
  AND3_X1   g542(.A1(new_n724), .A2(new_n728), .A3(KEYINPUT108), .ZN(new_n729));
  AOI21_X1  g543(.A(KEYINPUT108), .B1(new_n724), .B2(new_n728), .ZN(new_n730));
  OAI211_X1 g544(.A(new_n541), .B(new_n471), .C1(new_n729), .C2(new_n730), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n721), .B1(new_n731), .B2(new_n669), .ZN(new_n732));
  AND2_X1   g546(.A1(new_n541), .A2(new_n471), .ZN(new_n733));
  INV_X1    g547(.A(new_n669), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n724), .A2(new_n728), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT108), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n724), .A2(new_n728), .A3(KEYINPUT108), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n733), .A2(KEYINPUT42), .A3(new_n734), .A4(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n732), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G131), .ZN(G33));
  OR2_X1    g556(.A1(new_n731), .A2(new_n649), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G134), .ZN(G36));
  AND2_X1   g558(.A1(new_n610), .A2(new_n441), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT43), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n746), .B1(new_n613), .B2(KEYINPUT110), .ZN(new_n747));
  OR2_X1    g561(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n745), .A2(new_n747), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(new_n595), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n750), .A2(new_n751), .A3(new_n639), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT44), .ZN(new_n753));
  OR2_X1    g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(new_n722), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n725), .A2(KEYINPUT45), .A3(new_n582), .A4(new_n726), .ZN(new_n756));
  OAI211_X1 g570(.A(new_n756), .B(G469), .C1(KEYINPUT45), .C2(new_n584), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n757), .A2(KEYINPUT46), .A3(new_n586), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(new_n580), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(KEYINPUT109), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n757), .A2(new_n586), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT46), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT109), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n758), .A2(new_n764), .A3(new_n580), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n760), .A2(new_n763), .A3(new_n765), .ZN(new_n766));
  AND3_X1   g580(.A1(new_n766), .A2(new_n588), .A3(new_n655), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n752), .A2(new_n753), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n754), .A2(new_n755), .A3(new_n767), .A4(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G137), .ZN(G39));
  NAND2_X1  g584(.A1(new_n766), .A2(new_n588), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(KEYINPUT47), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT47), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n766), .A2(new_n773), .A3(new_n588), .ZN(new_n774));
  NOR3_X1   g588(.A1(new_n541), .A2(new_n471), .A3(new_n722), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n772), .A2(new_n734), .A3(new_n774), .A4(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G140), .ZN(G42));
  NAND4_X1  g591(.A1(new_n745), .A2(new_n471), .A3(new_n588), .A4(new_n300), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT111), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n780), .A2(new_n664), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n665), .B1(new_n778), .B2(new_n779), .ZN(new_n782));
  AND2_X1   g596(.A1(new_n676), .A2(new_n677), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(KEYINPUT49), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n781), .A2(new_n782), .A3(new_n784), .ZN(new_n785));
  XOR2_X1   g599(.A(new_n785), .B(KEYINPUT112), .Z(new_n786));
  INV_X1    g600(.A(new_n471), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n678), .A2(new_n755), .ZN(new_n788));
  OR4_X1    g602(.A1(new_n787), .A2(new_n664), .A3(new_n788), .A4(new_n385), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n789), .A2(new_n614), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n320), .A2(G952), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n695), .A2(new_n471), .ZN(new_n792));
  AOI211_X1 g606(.A(new_n385), .B(new_n792), .C1(new_n748), .C2(new_n749), .ZN(new_n793));
  INV_X1    g607(.A(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n772), .A2(new_n774), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n783), .A2(new_n723), .ZN(new_n796));
  AOI211_X1 g610(.A(new_n722), .B(new_n794), .C1(new_n795), .C2(new_n796), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n385), .B1(new_n748), .B2(new_n749), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n678), .A2(new_n615), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n665), .B1(new_n799), .B2(KEYINPUT117), .ZN(new_n800));
  INV_X1    g614(.A(new_n792), .ZN(new_n801));
  OR2_X1    g615(.A1(new_n799), .A2(KEYINPUT117), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n798), .A2(new_n800), .A3(new_n801), .A4(new_n802), .ZN(new_n803));
  NOR2_X1   g617(.A1(KEYINPUT118), .A2(KEYINPUT50), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(new_n804), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n793), .A2(new_n806), .A3(new_n802), .A4(new_n800), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(new_n788), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n798), .A2(new_n639), .A3(new_n695), .A4(new_n809), .ZN(new_n810));
  OR3_X1    g624(.A1(new_n789), .A2(new_n613), .A3(new_n610), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n808), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n797), .B1(KEYINPUT119), .B2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT119), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n808), .A2(new_n814), .A3(new_n810), .A4(new_n811), .ZN(new_n815));
  AND2_X1   g629(.A1(new_n815), .A2(KEYINPUT51), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n791), .B1(new_n813), .B2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT51), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n795), .A2(new_n796), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT116), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n819), .A2(new_n820), .A3(new_n755), .A4(new_n793), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n821), .A2(new_n810), .A3(new_n808), .A4(new_n811), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n797), .A2(new_n820), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n818), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n798), .A2(new_n733), .A3(new_n809), .ZN(new_n825));
  XNOR2_X1  g639(.A(new_n825), .B(KEYINPUT48), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n793), .A2(new_n618), .A3(new_n678), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n817), .A2(new_n824), .A3(new_n826), .A4(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT52), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT114), .ZN(new_n830));
  OAI211_X1 g644(.A(new_n541), .B(new_n618), .C1(new_n650), .C2(new_n670), .ZN(new_n831));
  AND3_X1   g645(.A1(new_n713), .A2(new_n717), .A3(new_n716), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n717), .B1(new_n713), .B2(new_n716), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n831), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(new_n648), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n639), .A2(new_n835), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n664), .A2(new_n588), .A3(new_n728), .A4(new_n836), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n837), .B1(new_n704), .B2(new_n702), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n830), .B1(new_n834), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n702), .A2(new_n704), .ZN(new_n840));
  INV_X1    g654(.A(new_n837), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n842), .A2(new_n719), .A3(KEYINPUT114), .A4(new_n831), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n829), .B1(new_n839), .B2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(new_n844), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n713), .B1(new_n729), .B2(new_n730), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n722), .A2(new_n628), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT113), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n699), .A2(new_n835), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n847), .A2(new_n627), .A3(new_n848), .A4(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n541), .A2(new_n589), .A3(new_n850), .ZN(new_n851));
  AND2_X1   g665(.A1(new_n627), .A2(new_n849), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n848), .B1(new_n852), .B2(new_n847), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n846), .B1(new_n851), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(new_n639), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n741), .A2(new_n743), .A3(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n684), .A2(new_n679), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n705), .A2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(new_n689), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n299), .A2(new_n300), .A3(new_n389), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n441), .A2(new_n699), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n861), .B1(new_n614), .B2(new_n862), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n595), .A2(new_n863), .A3(new_n471), .A4(new_n589), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n864), .A2(new_n590), .A3(new_n642), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n856), .A2(new_n860), .A3(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n839), .A2(new_n829), .A3(new_n843), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n845), .A2(new_n866), .A3(KEYINPUT53), .A4(new_n867), .ZN(new_n868));
  OAI21_X1  g682(.A(KEYINPUT52), .B1(new_n834), .B2(new_n838), .ZN(new_n869));
  AND3_X1   g683(.A1(new_n866), .A2(new_n867), .A3(new_n869), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n868), .B1(new_n870), .B2(KEYINPUT53), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n871), .A2(KEYINPUT54), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT53), .ZN(new_n873));
  AND3_X1   g687(.A1(new_n741), .A2(new_n743), .A3(new_n855), .ZN(new_n874));
  NOR4_X1   g688(.A1(new_n865), .A2(new_n705), .A3(new_n857), .A4(new_n689), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n867), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n873), .B1(new_n876), .B2(new_n844), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT54), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n866), .A2(KEYINPUT53), .A3(new_n869), .A4(new_n867), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n872), .A2(KEYINPUT115), .A3(new_n880), .ZN(new_n881));
  OR2_X1    g695(.A1(new_n880), .A2(KEYINPUT115), .ZN(new_n882));
  AOI211_X1 g696(.A(new_n790), .B(new_n828), .C1(new_n881), .C2(new_n882), .ZN(new_n883));
  NOR2_X1   g697(.A1(G952), .A2(G953), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n786), .B1(new_n883), .B2(new_n884), .ZN(G75));
  NAND2_X1  g699(.A1(new_n295), .A2(new_n296), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n886), .A2(new_n287), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n887), .B(KEYINPUT55), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n888), .A2(KEYINPUT56), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n877), .A2(new_n879), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n890), .A2(new_n387), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n889), .B1(new_n891), .B2(new_n289), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n320), .A2(G952), .ZN(new_n893));
  XOR2_X1   g707(.A(new_n893), .B(KEYINPUT120), .Z(new_n894));
  INV_X1    g708(.A(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(new_n888), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n426), .B1(new_n877), .B2(new_n879), .ZN(new_n897));
  AOI21_X1  g711(.A(KEYINPUT56), .B1(new_n897), .B2(new_n616), .ZN(new_n898));
  OAI211_X1 g712(.A(new_n892), .B(new_n895), .C1(new_n896), .C2(new_n898), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n899), .B(KEYINPUT121), .ZN(G51));
  XOR2_X1   g714(.A(new_n586), .B(KEYINPUT57), .Z(new_n901));
  INV_X1    g715(.A(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n890), .A2(KEYINPUT54), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n902), .B1(new_n903), .B2(new_n880), .ZN(new_n904));
  INV_X1    g718(.A(new_n578), .ZN(new_n905));
  OAI21_X1  g719(.A(KEYINPUT122), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  OR2_X1    g720(.A1(new_n891), .A2(new_n757), .ZN(new_n907));
  AND3_X1   g721(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n878), .B1(new_n877), .B2(new_n879), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n901), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT122), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n910), .A2(new_n911), .A3(new_n578), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n906), .A2(new_n907), .A3(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(new_n893), .ZN(new_n914));
  AND2_X1   g728(.A1(new_n913), .A2(new_n914), .ZN(G54));
  NAND3_X1  g729(.A1(new_n897), .A2(KEYINPUT58), .A3(G475), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n916), .B(new_n368), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n917), .A2(new_n893), .ZN(G60));
  NAND2_X1  g732(.A1(G478), .A2(G902), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n919), .B(KEYINPUT59), .ZN(new_n920));
  OAI211_X1 g734(.A(new_n600), .B(new_n920), .C1(new_n908), .C2(new_n909), .ZN(new_n921));
  INV_X1    g735(.A(new_n921), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n881), .A2(new_n882), .A3(new_n920), .ZN(new_n923));
  INV_X1    g737(.A(new_n600), .ZN(new_n924));
  AOI211_X1 g738(.A(new_n894), .B(new_n922), .C1(new_n923), .C2(new_n924), .ZN(G63));
  NAND2_X1  g739(.A1(G217), .A2(G902), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n926), .B(KEYINPUT123), .Z(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(KEYINPUT60), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n928), .B1(new_n877), .B2(new_n879), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n894), .B1(new_n929), .B2(new_n637), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n930), .B1(new_n463), .B2(new_n929), .ZN(new_n931));
  XOR2_X1   g745(.A(KEYINPUT124), .B(KEYINPUT61), .Z(new_n932));
  XNOR2_X1  g746(.A(new_n931), .B(new_n932), .ZN(G66));
  INV_X1    g747(.A(new_n386), .ZN(new_n934));
  OAI21_X1  g748(.A(G953), .B1(new_n225), .B2(new_n934), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n935), .B1(new_n875), .B2(G953), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(KEYINPUT125), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n296), .B1(G898), .B2(new_n320), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n937), .B(new_n938), .ZN(G69));
  INV_X1    g753(.A(new_n834), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n667), .A2(new_n940), .ZN(new_n941));
  XOR2_X1   g755(.A(new_n941), .B(KEYINPUT62), .Z(new_n942));
  NAND2_X1  g756(.A1(new_n614), .A2(new_n862), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n733), .A2(new_n943), .ZN(new_n944));
  OR3_X1    g758(.A1(new_n944), .A2(new_n656), .A3(new_n722), .ZN(new_n945));
  AND2_X1   g759(.A1(new_n769), .A2(new_n945), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n942), .A2(new_n946), .A3(new_n776), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(KEYINPUT126), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT126), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n942), .A2(new_n946), .A3(new_n949), .A4(new_n776), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n511), .B(new_n339), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n951), .A2(new_n320), .A3(new_n952), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n952), .B1(new_n566), .B2(G953), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n954), .B1(new_n566), .B2(new_n952), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n320), .B1(new_n955), .B2(G900), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n741), .A2(new_n743), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n776), .A2(new_n940), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n754), .A2(new_n755), .A3(new_n768), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n840), .A2(new_n733), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  AOI211_X1 g775(.A(new_n957), .B(new_n958), .C1(new_n961), .C2(new_n767), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n956), .B1(new_n962), .B2(new_n954), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n953), .A2(new_n963), .ZN(G72));
  INV_X1    g778(.A(new_n660), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n948), .A2(new_n875), .A3(new_n950), .ZN(new_n966));
  NAND2_X1  g780(.A1(G472), .A2(G902), .ZN(new_n967));
  XOR2_X1   g781(.A(new_n967), .B(KEYINPUT63), .Z(new_n968));
  XOR2_X1   g782(.A(new_n968), .B(KEYINPUT127), .Z(new_n969));
  AOI21_X1  g783(.A(new_n965), .B1(new_n966), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n512), .A2(new_n506), .ZN(new_n971));
  AND4_X1   g785(.A1(new_n965), .A2(new_n871), .A3(new_n968), .A4(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n962), .A2(new_n875), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n971), .B1(new_n973), .B2(new_n969), .ZN(new_n974));
  NOR4_X1   g788(.A1(new_n970), .A2(new_n893), .A3(new_n972), .A4(new_n974), .ZN(G57));
endmodule


