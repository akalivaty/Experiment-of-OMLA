

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761;

  INV_X1 U375 ( .A(n532), .ZN(n680) );
  NOR2_X1 U376 ( .A1(n723), .A2(G902), .ZN(n512) );
  XNOR2_X1 U377 ( .A(n352), .B(n401), .ZN(n399) );
  NAND2_X1 U378 ( .A1(n606), .A2(n366), .ZN(n352) );
  NOR2_X2 U379 ( .A1(n588), .A2(n587), .ZN(n593) );
  XNOR2_X1 U380 ( .A(n388), .B(KEYINPUT19), .ZN(n457) );
  XNOR2_X1 U381 ( .A(n497), .B(n432), .ZN(n740) );
  XNOR2_X2 U382 ( .A(G119), .B(KEYINPUT71), .ZN(n405) );
  XNOR2_X2 U383 ( .A(n398), .B(n364), .ZN(n629) );
  NAND2_X1 U384 ( .A1(n457), .A2(n357), .ZN(n429) );
  XNOR2_X2 U385 ( .A(G113), .B(KEYINPUT94), .ZN(n426) );
  XNOR2_X2 U386 ( .A(KEYINPUT72), .B(KEYINPUT3), .ZN(n404) );
  XNOR2_X2 U387 ( .A(n554), .B(KEYINPUT33), .ZN(n702) );
  NOR2_X2 U388 ( .A1(n564), .A2(n553), .ZN(n554) );
  XNOR2_X2 U389 ( .A(n447), .B(n446), .ZN(n542) );
  NOR2_X1 U390 ( .A1(n670), .A2(n673), .ZN(n698) );
  XNOR2_X1 U391 ( .A(n462), .B(n461), .ZN(n494) );
  XNOR2_X1 U392 ( .A(n373), .B(G143), .ZN(n462) );
  AND2_X1 U393 ( .A1(n380), .A2(n379), .ZN(n676) );
  XNOR2_X1 U394 ( .A(n605), .B(KEYINPUT42), .ZN(n760) );
  XNOR2_X1 U395 ( .A(n396), .B(n599), .ZN(n699) );
  NAND2_X1 U396 ( .A1(n694), .A2(n693), .ZN(n396) );
  XNOR2_X1 U397 ( .A(n375), .B(n374), .ZN(n496) );
  XNOR2_X1 U398 ( .A(G146), .B(KEYINPUT69), .ZN(n375) );
  XNOR2_X1 U399 ( .A(G128), .B(KEYINPUT65), .ZN(n373) );
  XNOR2_X1 U400 ( .A(n505), .B(n376), .ZN(n640) );
  NOR2_X2 U401 ( .A1(n719), .A2(n612), .ZN(n605) );
  XOR2_X1 U402 ( .A(G137), .B(KEYINPUT70), .Z(n518) );
  OR2_X1 U403 ( .A1(n565), .A2(KEYINPUT34), .ZN(n353) );
  XNOR2_X1 U404 ( .A(n494), .B(n425), .ZN(n505) );
  XNOR2_X1 U405 ( .A(n496), .B(G131), .ZN(n425) );
  AND2_X1 U406 ( .A1(n408), .A2(n410), .ZN(n372) );
  AND2_X1 U407 ( .A1(n746), .A2(n409), .ZN(n408) );
  NOR2_X1 U408 ( .A1(n601), .A2(n600), .ZN(n602) );
  NAND2_X1 U409 ( .A1(n394), .A2(n393), .ZN(n392) );
  NOR2_X1 U410 ( .A1(n620), .A2(n759), .ZN(n621) );
  XNOR2_X1 U411 ( .A(n397), .B(KEYINPUT38), .ZN(n598) );
  XNOR2_X1 U412 ( .A(n501), .B(KEYINPUT5), .ZN(n378) );
  XNOR2_X1 U413 ( .A(G137), .B(G101), .ZN(n501) );
  INV_X1 U414 ( .A(KEYINPUT78), .ZN(n516) );
  XNOR2_X1 U415 ( .A(KEYINPUT24), .B(KEYINPUT73), .ZN(n517) );
  XNOR2_X1 U416 ( .A(G128), .B(G110), .ZN(n514) );
  NAND2_X1 U417 ( .A1(n407), .A2(n406), .ZN(n371) );
  NAND2_X1 U418 ( .A1(n415), .A2(n616), .ZN(n414) );
  NAND2_X1 U419 ( .A1(n565), .A2(KEYINPUT34), .ZN(n415) );
  BUF_X2 U420 ( .A(n542), .Z(n397) );
  NAND2_X1 U421 ( .A1(n640), .A2(n525), .ZN(n503) );
  NOR2_X1 U422 ( .A1(n717), .A2(n421), .ZN(n418) );
  NAND2_X1 U423 ( .A1(n355), .A2(n757), .ZN(n563) );
  INV_X1 U424 ( .A(KEYINPUT75), .ZN(n561) );
  INV_X1 U425 ( .A(KEYINPUT46), .ZN(n401) );
  INV_X1 U426 ( .A(KEYINPUT4), .ZN(n374) );
  XNOR2_X1 U427 ( .A(G143), .B(G113), .ZN(n475) );
  XNOR2_X1 U428 ( .A(KEYINPUT18), .B(G125), .ZN(n437) );
  XNOR2_X1 U429 ( .A(n603), .B(n513), .ZN(n532) );
  NOR2_X1 U430 ( .A1(n696), .A2(n552), .ZN(n427) );
  XNOR2_X1 U431 ( .A(G122), .B(G104), .ZN(n476) );
  INV_X1 U432 ( .A(G953), .ZN(n734) );
  XNOR2_X1 U433 ( .A(G107), .B(G116), .ZN(n458) );
  XOR2_X1 U434 ( .A(KEYINPUT109), .B(G122), .Z(n459) );
  NOR2_X1 U435 ( .A1(n618), .A2(n598), .ZN(n594) );
  NAND2_X1 U436 ( .A1(n608), .A2(KEYINPUT36), .ZN(n382) );
  NOR2_X1 U437 ( .A1(n609), .A2(n384), .ZN(n383) );
  NAND2_X1 U438 ( .A1(n397), .A2(n385), .ZN(n384) );
  OR2_X1 U439 ( .A1(n612), .A2(n611), .ZN(n622) );
  INV_X1 U440 ( .A(KEYINPUT0), .ZN(n428) );
  XNOR2_X1 U441 ( .A(n570), .B(n569), .ZN(n587) );
  INV_X1 U442 ( .A(KEYINPUT103), .ZN(n569) );
  XNOR2_X1 U443 ( .A(n498), .B(n377), .ZN(n376) );
  XNOR2_X1 U444 ( .A(n378), .B(n500), .ZN(n377) );
  INV_X1 U445 ( .A(KEYINPUT64), .ZN(n436) );
  XNOR2_X1 U446 ( .A(G110), .B(G107), .ZN(n433) );
  XNOR2_X1 U447 ( .A(n522), .B(n365), .ZN(n524) );
  XNOR2_X1 U448 ( .A(n520), .B(n358), .ZN(n365) );
  AND2_X2 U449 ( .A1(n369), .A2(n367), .ZN(n728) );
  OR2_X1 U450 ( .A1(n751), .A2(G952), .ZN(n722) );
  NAND2_X1 U451 ( .A1(n422), .A2(n354), .ZN(n416) );
  NOR2_X1 U452 ( .A1(n713), .A2(n712), .ZN(n714) );
  NAND2_X1 U453 ( .A1(n609), .A2(KEYINPUT36), .ZN(n379) );
  NOR2_X1 U454 ( .A1(n383), .A2(n381), .ZN(n380) );
  NAND2_X1 U455 ( .A1(n680), .A2(n382), .ZN(n381) );
  NAND2_X1 U456 ( .A1(n616), .A2(n397), .ZN(n617) );
  XNOR2_X1 U457 ( .A(n387), .B(n363), .ZN(n550) );
  INV_X1 U458 ( .A(n550), .ZN(n393) );
  NAND2_X1 U459 ( .A1(n424), .A2(KEYINPUT53), .ZN(n354) );
  AND2_X1 U460 ( .A1(n393), .A2(n390), .ZN(n355) );
  NOR2_X1 U461 ( .A1(n626), .A2(n625), .ZN(n356) );
  XOR2_X1 U462 ( .A(n456), .B(KEYINPUT99), .Z(n357) );
  XOR2_X1 U463 ( .A(n515), .B(n514), .Z(n358) );
  AND2_X1 U464 ( .A1(n583), .A2(n582), .ZN(n359) );
  AND2_X1 U465 ( .A1(n667), .A2(n624), .ZN(n360) );
  BUF_X1 U466 ( .A(n532), .Z(n610) );
  INV_X1 U467 ( .A(n397), .ZN(n608) );
  INV_X1 U468 ( .A(n422), .ZN(n421) );
  OR2_X1 U469 ( .A1(n424), .A2(KEYINPUT53), .ZN(n422) );
  AND2_X1 U470 ( .A1(n367), .A2(n423), .ZN(n361) );
  NAND2_X1 U471 ( .A1(n721), .A2(n734), .ZN(n362) );
  INV_X1 U472 ( .A(KEYINPUT36), .ZN(n385) );
  XNOR2_X1 U473 ( .A(KEYINPUT79), .B(KEYINPUT32), .ZN(n363) );
  XNOR2_X1 U474 ( .A(n505), .B(n518), .ZN(n747) );
  XOR2_X1 U475 ( .A(KEYINPUT90), .B(KEYINPUT48), .Z(n364) );
  INV_X1 U476 ( .A(KEYINPUT53), .ZN(n423) );
  XNOR2_X1 U477 ( .A(n517), .B(n516), .ZN(n519) );
  XNOR2_X1 U478 ( .A(n368), .B(n633), .ZN(n716) );
  INV_X1 U479 ( .A(n760), .ZN(n366) );
  NAND2_X1 U480 ( .A1(n392), .A2(n391), .ZN(n560) );
  NAND2_X1 U481 ( .A1(n716), .A2(n407), .ZN(n367) );
  NAND2_X1 U482 ( .A1(n746), .A2(KEYINPUT2), .ZN(n368) );
  NAND2_X1 U483 ( .A1(n370), .A2(n632), .ZN(n369) );
  NAND2_X1 U484 ( .A1(n372), .A2(n371), .ZN(n370) );
  INV_X1 U485 ( .A(n496), .ZN(n495) );
  NAND2_X1 U486 ( .A1(n540), .A2(n693), .ZN(n609) );
  AND2_X1 U487 ( .A1(n546), .A2(n553), .ZN(n545) );
  NAND2_X1 U488 ( .A1(n546), .A2(n386), .ZN(n387) );
  AND2_X1 U489 ( .A1(n544), .A2(n553), .ZN(n386) );
  XNOR2_X2 U490 ( .A(n493), .B(n492), .ZN(n546) );
  NAND2_X1 U491 ( .A1(n542), .A2(n693), .ZN(n388) );
  NAND2_X1 U492 ( .A1(n389), .A2(KEYINPUT91), .ZN(n391) );
  NAND2_X1 U493 ( .A1(n393), .A2(n390), .ZN(n389) );
  INV_X1 U494 ( .A(n638), .ZN(n390) );
  NOR2_X1 U495 ( .A1(n638), .A2(KEYINPUT91), .ZN(n394) );
  XNOR2_X2 U496 ( .A(n395), .B(KEYINPUT41), .ZN(n719) );
  NOR2_X2 U497 ( .A1(n699), .A2(n696), .ZN(n395) );
  NAND2_X1 U498 ( .A1(n400), .A2(n399), .ZN(n398) );
  AND2_X1 U499 ( .A1(n403), .A2(n402), .ZN(n400) );
  NOR2_X1 U500 ( .A1(n676), .A2(n360), .ZN(n403) );
  XNOR2_X1 U501 ( .A(n621), .B(KEYINPUT82), .ZN(n402) );
  XNOR2_X1 U502 ( .A(n405), .B(n404), .ZN(n431) );
  NAND2_X1 U503 ( .A1(n710), .A2(KEYINPUT86), .ZN(n410) );
  XNOR2_X2 U504 ( .A(n586), .B(n585), .ZN(n710) );
  NOR2_X1 U505 ( .A1(n630), .A2(KEYINPUT86), .ZN(n406) );
  INV_X1 U506 ( .A(n710), .ZN(n407) );
  NAND2_X1 U507 ( .A1(n630), .A2(KEYINPUT86), .ZN(n409) );
  INV_X1 U508 ( .A(n457), .ZN(n611) );
  AND2_X2 U509 ( .A1(n549), .A2(n548), .ZN(n638) );
  NAND2_X1 U510 ( .A1(n412), .A2(n411), .ZN(n557) );
  NAND2_X1 U511 ( .A1(n702), .A2(KEYINPUT34), .ZN(n411) );
  NOR2_X1 U512 ( .A1(n413), .A2(n414), .ZN(n412) );
  NOR2_X1 U513 ( .A1(n702), .A2(n353), .ZN(n413) );
  NAND2_X1 U514 ( .A1(n417), .A2(n416), .ZN(n420) );
  NAND2_X1 U515 ( .A1(n715), .A2(n418), .ZN(n417) );
  NAND2_X1 U516 ( .A1(n420), .A2(n419), .ZN(G75) );
  NAND2_X1 U517 ( .A1(n715), .A2(n361), .ZN(n419) );
  NOR2_X1 U518 ( .A1(n718), .A2(n362), .ZN(n424) );
  XNOR2_X1 U519 ( .A(n426), .B(G116), .ZN(n430) );
  INV_X1 U520 ( .A(n571), .ZN(n565) );
  NAND2_X1 U521 ( .A1(n571), .A2(n427), .ZN(n493) );
  NAND2_X1 U522 ( .A1(n574), .A2(n555), .ZN(n696) );
  XNOR2_X2 U523 ( .A(n429), .B(n428), .ZN(n571) );
  AND2_X1 U524 ( .A1(n757), .A2(n558), .ZN(n559) );
  INV_X1 U525 ( .A(G134), .ZN(n461) );
  XNOR2_X1 U526 ( .A(n519), .B(n518), .ZN(n520) );
  INV_X1 U527 ( .A(KEYINPUT117), .ZN(n599) );
  XNOR2_X1 U528 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U529 ( .A(n723), .B(n724), .ZN(n725) );
  XNOR2_X1 U530 ( .A(n726), .B(n725), .ZN(n727) );
  XNOR2_X1 U531 ( .A(n431), .B(n430), .ZN(n497) );
  XNOR2_X1 U532 ( .A(n476), .B(KEYINPUT16), .ZN(n432) );
  XOR2_X1 U533 ( .A(G101), .B(KEYINPUT93), .Z(n434) );
  XNOR2_X1 U534 ( .A(n434), .B(n433), .ZN(n741) );
  INV_X1 U535 ( .A(KEYINPUT74), .ZN(n435) );
  XNOR2_X1 U536 ( .A(n741), .B(n435), .ZN(n508) );
  XNOR2_X1 U537 ( .A(n740), .B(n508), .ZN(n444) );
  XNOR2_X1 U538 ( .A(n495), .B(n462), .ZN(n442) );
  XNOR2_X2 U539 ( .A(n436), .B(G953), .ZN(n751) );
  NAND2_X1 U540 ( .A1(n751), .A2(G224), .ZN(n440) );
  XNOR2_X1 U541 ( .A(KEYINPUT95), .B(KEYINPUT17), .ZN(n438) );
  XNOR2_X1 U542 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U543 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U544 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U545 ( .A(n444), .B(n443), .ZN(n652) );
  XNOR2_X1 U546 ( .A(G902), .B(KEYINPUT15), .ZN(n630) );
  NAND2_X1 U547 ( .A1(n652), .A2(n630), .ZN(n447) );
  INV_X1 U548 ( .A(G902), .ZN(n525) );
  INV_X1 U549 ( .A(G237), .ZN(n445) );
  NAND2_X1 U550 ( .A1(n525), .A2(n445), .ZN(n448) );
  AND2_X1 U551 ( .A1(n448), .A2(G210), .ZN(n446) );
  NAND2_X1 U552 ( .A1(n448), .A2(G214), .ZN(n693) );
  XOR2_X1 U553 ( .A(KEYINPUT77), .B(KEYINPUT14), .Z(n450) );
  NAND2_X1 U554 ( .A1(G237), .A2(G234), .ZN(n449) );
  XNOR2_X1 U555 ( .A(n450), .B(n449), .ZN(n453) );
  NAND2_X1 U556 ( .A1(n453), .A2(G952), .ZN(n451) );
  XNOR2_X1 U557 ( .A(n451), .B(KEYINPUT96), .ZN(n708) );
  NOR2_X1 U558 ( .A1(G953), .A2(n708), .ZN(n536) );
  NOR2_X1 U559 ( .A1(n734), .A2(G898), .ZN(n452) );
  XNOR2_X1 U560 ( .A(n452), .B(KEYINPUT97), .ZN(n742) );
  NAND2_X1 U561 ( .A1(G902), .A2(n453), .ZN(n533) );
  NOR2_X1 U562 ( .A1(n742), .A2(n533), .ZN(n454) );
  XNOR2_X1 U563 ( .A(n454), .B(KEYINPUT98), .ZN(n455) );
  OR2_X1 U564 ( .A1(n536), .A2(n455), .ZN(n456) );
  XNOR2_X1 U565 ( .A(n459), .B(n458), .ZN(n460) );
  XOR2_X1 U566 ( .A(n460), .B(KEYINPUT9), .Z(n464) );
  XNOR2_X1 U567 ( .A(n494), .B(KEYINPUT7), .ZN(n463) );
  XNOR2_X1 U568 ( .A(n464), .B(n463), .ZN(n468) );
  XOR2_X1 U569 ( .A(KEYINPUT84), .B(KEYINPUT8), .Z(n466) );
  NAND2_X1 U570 ( .A1(G234), .A2(n751), .ZN(n465) );
  XNOR2_X1 U571 ( .A(n466), .B(n465), .ZN(n521) );
  NAND2_X1 U572 ( .A1(G217), .A2(n521), .ZN(n467) );
  XOR2_X1 U573 ( .A(n468), .B(n467), .Z(n729) );
  NOR2_X1 U574 ( .A1(G902), .A2(n729), .ZN(n470) );
  XNOR2_X1 U575 ( .A(KEYINPUT110), .B(G478), .ZN(n469) );
  XNOR2_X1 U576 ( .A(n470), .B(n469), .ZN(n574) );
  XNOR2_X1 U577 ( .A(G125), .B(KEYINPUT10), .ZN(n471) );
  XNOR2_X1 U578 ( .A(n471), .B(G140), .ZN(n748) );
  XNOR2_X1 U579 ( .A(n748), .B(G146), .ZN(n523) );
  XOR2_X1 U580 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n473) );
  NOR2_X1 U581 ( .A1(G953), .A2(G237), .ZN(n499) );
  NAND2_X1 U582 ( .A1(n499), .A2(G214), .ZN(n472) );
  XNOR2_X1 U583 ( .A(n473), .B(n472), .ZN(n474) );
  XOR2_X1 U584 ( .A(n474), .B(KEYINPUT105), .Z(n480) );
  XNOR2_X1 U585 ( .A(n476), .B(n475), .ZN(n478) );
  XOR2_X1 U586 ( .A(KEYINPUT106), .B(G131), .Z(n477) );
  XNOR2_X1 U587 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U588 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U589 ( .A(n523), .B(n481), .ZN(n646) );
  NAND2_X1 U590 ( .A1(n646), .A2(n525), .ZN(n485) );
  XOR2_X1 U591 ( .A(KEYINPUT108), .B(KEYINPUT13), .Z(n483) );
  XNOR2_X1 U592 ( .A(KEYINPUT107), .B(G475), .ZN(n482) );
  XOR2_X1 U593 ( .A(n483), .B(n482), .Z(n484) );
  XNOR2_X1 U594 ( .A(n485), .B(n484), .ZN(n573) );
  INV_X1 U595 ( .A(n573), .ZN(n555) );
  XOR2_X1 U596 ( .A(KEYINPUT101), .B(KEYINPUT20), .Z(n487) );
  NAND2_X1 U597 ( .A1(G234), .A2(n630), .ZN(n486) );
  XNOR2_X1 U598 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U599 ( .A(KEYINPUT100), .B(n488), .ZN(n526) );
  NAND2_X1 U600 ( .A1(n526), .A2(G221), .ZN(n490) );
  INV_X1 U601 ( .A(KEYINPUT21), .ZN(n489) );
  XNOR2_X1 U602 ( .A(n490), .B(n489), .ZN(n683) );
  INV_X1 U603 ( .A(n683), .ZN(n552) );
  INV_X1 U604 ( .A(KEYINPUT66), .ZN(n491) );
  XNOR2_X1 U605 ( .A(n491), .B(KEYINPUT22), .ZN(n492) );
  BUF_X1 U606 ( .A(n497), .Z(n498) );
  NAND2_X1 U607 ( .A1(G210), .A2(n499), .ZN(n500) );
  INV_X1 U608 ( .A(G472), .ZN(n502) );
  XNOR2_X1 U609 ( .A(n503), .B(n502), .ZN(n601) );
  INV_X1 U610 ( .A(KEYINPUT6), .ZN(n504) );
  XNOR2_X1 U611 ( .A(n601), .B(n504), .ZN(n553) );
  XOR2_X1 U612 ( .A(G104), .B(G140), .Z(n507) );
  NAND2_X1 U613 ( .A1(G227), .A2(n751), .ZN(n506) );
  XNOR2_X1 U614 ( .A(n507), .B(n506), .ZN(n509) );
  XNOR2_X1 U615 ( .A(n747), .B(n510), .ZN(n723) );
  INV_X1 U616 ( .A(G469), .ZN(n511) );
  XNOR2_X2 U617 ( .A(n512), .B(n511), .ZN(n603) );
  INV_X1 U618 ( .A(KEYINPUT1), .ZN(n513) );
  XOR2_X1 U619 ( .A(KEYINPUT23), .B(G119), .Z(n515) );
  NAND2_X1 U620 ( .A1(G221), .A2(n521), .ZN(n522) );
  XNOR2_X1 U621 ( .A(n524), .B(n523), .ZN(n634) );
  NAND2_X1 U622 ( .A1(n634), .A2(n525), .ZN(n530) );
  NAND2_X1 U623 ( .A1(n526), .A2(G217), .ZN(n528) );
  XNOR2_X1 U624 ( .A(KEYINPUT25), .B(KEYINPUT102), .ZN(n527) );
  XNOR2_X1 U625 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X2 U626 ( .A(n530), .B(n529), .ZN(n551) );
  INV_X1 U627 ( .A(n551), .ZN(n684) );
  AND2_X1 U628 ( .A1(n610), .A2(n684), .ZN(n531) );
  NAND2_X1 U629 ( .A1(n545), .A2(n531), .ZN(n578) );
  XNOR2_X1 U630 ( .A(n578), .B(G101), .ZN(G3) );
  AND2_X1 U631 ( .A1(n574), .A2(n573), .ZN(n670) );
  INV_X1 U632 ( .A(n670), .ZN(n595) );
  OR2_X1 U633 ( .A1(n533), .A2(n751), .ZN(n534) );
  NOR2_X1 U634 ( .A1(G900), .A2(n534), .ZN(n535) );
  NOR2_X1 U635 ( .A1(n536), .A2(n535), .ZN(n588) );
  NOR2_X1 U636 ( .A1(n552), .A2(n588), .ZN(n537) );
  NAND2_X1 U637 ( .A1(n537), .A2(n551), .ZN(n600) );
  NOR2_X1 U638 ( .A1(n553), .A2(n600), .ZN(n538) );
  XOR2_X1 U639 ( .A(KEYINPUT114), .B(n538), .Z(n539) );
  NOR2_X1 U640 ( .A1(n595), .A2(n539), .ZN(n540) );
  OR2_X1 U641 ( .A1(n680), .A2(n609), .ZN(n541) );
  XNOR2_X1 U642 ( .A(n541), .B(KEYINPUT43), .ZN(n543) );
  AND2_X1 U643 ( .A1(n543), .A2(n608), .ZN(n627) );
  XOR2_X1 U644 ( .A(n627), .B(G140), .Z(G42) );
  NOR2_X1 U645 ( .A1(n610), .A2(n684), .ZN(n544) );
  XOR2_X1 U646 ( .A(n550), .B(G119), .Z(G21) );
  NAND2_X1 U647 ( .A1(n546), .A2(n610), .ZN(n547) );
  XNOR2_X1 U648 ( .A(n547), .B(KEYINPUT113), .ZN(n549) );
  INV_X1 U649 ( .A(n601), .ZN(n589) );
  AND2_X1 U650 ( .A1(n601), .A2(n551), .ZN(n548) );
  NOR2_X2 U651 ( .A1(n552), .A2(n551), .ZN(n679) );
  NAND2_X1 U652 ( .A1(n680), .A2(n679), .ZN(n564) );
  NOR2_X1 U653 ( .A1(n574), .A2(n555), .ZN(n616) );
  INV_X1 U654 ( .A(KEYINPUT35), .ZN(n556) );
  XNOR2_X2 U655 ( .A(n557), .B(n556), .ZN(n757) );
  INV_X1 U656 ( .A(KEYINPUT44), .ZN(n558) );
  NAND2_X1 U657 ( .A1(n560), .A2(n559), .ZN(n562) );
  XNOR2_X1 U658 ( .A(n562), .B(n561), .ZN(n584) );
  NAND2_X1 U659 ( .A1(n563), .A2(KEYINPUT44), .ZN(n583) );
  OR2_X1 U660 ( .A1(n564), .A2(n601), .ZN(n689) );
  NOR2_X1 U661 ( .A1(n689), .A2(n565), .ZN(n568) );
  INV_X1 U662 ( .A(KEYINPUT104), .ZN(n566) );
  XNOR2_X1 U663 ( .A(n566), .B(KEYINPUT31), .ZN(n567) );
  XNOR2_X1 U664 ( .A(n568), .B(n567), .ZN(n672) );
  NAND2_X1 U665 ( .A1(n679), .A2(n603), .ZN(n570) );
  NOR2_X1 U666 ( .A1(n587), .A2(n589), .ZN(n572) );
  AND2_X1 U667 ( .A1(n571), .A2(n572), .ZN(n661) );
  OR2_X1 U668 ( .A1(n672), .A2(n661), .ZN(n577) );
  NOR2_X1 U669 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U670 ( .A(KEYINPUT111), .B(n575), .ZN(n625) );
  INV_X1 U671 ( .A(n625), .ZN(n673) );
  INV_X1 U672 ( .A(n698), .ZN(n576) );
  NAND2_X1 U673 ( .A1(n577), .A2(n576), .ZN(n579) );
  NAND2_X1 U674 ( .A1(n579), .A2(n578), .ZN(n581) );
  INV_X1 U675 ( .A(KEYINPUT112), .ZN(n580) );
  XNOR2_X1 U676 ( .A(n581), .B(n580), .ZN(n582) );
  NAND2_X1 U677 ( .A1(n584), .A2(n359), .ZN(n586) );
  INV_X1 U678 ( .A(KEYINPUT45), .ZN(n585) );
  INV_X1 U679 ( .A(KEYINPUT30), .ZN(n591) );
  NAND2_X1 U680 ( .A1(n589), .A2(n693), .ZN(n590) );
  XNOR2_X1 U681 ( .A(n591), .B(n590), .ZN(n592) );
  NAND2_X1 U682 ( .A1(n593), .A2(n592), .ZN(n618) );
  XNOR2_X1 U683 ( .A(n594), .B(KEYINPUT39), .ZN(n626) );
  NOR2_X1 U684 ( .A1(n595), .A2(n626), .ZN(n597) );
  XNOR2_X1 U685 ( .A(KEYINPUT40), .B(KEYINPUT116), .ZN(n596) );
  XNOR2_X1 U686 ( .A(n597), .B(n596), .ZN(n758) );
  INV_X1 U687 ( .A(n758), .ZN(n606) );
  INV_X1 U688 ( .A(n598), .ZN(n694) );
  XNOR2_X1 U689 ( .A(KEYINPUT28), .B(n602), .ZN(n604) );
  NAND2_X1 U690 ( .A1(n604), .A2(n603), .ZN(n612) );
  NAND2_X1 U691 ( .A1(n622), .A2(KEYINPUT47), .ZN(n613) );
  XOR2_X1 U692 ( .A(n613), .B(KEYINPUT83), .Z(n615) );
  NAND2_X1 U693 ( .A1(n698), .A2(KEYINPUT47), .ZN(n614) );
  NAND2_X1 U694 ( .A1(n615), .A2(n614), .ZN(n620) );
  OR2_X1 U695 ( .A1(n618), .A2(n617), .ZN(n619) );
  XNOR2_X1 U696 ( .A(KEYINPUT115), .B(n619), .ZN(n759) );
  INV_X1 U697 ( .A(n622), .ZN(n667) );
  NOR2_X1 U698 ( .A1(n698), .A2(KEYINPUT47), .ZN(n623) );
  XNOR2_X1 U699 ( .A(KEYINPUT76), .B(n623), .ZN(n624) );
  NOR2_X1 U700 ( .A1(n627), .A2(n356), .ZN(n628) );
  AND2_X2 U701 ( .A1(n629), .A2(n628), .ZN(n746) );
  XNOR2_X1 U702 ( .A(n630), .B(KEYINPUT87), .ZN(n631) );
  NAND2_X1 U703 ( .A1(n631), .A2(KEYINPUT2), .ZN(n632) );
  INV_X1 U704 ( .A(KEYINPUT88), .ZN(n633) );
  NAND2_X1 U705 ( .A1(n728), .A2(G217), .ZN(n635) );
  XNOR2_X1 U706 ( .A(n635), .B(n634), .ZN(n636) );
  NAND2_X1 U707 ( .A1(n636), .A2(n722), .ZN(n637) );
  XNOR2_X1 U708 ( .A(n637), .B(KEYINPUT125), .ZN(G66) );
  XOR2_X1 U709 ( .A(G110), .B(n638), .Z(G12) );
  NAND2_X1 U710 ( .A1(n728), .A2(G472), .ZN(n642) );
  XNOR2_X1 U711 ( .A(KEYINPUT92), .B(KEYINPUT62), .ZN(n639) );
  XNOR2_X1 U712 ( .A(n640), .B(n639), .ZN(n641) );
  XNOR2_X1 U713 ( .A(n642), .B(n641), .ZN(n643) );
  NAND2_X1 U714 ( .A1(n643), .A2(n722), .ZN(n644) );
  XNOR2_X1 U715 ( .A(n644), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U716 ( .A1(n728), .A2(G475), .ZN(n648) );
  XNOR2_X1 U717 ( .A(KEYINPUT67), .B(KEYINPUT59), .ZN(n645) );
  XNOR2_X1 U718 ( .A(n646), .B(n645), .ZN(n647) );
  XNOR2_X1 U719 ( .A(n648), .B(n647), .ZN(n649) );
  NAND2_X1 U720 ( .A1(n649), .A2(n722), .ZN(n651) );
  XOR2_X1 U721 ( .A(KEYINPUT68), .B(KEYINPUT60), .Z(n650) );
  XNOR2_X1 U722 ( .A(n651), .B(n650), .ZN(G60) );
  NAND2_X1 U723 ( .A1(n728), .A2(G210), .ZN(n656) );
  XNOR2_X1 U724 ( .A(KEYINPUT81), .B(KEYINPUT54), .ZN(n653) );
  XNOR2_X1 U725 ( .A(n653), .B(KEYINPUT55), .ZN(n654) );
  XNOR2_X1 U726 ( .A(n652), .B(n654), .ZN(n655) );
  XNOR2_X1 U727 ( .A(n656), .B(n655), .ZN(n657) );
  NAND2_X1 U728 ( .A1(n657), .A2(n722), .ZN(n659) );
  XNOR2_X1 U729 ( .A(KEYINPUT89), .B(KEYINPUT56), .ZN(n658) );
  XNOR2_X1 U730 ( .A(n659), .B(n658), .ZN(G51) );
  NAND2_X1 U731 ( .A1(n661), .A2(n670), .ZN(n660) );
  XNOR2_X1 U732 ( .A(n660), .B(G104), .ZN(G6) );
  XOR2_X1 U733 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n663) );
  NAND2_X1 U734 ( .A1(n661), .A2(n673), .ZN(n662) );
  XNOR2_X1 U735 ( .A(n663), .B(n662), .ZN(n664) );
  XNOR2_X1 U736 ( .A(G107), .B(n664), .ZN(G9) );
  XOR2_X1 U737 ( .A(G128), .B(KEYINPUT29), .Z(n666) );
  NAND2_X1 U738 ( .A1(n667), .A2(n673), .ZN(n665) );
  XNOR2_X1 U739 ( .A(n666), .B(n665), .ZN(G30) );
  NAND2_X1 U740 ( .A1(n667), .A2(n670), .ZN(n668) );
  XNOR2_X1 U741 ( .A(n668), .B(KEYINPUT118), .ZN(n669) );
  XNOR2_X1 U742 ( .A(G146), .B(n669), .ZN(G48) );
  NAND2_X1 U743 ( .A1(n672), .A2(n670), .ZN(n671) );
  XNOR2_X1 U744 ( .A(n671), .B(G113), .ZN(G15) );
  XOR2_X1 U745 ( .A(G116), .B(KEYINPUT119), .Z(n675) );
  NAND2_X1 U746 ( .A1(n673), .A2(n672), .ZN(n674) );
  XNOR2_X1 U747 ( .A(n675), .B(n674), .ZN(G18) );
  XNOR2_X1 U748 ( .A(G125), .B(n676), .ZN(n677) );
  XNOR2_X1 U749 ( .A(n677), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U750 ( .A(G134), .B(n356), .Z(n678) );
  XNOR2_X1 U751 ( .A(KEYINPUT120), .B(n678), .ZN(G36) );
  NOR2_X1 U752 ( .A1(n680), .A2(n679), .ZN(n681) );
  XNOR2_X1 U753 ( .A(n681), .B(KEYINPUT121), .ZN(n682) );
  XNOR2_X1 U754 ( .A(n682), .B(KEYINPUT50), .ZN(n688) );
  NOR2_X1 U755 ( .A1(n684), .A2(n683), .ZN(n685) );
  XOR2_X1 U756 ( .A(KEYINPUT49), .B(n685), .Z(n686) );
  NOR2_X1 U757 ( .A1(n589), .A2(n686), .ZN(n687) );
  NAND2_X1 U758 ( .A1(n688), .A2(n687), .ZN(n690) );
  NAND2_X1 U759 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U760 ( .A(KEYINPUT51), .B(n691), .ZN(n692) );
  NOR2_X1 U761 ( .A1(n719), .A2(n692), .ZN(n705) );
  NOR2_X1 U762 ( .A1(n694), .A2(n693), .ZN(n695) );
  NOR2_X1 U763 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U764 ( .A(n697), .B(KEYINPUT122), .ZN(n701) );
  NOR2_X1 U765 ( .A1(n699), .A2(n698), .ZN(n700) );
  NOR2_X1 U766 ( .A1(n701), .A2(n700), .ZN(n703) );
  NOR2_X1 U767 ( .A1(n703), .A2(n702), .ZN(n704) );
  NOR2_X1 U768 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U769 ( .A(n706), .B(KEYINPUT52), .ZN(n707) );
  NOR2_X1 U770 ( .A1(n708), .A2(n707), .ZN(n718) );
  INV_X1 U771 ( .A(KEYINPUT2), .ZN(n709) );
  NAND2_X1 U772 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U773 ( .A(n711), .B(KEYINPUT85), .ZN(n713) );
  NOR2_X1 U774 ( .A1(n746), .A2(KEYINPUT2), .ZN(n712) );
  XNOR2_X1 U775 ( .A(n714), .B(KEYINPUT80), .ZN(n715) );
  AND2_X1 U776 ( .A1(n716), .A2(n407), .ZN(n717) );
  NOR2_X1 U777 ( .A1(n719), .A2(n702), .ZN(n720) );
  XNOR2_X1 U778 ( .A(n720), .B(KEYINPUT123), .ZN(n721) );
  INV_X1 U779 ( .A(n722), .ZN(n733) );
  NAND2_X1 U780 ( .A1(n728), .A2(G469), .ZN(n726) );
  XOR2_X1 U781 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n724) );
  NOR2_X1 U782 ( .A1(n733), .A2(n727), .ZN(G54) );
  NAND2_X1 U783 ( .A1(n728), .A2(G478), .ZN(n731) );
  XNOR2_X1 U784 ( .A(n729), .B(KEYINPUT124), .ZN(n730) );
  XNOR2_X1 U785 ( .A(n731), .B(n730), .ZN(n732) );
  NOR2_X1 U786 ( .A1(n733), .A2(n732), .ZN(G63) );
  NAND2_X1 U787 ( .A1(n407), .A2(n734), .ZN(n739) );
  NAND2_X1 U788 ( .A1(G224), .A2(G953), .ZN(n735) );
  XNOR2_X1 U789 ( .A(n735), .B(KEYINPUT126), .ZN(n736) );
  XNOR2_X1 U790 ( .A(KEYINPUT61), .B(n736), .ZN(n737) );
  NAND2_X1 U791 ( .A1(G898), .A2(n737), .ZN(n738) );
  NAND2_X1 U792 ( .A1(n739), .A2(n738), .ZN(n745) );
  XNOR2_X1 U793 ( .A(n740), .B(n741), .ZN(n743) );
  NAND2_X1 U794 ( .A1(n743), .A2(n742), .ZN(n744) );
  XOR2_X1 U795 ( .A(n745), .B(n744), .Z(G69) );
  INV_X1 U796 ( .A(n746), .ZN(n749) );
  XOR2_X1 U797 ( .A(n748), .B(n747), .Z(n752) );
  XOR2_X1 U798 ( .A(n749), .B(n752), .Z(n750) );
  NAND2_X1 U799 ( .A1(n751), .A2(n750), .ZN(n756) );
  XOR2_X1 U800 ( .A(G227), .B(n752), .Z(n753) );
  NAND2_X1 U801 ( .A1(n753), .A2(G900), .ZN(n754) );
  NAND2_X1 U802 ( .A1(G953), .A2(n754), .ZN(n755) );
  NAND2_X1 U803 ( .A1(n756), .A2(n755), .ZN(G72) );
  XNOR2_X1 U804 ( .A(n757), .B(G122), .ZN(G24) );
  XOR2_X1 U805 ( .A(n758), .B(G131), .Z(G33) );
  XOR2_X1 U806 ( .A(G143), .B(n759), .Z(G45) );
  XNOR2_X1 U807 ( .A(G137), .B(KEYINPUT127), .ZN(n761) );
  XNOR2_X1 U808 ( .A(n761), .B(n760), .ZN(G39) );
endmodule

