//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 0 1 1 1 1 1 0 0 1 0 1 0 0 1 0 1 0 1 1 0 0 1 0 1 1 1 1 1 0 1 1 1 1 0 0 0 0 1 0 0 1 0 0 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:05 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n736, new_n737, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n760, new_n761, new_n762, new_n763, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n781, new_n782, new_n783, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  XOR2_X1   g001(.A(new_n187), .B(KEYINPUT82), .Z(new_n188));
  INV_X1    g002(.A(G143), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n189), .A2(G146), .ZN(new_n190));
  OR2_X1    g004(.A1(KEYINPUT64), .A2(G146), .ZN(new_n191));
  NAND2_X1  g005(.A1(KEYINPUT64), .A2(G146), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  AOI21_X1  g007(.A(new_n190), .B1(new_n193), .B2(new_n189), .ZN(new_n194));
  XNOR2_X1  g008(.A(KEYINPUT0), .B(G128), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n191), .A2(G143), .A3(new_n192), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n189), .A2(G146), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(KEYINPUT0), .A2(G128), .ZN(new_n199));
  OAI22_X1  g013(.A1(new_n194), .A2(new_n195), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G125), .ZN(new_n201));
  INV_X1    g015(.A(G128), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n202), .A2(KEYINPUT1), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n196), .A2(new_n197), .A3(new_n203), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n202), .B1(new_n196), .B2(KEYINPUT1), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n204), .B1(new_n205), .B2(new_n194), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n201), .B1(G125), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G224), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n208), .A2(G953), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  OAI221_X1 g024(.A(new_n201), .B1(G125), .B2(new_n206), .C1(new_n208), .C2(G953), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  XNOR2_X1  g026(.A(G110), .B(G122), .ZN(new_n213));
  AND2_X1   g027(.A1(KEYINPUT3), .A2(G107), .ZN(new_n214));
  NOR2_X1   g028(.A1(KEYINPUT3), .A2(G107), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n214), .B1(G104), .B2(new_n215), .ZN(new_n216));
  OR2_X1    g030(.A1(KEYINPUT3), .A2(G107), .ZN(new_n217));
  INV_X1    g031(.A(G104), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(KEYINPUT80), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT80), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G104), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n217), .A2(new_n219), .A3(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n216), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(G101), .ZN(new_n224));
  INV_X1    g038(.A(G101), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n216), .A2(new_n222), .A3(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n224), .A2(KEYINPUT4), .A3(new_n226), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n225), .B1(new_n216), .B2(new_n222), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT4), .ZN(new_n229));
  XOR2_X1   g043(.A(G116), .B(G119), .Z(new_n230));
  XNOR2_X1  g044(.A(KEYINPUT2), .B(G113), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  XOR2_X1   g046(.A(KEYINPUT2), .B(G113), .Z(new_n233));
  XNOR2_X1  g047(.A(G116), .B(G119), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  AOI22_X1  g049(.A1(new_n228), .A2(new_n229), .B1(new_n232), .B2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n227), .A2(new_n236), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n230), .A2(new_n231), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT5), .ZN(new_n239));
  INV_X1    g053(.A(G119), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n239), .A2(new_n240), .A3(G116), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT83), .ZN(new_n242));
  XNOR2_X1  g056(.A(new_n241), .B(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(G113), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n244), .B1(new_n234), .B2(KEYINPUT5), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n238), .B1(new_n243), .B2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(G107), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n219), .A2(new_n221), .A3(new_n247), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n225), .B1(G104), .B2(G107), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  AND2_X1   g064(.A1(new_n226), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n246), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n237), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT84), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n213), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  AOI22_X1  g069(.A1(new_n227), .A2(new_n236), .B1(new_n246), .B2(new_n251), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(KEYINPUT84), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n255), .A2(KEYINPUT6), .A3(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n256), .A2(new_n213), .ZN(new_n260));
  AOI22_X1  g074(.A1(new_n255), .A2(new_n257), .B1(KEYINPUT6), .B2(new_n260), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n212), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(G902), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n209), .A2(KEYINPUT7), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n264), .B1(new_n210), .B2(new_n211), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n207), .A2(new_n264), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT85), .ZN(new_n267));
  AND2_X1   g081(.A1(new_n243), .A2(new_n245), .ZN(new_n268));
  OAI211_X1 g082(.A(new_n267), .B(new_n251), .C1(new_n268), .C2(new_n238), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n226), .A2(new_n250), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n246), .B1(KEYINPUT85), .B2(new_n270), .ZN(new_n271));
  XNOR2_X1  g085(.A(new_n213), .B(KEYINPUT8), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n269), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n260), .A2(new_n266), .A3(new_n273), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n263), .B1(new_n265), .B2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  OAI21_X1  g090(.A(G210), .B1(G237), .B2(G902), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n262), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n277), .ZN(new_n279));
  INV_X1    g093(.A(new_n212), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n260), .A2(KEYINPUT6), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n253), .A2(new_n254), .ZN(new_n282));
  INV_X1    g096(.A(new_n213), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n283), .B1(new_n256), .B2(KEYINPUT84), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n281), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n280), .B1(new_n285), .B2(new_n258), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n279), .B1(new_n286), .B2(new_n275), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n188), .B1(new_n278), .B2(new_n287), .ZN(new_n288));
  XNOR2_X1  g102(.A(KEYINPUT22), .B(G137), .ZN(new_n289));
  INV_X1    g103(.A(G953), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n290), .A2(G221), .A3(G234), .ZN(new_n291));
  XNOR2_X1  g105(.A(new_n289), .B(new_n291), .ZN(new_n292));
  XOR2_X1   g106(.A(G119), .B(G128), .Z(new_n293));
  XNOR2_X1  g107(.A(KEYINPUT24), .B(G110), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT23), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n296), .B1(new_n240), .B2(G128), .ZN(new_n297));
  OAI21_X1  g111(.A(KEYINPUT74), .B1(new_n240), .B2(G128), .ZN(new_n298));
  XNOR2_X1  g112(.A(new_n297), .B(new_n298), .ZN(new_n299));
  XNOR2_X1  g113(.A(KEYINPUT77), .B(G110), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n295), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(new_n193), .ZN(new_n302));
  XNOR2_X1  g116(.A(G125), .B(G140), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(G125), .ZN(new_n305));
  NOR3_X1   g119(.A1(new_n305), .A2(KEYINPUT16), .A3(G140), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT75), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  AOI21_X1  g122(.A(KEYINPUT75), .B1(new_n303), .B2(KEYINPUT16), .ZN(new_n309));
  OAI211_X1 g123(.A(G146), .B(new_n308), .C1(new_n309), .C2(new_n306), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n301), .A2(new_n304), .A3(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(G146), .ZN(new_n313));
  INV_X1    g127(.A(G140), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(G125), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n305), .A2(G140), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n315), .A2(new_n316), .A3(KEYINPUT16), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n306), .B1(new_n317), .B2(new_n307), .ZN(new_n318));
  INV_X1    g132(.A(new_n308), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n313), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(new_n310), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n293), .A2(new_n294), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n322), .B1(new_n299), .B2(G110), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT76), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n321), .A2(KEYINPUT76), .A3(new_n323), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n312), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT78), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n292), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  AND3_X1   g144(.A1(new_n321), .A2(KEYINPUT76), .A3(new_n323), .ZN(new_n331));
  AOI21_X1  g145(.A(KEYINPUT76), .B1(new_n321), .B2(new_n323), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n311), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(KEYINPUT78), .ZN(new_n334));
  OAI211_X1 g148(.A(new_n329), .B(new_n311), .C1(new_n331), .C2(new_n332), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n330), .B1(new_n336), .B2(new_n292), .ZN(new_n337));
  XOR2_X1   g151(.A(KEYINPUT73), .B(G217), .Z(new_n338));
  XOR2_X1   g152(.A(KEYINPUT72), .B(G902), .Z(new_n339));
  AOI21_X1  g153(.A(new_n338), .B1(G234), .B2(new_n339), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n340), .A2(G902), .ZN(new_n341));
  AND2_X1   g155(.A1(new_n337), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n326), .A2(new_n327), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n329), .B1(new_n343), .B2(new_n311), .ZN(new_n344));
  INV_X1    g158(.A(new_n335), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n292), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(new_n330), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n346), .A2(new_n339), .A3(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT25), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n337), .A2(KEYINPUT25), .A3(new_n339), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n342), .B1(new_n352), .B2(new_n340), .ZN(new_n353));
  OR2_X1    g167(.A1(new_n251), .A2(new_n206), .ZN(new_n354));
  INV_X1    g168(.A(new_n204), .ZN(new_n355));
  OAI21_X1  g169(.A(KEYINPUT1), .B1(new_n189), .B2(G146), .ZN(new_n356));
  AOI22_X1  g170(.A1(new_n196), .A2(new_n197), .B1(G128), .B2(new_n356), .ZN(new_n357));
  OAI211_X1 g171(.A(new_n226), .B(new_n250), .C1(new_n355), .C2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n354), .A2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT65), .ZN(new_n360));
  INV_X1    g174(.A(G134), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(KEYINPUT65), .A2(G134), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n362), .A2(G137), .A3(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(G137), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n365), .A2(KEYINPUT11), .A3(G134), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  AND2_X1   g182(.A1(KEYINPUT65), .A2(G134), .ZN(new_n369));
  NOR2_X1   g183(.A1(KEYINPUT65), .A2(G134), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n365), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT11), .ZN(new_n372));
  AND3_X1   g186(.A1(new_n371), .A2(KEYINPUT66), .A3(new_n372), .ZN(new_n373));
  AOI21_X1  g187(.A(KEYINPUT66), .B1(new_n371), .B2(new_n372), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n368), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(G131), .ZN(new_n376));
  INV_X1    g190(.A(G131), .ZN(new_n377));
  OAI211_X1 g191(.A(new_n377), .B(new_n368), .C1(new_n373), .C2(new_n374), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n359), .A2(KEYINPUT12), .A3(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT67), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT66), .ZN(new_n382));
  AOI21_X1  g196(.A(G137), .B1(new_n362), .B2(new_n363), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n382), .B1(new_n383), .B2(KEYINPUT11), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n371), .A2(KEYINPUT66), .A3(new_n372), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n377), .B1(new_n386), .B2(new_n368), .ZN(new_n387));
  AOI211_X1 g201(.A(G131), .B(new_n367), .C1(new_n384), .C2(new_n385), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n381), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n376), .A2(KEYINPUT67), .A3(new_n378), .ZN(new_n390));
  AOI22_X1  g204(.A1(new_n389), .A2(new_n390), .B1(new_n358), .B2(new_n354), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n380), .B1(new_n391), .B2(KEYINPUT12), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT10), .ZN(new_n393));
  AND3_X1   g207(.A1(new_n226), .A2(KEYINPUT10), .A3(new_n250), .ZN(new_n394));
  AOI22_X1  g208(.A1(new_n358), .A2(new_n393), .B1(new_n394), .B2(new_n206), .ZN(new_n395));
  INV_X1    g209(.A(new_n200), .ZN(new_n396));
  OAI211_X1 g210(.A(new_n396), .B(new_n227), .C1(KEYINPUT4), .C2(new_n224), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n389), .A2(new_n390), .A3(new_n395), .A4(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n392), .A2(new_n398), .ZN(new_n399));
  XNOR2_X1  g213(.A(G110), .B(G140), .ZN(new_n400));
  INV_X1    g214(.A(G227), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n401), .A2(G953), .ZN(new_n402));
  XNOR2_X1  g216(.A(new_n400), .B(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  AND2_X1   g218(.A1(new_n398), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n389), .A2(new_n390), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n395), .A2(new_n397), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  AOI22_X1  g222(.A1(new_n399), .A2(new_n403), .B1(new_n405), .B2(new_n408), .ZN(new_n409));
  OAI21_X1  g223(.A(G469), .B1(new_n409), .B2(G902), .ZN(new_n410));
  INV_X1    g224(.A(new_n339), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n392), .A2(new_n405), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n408), .A2(new_n398), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(new_n403), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n411), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(G469), .ZN(new_n416));
  AOI21_X1  g230(.A(KEYINPUT81), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  AOI22_X1  g231(.A1(new_n392), .A2(new_n405), .B1(new_n413), .B2(new_n403), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT81), .ZN(new_n419));
  NOR4_X1   g233(.A1(new_n418), .A2(new_n419), .A3(G469), .A4(new_n411), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n410), .B1(new_n417), .B2(new_n420), .ZN(new_n421));
  XNOR2_X1  g235(.A(KEYINPUT9), .B(G234), .ZN(new_n422));
  OAI21_X1  g236(.A(G221), .B1(new_n422), .B2(G902), .ZN(new_n423));
  XOR2_X1   g237(.A(new_n423), .B(KEYINPUT79), .Z(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  AND4_X1   g239(.A1(new_n288), .A2(new_n353), .A3(new_n421), .A4(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(G475), .ZN(new_n427));
  NOR2_X1   g241(.A1(G237), .A2(G953), .ZN(new_n428));
  AND3_X1   g242(.A1(new_n428), .A2(G143), .A3(G214), .ZN(new_n429));
  AOI21_X1  g243(.A(G143), .B1(new_n428), .B2(G214), .ZN(new_n430));
  OAI21_X1  g244(.A(G131), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT87), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(G237), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n434), .A2(new_n290), .A3(G214), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(new_n189), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n428), .A2(G143), .A3(G214), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n438), .A2(KEYINPUT87), .A3(G131), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n433), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(KEYINPUT17), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT17), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n436), .A2(new_n377), .A3(new_n437), .ZN(new_n443));
  NAND4_X1  g257(.A1(new_n433), .A2(new_n439), .A3(new_n442), .A4(new_n443), .ZN(new_n444));
  NAND4_X1  g258(.A1(new_n441), .A2(new_n444), .A3(new_n320), .A4(new_n310), .ZN(new_n445));
  NAND2_X1  g259(.A1(KEYINPUT18), .A2(G131), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  OAI21_X1  g261(.A(KEYINPUT86), .B1(new_n438), .B2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT86), .ZN(new_n449));
  NAND4_X1  g263(.A1(new_n436), .A2(new_n449), .A3(new_n437), .A4(new_n446), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n315), .A2(new_n316), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(G146), .ZN(new_n453));
  AOI22_X1  g267(.A1(new_n304), .A2(new_n453), .B1(new_n438), .B2(new_n447), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n451), .A2(new_n454), .ZN(new_n455));
  XNOR2_X1  g269(.A(G113), .B(G122), .ZN(new_n456));
  XNOR2_X1  g270(.A(KEYINPUT89), .B(G104), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n456), .B(new_n457), .ZN(new_n458));
  XNOR2_X1  g272(.A(new_n458), .B(KEYINPUT90), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n445), .A2(new_n455), .A3(new_n459), .ZN(new_n460));
  AND2_X1   g274(.A1(new_n451), .A2(new_n454), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n442), .B1(new_n433), .B2(new_n439), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n462), .A2(new_n321), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n461), .B1(new_n463), .B2(new_n444), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n460), .B1(new_n464), .B2(new_n458), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n427), .B1(new_n465), .B2(new_n263), .ZN(new_n466));
  AND3_X1   g280(.A1(new_n433), .A2(new_n439), .A3(new_n443), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT19), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n452), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n303), .A2(KEYINPUT19), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n193), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(new_n310), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n455), .B1(new_n467), .B2(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n458), .B1(new_n474), .B2(KEYINPUT88), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n318), .A2(new_n319), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n471), .B1(new_n476), .B2(G146), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n433), .A2(new_n439), .A3(new_n443), .ZN(new_n478));
  AOI22_X1  g292(.A1(new_n477), .A2(new_n478), .B1(new_n451), .B2(new_n454), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT88), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  AOI22_X1  g295(.A1(new_n475), .A2(new_n481), .B1(new_n464), .B2(new_n459), .ZN(new_n482));
  NOR2_X1   g296(.A1(G475), .A2(G902), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(KEYINPUT20), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n458), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n486), .B1(new_n479), .B2(new_n480), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n474), .A2(KEYINPUT88), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n460), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT20), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n489), .A2(new_n490), .A3(new_n483), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n466), .B1(new_n485), .B2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(G478), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n493), .A2(KEYINPUT15), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  XNOR2_X1  g309(.A(G116), .B(G122), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(new_n247), .ZN(new_n497));
  XNOR2_X1  g311(.A(new_n497), .B(KEYINPUT92), .ZN(new_n498));
  XOR2_X1   g312(.A(G128), .B(G143), .Z(new_n499));
  NAND2_X1  g313(.A1(new_n362), .A2(new_n363), .ZN(new_n500));
  XNOR2_X1  g314(.A(new_n499), .B(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(G116), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n502), .A2(KEYINPUT14), .A3(G122), .ZN(new_n503));
  INV_X1    g317(.A(new_n496), .ZN(new_n504));
  OAI211_X1 g318(.A(G107), .B(new_n503), .C1(new_n504), .C2(KEYINPUT14), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n498), .A2(new_n501), .A3(new_n505), .ZN(new_n506));
  XNOR2_X1  g320(.A(KEYINPUT91), .B(KEYINPUT13), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n507), .A2(G128), .A3(new_n189), .ZN(new_n508));
  OAI211_X1 g322(.A(new_n508), .B(G134), .C1(new_n499), .C2(new_n507), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n496), .B(new_n247), .ZN(new_n510));
  OAI211_X1 g324(.A(new_n509), .B(new_n510), .C1(new_n499), .C2(new_n500), .ZN(new_n511));
  NOR3_X1   g325(.A1(new_n338), .A2(G953), .A3(new_n422), .ZN(new_n512));
  AND3_X1   g326(.A1(new_n506), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n512), .B1(new_n506), .B2(new_n511), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n495), .B1(new_n516), .B2(new_n339), .ZN(new_n517));
  OAI211_X1 g331(.A(new_n339), .B(new_n495), .C1(new_n513), .C2(new_n514), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n492), .A2(new_n520), .ZN(new_n521));
  OR2_X1    g335(.A1(KEYINPUT93), .A2(G952), .ZN(new_n522));
  NAND2_X1  g336(.A1(KEYINPUT93), .A2(G952), .ZN(new_n523));
  AOI21_X1  g337(.A(G953), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(G234), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n524), .B1(new_n525), .B2(new_n434), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  AOI211_X1 g341(.A(new_n290), .B(new_n339), .C1(G234), .C2(G237), .ZN(new_n528));
  XNOR2_X1  g342(.A(KEYINPUT21), .B(G898), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n521), .A2(new_n530), .ZN(new_n531));
  NOR3_X1   g345(.A1(new_n387), .A2(new_n388), .A3(new_n381), .ZN(new_n532));
  AOI21_X1  g346(.A(KEYINPUT67), .B1(new_n376), .B2(new_n378), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n396), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n365), .A2(G134), .ZN(new_n535));
  OAI21_X1  g349(.A(G131), .B1(new_n383), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n378), .A2(new_n536), .A3(new_n206), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n232), .A2(new_n235), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(KEYINPUT28), .B1(new_n534), .B2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n428), .A2(G210), .ZN(new_n544));
  XOR2_X1   g358(.A(new_n544), .B(KEYINPUT27), .Z(new_n545));
  XNOR2_X1  g359(.A(KEYINPUT26), .B(G101), .ZN(new_n546));
  XNOR2_X1  g360(.A(new_n545), .B(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT29), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n540), .B1(new_n406), .B2(new_n396), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n534), .A2(new_n537), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n550), .B1(new_n551), .B2(new_n538), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT28), .ZN(new_n553));
  OAI211_X1 g367(.A(new_n543), .B(new_n549), .C1(new_n552), .C2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT71), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n200), .B1(new_n389), .B2(new_n390), .ZN(new_n557));
  INV_X1    g371(.A(new_n537), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n538), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n534), .A2(new_n541), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(KEYINPUT28), .ZN(new_n562));
  NAND4_X1  g376(.A1(new_n562), .A2(KEYINPUT71), .A3(new_n543), .A4(new_n549), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n556), .A2(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n200), .B1(new_n376), .B2(new_n378), .ZN(new_n565));
  OAI211_X1 g379(.A(KEYINPUT70), .B(new_n538), .C1(new_n565), .C2(new_n558), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n538), .B1(new_n565), .B2(new_n558), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT70), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n560), .A2(new_n566), .A3(new_n569), .ZN(new_n570));
  AOI211_X1 g384(.A(new_n547), .B(new_n542), .C1(new_n570), .C2(KEYINPUT28), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n534), .A2(KEYINPUT30), .A3(new_n537), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n379), .A2(new_n396), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(new_n537), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT30), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n539), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n550), .B1(new_n572), .B2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(new_n547), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n548), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n339), .B1(new_n571), .B2(new_n579), .ZN(new_n580));
  OAI21_X1  g394(.A(G472), .B1(new_n564), .B2(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n547), .B1(new_n534), .B2(new_n541), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n575), .B1(new_n565), .B2(new_n558), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n537), .A2(KEYINPUT30), .ZN(new_n584));
  OAI211_X1 g398(.A(new_n538), .B(new_n583), .C1(new_n557), .C2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT31), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n582), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n542), .B1(new_n570), .B2(KEYINPUT28), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n587), .B1(new_n588), .B2(new_n578), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n582), .A2(new_n585), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(KEYINPUT68), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT68), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n582), .A2(new_n585), .A3(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n591), .A2(KEYINPUT31), .A3(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT69), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n591), .A2(KEYINPUT69), .A3(KEYINPUT31), .A4(new_n593), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n589), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NOR2_X1   g412(.A1(G472), .A2(G902), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT32), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n581), .B1(new_n598), .B2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n589), .ZN(new_n605));
  AND3_X1   g419(.A1(new_n582), .A2(new_n585), .A3(new_n592), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n592), .B1(new_n582), .B2(new_n585), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  AOI21_X1  g422(.A(KEYINPUT69), .B1(new_n608), .B2(KEYINPUT31), .ZN(new_n609));
  INV_X1    g423(.A(new_n597), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n605), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  AOI21_X1  g425(.A(KEYINPUT32), .B1(new_n611), .B2(new_n599), .ZN(new_n612));
  OAI211_X1 g426(.A(new_n426), .B(new_n531), .C1(new_n604), .C2(new_n612), .ZN(new_n613));
  XNOR2_X1  g427(.A(KEYINPUT94), .B(G101), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n613), .B(new_n614), .ZN(G3));
  NAND2_X1  g429(.A1(new_n421), .A2(new_n425), .ZN(new_n616));
  INV_X1    g430(.A(new_n353), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n611), .A2(new_n599), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n516), .A2(new_n339), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(new_n493), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(KEYINPUT96), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT96), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n620), .A2(new_n623), .A3(new_n493), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT33), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n625), .A2(KEYINPUT95), .ZN(new_n626));
  OR2_X1    g440(.A1(new_n625), .A2(KEYINPUT95), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n516), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n515), .A2(KEYINPUT95), .A3(new_n625), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n411), .A2(new_n493), .ZN(new_n631));
  AOI22_X1  g445(.A1(new_n622), .A2(new_n624), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n465), .A2(new_n263), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(G475), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n474), .A2(KEYINPUT88), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n636), .A2(new_n481), .A3(new_n486), .ZN(new_n637));
  AOI211_X1 g451(.A(KEYINPUT20), .B(new_n484), .C1(new_n637), .C2(new_n460), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n490), .B1(new_n489), .B2(new_n483), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n635), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n633), .A2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n530), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n288), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  OAI21_X1  g458(.A(G472), .B1(new_n598), .B2(new_n411), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n618), .A2(new_n619), .A3(new_n644), .A4(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(G104), .ZN(new_n647));
  XNOR2_X1  g461(.A(KEYINPUT97), .B(KEYINPUT34), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G6));
  INV_X1    g463(.A(new_n520), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n492), .A2(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n643), .A2(new_n651), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n618), .A2(new_n619), .A3(new_n645), .A4(new_n652), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT35), .B(G107), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G9));
  NAND2_X1  g469(.A1(new_n398), .A2(new_n404), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n359), .B1(new_n532), .B2(new_n533), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT12), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n656), .B1(new_n659), .B2(new_n380), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n404), .B1(new_n408), .B2(new_n398), .ZN(new_n661));
  OAI211_X1 g475(.A(new_n416), .B(new_n339), .C1(new_n660), .C2(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(new_n419), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n415), .A2(KEYINPUT81), .A3(new_n416), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n424), .B1(new_n665), .B2(new_n410), .ZN(new_n666));
  INV_X1    g480(.A(new_n188), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n277), .B1(new_n262), .B2(new_n276), .ZN(new_n668));
  NOR3_X1   g482(.A1(new_n286), .A2(new_n279), .A3(new_n275), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n667), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  AOI21_X1  g484(.A(KEYINPUT25), .B1(new_n337), .B2(new_n339), .ZN(new_n671));
  INV_X1    g485(.A(new_n292), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n672), .B1(new_n334), .B2(new_n335), .ZN(new_n673));
  NOR4_X1   g487(.A1(new_n673), .A2(new_n330), .A3(new_n349), .A4(new_n411), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n340), .B1(new_n671), .B2(new_n674), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n672), .A2(KEYINPUT36), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n333), .B(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(new_n341), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n670), .B1(new_n675), .B2(new_n678), .ZN(new_n679));
  AND2_X1   g493(.A1(new_n666), .A2(new_n679), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n680), .A2(new_n531), .A3(new_n619), .A4(new_n645), .ZN(new_n681));
  XOR2_X1   g495(.A(KEYINPUT37), .B(G110), .Z(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G12));
  INV_X1    g497(.A(new_n528), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n526), .B1(new_n684), .B2(G900), .ZN(new_n685));
  XOR2_X1   g499(.A(new_n685), .B(KEYINPUT98), .Z(new_n686));
  NOR2_X1   g500(.A1(new_n651), .A2(new_n686), .ZN(new_n687));
  AND3_X1   g501(.A1(new_n666), .A2(new_n679), .A3(new_n687), .ZN(new_n688));
  OAI21_X1  g502(.A(new_n688), .B1(new_n612), .B2(new_n604), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G128), .ZN(G30));
  XOR2_X1   g504(.A(new_n686), .B(KEYINPUT39), .Z(new_n691));
  NAND2_X1  g505(.A1(new_n666), .A2(new_n691), .ZN(new_n692));
  XOR2_X1   g506(.A(new_n692), .B(KEYINPUT40), .Z(new_n693));
  NAND2_X1  g507(.A1(new_n675), .A2(new_n678), .ZN(new_n694));
  NOR4_X1   g508(.A1(new_n694), .A2(new_n520), .A3(new_n492), .A4(new_n188), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(KEYINPUT100), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n601), .B1(new_n598), .B2(new_n600), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n611), .A2(new_n602), .ZN(new_n698));
  AOI211_X1 g512(.A(new_n607), .B(new_n606), .C1(new_n547), .C2(new_n561), .ZN(new_n699));
  OAI21_X1  g513(.A(G472), .B1(new_n699), .B2(G902), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n697), .A2(new_n698), .A3(new_n700), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n668), .A2(new_n669), .ZN(new_n702));
  XNOR2_X1  g516(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n702), .B(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n693), .A2(new_n696), .A3(new_n701), .A4(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G143), .ZN(G45));
  NOR3_X1   g521(.A1(new_n632), .A2(new_n492), .A3(new_n686), .ZN(new_n708));
  AND3_X1   g522(.A1(new_n666), .A2(new_n679), .A3(new_n708), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n709), .B1(new_n612), .B2(new_n604), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(KEYINPUT101), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n697), .A2(new_n698), .A3(new_n581), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT101), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n712), .A2(new_n713), .A3(new_n709), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n711), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G146), .ZN(G48));
  NOR2_X1   g530(.A1(new_n415), .A2(new_n416), .ZN(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n665), .A2(new_n425), .A3(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(new_n719), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n712), .A2(new_n720), .A3(new_n353), .A4(new_n644), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT102), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n588), .A2(new_n578), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n585), .A2(new_n560), .ZN(new_n725));
  AOI21_X1  g539(.A(KEYINPUT29), .B1(new_n725), .B2(new_n547), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n411), .B1(new_n724), .B2(new_n726), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n727), .A2(new_n556), .A3(new_n563), .ZN(new_n728));
  AOI22_X1  g542(.A1(new_n611), .A2(new_n602), .B1(new_n728), .B2(G472), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n617), .B1(new_n729), .B2(new_n697), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n730), .A2(KEYINPUT102), .A3(new_n644), .A4(new_n720), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n723), .A2(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(KEYINPUT41), .B(G113), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n732), .B(new_n733), .ZN(G15));
  NAND4_X1  g548(.A1(new_n712), .A2(new_n720), .A3(new_n353), .A4(new_n652), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT103), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n730), .A2(KEYINPUT103), .A3(new_n652), .A4(new_n720), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G116), .ZN(G18));
  NAND4_X1  g554(.A1(new_n665), .A2(new_n288), .A3(new_n425), .A4(new_n718), .ZN(new_n741));
  AOI22_X1  g555(.A1(new_n352), .A2(new_n340), .B1(new_n341), .B2(new_n677), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  OAI211_X1 g557(.A(new_n531), .B(new_n743), .C1(new_n604), .C2(new_n612), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G119), .ZN(G21));
  NAND4_X1  g559(.A1(new_n665), .A2(new_n642), .A3(new_n425), .A4(new_n718), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT104), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n747), .B1(new_n492), .B2(new_n520), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n640), .A2(KEYINPUT104), .A3(new_n650), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n748), .A2(new_n749), .A3(new_n288), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(KEYINPUT105), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT105), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n748), .A2(new_n749), .A3(new_n288), .A4(new_n752), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n746), .B1(new_n751), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n594), .A2(new_n587), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n578), .B1(new_n562), .B2(new_n543), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n599), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n754), .A2(new_n353), .A3(new_n645), .A4(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G122), .ZN(G24));
  INV_X1    g573(.A(new_n686), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n633), .A2(new_n640), .A3(new_n760), .ZN(new_n761));
  NOR3_X1   g575(.A1(new_n741), .A2(new_n742), .A3(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n762), .A2(new_n645), .A3(new_n757), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G125), .ZN(G27));
  NOR2_X1   g578(.A1(new_n598), .A2(new_n603), .ZN(new_n765));
  OAI21_X1  g579(.A(KEYINPUT106), .B1(new_n612), .B2(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT106), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n697), .A2(new_n767), .A3(new_n698), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n766), .A2(new_n581), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n702), .A2(new_n667), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n616), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(new_n708), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT42), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n769), .A2(new_n353), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n712), .A2(new_n353), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n773), .B1(new_n776), .B2(new_n772), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  XOR2_X1   g592(.A(KEYINPUT107), .B(G131), .Z(new_n779));
  XNOR2_X1  g593(.A(new_n778), .B(new_n779), .ZN(G33));
  AND2_X1   g594(.A1(new_n712), .A2(new_n771), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n781), .A2(new_n353), .A3(new_n687), .ZN(new_n782));
  XOR2_X1   g596(.A(KEYINPUT108), .B(G134), .Z(new_n783));
  XNOR2_X1  g597(.A(new_n782), .B(new_n783), .ZN(G36));
  INV_X1    g598(.A(KEYINPUT110), .ZN(new_n785));
  AND2_X1   g599(.A1(new_n409), .A2(KEYINPUT45), .ZN(new_n786));
  OR2_X1    g600(.A1(new_n409), .A2(KEYINPUT45), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n787), .A2(G469), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n786), .B1(new_n788), .B2(KEYINPUT109), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT109), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n787), .A2(new_n790), .A3(G469), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(G469), .A2(G902), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT46), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n785), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  AOI22_X1  g610(.A1(new_n789), .A2(new_n791), .B1(G469), .B2(G902), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n797), .A2(KEYINPUT110), .A3(KEYINPUT46), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(new_n665), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n800), .B1(new_n794), .B2(new_n795), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n424), .B1(new_n799), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n802), .A2(new_n691), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n645), .A2(new_n619), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n633), .A2(new_n492), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n805), .A2(KEYINPUT43), .ZN(new_n806));
  OR2_X1    g620(.A1(new_n805), .A2(KEYINPUT43), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n804), .A2(new_n694), .A3(new_n806), .A4(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT44), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n770), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n810), .B1(new_n809), .B2(new_n808), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n803), .A2(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(new_n365), .ZN(G39));
  AND3_X1   g627(.A1(new_n797), .A2(KEYINPUT110), .A3(KEYINPUT46), .ZN(new_n814));
  AOI21_X1  g628(.A(KEYINPUT110), .B1(new_n797), .B2(KEYINPUT46), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n801), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  XOR2_X1   g630(.A(KEYINPUT111), .B(KEYINPUT47), .Z(new_n817));
  INV_X1    g631(.A(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n816), .A2(new_n425), .A3(new_n818), .ZN(new_n819));
  NOR2_X1   g633(.A1(KEYINPUT111), .A2(KEYINPUT47), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n819), .B1(new_n802), .B2(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(new_n770), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n617), .A2(new_n708), .A3(new_n822), .ZN(new_n823));
  OR3_X1    g637(.A1(new_n821), .A2(new_n712), .A3(new_n823), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n824), .B(G140), .ZN(G42));
  INV_X1    g639(.A(KEYINPUT113), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n697), .A2(new_n698), .A3(new_n700), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n751), .A2(new_n753), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n694), .A2(new_n686), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n828), .A2(new_n666), .A3(new_n829), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n826), .B1(new_n827), .B2(new_n830), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n616), .A2(new_n694), .A3(new_n686), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n701), .A2(KEYINPUT113), .A3(new_n832), .A4(new_n828), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  AND2_X1   g648(.A1(new_n645), .A2(new_n757), .ZN(new_n835));
  AOI22_X1  g649(.A1(new_n835), .A2(new_n762), .B1(new_n712), .B2(new_n688), .ZN(new_n836));
  AND3_X1   g650(.A1(new_n712), .A2(new_n713), .A3(new_n709), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n713), .B1(new_n712), .B2(new_n709), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n836), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  OAI21_X1  g653(.A(KEYINPUT52), .B1(new_n834), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n689), .A2(new_n763), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n841), .B1(new_n714), .B2(new_n711), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT52), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n831), .A2(new_n833), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n842), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n840), .A2(new_n845), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n758), .A2(new_n744), .A3(new_n653), .A4(new_n681), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT112), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n848), .B1(new_n613), .B2(new_n646), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n613), .A2(new_n646), .A3(new_n848), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n850), .A2(new_n732), .A3(new_n739), .A4(new_n851), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n742), .A2(new_n521), .A3(new_n686), .ZN(new_n853));
  INV_X1    g667(.A(new_n772), .ZN(new_n854));
  AND3_X1   g668(.A1(new_n645), .A2(new_n694), .A3(new_n757), .ZN(new_n855));
  AOI22_X1  g669(.A1(new_n781), .A2(new_n853), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n778), .A2(new_n782), .A3(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT53), .ZN(new_n858));
  NOR4_X1   g672(.A1(new_n846), .A2(new_n852), .A3(new_n857), .A4(new_n858), .ZN(new_n859));
  AND4_X1   g673(.A1(new_n843), .A2(new_n844), .A3(new_n715), .A4(new_n836), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n843), .B1(new_n842), .B2(new_n844), .ZN(new_n861));
  OAI21_X1  g675(.A(KEYINPUT114), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n852), .A2(new_n857), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT114), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n840), .A2(new_n864), .A3(new_n845), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n862), .A2(new_n863), .A3(new_n865), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n859), .B1(new_n858), .B2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT54), .ZN(new_n868));
  OAI21_X1  g682(.A(KEYINPUT115), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n866), .A2(new_n858), .ZN(new_n870));
  INV_X1    g684(.A(new_n846), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n871), .A2(new_n863), .A3(KEYINPUT53), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT115), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n873), .A2(new_n874), .A3(KEYINPUT54), .ZN(new_n875));
  OR2_X1    g689(.A1(new_n866), .A2(new_n858), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n871), .A2(new_n863), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n877), .A2(new_n858), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n876), .A2(new_n868), .A3(new_n878), .ZN(new_n879));
  AND3_X1   g693(.A1(new_n807), .A2(new_n527), .A3(new_n806), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n880), .A2(new_n353), .A3(new_n835), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n524), .B1(new_n881), .B2(new_n741), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n827), .A2(new_n353), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n719), .A2(new_n770), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n884), .A2(new_n527), .ZN(new_n885));
  NOR3_X1   g699(.A1(new_n883), .A2(new_n641), .A3(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT120), .ZN(new_n887));
  OR3_X1    g701(.A1(new_n882), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n887), .B1(new_n882), .B2(new_n886), .ZN(new_n889));
  AND2_X1   g703(.A1(new_n880), .A2(new_n884), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n890), .A2(new_n353), .A3(new_n769), .ZN(new_n891));
  OR2_X1    g705(.A1(new_n891), .A2(KEYINPUT48), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n891), .A2(KEYINPUT48), .ZN(new_n893));
  AOI22_X1  g707(.A1(new_n888), .A2(new_n889), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  OR4_X1    g708(.A1(new_n640), .A2(new_n883), .A3(new_n633), .A4(new_n885), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n890), .A2(new_n855), .ZN(new_n896));
  AND2_X1   g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT118), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n898), .B1(new_n720), .B2(new_n188), .ZN(new_n899));
  NOR3_X1   g713(.A1(new_n719), .A2(KEYINPUT118), .A3(new_n667), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n899), .A2(new_n705), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n881), .B1(new_n901), .B2(KEYINPUT119), .ZN(new_n902));
  OR2_X1    g716(.A1(new_n901), .A2(KEYINPUT119), .ZN(new_n903));
  AOI21_X1  g717(.A(KEYINPUT50), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  AND3_X1   g718(.A1(new_n902), .A2(KEYINPUT50), .A3(new_n903), .ZN(new_n905));
  OAI211_X1 g719(.A(new_n897), .B(KEYINPUT51), .C1(new_n904), .C2(new_n905), .ZN(new_n906));
  OR2_X1    g720(.A1(new_n881), .A2(new_n770), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n800), .A2(new_n717), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(new_n424), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n907), .B1(new_n821), .B2(new_n909), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n894), .B1(new_n906), .B2(new_n910), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n905), .A2(new_n904), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n895), .A2(new_n896), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT117), .ZN(new_n915));
  AND3_X1   g729(.A1(new_n816), .A2(new_n425), .A3(new_n818), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n820), .B1(new_n816), .B2(new_n425), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n915), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  OAI211_X1 g732(.A(new_n819), .B(KEYINPUT117), .C1(new_n802), .C2(new_n820), .ZN(new_n919));
  AND3_X1   g733(.A1(new_n918), .A2(new_n919), .A3(new_n909), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n914), .B1(new_n920), .B2(new_n907), .ZN(new_n921));
  XOR2_X1   g735(.A(KEYINPUT116), .B(KEYINPUT51), .Z(new_n922));
  AOI21_X1  g736(.A(new_n911), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n869), .A2(new_n875), .A3(new_n879), .A4(new_n923), .ZN(new_n924));
  OR2_X1    g738(.A1(G952), .A2(G953), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NOR3_X1   g740(.A1(new_n800), .A2(KEYINPUT49), .A3(new_n717), .ZN(new_n927));
  NOR3_X1   g741(.A1(new_n805), .A2(new_n188), .A3(new_n424), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT49), .ZN(new_n929));
  OAI211_X1 g743(.A(new_n928), .B(new_n704), .C1(new_n929), .C2(new_n908), .ZN(new_n930));
  OR3_X1    g744(.A1(new_n883), .A2(new_n927), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n926), .A2(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT121), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n926), .A2(KEYINPUT121), .A3(new_n931), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n934), .A2(new_n935), .ZN(G75));
  NOR2_X1   g750(.A1(new_n290), .A2(G952), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n339), .B1(new_n876), .B2(new_n878), .ZN(new_n938));
  AOI21_X1  g752(.A(KEYINPUT56), .B1(new_n938), .B2(new_n279), .ZN(new_n939));
  NOR3_X1   g753(.A1(new_n259), .A2(new_n261), .A3(new_n212), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n940), .A2(new_n286), .ZN(new_n941));
  XNOR2_X1  g755(.A(KEYINPUT122), .B(KEYINPUT55), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n941), .B(new_n942), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n939), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n938), .A2(new_n279), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT56), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n945), .A2(new_n946), .A3(new_n943), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT123), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n939), .A2(KEYINPUT123), .A3(new_n943), .ZN(new_n950));
  AOI211_X1 g764(.A(new_n937), .B(new_n944), .C1(new_n949), .C2(new_n950), .ZN(G51));
  NAND2_X1  g765(.A1(new_n876), .A2(new_n878), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n952), .A2(KEYINPUT54), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n953), .A2(new_n879), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n793), .B(KEYINPUT57), .Z(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n956), .B1(new_n660), .B2(new_n661), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n938), .A2(new_n791), .A3(new_n789), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n937), .B1(new_n957), .B2(new_n958), .ZN(G54));
  AND3_X1   g773(.A1(new_n938), .A2(KEYINPUT58), .A3(G475), .ZN(new_n960));
  AND2_X1   g774(.A1(new_n960), .A2(new_n489), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n960), .A2(new_n489), .ZN(new_n962));
  NOR3_X1   g776(.A1(new_n961), .A2(new_n962), .A3(new_n937), .ZN(G60));
  NAND2_X1  g777(.A1(G478), .A2(G902), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n964), .B(KEYINPUT59), .Z(new_n965));
  INV_X1    g779(.A(new_n965), .ZN(new_n966));
  AND3_X1   g780(.A1(new_n954), .A2(new_n630), .A3(new_n966), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n869), .A2(new_n875), .A3(new_n879), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n630), .B1(new_n968), .B2(new_n966), .ZN(new_n969));
  NOR3_X1   g783(.A1(new_n967), .A2(new_n969), .A3(new_n937), .ZN(G63));
  NAND2_X1  g784(.A1(G217), .A2(G902), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n971), .B(KEYINPUT60), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n972), .B1(new_n876), .B2(new_n878), .ZN(new_n973));
  INV_X1    g787(.A(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(new_n337), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n937), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  AND3_X1   g790(.A1(new_n973), .A2(KEYINPUT124), .A3(new_n677), .ZN(new_n977));
  AOI21_X1  g791(.A(KEYINPUT124), .B1(new_n973), .B2(new_n677), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n976), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(KEYINPUT61), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  OAI211_X1 g795(.A(new_n976), .B(KEYINPUT61), .C1(new_n977), .C2(new_n978), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n981), .A2(new_n982), .ZN(G66));
  OAI21_X1  g797(.A(G953), .B1(new_n529), .B2(new_n208), .ZN(new_n984));
  INV_X1    g798(.A(new_n852), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n984), .B1(new_n985), .B2(G953), .ZN(new_n986));
  OAI211_X1 g800(.A(new_n285), .B(new_n258), .C1(G898), .C2(new_n290), .ZN(new_n987));
  XOR2_X1   g801(.A(new_n987), .B(KEYINPUT125), .Z(new_n988));
  XNOR2_X1  g802(.A(new_n986), .B(new_n988), .ZN(G69));
  NAND2_X1  g803(.A1(new_n572), .A2(new_n583), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n469), .A2(new_n470), .ZN(new_n991));
  XOR2_X1   g805(.A(new_n990), .B(new_n991), .Z(new_n992));
  AOI21_X1  g806(.A(new_n290), .B1(G227), .B2(G900), .ZN(new_n993));
  AOI211_X1 g807(.A(new_n770), .B(new_n692), .C1(new_n641), .C2(new_n651), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n812), .B1(new_n730), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n842), .A2(new_n706), .ZN(new_n996));
  XOR2_X1   g810(.A(new_n996), .B(KEYINPUT62), .Z(new_n997));
  NAND3_X1  g811(.A1(new_n995), .A2(new_n824), .A3(new_n997), .ZN(new_n998));
  AOI211_X1 g812(.A(new_n992), .B(new_n993), .C1(new_n998), .C2(new_n290), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n401), .A2(G900), .A3(G953), .ZN(new_n1000));
  AND2_X1   g814(.A1(new_n778), .A2(new_n782), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n769), .A2(new_n353), .A3(new_n828), .ZN(new_n1002));
  OR2_X1    g816(.A1(new_n803), .A2(new_n1002), .ZN(new_n1003));
  AND3_X1   g817(.A1(new_n824), .A2(new_n1001), .A3(new_n1003), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n842), .B1(new_n803), .B2(new_n811), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n1005), .B(KEYINPUT126), .ZN(new_n1006));
  AND2_X1   g820(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n1000), .B1(new_n1007), .B2(G953), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n999), .B1(new_n1008), .B2(new_n992), .ZN(G72));
  NAND3_X1  g823(.A1(new_n1004), .A2(new_n1006), .A3(new_n985), .ZN(new_n1010));
  NAND2_X1  g824(.A1(G472), .A2(G902), .ZN(new_n1011));
  XOR2_X1   g825(.A(new_n1011), .B(KEYINPUT63), .Z(new_n1012));
  NAND2_X1  g826(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n1013), .A2(new_n547), .A3(new_n577), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n608), .B1(new_n578), .B2(new_n577), .ZN(new_n1015));
  NAND3_X1  g829(.A1(new_n873), .A2(new_n1012), .A3(new_n1015), .ZN(new_n1016));
  OAI21_X1  g830(.A(new_n1012), .B1(new_n998), .B2(new_n852), .ZN(new_n1017));
  NOR2_X1   g831(.A1(new_n577), .A2(new_n547), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n937), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  NAND3_X1  g833(.A1(new_n1014), .A2(new_n1016), .A3(new_n1019), .ZN(new_n1020));
  XNOR2_X1  g834(.A(new_n1020), .B(KEYINPUT127), .ZN(G57));
endmodule


