

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590;

  NOR2_X1 U324 ( .A1(n588), .A2(n491), .ZN(n492) );
  NAND2_X1 U325 ( .A1(n570), .A2(n569), .ZN(n292) );
  XNOR2_X1 U326 ( .A(n301), .B(KEYINPUT79), .ZN(n302) );
  INV_X1 U327 ( .A(KEYINPUT54), .ZN(n425) );
  XNOR2_X1 U328 ( .A(n303), .B(n302), .ZN(n305) );
  XNOR2_X1 U329 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U330 ( .A(n414), .B(n308), .ZN(n309) );
  XNOR2_X1 U331 ( .A(n428), .B(n427), .ZN(n452) );
  XNOR2_X1 U332 ( .A(KEYINPUT97), .B(KEYINPUT26), .ZN(n464) );
  XNOR2_X1 U333 ( .A(n435), .B(n309), .ZN(n310) );
  XNOR2_X1 U334 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U335 ( .A(n465), .B(n464), .ZN(n575) );
  XNOR2_X1 U336 ( .A(n383), .B(n382), .ZN(n403) );
  NOR2_X1 U337 ( .A1(n532), .A2(n571), .ZN(n565) );
  NOR2_X1 U338 ( .A1(n532), .A2(n502), .ZN(n500) );
  XNOR2_X1 U339 ( .A(KEYINPUT38), .B(n494), .ZN(n502) );
  XNOR2_X1 U340 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U341 ( .A(n459), .B(n458), .ZN(G1349GAT) );
  NAND2_X1 U342 ( .A1(G227GAT), .A2(G233GAT), .ZN(n298) );
  XOR2_X1 U343 ( .A(KEYINPUT81), .B(KEYINPUT83), .Z(n294) );
  XNOR2_X1 U344 ( .A(G183GAT), .B(KEYINPUT82), .ZN(n293) );
  XNOR2_X1 U345 ( .A(n294), .B(n293), .ZN(n296) );
  XOR2_X1 U346 ( .A(G43GAT), .B(G99GAT), .Z(n295) );
  XNOR2_X1 U347 ( .A(n296), .B(n295), .ZN(n297) );
  XNOR2_X1 U348 ( .A(n298), .B(n297), .ZN(n313) );
  XOR2_X1 U349 ( .A(G176GAT), .B(KEYINPUT20), .Z(n300) );
  XNOR2_X1 U350 ( .A(G169GAT), .B(G15GAT), .ZN(n299) );
  XNOR2_X1 U351 ( .A(n300), .B(n299), .ZN(n311) );
  XNOR2_X1 U352 ( .A(G120GAT), .B(KEYINPUT80), .ZN(n303) );
  INV_X1 U353 ( .A(KEYINPUT0), .ZN(n301) );
  XNOR2_X1 U354 ( .A(G113GAT), .B(G134GAT), .ZN(n304) );
  XNOR2_X1 U355 ( .A(n305), .B(n304), .ZN(n435) );
  XOR2_X1 U356 ( .A(KEYINPUT17), .B(KEYINPUT19), .Z(n307) );
  XNOR2_X1 U357 ( .A(G190GAT), .B(KEYINPUT18), .ZN(n306) );
  XNOR2_X1 U358 ( .A(n307), .B(n306), .ZN(n414) );
  XOR2_X1 U359 ( .A(G71GAT), .B(G127GAT), .Z(n308) );
  XOR2_X1 U360 ( .A(n311), .B(n310), .Z(n312) );
  XOR2_X1 U361 ( .A(n313), .B(n312), .Z(n570) );
  INV_X1 U362 ( .A(n570), .ZN(n532) );
  XOR2_X1 U363 ( .A(G197GAT), .B(KEYINPUT21), .Z(n418) );
  XOR2_X1 U364 ( .A(G211GAT), .B(n418), .Z(n315) );
  XOR2_X1 U365 ( .A(G218GAT), .B(G162GAT), .Z(n395) );
  XNOR2_X1 U366 ( .A(G50GAT), .B(n395), .ZN(n314) );
  XNOR2_X1 U367 ( .A(n315), .B(n314), .ZN(n319) );
  XOR2_X1 U368 ( .A(KEYINPUT22), .B(G204GAT), .Z(n317) );
  NAND2_X1 U369 ( .A1(G228GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U370 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U371 ( .A(n319), .B(n318), .Z(n321) );
  XOR2_X1 U372 ( .A(G141GAT), .B(G22GAT), .Z(n359) );
  XNOR2_X1 U373 ( .A(n359), .B(KEYINPUT23), .ZN(n320) );
  XNOR2_X1 U374 ( .A(n321), .B(n320), .ZN(n325) );
  XOR2_X1 U375 ( .A(KEYINPUT86), .B(G155GAT), .Z(n323) );
  XNOR2_X1 U376 ( .A(KEYINPUT24), .B(KEYINPUT87), .ZN(n322) );
  XNOR2_X1 U377 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U378 ( .A(n325), .B(n324), .Z(n330) );
  XOR2_X1 U379 ( .A(G106GAT), .B(G78GAT), .Z(n326) );
  XOR2_X1 U380 ( .A(G148GAT), .B(n326), .Z(n376) );
  XOR2_X1 U381 ( .A(KEYINPUT2), .B(KEYINPUT84), .Z(n328) );
  XNOR2_X1 U382 ( .A(KEYINPUT85), .B(KEYINPUT3), .ZN(n327) );
  XNOR2_X1 U383 ( .A(n328), .B(n327), .ZN(n443) );
  XNOR2_X1 U384 ( .A(n376), .B(n443), .ZN(n329) );
  XNOR2_X1 U385 ( .A(n330), .B(n329), .ZN(n471) );
  XOR2_X1 U386 ( .A(KEYINPUT77), .B(KEYINPUT12), .Z(n332) );
  XNOR2_X1 U387 ( .A(KEYINPUT78), .B(KEYINPUT76), .ZN(n331) );
  XOR2_X1 U388 ( .A(n332), .B(n331), .Z(n336) );
  XOR2_X1 U389 ( .A(G183GAT), .B(G211GAT), .Z(n411) );
  XOR2_X1 U390 ( .A(G127GAT), .B(G155GAT), .Z(n442) );
  XOR2_X1 U391 ( .A(n411), .B(n442), .Z(n334) );
  XNOR2_X1 U392 ( .A(G22GAT), .B(G78GAT), .ZN(n333) );
  XNOR2_X1 U393 ( .A(n334), .B(n333), .ZN(n335) );
  XNOR2_X1 U394 ( .A(n336), .B(n335), .ZN(n338) );
  NAND2_X1 U395 ( .A1(G231GAT), .A2(G233GAT), .ZN(n337) );
  XNOR2_X1 U396 ( .A(n338), .B(n337), .ZN(n342) );
  XOR2_X1 U397 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n340) );
  XNOR2_X1 U398 ( .A(G8GAT), .B(G64GAT), .ZN(n339) );
  XNOR2_X1 U399 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U400 ( .A(n342), .B(n341), .Z(n347) );
  XOR2_X1 U401 ( .A(KEYINPUT66), .B(KEYINPUT67), .Z(n344) );
  XNOR2_X1 U402 ( .A(G15GAT), .B(G1GAT), .ZN(n343) );
  XNOR2_X1 U403 ( .A(n344), .B(n343), .ZN(n352) );
  XNOR2_X1 U404 ( .A(G71GAT), .B(G57GAT), .ZN(n345) );
  XNOR2_X1 U405 ( .A(n345), .B(KEYINPUT13), .ZN(n363) );
  XNOR2_X1 U406 ( .A(n352), .B(n363), .ZN(n346) );
  XOR2_X1 U407 ( .A(n347), .B(n346), .Z(n559) );
  XOR2_X1 U408 ( .A(n559), .B(KEYINPUT109), .Z(n566) );
  XNOR2_X1 U409 ( .A(G36GAT), .B(KEYINPUT7), .ZN(n348) );
  XNOR2_X1 U410 ( .A(n348), .B(G29GAT), .ZN(n349) );
  XOR2_X1 U411 ( .A(n349), .B(KEYINPUT8), .Z(n351) );
  XNOR2_X1 U412 ( .A(G43GAT), .B(G50GAT), .ZN(n350) );
  XNOR2_X1 U413 ( .A(n351), .B(n350), .ZN(n399) );
  XOR2_X1 U414 ( .A(n352), .B(KEYINPUT65), .Z(n354) );
  NAND2_X1 U415 ( .A1(G229GAT), .A2(G233GAT), .ZN(n353) );
  XNOR2_X1 U416 ( .A(n354), .B(n353), .ZN(n358) );
  XOR2_X1 U417 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n356) );
  XNOR2_X1 U418 ( .A(G197GAT), .B(G113GAT), .ZN(n355) );
  XNOR2_X1 U419 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U420 ( .A(n358), .B(n357), .Z(n361) );
  XOR2_X1 U421 ( .A(G169GAT), .B(G8GAT), .Z(n412) );
  XNOR2_X1 U422 ( .A(n359), .B(n412), .ZN(n360) );
  XNOR2_X1 U423 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U424 ( .A(n399), .B(n362), .Z(n578) );
  XNOR2_X1 U425 ( .A(n363), .B(KEYINPUT33), .ZN(n365) );
  XOR2_X1 U426 ( .A(G99GAT), .B(G85GAT), .Z(n388) );
  XOR2_X1 U427 ( .A(G120GAT), .B(n388), .Z(n364) );
  XNOR2_X1 U428 ( .A(n365), .B(n364), .ZN(n368) );
  XOR2_X1 U429 ( .A(KEYINPUT31), .B(KEYINPUT32), .Z(n367) );
  NAND2_X1 U430 ( .A1(G230GAT), .A2(G233GAT), .ZN(n366) );
  XNOR2_X1 U431 ( .A(n367), .B(n366), .ZN(n369) );
  NAND2_X1 U432 ( .A1(n368), .A2(n369), .ZN(n373) );
  INV_X1 U433 ( .A(n368), .ZN(n371) );
  INV_X1 U434 ( .A(n369), .ZN(n370) );
  NAND2_X1 U435 ( .A1(n371), .A2(n370), .ZN(n372) );
  NAND2_X1 U436 ( .A1(n373), .A2(n372), .ZN(n383) );
  XOR2_X1 U437 ( .A(G64GAT), .B(G92GAT), .Z(n375) );
  XNOR2_X1 U438 ( .A(G176GAT), .B(G204GAT), .ZN(n374) );
  XNOR2_X1 U439 ( .A(n375), .B(n374), .ZN(n413) );
  XOR2_X1 U440 ( .A(n413), .B(n376), .Z(n381) );
  XOR2_X1 U441 ( .A(KEYINPUT69), .B(KEYINPUT70), .Z(n378) );
  XNOR2_X1 U442 ( .A(KEYINPUT73), .B(KEYINPUT71), .ZN(n377) );
  XNOR2_X1 U443 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X1 U444 ( .A(n379), .B(KEYINPUT72), .Z(n380) );
  XOR2_X1 U445 ( .A(KEYINPUT41), .B(n403), .Z(n554) );
  INV_X1 U446 ( .A(n554), .ZN(n504) );
  NOR2_X1 U447 ( .A1(n578), .A2(n504), .ZN(n384) );
  XNOR2_X1 U448 ( .A(n384), .B(KEYINPUT46), .ZN(n385) );
  NOR2_X1 U449 ( .A1(n566), .A2(n385), .ZN(n400) );
  XOR2_X1 U450 ( .A(KEYINPUT75), .B(KEYINPUT11), .Z(n387) );
  XNOR2_X1 U451 ( .A(G190GAT), .B(G106GAT), .ZN(n386) );
  XNOR2_X1 U452 ( .A(n387), .B(n386), .ZN(n389) );
  XNOR2_X1 U453 ( .A(n389), .B(n388), .ZN(n393) );
  XOR2_X1 U454 ( .A(KEYINPUT10), .B(KEYINPUT9), .Z(n391) );
  NAND2_X1 U455 ( .A1(G232GAT), .A2(G233GAT), .ZN(n390) );
  XNOR2_X1 U456 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U457 ( .A(n393), .B(n392), .ZN(n394) );
  XOR2_X1 U458 ( .A(n394), .B(G92GAT), .Z(n397) );
  XNOR2_X1 U459 ( .A(G134GAT), .B(n395), .ZN(n396) );
  XNOR2_X1 U460 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U461 ( .A(n399), .B(n398), .ZN(n476) );
  NAND2_X1 U462 ( .A1(n400), .A2(n476), .ZN(n402) );
  XOR2_X1 U463 ( .A(KEYINPUT110), .B(KEYINPUT47), .Z(n401) );
  XNOR2_X1 U464 ( .A(n402), .B(n401), .ZN(n409) );
  XOR2_X1 U465 ( .A(KEYINPUT68), .B(n578), .Z(n563) );
  INV_X1 U466 ( .A(n563), .ZN(n479) );
  XOR2_X1 U467 ( .A(KEYINPUT45), .B(KEYINPUT111), .Z(n405) );
  INV_X1 U468 ( .A(n476), .ZN(n569) );
  XOR2_X1 U469 ( .A(KEYINPUT36), .B(n569), .Z(n588) );
  INV_X1 U470 ( .A(n559), .ZN(n585) );
  NOR2_X1 U471 ( .A1(n588), .A2(n585), .ZN(n404) );
  XOR2_X1 U472 ( .A(n405), .B(n404), .Z(n406) );
  NOR2_X1 U473 ( .A1(n403), .A2(n406), .ZN(n407) );
  NAND2_X1 U474 ( .A1(n479), .A2(n407), .ZN(n408) );
  NAND2_X1 U475 ( .A1(n409), .A2(n408), .ZN(n410) );
  XNOR2_X1 U476 ( .A(n410), .B(KEYINPUT48), .ZN(n529) );
  XNOR2_X1 U477 ( .A(n412), .B(n411), .ZN(n424) );
  XNOR2_X1 U478 ( .A(n414), .B(n413), .ZN(n422) );
  XOR2_X1 U479 ( .A(KEYINPUT95), .B(KEYINPUT94), .Z(n416) );
  XNOR2_X1 U480 ( .A(G36GAT), .B(G218GAT), .ZN(n415) );
  XNOR2_X1 U481 ( .A(n416), .B(n415), .ZN(n417) );
  XOR2_X1 U482 ( .A(n418), .B(n417), .Z(n420) );
  NAND2_X1 U483 ( .A1(G226GAT), .A2(G233GAT), .ZN(n419) );
  XNOR2_X1 U484 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U485 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U486 ( .A(n424), .B(n423), .Z(n522) );
  INV_X1 U487 ( .A(n522), .ZN(n460) );
  NAND2_X1 U488 ( .A1(n529), .A2(n460), .ZN(n428) );
  XOR2_X1 U489 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n426) );
  XOR2_X1 U490 ( .A(G57GAT), .B(KEYINPUT93), .Z(n430) );
  XNOR2_X1 U491 ( .A(KEYINPUT90), .B(KEYINPUT92), .ZN(n429) );
  XNOR2_X1 U492 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U493 ( .A(G1GAT), .B(n431), .Z(n433) );
  NAND2_X1 U494 ( .A1(G225GAT), .A2(G233GAT), .ZN(n432) );
  XNOR2_X1 U495 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U496 ( .A(n434), .B(KEYINPUT91), .Z(n437) );
  XNOR2_X1 U497 ( .A(n435), .B(KEYINPUT6), .ZN(n436) );
  XNOR2_X1 U498 ( .A(n437), .B(n436), .ZN(n441) );
  XOR2_X1 U499 ( .A(KEYINPUT4), .B(G162GAT), .Z(n439) );
  XNOR2_X1 U500 ( .A(G141GAT), .B(G148GAT), .ZN(n438) );
  XNOR2_X1 U501 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U502 ( .A(n441), .B(n440), .Z(n451) );
  XOR2_X1 U503 ( .A(n442), .B(G85GAT), .Z(n445) );
  XNOR2_X1 U504 ( .A(G29GAT), .B(n443), .ZN(n444) );
  XNOR2_X1 U505 ( .A(n445), .B(n444), .ZN(n449) );
  XOR2_X1 U506 ( .A(KEYINPUT5), .B(KEYINPUT1), .Z(n447) );
  XNOR2_X1 U507 ( .A(KEYINPUT88), .B(KEYINPUT89), .ZN(n446) );
  XNOR2_X1 U508 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U509 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U510 ( .A(n451), .B(n450), .ZN(n519) );
  NAND2_X1 U511 ( .A1(n452), .A2(n519), .ZN(n453) );
  XOR2_X1 U512 ( .A(KEYINPUT64), .B(n453), .Z(n577) );
  NAND2_X1 U513 ( .A1(n471), .A2(n577), .ZN(n455) );
  XOR2_X1 U514 ( .A(KEYINPUT55), .B(KEYINPUT124), .Z(n454) );
  XNOR2_X1 U515 ( .A(n455), .B(n454), .ZN(n571) );
  NAND2_X1 U516 ( .A1(n565), .A2(n554), .ZN(n459) );
  XOR2_X1 U517 ( .A(G176GAT), .B(KEYINPUT125), .Z(n457) );
  XOR2_X1 U518 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n456) );
  NAND2_X1 U519 ( .A1(n460), .A2(n570), .ZN(n461) );
  XNOR2_X1 U520 ( .A(KEYINPUT98), .B(n461), .ZN(n462) );
  NAND2_X1 U521 ( .A1(n462), .A2(n471), .ZN(n463) );
  XNOR2_X1 U522 ( .A(n463), .B(KEYINPUT25), .ZN(n467) );
  XNOR2_X1 U523 ( .A(n522), .B(KEYINPUT27), .ZN(n470) );
  NOR2_X1 U524 ( .A1(n471), .A2(n570), .ZN(n465) );
  NOR2_X1 U525 ( .A1(n470), .A2(n575), .ZN(n466) );
  NOR2_X1 U526 ( .A1(n467), .A2(n466), .ZN(n468) );
  XNOR2_X1 U527 ( .A(n468), .B(KEYINPUT99), .ZN(n469) );
  NAND2_X1 U528 ( .A1(n469), .A2(n519), .ZN(n475) );
  NOR2_X1 U529 ( .A1(n519), .A2(n470), .ZN(n530) );
  XNOR2_X1 U530 ( .A(n471), .B(KEYINPUT28), .ZN(n528) );
  NAND2_X1 U531 ( .A1(n530), .A2(n528), .ZN(n472) );
  XOR2_X1 U532 ( .A(KEYINPUT96), .B(n472), .Z(n473) );
  NAND2_X1 U533 ( .A1(n532), .A2(n473), .ZN(n474) );
  NAND2_X1 U534 ( .A1(n475), .A2(n474), .ZN(n490) );
  NAND2_X1 U535 ( .A1(n476), .A2(n559), .ZN(n477) );
  XOR2_X1 U536 ( .A(KEYINPUT16), .B(n477), .Z(n478) );
  AND2_X1 U537 ( .A1(n490), .A2(n478), .ZN(n506) );
  NOR2_X1 U538 ( .A1(n403), .A2(n479), .ZN(n480) );
  XNOR2_X1 U539 ( .A(n480), .B(KEYINPUT74), .ZN(n493) );
  NAND2_X1 U540 ( .A1(n506), .A2(n493), .ZN(n487) );
  NOR2_X1 U541 ( .A1(n519), .A2(n487), .ZN(n482) );
  XNOR2_X1 U542 ( .A(KEYINPUT100), .B(KEYINPUT34), .ZN(n481) );
  XNOR2_X1 U543 ( .A(n482), .B(n481), .ZN(n483) );
  XOR2_X1 U544 ( .A(G1GAT), .B(n483), .Z(G1324GAT) );
  NOR2_X1 U545 ( .A1(n522), .A2(n487), .ZN(n484) );
  XOR2_X1 U546 ( .A(G8GAT), .B(n484), .Z(G1325GAT) );
  NOR2_X1 U547 ( .A1(n532), .A2(n487), .ZN(n486) );
  XNOR2_X1 U548 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n485) );
  XNOR2_X1 U549 ( .A(n486), .B(n485), .ZN(G1326GAT) );
  NOR2_X1 U550 ( .A1(n528), .A2(n487), .ZN(n489) );
  XNOR2_X1 U551 ( .A(G22GAT), .B(KEYINPUT101), .ZN(n488) );
  XNOR2_X1 U552 ( .A(n489), .B(n488), .ZN(G1327GAT) );
  XNOR2_X1 U553 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n496) );
  NAND2_X1 U554 ( .A1(n585), .A2(n490), .ZN(n491) );
  XOR2_X1 U555 ( .A(KEYINPUT37), .B(n492), .Z(n518) );
  NAND2_X1 U556 ( .A1(n518), .A2(n493), .ZN(n494) );
  NOR2_X1 U557 ( .A1(n519), .A2(n502), .ZN(n495) );
  XNOR2_X1 U558 ( .A(n496), .B(n495), .ZN(G1328GAT) );
  NOR2_X1 U559 ( .A1(n502), .A2(n522), .ZN(n498) );
  XNOR2_X1 U560 ( .A(KEYINPUT102), .B(KEYINPUT103), .ZN(n497) );
  XNOR2_X1 U561 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U562 ( .A(G36GAT), .B(n499), .ZN(G1329GAT) );
  XOR2_X1 U563 ( .A(KEYINPUT40), .B(n500), .Z(n501) );
  XNOR2_X1 U564 ( .A(G43GAT), .B(n501), .ZN(G1330GAT) );
  NOR2_X1 U565 ( .A1(n502), .A2(n528), .ZN(n503) );
  XOR2_X1 U566 ( .A(G50GAT), .B(n503), .Z(G1331GAT) );
  INV_X1 U567 ( .A(n578), .ZN(n549) );
  NOR2_X1 U568 ( .A1(n549), .A2(n504), .ZN(n505) );
  XNOR2_X1 U569 ( .A(n505), .B(KEYINPUT104), .ZN(n517) );
  NAND2_X1 U570 ( .A1(n506), .A2(n517), .ZN(n513) );
  NOR2_X1 U571 ( .A1(n519), .A2(n513), .ZN(n507) );
  XOR2_X1 U572 ( .A(G57GAT), .B(n507), .Z(n508) );
  XNOR2_X1 U573 ( .A(KEYINPUT42), .B(n508), .ZN(G1332GAT) );
  NOR2_X1 U574 ( .A1(n522), .A2(n513), .ZN(n509) );
  XOR2_X1 U575 ( .A(G64GAT), .B(n509), .Z(G1333GAT) );
  NOR2_X1 U576 ( .A1(n532), .A2(n513), .ZN(n511) );
  XNOR2_X1 U577 ( .A(KEYINPUT105), .B(KEYINPUT106), .ZN(n510) );
  XNOR2_X1 U578 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U579 ( .A(G71GAT), .B(n512), .ZN(G1334GAT) );
  NOR2_X1 U580 ( .A1(n528), .A2(n513), .ZN(n515) );
  XNOR2_X1 U581 ( .A(KEYINPUT107), .B(KEYINPUT43), .ZN(n514) );
  XNOR2_X1 U582 ( .A(n515), .B(n514), .ZN(n516) );
  XOR2_X1 U583 ( .A(G78GAT), .B(n516), .Z(G1335GAT) );
  NAND2_X1 U584 ( .A1(n518), .A2(n517), .ZN(n525) );
  NOR2_X1 U585 ( .A1(n519), .A2(n525), .ZN(n520) );
  XOR2_X1 U586 ( .A(n520), .B(KEYINPUT108), .Z(n521) );
  XNOR2_X1 U587 ( .A(G85GAT), .B(n521), .ZN(G1336GAT) );
  NOR2_X1 U588 ( .A1(n522), .A2(n525), .ZN(n523) );
  XOR2_X1 U589 ( .A(G92GAT), .B(n523), .Z(G1337GAT) );
  NOR2_X1 U590 ( .A1(n532), .A2(n525), .ZN(n524) );
  XOR2_X1 U591 ( .A(G99GAT), .B(n524), .Z(G1338GAT) );
  NOR2_X1 U592 ( .A1(n528), .A2(n525), .ZN(n526) );
  XOR2_X1 U593 ( .A(KEYINPUT44), .B(n526), .Z(n527) );
  XNOR2_X1 U594 ( .A(G106GAT), .B(n527), .ZN(G1339GAT) );
  INV_X1 U595 ( .A(n528), .ZN(n535) );
  NAND2_X1 U596 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U597 ( .A(n531), .B(KEYINPUT112), .ZN(n547) );
  NOR2_X1 U598 ( .A1(n532), .A2(n547), .ZN(n533) );
  XNOR2_X1 U599 ( .A(n533), .B(KEYINPUT113), .ZN(n534) );
  NOR2_X1 U600 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U601 ( .A(KEYINPUT114), .B(n536), .ZN(n544) );
  NAND2_X1 U602 ( .A1(n544), .A2(n563), .ZN(n537) );
  XNOR2_X1 U603 ( .A(n537), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT115), .B(KEYINPUT49), .Z(n539) );
  NAND2_X1 U605 ( .A1(n544), .A2(n554), .ZN(n538) );
  XNOR2_X1 U606 ( .A(n539), .B(n538), .ZN(n540) );
  XOR2_X1 U607 ( .A(G120GAT), .B(n540), .Z(G1341GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n542) );
  NAND2_X1 U609 ( .A1(n544), .A2(n566), .ZN(n541) );
  XNOR2_X1 U610 ( .A(n542), .B(n541), .ZN(n543) );
  XOR2_X1 U611 ( .A(G127GAT), .B(n543), .Z(G1342GAT) );
  XOR2_X1 U612 ( .A(G134GAT), .B(KEYINPUT51), .Z(n546) );
  NAND2_X1 U613 ( .A1(n569), .A2(n544), .ZN(n545) );
  XNOR2_X1 U614 ( .A(n546), .B(n545), .ZN(G1343GAT) );
  XNOR2_X1 U615 ( .A(G141GAT), .B(KEYINPUT118), .ZN(n551) );
  NOR2_X1 U616 ( .A1(n547), .A2(n575), .ZN(n548) );
  XOR2_X1 U617 ( .A(KEYINPUT117), .B(n548), .Z(n561) );
  NAND2_X1 U618 ( .A1(n561), .A2(n549), .ZN(n550) );
  XNOR2_X1 U619 ( .A(n551), .B(n550), .ZN(G1344GAT) );
  XOR2_X1 U620 ( .A(KEYINPUT121), .B(KEYINPUT53), .Z(n553) );
  XNOR2_X1 U621 ( .A(KEYINPUT119), .B(KEYINPUT120), .ZN(n552) );
  XNOR2_X1 U622 ( .A(n553), .B(n552), .ZN(n558) );
  XNOR2_X1 U623 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n556) );
  NAND2_X1 U624 ( .A1(n561), .A2(n554), .ZN(n555) );
  XNOR2_X1 U625 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U626 ( .A(n558), .B(n557), .ZN(G1345GAT) );
  NAND2_X1 U627 ( .A1(n561), .A2(n559), .ZN(n560) );
  XNOR2_X1 U628 ( .A(G155GAT), .B(n560), .ZN(G1346GAT) );
  NAND2_X1 U629 ( .A1(n561), .A2(n569), .ZN(n562) );
  XNOR2_X1 U630 ( .A(n562), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U631 ( .A1(n563), .A2(n565), .ZN(n564) );
  XNOR2_X1 U632 ( .A(G169GAT), .B(n564), .ZN(G1348GAT) );
  NAND2_X1 U633 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n567), .B(KEYINPUT126), .ZN(n568) );
  XNOR2_X1 U635 ( .A(G183GAT), .B(n568), .ZN(G1350GAT) );
  XOR2_X1 U636 ( .A(KEYINPUT127), .B(KEYINPUT58), .Z(n573) );
  OR2_X1 U637 ( .A1(n292), .A2(n571), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(n574) );
  XNOR2_X1 U639 ( .A(G190GAT), .B(n574), .ZN(G1351GAT) );
  INV_X1 U640 ( .A(n575), .ZN(n576) );
  NAND2_X1 U641 ( .A1(n577), .A2(n576), .ZN(n587) );
  NOR2_X1 U642 ( .A1(n578), .A2(n587), .ZN(n580) );
  XNOR2_X1 U643 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U645 ( .A(G197GAT), .B(n581), .ZN(G1352GAT) );
  XOR2_X1 U646 ( .A(G204GAT), .B(KEYINPUT61), .Z(n584) );
  INV_X1 U647 ( .A(n587), .ZN(n582) );
  NAND2_X1 U648 ( .A1(n582), .A2(n403), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(G1353GAT) );
  NOR2_X1 U650 ( .A1(n585), .A2(n587), .ZN(n586) );
  XOR2_X1 U651 ( .A(G211GAT), .B(n586), .Z(G1354GAT) );
  NOR2_X1 U652 ( .A1(n588), .A2(n587), .ZN(n589) );
  XOR2_X1 U653 ( .A(KEYINPUT62), .B(n589), .Z(n590) );
  XNOR2_X1 U654 ( .A(G218GAT), .B(n590), .ZN(G1355GAT) );
endmodule

