

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583;

  XNOR2_X1 U322 ( .A(G148GAT), .B(KEYINPUT72), .ZN(n331) );
  XNOR2_X1 U323 ( .A(KEYINPUT113), .B(KEYINPUT47), .ZN(n381) );
  INV_X1 U324 ( .A(KEYINPUT65), .ZN(n340) );
  XNOR2_X1 U325 ( .A(n382), .B(n381), .ZN(n387) );
  XNOR2_X1 U326 ( .A(n340), .B(KEYINPUT41), .ZN(n341) );
  XNOR2_X1 U327 ( .A(n573), .B(n341), .ZN(n495) );
  INV_X1 U328 ( .A(G183GAT), .ZN(n450) );
  XOR2_X1 U329 ( .A(n360), .B(n359), .Z(n538) );
  XNOR2_X1 U330 ( .A(n450), .B(KEYINPUT124), .ZN(n451) );
  XNOR2_X1 U331 ( .A(n452), .B(n451), .ZN(G1350GAT) );
  XOR2_X1 U332 ( .A(G64GAT), .B(G78GAT), .Z(n291) );
  XNOR2_X1 U333 ( .A(G1GAT), .B(G8GAT), .ZN(n290) );
  XNOR2_X1 U334 ( .A(n291), .B(n290), .ZN(n306) );
  XOR2_X1 U335 ( .A(KEYINPUT12), .B(KEYINPUT81), .Z(n293) );
  XNOR2_X1 U336 ( .A(KEYINPUT83), .B(KEYINPUT82), .ZN(n292) );
  XNOR2_X1 U337 ( .A(n293), .B(n292), .ZN(n297) );
  XOR2_X1 U338 ( .A(G22GAT), .B(G155GAT), .Z(n416) );
  XOR2_X1 U339 ( .A(n416), .B(G211GAT), .Z(n295) );
  XOR2_X1 U340 ( .A(G15GAT), .B(G127GAT), .Z(n432) );
  XNOR2_X1 U341 ( .A(n432), .B(G183GAT), .ZN(n294) );
  XNOR2_X1 U342 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U343 ( .A(n297), .B(n296), .Z(n299) );
  NAND2_X1 U344 ( .A1(G231GAT), .A2(G233GAT), .ZN(n298) );
  XNOR2_X1 U345 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U346 ( .A(n300), .B(KEYINPUT15), .Z(n304) );
  XOR2_X1 U347 ( .A(KEYINPUT70), .B(KEYINPUT13), .Z(n302) );
  XNOR2_X1 U348 ( .A(G71GAT), .B(G57GAT), .ZN(n301) );
  XNOR2_X1 U349 ( .A(n302), .B(n301), .ZN(n321) );
  XNOR2_X1 U350 ( .A(n321), .B(KEYINPUT14), .ZN(n303) );
  XNOR2_X1 U351 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U352 ( .A(n306), .B(n305), .ZN(n576) );
  XOR2_X1 U353 ( .A(G36GAT), .B(G190GAT), .Z(n371) );
  XOR2_X1 U354 ( .A(G176GAT), .B(G64GAT), .Z(n322) );
  XNOR2_X1 U355 ( .A(n371), .B(n322), .ZN(n320) );
  XOR2_X1 U356 ( .A(KEYINPUT95), .B(KEYINPUT96), .Z(n308) );
  NAND2_X1 U357 ( .A1(G226GAT), .A2(G233GAT), .ZN(n307) );
  XNOR2_X1 U358 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U359 ( .A(n309), .B(KEYINPUT94), .Z(n315) );
  XOR2_X1 U360 ( .A(G183GAT), .B(KEYINPUT19), .Z(n311) );
  XNOR2_X1 U361 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n310) );
  XNOR2_X1 U362 ( .A(n311), .B(n310), .ZN(n433) );
  XOR2_X1 U363 ( .A(G211GAT), .B(KEYINPUT21), .Z(n313) );
  XNOR2_X1 U364 ( .A(G197GAT), .B(G218GAT), .ZN(n312) );
  XNOR2_X1 U365 ( .A(n313), .B(n312), .ZN(n415) );
  XNOR2_X1 U366 ( .A(n433), .B(n415), .ZN(n314) );
  XNOR2_X1 U367 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U368 ( .A(n316), .B(G92GAT), .Z(n318) );
  XOR2_X1 U369 ( .A(G169GAT), .B(G8GAT), .Z(n347) );
  XNOR2_X1 U370 ( .A(n347), .B(G204GAT), .ZN(n317) );
  XNOR2_X1 U371 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U372 ( .A(n320), .B(n319), .Z(n512) );
  INV_X1 U373 ( .A(n512), .ZN(n391) );
  INV_X1 U374 ( .A(n576), .ZN(n548) );
  XOR2_X1 U375 ( .A(KEYINPUT31), .B(n321), .Z(n324) );
  XNOR2_X1 U376 ( .A(G120GAT), .B(n322), .ZN(n323) );
  XNOR2_X1 U377 ( .A(n324), .B(n323), .ZN(n330) );
  XOR2_X1 U378 ( .A(KEYINPUT74), .B(G92GAT), .Z(n326) );
  XNOR2_X1 U379 ( .A(G99GAT), .B(G85GAT), .ZN(n325) );
  XNOR2_X1 U380 ( .A(n326), .B(n325), .ZN(n368) );
  XOR2_X1 U381 ( .A(n368), .B(KEYINPUT76), .Z(n328) );
  NAND2_X1 U382 ( .A1(G230GAT), .A2(G233GAT), .ZN(n327) );
  XNOR2_X1 U383 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U384 ( .A(n330), .B(n329), .ZN(n339) );
  XNOR2_X1 U385 ( .A(n331), .B(KEYINPUT73), .ZN(n332) );
  XOR2_X1 U386 ( .A(G204GAT), .B(n332), .Z(n334) );
  XNOR2_X1 U387 ( .A(G78GAT), .B(G106GAT), .ZN(n333) );
  XOR2_X1 U388 ( .A(n334), .B(n333), .Z(n428) );
  XOR2_X1 U389 ( .A(KEYINPUT71), .B(KEYINPUT33), .Z(n336) );
  XNOR2_X1 U390 ( .A(KEYINPUT32), .B(KEYINPUT75), .ZN(n335) );
  XNOR2_X1 U391 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U392 ( .A(n428), .B(n337), .ZN(n338) );
  XNOR2_X1 U393 ( .A(n339), .B(n338), .ZN(n573) );
  XOR2_X1 U394 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n343) );
  XNOR2_X1 U395 ( .A(G22GAT), .B(G1GAT), .ZN(n342) );
  XNOR2_X1 U396 ( .A(n343), .B(n342), .ZN(n360) );
  XOR2_X1 U397 ( .A(G197GAT), .B(G141GAT), .Z(n345) );
  XNOR2_X1 U398 ( .A(G113GAT), .B(G15GAT), .ZN(n344) );
  XNOR2_X1 U399 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U400 ( .A(n346), .B(G36GAT), .Z(n349) );
  XNOR2_X1 U401 ( .A(n347), .B(G50GAT), .ZN(n348) );
  XNOR2_X1 U402 ( .A(n349), .B(n348), .ZN(n353) );
  XOR2_X1 U403 ( .A(KEYINPUT69), .B(KEYINPUT67), .Z(n351) );
  NAND2_X1 U404 ( .A1(G229GAT), .A2(G233GAT), .ZN(n350) );
  XNOR2_X1 U405 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U406 ( .A(n353), .B(n352), .Z(n358) );
  XOR2_X1 U407 ( .A(KEYINPUT68), .B(KEYINPUT8), .Z(n355) );
  XNOR2_X1 U408 ( .A(G43GAT), .B(G29GAT), .ZN(n354) );
  XNOR2_X1 U409 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U410 ( .A(KEYINPUT7), .B(n356), .Z(n379) );
  XNOR2_X1 U411 ( .A(n379), .B(KEYINPUT66), .ZN(n357) );
  XNOR2_X1 U412 ( .A(n358), .B(n357), .ZN(n359) );
  AND2_X1 U413 ( .A1(n495), .A2(n538), .ZN(n361) );
  XNOR2_X1 U414 ( .A(n361), .B(KEYINPUT46), .ZN(n362) );
  NOR2_X1 U415 ( .A1(n548), .A2(n362), .ZN(n363) );
  XNOR2_X1 U416 ( .A(KEYINPUT112), .B(n363), .ZN(n380) );
  XOR2_X1 U417 ( .A(KEYINPUT11), .B(KEYINPUT10), .Z(n365) );
  NAND2_X1 U418 ( .A1(G232GAT), .A2(G233GAT), .ZN(n364) );
  XNOR2_X1 U419 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U420 ( .A(n366), .B(KEYINPUT80), .Z(n370) );
  XNOR2_X1 U421 ( .A(G50GAT), .B(KEYINPUT77), .ZN(n367) );
  XNOR2_X1 U422 ( .A(n367), .B(G162GAT), .ZN(n423) );
  XNOR2_X1 U423 ( .A(n423), .B(n368), .ZN(n369) );
  XNOR2_X1 U424 ( .A(n370), .B(n369), .ZN(n375) );
  XOR2_X1 U425 ( .A(KEYINPUT78), .B(n371), .Z(n373) );
  XOR2_X1 U426 ( .A(G134GAT), .B(KEYINPUT79), .Z(n406) );
  XNOR2_X1 U427 ( .A(G218GAT), .B(n406), .ZN(n372) );
  XNOR2_X1 U428 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U429 ( .A(n375), .B(n374), .Z(n377) );
  XNOR2_X1 U430 ( .A(G106GAT), .B(KEYINPUT9), .ZN(n376) );
  XNOR2_X1 U431 ( .A(n377), .B(n376), .ZN(n378) );
  XOR2_X1 U432 ( .A(n379), .B(n378), .Z(n551) );
  INV_X1 U433 ( .A(n551), .ZN(n560) );
  NAND2_X1 U434 ( .A1(n380), .A2(n560), .ZN(n382) );
  XOR2_X1 U435 ( .A(KEYINPUT36), .B(n551), .Z(n580) );
  NOR2_X1 U436 ( .A1(n580), .A2(n576), .ZN(n383) );
  XOR2_X1 U437 ( .A(KEYINPUT45), .B(n383), .Z(n384) );
  NOR2_X1 U438 ( .A1(n538), .A2(n384), .ZN(n385) );
  NAND2_X1 U439 ( .A1(n385), .A2(n573), .ZN(n386) );
  NAND2_X1 U440 ( .A1(n387), .A2(n386), .ZN(n390) );
  XOR2_X1 U441 ( .A(KEYINPUT64), .B(KEYINPUT114), .Z(n388) );
  XNOR2_X1 U442 ( .A(KEYINPUT48), .B(n388), .ZN(n389) );
  XNOR2_X1 U443 ( .A(n390), .B(n389), .ZN(n535) );
  NOR2_X1 U444 ( .A1(n391), .A2(n535), .ZN(n392) );
  XNOR2_X1 U445 ( .A(n392), .B(KEYINPUT54), .ZN(n565) );
  XOR2_X1 U446 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n394) );
  XNOR2_X1 U447 ( .A(KEYINPUT1), .B(KEYINPUT91), .ZN(n393) );
  XNOR2_X1 U448 ( .A(n394), .B(n393), .ZN(n414) );
  XOR2_X1 U449 ( .A(G85GAT), .B(G155GAT), .Z(n396) );
  XNOR2_X1 U450 ( .A(G127GAT), .B(G148GAT), .ZN(n395) );
  XNOR2_X1 U451 ( .A(n396), .B(n395), .ZN(n400) );
  XOR2_X1 U452 ( .A(KEYINPUT92), .B(KEYINPUT93), .Z(n398) );
  XNOR2_X1 U453 ( .A(G1GAT), .B(G57GAT), .ZN(n397) );
  XNOR2_X1 U454 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U455 ( .A(n400), .B(n399), .Z(n412) );
  XNOR2_X1 U456 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n401) );
  XNOR2_X1 U457 ( .A(n401), .B(G120GAT), .ZN(n436) );
  XOR2_X1 U458 ( .A(n436), .B(KEYINPUT6), .Z(n403) );
  NAND2_X1 U459 ( .A1(G225GAT), .A2(G233GAT), .ZN(n402) );
  XNOR2_X1 U460 ( .A(n403), .B(n402), .ZN(n410) );
  XOR2_X1 U461 ( .A(KEYINPUT88), .B(KEYINPUT3), .Z(n405) );
  XNOR2_X1 U462 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n404) );
  XNOR2_X1 U463 ( .A(n405), .B(n404), .ZN(n422) );
  XOR2_X1 U464 ( .A(n406), .B(n422), .Z(n408) );
  XNOR2_X1 U465 ( .A(G29GAT), .B(G162GAT), .ZN(n407) );
  XNOR2_X1 U466 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U467 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U468 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U469 ( .A(n414), .B(n413), .ZN(n564) );
  XOR2_X1 U470 ( .A(n416), .B(n415), .Z(n418) );
  XNOR2_X1 U471 ( .A(KEYINPUT24), .B(KEYINPUT22), .ZN(n417) );
  XNOR2_X1 U472 ( .A(n418), .B(n417), .ZN(n427) );
  XOR2_X1 U473 ( .A(KEYINPUT23), .B(KEYINPUT90), .Z(n420) );
  NAND2_X1 U474 ( .A1(G228GAT), .A2(G233GAT), .ZN(n419) );
  XNOR2_X1 U475 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U476 ( .A(n421), .B(KEYINPUT89), .Z(n425) );
  XNOR2_X1 U477 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U478 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U479 ( .A(n427), .B(n426), .ZN(n429) );
  XNOR2_X1 U480 ( .A(n429), .B(n428), .ZN(n464) );
  AND2_X1 U481 ( .A1(n564), .A2(n464), .ZN(n430) );
  NAND2_X1 U482 ( .A1(n565), .A2(n430), .ZN(n431) );
  XNOR2_X1 U483 ( .A(n431), .B(KEYINPUT55), .ZN(n449) );
  XOR2_X1 U484 ( .A(n433), .B(n432), .Z(n435) );
  XNOR2_X1 U485 ( .A(G134GAT), .B(G190GAT), .ZN(n434) );
  XNOR2_X1 U486 ( .A(n435), .B(n434), .ZN(n440) );
  XOR2_X1 U487 ( .A(n436), .B(G169GAT), .Z(n438) );
  NAND2_X1 U488 ( .A1(G227GAT), .A2(G233GAT), .ZN(n437) );
  XNOR2_X1 U489 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U490 ( .A(n440), .B(n439), .Z(n448) );
  XOR2_X1 U491 ( .A(KEYINPUT20), .B(KEYINPUT86), .Z(n442) );
  XNOR2_X1 U492 ( .A(G43GAT), .B(G99GAT), .ZN(n441) );
  XNOR2_X1 U493 ( .A(n442), .B(n441), .ZN(n446) );
  XOR2_X1 U494 ( .A(KEYINPUT87), .B(G71GAT), .Z(n444) );
  XNOR2_X1 U495 ( .A(KEYINPUT85), .B(G176GAT), .ZN(n443) );
  XNOR2_X1 U496 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U497 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U498 ( .A(n448), .B(n447), .ZN(n522) );
  NAND2_X1 U499 ( .A1(n449), .A2(n522), .ZN(n559) );
  NOR2_X1 U500 ( .A1(n576), .A2(n559), .ZN(n452) );
  XNOR2_X1 U501 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n471) );
  INV_X1 U502 ( .A(n564), .ZN(n510) );
  NAND2_X1 U503 ( .A1(n538), .A2(n573), .ZN(n482) );
  XOR2_X1 U504 ( .A(KEYINPUT84), .B(KEYINPUT16), .Z(n454) );
  NAND2_X1 U505 ( .A1(n548), .A2(n560), .ZN(n453) );
  XNOR2_X1 U506 ( .A(n454), .B(n453), .ZN(n469) );
  NAND2_X1 U507 ( .A1(n512), .A2(n522), .ZN(n455) );
  NAND2_X1 U508 ( .A1(n455), .A2(n464), .ZN(n456) );
  XNOR2_X1 U509 ( .A(n456), .B(KEYINPUT98), .ZN(n457) );
  XOR2_X1 U510 ( .A(KEYINPUT25), .B(n457), .Z(n460) );
  XNOR2_X1 U511 ( .A(n512), .B(KEYINPUT27), .ZN(n463) );
  NOR2_X1 U512 ( .A1(n464), .A2(n522), .ZN(n458) );
  XNOR2_X1 U513 ( .A(n458), .B(KEYINPUT26), .ZN(n566) );
  NAND2_X1 U514 ( .A1(n463), .A2(n566), .ZN(n459) );
  NAND2_X1 U515 ( .A1(n460), .A2(n459), .ZN(n461) );
  NAND2_X1 U516 ( .A1(n564), .A2(n461), .ZN(n462) );
  XNOR2_X1 U517 ( .A(n462), .B(KEYINPUT99), .ZN(n467) );
  NAND2_X1 U518 ( .A1(n510), .A2(n463), .ZN(n534) );
  XOR2_X1 U519 ( .A(KEYINPUT28), .B(n464), .Z(n516) );
  NOR2_X1 U520 ( .A1(n534), .A2(n516), .ZN(n521) );
  XNOR2_X1 U521 ( .A(n521), .B(KEYINPUT97), .ZN(n465) );
  NOR2_X1 U522 ( .A1(n465), .A2(n522), .ZN(n466) );
  NOR2_X1 U523 ( .A1(n467), .A2(n466), .ZN(n478) );
  INV_X1 U524 ( .A(n478), .ZN(n468) );
  NAND2_X1 U525 ( .A1(n469), .A2(n468), .ZN(n496) );
  NOR2_X1 U526 ( .A1(n482), .A2(n496), .ZN(n475) );
  NAND2_X1 U527 ( .A1(n510), .A2(n475), .ZN(n470) );
  XNOR2_X1 U528 ( .A(n471), .B(n470), .ZN(G1324GAT) );
  NAND2_X1 U529 ( .A1(n512), .A2(n475), .ZN(n472) );
  XNOR2_X1 U530 ( .A(n472), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U531 ( .A(G15GAT), .B(KEYINPUT35), .Z(n474) );
  NAND2_X1 U532 ( .A1(n475), .A2(n522), .ZN(n473) );
  XNOR2_X1 U533 ( .A(n474), .B(n473), .ZN(G1326GAT) );
  NAND2_X1 U534 ( .A1(n516), .A2(n475), .ZN(n476) );
  XNOR2_X1 U535 ( .A(n476), .B(KEYINPUT100), .ZN(n477) );
  XNOR2_X1 U536 ( .A(G22GAT), .B(n477), .ZN(G1327GAT) );
  XOR2_X1 U537 ( .A(KEYINPUT39), .B(KEYINPUT103), .Z(n486) );
  NOR2_X1 U538 ( .A1(n580), .A2(n478), .ZN(n479) );
  NAND2_X1 U539 ( .A1(n576), .A2(n479), .ZN(n480) );
  XNOR2_X1 U540 ( .A(n480), .B(KEYINPUT101), .ZN(n481) );
  XNOR2_X1 U541 ( .A(KEYINPUT37), .B(n481), .ZN(n509) );
  NOR2_X1 U542 ( .A1(n509), .A2(n482), .ZN(n484) );
  XNOR2_X1 U543 ( .A(KEYINPUT102), .B(KEYINPUT38), .ZN(n483) );
  XNOR2_X1 U544 ( .A(n484), .B(n483), .ZN(n493) );
  NAND2_X1 U545 ( .A1(n493), .A2(n510), .ZN(n485) );
  XNOR2_X1 U546 ( .A(n486), .B(n485), .ZN(n487) );
  XOR2_X1 U547 ( .A(G29GAT), .B(n487), .Z(G1328GAT) );
  NAND2_X1 U548 ( .A1(n512), .A2(n493), .ZN(n488) );
  XNOR2_X1 U549 ( .A(n488), .B(KEYINPUT104), .ZN(n489) );
  XNOR2_X1 U550 ( .A(G36GAT), .B(n489), .ZN(G1329GAT) );
  XOR2_X1 U551 ( .A(KEYINPUT40), .B(KEYINPUT105), .Z(n491) );
  NAND2_X1 U552 ( .A1(n493), .A2(n522), .ZN(n490) );
  XNOR2_X1 U553 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U554 ( .A(G43GAT), .B(n492), .ZN(G1330GAT) );
  NAND2_X1 U555 ( .A1(n516), .A2(n493), .ZN(n494) );
  XNOR2_X1 U556 ( .A(n494), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U557 ( .A(KEYINPUT106), .B(KEYINPUT42), .Z(n498) );
  INV_X1 U558 ( .A(n538), .ZN(n568) );
  INV_X1 U559 ( .A(n495), .ZN(n554) );
  NAND2_X1 U560 ( .A1(n568), .A2(n495), .ZN(n508) );
  NOR2_X1 U561 ( .A1(n508), .A2(n496), .ZN(n504) );
  NAND2_X1 U562 ( .A1(n504), .A2(n510), .ZN(n497) );
  XNOR2_X1 U563 ( .A(n498), .B(n497), .ZN(n499) );
  XOR2_X1 U564 ( .A(G57GAT), .B(n499), .Z(G1332GAT) );
  XOR2_X1 U565 ( .A(G64GAT), .B(KEYINPUT107), .Z(n501) );
  NAND2_X1 U566 ( .A1(n504), .A2(n512), .ZN(n500) );
  XNOR2_X1 U567 ( .A(n501), .B(n500), .ZN(G1333GAT) );
  NAND2_X1 U568 ( .A1(n504), .A2(n522), .ZN(n502) );
  XNOR2_X1 U569 ( .A(n502), .B(KEYINPUT108), .ZN(n503) );
  XNOR2_X1 U570 ( .A(G71GAT), .B(n503), .ZN(G1334GAT) );
  XOR2_X1 U571 ( .A(KEYINPUT43), .B(KEYINPUT109), .Z(n506) );
  NAND2_X1 U572 ( .A1(n504), .A2(n516), .ZN(n505) );
  XNOR2_X1 U573 ( .A(n506), .B(n505), .ZN(n507) );
  XOR2_X1 U574 ( .A(G78GAT), .B(n507), .Z(G1335GAT) );
  NOR2_X1 U575 ( .A1(n509), .A2(n508), .ZN(n517) );
  NAND2_X1 U576 ( .A1(n510), .A2(n517), .ZN(n511) );
  XNOR2_X1 U577 ( .A(G85GAT), .B(n511), .ZN(G1336GAT) );
  NAND2_X1 U578 ( .A1(n512), .A2(n517), .ZN(n513) );
  XNOR2_X1 U579 ( .A(n513), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U580 ( .A1(n517), .A2(n522), .ZN(n514) );
  XNOR2_X1 U581 ( .A(n514), .B(KEYINPUT110), .ZN(n515) );
  XNOR2_X1 U582 ( .A(G99GAT), .B(n515), .ZN(G1338GAT) );
  XOR2_X1 U583 ( .A(KEYINPUT44), .B(KEYINPUT111), .Z(n519) );
  NAND2_X1 U584 ( .A1(n517), .A2(n516), .ZN(n518) );
  XNOR2_X1 U585 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U586 ( .A(G106GAT), .B(n520), .ZN(G1339GAT) );
  NAND2_X1 U587 ( .A1(n522), .A2(n521), .ZN(n523) );
  NOR2_X1 U588 ( .A1(n535), .A2(n523), .ZN(n530) );
  NAND2_X1 U589 ( .A1(n530), .A2(n538), .ZN(n524) );
  XNOR2_X1 U590 ( .A(n524), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U591 ( .A(G120GAT), .B(KEYINPUT49), .Z(n526) );
  NAND2_X1 U592 ( .A1(n530), .A2(n495), .ZN(n525) );
  XNOR2_X1 U593 ( .A(n526), .B(n525), .ZN(G1341GAT) );
  XOR2_X1 U594 ( .A(KEYINPUT115), .B(KEYINPUT50), .Z(n528) );
  NAND2_X1 U595 ( .A1(n530), .A2(n548), .ZN(n527) );
  XNOR2_X1 U596 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U597 ( .A(G127GAT), .B(n529), .ZN(G1342GAT) );
  XOR2_X1 U598 ( .A(KEYINPUT116), .B(KEYINPUT51), .Z(n532) );
  NAND2_X1 U599 ( .A1(n530), .A2(n551), .ZN(n531) );
  XNOR2_X1 U600 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U601 ( .A(G134GAT), .B(n533), .ZN(G1343GAT) );
  XOR2_X1 U602 ( .A(KEYINPUT118), .B(KEYINPUT119), .Z(n540) );
  NOR2_X1 U603 ( .A1(n535), .A2(n534), .ZN(n536) );
  NAND2_X1 U604 ( .A1(n566), .A2(n536), .ZN(n537) );
  XNOR2_X1 U605 ( .A(n537), .B(KEYINPUT117), .ZN(n550) );
  NAND2_X1 U606 ( .A1(n550), .A2(n538), .ZN(n539) );
  XNOR2_X1 U607 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U608 ( .A(G141GAT), .B(n541), .ZN(G1344GAT) );
  XOR2_X1 U609 ( .A(KEYINPUT122), .B(KEYINPUT53), .Z(n543) );
  XNOR2_X1 U610 ( .A(KEYINPUT120), .B(KEYINPUT121), .ZN(n542) );
  XNOR2_X1 U611 ( .A(n543), .B(n542), .ZN(n547) );
  XOR2_X1 U612 ( .A(G148GAT), .B(KEYINPUT52), .Z(n545) );
  NAND2_X1 U613 ( .A1(n550), .A2(n495), .ZN(n544) );
  XNOR2_X1 U614 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U615 ( .A(n547), .B(n546), .ZN(G1345GAT) );
  NAND2_X1 U616 ( .A1(n550), .A2(n548), .ZN(n549) );
  XNOR2_X1 U617 ( .A(n549), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U618 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U619 ( .A(G162GAT), .B(n552), .ZN(G1347GAT) );
  NOR2_X1 U620 ( .A1(n568), .A2(n559), .ZN(n553) );
  XOR2_X1 U621 ( .A(G169GAT), .B(n553), .Z(G1348GAT) );
  NOR2_X1 U622 ( .A1(n559), .A2(n554), .ZN(n558) );
  XOR2_X1 U623 ( .A(KEYINPUT123), .B(KEYINPUT56), .Z(n556) );
  XNOR2_X1 U624 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n555) );
  XNOR2_X1 U625 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U626 ( .A(n558), .B(n557), .ZN(G1349GAT) );
  INV_X1 U627 ( .A(KEYINPUT58), .ZN(n562) );
  NOR2_X1 U628 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U629 ( .A(n562), .B(n561), .ZN(n563) );
  XNOR2_X1 U630 ( .A(G190GAT), .B(n563), .ZN(G1351GAT) );
  AND2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n567) );
  NAND2_X1 U632 ( .A1(n567), .A2(n566), .ZN(n579) );
  NOR2_X1 U633 ( .A1(n579), .A2(n568), .ZN(n572) );
  XOR2_X1 U634 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n570) );
  XNOR2_X1 U635 ( .A(G197GAT), .B(KEYINPUT125), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(G1352GAT) );
  NOR2_X1 U638 ( .A1(n573), .A2(n579), .ZN(n575) );
  XNOR2_X1 U639 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(G1353GAT) );
  NOR2_X1 U641 ( .A1(n576), .A2(n579), .ZN(n577) );
  XOR2_X1 U642 ( .A(KEYINPUT126), .B(n577), .Z(n578) );
  XNOR2_X1 U643 ( .A(G211GAT), .B(n578), .ZN(G1354GAT) );
  NOR2_X1 U644 ( .A1(n580), .A2(n579), .ZN(n582) );
  XNOR2_X1 U645 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U647 ( .A(G218GAT), .B(n583), .ZN(G1355GAT) );
endmodule

