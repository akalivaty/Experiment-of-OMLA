//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 1 1 0 0 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 0 0 0 0 1 1 0 0 0 0 0 1 0 0 0 1 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 1 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:49 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1289, new_n1290,
    new_n1291, new_n1292, new_n1293, new_n1295, new_n1296, new_n1297,
    new_n1298, new_n1299, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1356, new_n1357, new_n1358, new_n1359,
    new_n1360, new_n1361, new_n1362, new_n1363, new_n1364, new_n1365,
    new_n1366, new_n1367, new_n1368, new_n1369, new_n1370;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  INV_X1    g0002(.A(G77), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  XOR2_X1   g0004(.A(new_n204), .B(KEYINPUT64), .Z(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n209), .B(KEYINPUT0), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G13), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(new_n201), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(G50), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n217));
  INV_X1    g0017(.A(G244), .ZN(new_n218));
  INV_X1    g0018(.A(G107), .ZN(new_n219));
  INV_X1    g0019(.A(G264), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n217), .B1(new_n203), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n207), .B1(new_n221), .B2(new_n224), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n210), .B1(new_n214), .B2(new_n216), .C1(KEYINPUT1), .C2(new_n225), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n225), .ZN(G361));
  XOR2_X1   g0027(.A(G238), .B(G244), .Z(new_n228));
  XNOR2_X1  g0028(.A(KEYINPUT65), .B(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT2), .B(G226), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(G264), .B(G270), .Z(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  XOR2_X1   g0036(.A(G87), .B(G97), .Z(new_n237));
  XOR2_X1   g0037(.A(G107), .B(G116), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G50), .B(G68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G58), .B(G77), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G351));
  INV_X1    g0043(.A(G1), .ZN(new_n244));
  OAI21_X1  g0044(.A(new_n244), .B1(G41), .B2(G45), .ZN(new_n245));
  INV_X1    g0045(.A(new_n245), .ZN(new_n246));
  AND2_X1   g0046(.A1(G1), .A2(G13), .ZN(new_n247));
  NAND2_X1  g0047(.A1(G33), .A2(G41), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n246), .A2(new_n249), .A3(G274), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n245), .A2(KEYINPUT66), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT66), .ZN(new_n252));
  OAI211_X1 g0052(.A(new_n252), .B(new_n244), .C1(G41), .C2(G45), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n251), .A2(new_n249), .A3(new_n253), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n250), .B1(new_n254), .B2(new_n218), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT68), .ZN(new_n256));
  AND2_X1   g0056(.A1(KEYINPUT3), .A2(G33), .ZN(new_n257));
  NOR2_X1   g0057(.A1(KEYINPUT3), .A2(G33), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n256), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT3), .ZN(new_n260));
  INV_X1    g0060(.A(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(KEYINPUT3), .A2(G33), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n262), .A2(KEYINPUT68), .A3(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n259), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G1698), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n266), .A2(G232), .A3(new_n267), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n266), .A2(G238), .A3(G1698), .ZN(new_n269));
  XNOR2_X1  g0069(.A(KEYINPUT71), .B(G107), .ZN(new_n270));
  OAI211_X1 g0070(.A(new_n268), .B(new_n269), .C1(new_n266), .C2(new_n270), .ZN(new_n271));
  AND2_X1   g0071(.A1(G33), .A2(G41), .ZN(new_n272));
  NOR3_X1   g0072(.A1(new_n272), .A2(KEYINPUT69), .A3(new_n211), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT69), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n274), .B1(new_n247), .B2(new_n248), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n255), .B1(new_n271), .B2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G179), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G13), .ZN(new_n281));
  NOR3_X1   g0081(.A1(new_n281), .A2(new_n212), .A3(G1), .ZN(new_n282));
  NAND3_X1  g0082(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(new_n211), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n212), .A2(G1), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n286), .A2(new_n203), .ZN(new_n287));
  AOI22_X1  g0087(.A1(new_n285), .A2(new_n287), .B1(new_n203), .B2(new_n282), .ZN(new_n288));
  XNOR2_X1  g0088(.A(KEYINPUT15), .B(G87), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT72), .ZN(new_n290));
  XNOR2_X1  g0090(.A(new_n289), .B(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n212), .A2(G33), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  XNOR2_X1  g0093(.A(KEYINPUT8), .B(G58), .ZN(new_n294));
  NOR2_X1   g0094(.A1(G20), .A2(G33), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  OAI22_X1  g0096(.A1(new_n294), .A2(new_n296), .B1(new_n212), .B2(new_n203), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n293), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(new_n284), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n288), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n300), .B1(new_n277), .B2(G169), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n280), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n277), .A2(G190), .ZN(new_n304));
  INV_X1    g0104(.A(new_n300), .ZN(new_n305));
  INV_X1    g0105(.A(G200), .ZN(new_n306));
  OAI211_X1 g0106(.A(new_n304), .B(new_n305), .C1(new_n306), .C2(new_n277), .ZN(new_n307));
  INV_X1    g0107(.A(G226), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n250), .B1(new_n254), .B2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT67), .ZN(new_n310));
  XNOR2_X1  g0110(.A(new_n309), .B(new_n310), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n259), .A2(new_n264), .A3(G222), .A4(new_n267), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n259), .A2(new_n264), .A3(G223), .A4(G1698), .ZN(new_n313));
  OAI211_X1 g0113(.A(new_n312), .B(new_n313), .C1(new_n266), .C2(new_n203), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(new_n276), .ZN(new_n315));
  AND2_X1   g0115(.A1(new_n311), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(new_n278), .ZN(new_n317));
  XNOR2_X1  g0117(.A(new_n284), .B(KEYINPUT70), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n318), .A2(new_n282), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n286), .A2(new_n202), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n212), .B1(new_n201), .B2(new_n202), .ZN(new_n322));
  INV_X1    g0122(.A(G150), .ZN(new_n323));
  OAI22_X1  g0123(.A1(new_n294), .A2(new_n292), .B1(new_n323), .B2(new_n296), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n318), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n282), .A2(new_n202), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n321), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  OAI211_X1 g0127(.A(new_n317), .B(new_n327), .C1(G169), .C2(new_n316), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n303), .A2(new_n307), .A3(new_n328), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n311), .A2(G190), .A3(new_n315), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT9), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n327), .A2(new_n331), .ZN(new_n332));
  NAND4_X1  g0132(.A1(new_n321), .A2(new_n325), .A3(KEYINPUT9), .A4(new_n326), .ZN(new_n333));
  AND3_X1   g0133(.A1(new_n330), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n311), .A2(new_n315), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(G200), .ZN(new_n336));
  OAI211_X1 g0136(.A(new_n334), .B(new_n336), .C1(KEYINPUT73), .C2(KEYINPUT10), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT10), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n330), .A2(new_n332), .A3(KEYINPUT73), .A4(new_n333), .ZN(new_n339));
  INV_X1    g0139(.A(new_n336), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n330), .A2(new_n332), .A3(new_n333), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n338), .B(new_n339), .C1(new_n340), .C2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n337), .A2(new_n342), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n329), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n295), .A2(G50), .ZN(new_n345));
  INV_X1    g0145(.A(G68), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(G20), .ZN(new_n347));
  OAI211_X1 g0147(.A(new_n345), .B(new_n347), .C1(new_n203), .C2(new_n292), .ZN(new_n348));
  AOI21_X1  g0148(.A(KEYINPUT75), .B1(new_n318), .B2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT70), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n350), .B1(new_n283), .B2(new_n211), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n284), .A2(KEYINPUT70), .ZN(new_n352));
  OAI211_X1 g0152(.A(new_n348), .B(KEYINPUT75), .C1(new_n351), .C2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  OAI21_X1  g0154(.A(KEYINPUT11), .B1(new_n349), .B2(new_n354), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n348), .B1(new_n352), .B2(new_n351), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT75), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT11), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n358), .A2(new_n359), .A3(new_n353), .ZN(new_n360));
  INV_X1    g0160(.A(new_n282), .ZN(new_n361));
  OR3_X1    g0161(.A1(new_n361), .A2(KEYINPUT12), .A3(G68), .ZN(new_n362));
  OAI21_X1  g0162(.A(KEYINPUT12), .B1(new_n361), .B2(G68), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n286), .A2(new_n346), .ZN(new_n364));
  AOI22_X1  g0164(.A1(new_n362), .A2(new_n363), .B1(new_n285), .B2(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n355), .A2(new_n360), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(KEYINPUT76), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT76), .ZN(new_n368));
  NAND4_X1  g0168(.A1(new_n355), .A2(new_n368), .A3(new_n360), .A4(new_n365), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(G238), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n250), .B1(new_n254), .B2(new_n371), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n259), .A2(new_n264), .A3(G226), .A4(new_n267), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n259), .A2(new_n264), .A3(G232), .A4(G1698), .ZN(new_n374));
  NAND2_X1  g0174(.A1(G33), .A2(G97), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n373), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n372), .B1(new_n376), .B2(new_n276), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT13), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(KEYINPUT74), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT74), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n381), .B1(new_n377), .B2(new_n378), .ZN(new_n382));
  AOI211_X1 g0182(.A(KEYINPUT13), .B(new_n372), .C1(new_n376), .C2(new_n276), .ZN(new_n383));
  INV_X1    g0183(.A(new_n383), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n380), .A2(new_n382), .A3(G190), .A4(new_n384), .ZN(new_n385));
  OAI21_X1  g0185(.A(G200), .B1(new_n379), .B2(new_n383), .ZN(new_n386));
  AND3_X1   g0186(.A1(new_n370), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n370), .ZN(new_n388));
  OAI21_X1  g0188(.A(G169), .B1(new_n379), .B2(new_n383), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(KEYINPUT14), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n380), .A2(new_n382), .A3(G179), .A4(new_n384), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT14), .ZN(new_n392));
  OAI211_X1 g0192(.A(new_n392), .B(G169), .C1(new_n379), .C2(new_n383), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n390), .A2(new_n391), .A3(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n387), .B1(new_n388), .B2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(new_n254), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n249), .A2(G274), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  AOI22_X1  g0198(.A1(new_n396), .A2(G232), .B1(new_n246), .B2(new_n398), .ZN(new_n399));
  NOR2_X1   g0199(.A1(G223), .A2(G1698), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n400), .B1(new_n308), .B2(G1698), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n262), .A2(new_n263), .ZN(new_n402));
  AOI22_X1  g0202(.A1(new_n401), .A2(new_n402), .B1(G33), .B2(G87), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(KEYINPUT78), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n276), .B1(new_n403), .B2(KEYINPUT78), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n399), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  OAI21_X1  g0207(.A(KEYINPUT79), .B1(new_n407), .B2(G179), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n401), .A2(new_n402), .ZN(new_n409));
  NAND2_X1  g0209(.A1(G33), .A2(G87), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT78), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n413), .A2(new_n276), .A3(new_n404), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT79), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n414), .A2(new_n415), .A3(new_n278), .A4(new_n399), .ZN(new_n416));
  INV_X1    g0216(.A(G169), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n407), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n408), .A2(new_n416), .A3(new_n418), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n294), .A2(new_n286), .ZN(new_n420));
  XNOR2_X1  g0220(.A(new_n420), .B(KEYINPUT77), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(new_n319), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n294), .A2(new_n282), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(G58), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n425), .A2(new_n346), .ZN(new_n426));
  OAI21_X1  g0226(.A(G20), .B1(new_n426), .B2(new_n201), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n295), .A2(G159), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n257), .A2(new_n258), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n431), .A2(KEYINPUT7), .A3(new_n212), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  NOR3_X1   g0233(.A1(new_n257), .A2(new_n258), .A3(new_n256), .ZN(new_n434));
  AOI21_X1  g0234(.A(KEYINPUT68), .B1(new_n262), .B2(new_n263), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n212), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT7), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n433), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n430), .B1(new_n438), .B2(new_n346), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT16), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n437), .B1(new_n402), .B2(G20), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n346), .B1(new_n442), .B2(new_n432), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n443), .A2(new_n429), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n299), .B1(new_n444), .B2(KEYINPUT16), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n424), .B1(new_n441), .B2(new_n445), .ZN(new_n446));
  OAI21_X1  g0246(.A(KEYINPUT18), .B1(new_n419), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n407), .A2(G200), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n414), .A2(G190), .A3(new_n399), .ZN(new_n449));
  AND2_X1   g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(KEYINPUT80), .A2(KEYINPUT17), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT80), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT17), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n450), .A2(new_n446), .A3(new_n451), .A4(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(new_n443), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n456), .A2(KEYINPUT16), .A3(new_n430), .ZN(new_n457));
  AOI21_X1  g0257(.A(G20), .B1(new_n259), .B2(new_n264), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n432), .B1(new_n458), .B2(KEYINPUT7), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n429), .B1(new_n459), .B2(G68), .ZN(new_n460));
  OAI211_X1 g0260(.A(new_n457), .B(new_n284), .C1(new_n460), .C2(KEYINPUT16), .ZN(new_n461));
  AOI22_X1  g0261(.A1(new_n421), .A2(new_n319), .B1(new_n282), .B2(new_n294), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n461), .A2(new_n462), .A3(new_n449), .A4(new_n448), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n463), .A2(new_n452), .A3(new_n453), .ZN(new_n464));
  AND2_X1   g0264(.A1(new_n418), .A2(new_n416), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n461), .A2(new_n462), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT18), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n465), .A2(new_n466), .A3(new_n467), .A4(new_n408), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n447), .A2(new_n455), .A3(new_n464), .A4(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n344), .A2(new_n395), .A3(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(G87), .ZN(new_n472));
  NOR3_X1   g0272(.A1(new_n472), .A2(KEYINPUT22), .A3(G20), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n259), .A2(new_n264), .A3(new_n473), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n212), .B(G87), .C1(new_n257), .C2(new_n258), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(KEYINPUT22), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n219), .A2(G20), .ZN(new_n478));
  INV_X1    g0278(.A(G116), .ZN(new_n479));
  OAI22_X1  g0279(.A1(KEYINPUT23), .A2(new_n478), .B1(new_n292), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n270), .A2(G20), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n480), .B1(new_n481), .B2(KEYINPUT23), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n477), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(KEYINPUT86), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT86), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n477), .A2(new_n482), .A3(new_n485), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n484), .A2(KEYINPUT24), .A3(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n485), .B1(new_n477), .B2(new_n482), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT24), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n299), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n487), .A2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(new_n478), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n281), .A2(G1), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n492), .B(new_n493), .C1(KEYINPUT87), .C2(KEYINPUT25), .ZN(new_n494));
  NAND2_X1  g0294(.A1(KEYINPUT87), .A2(KEYINPUT25), .ZN(new_n495));
  OR2_X1    g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n494), .A2(new_n495), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n352), .A2(new_n351), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n244), .A2(G33), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n499), .A2(new_n361), .A3(new_n500), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n498), .B1(new_n501), .B2(new_n219), .ZN(new_n502));
  INV_X1    g0302(.A(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(G257), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(G1698), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n505), .B1(G250), .B2(G1698), .ZN(new_n506));
  INV_X1    g0306(.A(G294), .ZN(new_n507));
  OAI22_X1  g0307(.A1(new_n506), .A2(new_n431), .B1(new_n261), .B2(new_n507), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n272), .A2(new_n211), .ZN(new_n509));
  INV_X1    g0309(.A(G45), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n510), .A2(G1), .ZN(new_n511));
  XNOR2_X1  g0311(.A(KEYINPUT5), .B(G41), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n509), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  AOI22_X1  g0313(.A1(new_n276), .A2(new_n508), .B1(new_n513), .B2(G264), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT89), .ZN(new_n515));
  INV_X1    g0315(.A(G190), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n512), .A2(new_n249), .A3(G274), .A4(new_n511), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n514), .A2(new_n515), .A3(new_n516), .A4(new_n517), .ZN(new_n518));
  AND2_X1   g0318(.A1(KEYINPUT5), .A2(G41), .ZN(new_n519));
  NOR2_X1   g0319(.A1(KEYINPUT5), .A2(G41), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n511), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n521), .A2(G264), .A3(new_n249), .ZN(new_n522));
  NOR2_X1   g0322(.A1(G250), .A2(G1698), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n523), .B1(new_n504), .B2(G1698), .ZN(new_n524));
  AOI22_X1  g0324(.A1(new_n524), .A2(new_n402), .B1(G33), .B2(G294), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n249), .A2(KEYINPUT69), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n247), .A2(new_n274), .A3(new_n248), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n522), .B(new_n517), .C1(new_n525), .C2(new_n528), .ZN(new_n529));
  OAI21_X1  g0329(.A(KEYINPUT89), .B1(new_n529), .B2(G190), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n306), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n518), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n491), .A2(new_n503), .A3(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT90), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n502), .B1(new_n487), .B2(new_n490), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n536), .A2(KEYINPUT90), .A3(new_n532), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  AND3_X1   g0338(.A1(new_n477), .A2(new_n482), .A3(new_n485), .ZN(new_n539));
  NOR3_X1   g0339(.A1(new_n539), .A2(new_n488), .A3(new_n489), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n483), .A2(KEYINPUT86), .A3(new_n489), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(new_n284), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n503), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(KEYINPUT88), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT88), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n536), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n529), .A2(G169), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n547), .B1(new_n278), .B2(new_n529), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n544), .A2(new_n546), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n538), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n402), .A2(new_n212), .A3(G68), .ZN(new_n551));
  INV_X1    g0351(.A(G97), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n292), .A2(new_n552), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n551), .B1(KEYINPUT19), .B2(new_n553), .ZN(new_n554));
  NOR2_X1   g0354(.A1(G87), .A2(G97), .ZN(new_n555));
  NAND3_X1  g0355(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n270), .A2(new_n555), .B1(new_n212), .B2(new_n556), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n284), .B1(new_n554), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n291), .A2(new_n282), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n558), .B(new_n559), .C1(new_n501), .C2(new_n291), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n371), .A2(new_n267), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n218), .A2(G1698), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n561), .B(new_n562), .C1(new_n257), .C2(new_n258), .ZN(new_n563));
  NAND2_X1  g0363(.A1(G33), .A2(G116), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n276), .A2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT82), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n244), .A2(G45), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(G250), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n567), .B1(new_n509), .B2(new_n569), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n249), .A2(KEYINPUT82), .A3(G250), .A4(new_n568), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n398), .A2(new_n511), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n566), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n417), .ZN(new_n575));
  AOI22_X1  g0375(.A1(new_n276), .A2(new_n565), .B1(new_n398), .B2(new_n511), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n576), .A2(new_n278), .A3(new_n572), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n560), .A2(new_n575), .A3(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n566), .A2(new_n572), .A3(new_n573), .A4(G190), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(KEYINPUT83), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT83), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n576), .A2(new_n582), .A3(G190), .A4(new_n572), .ZN(new_n583));
  AOI21_X1  g0383(.A(KEYINPUT84), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n306), .B1(new_n576), .B2(new_n572), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n499), .A2(G87), .A3(new_n361), .A4(new_n500), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n558), .A2(new_n586), .A3(new_n559), .ZN(new_n587));
  NOR3_X1   g0387(.A1(new_n584), .A2(new_n585), .A3(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n581), .A2(KEYINPUT84), .A3(new_n583), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n579), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n220), .A2(G1698), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n402), .B(new_n591), .C1(G257), .C2(G1698), .ZN(new_n592));
  INV_X1    g0392(.A(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(G303), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n594), .B1(new_n259), .B2(new_n264), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n276), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n521), .A2(G270), .A3(new_n249), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT85), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n597), .A2(new_n598), .A3(new_n517), .ZN(new_n599));
  INV_X1    g0399(.A(new_n599), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n598), .B1(new_n597), .B2(new_n517), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n596), .B(G190), .C1(new_n600), .C2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(G33), .A2(G283), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n603), .B(new_n212), .C1(G33), .C2(new_n552), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n479), .A2(G20), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n604), .A2(new_n284), .A3(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT20), .ZN(new_n607));
  XNOR2_X1  g0407(.A(new_n606), .B(new_n607), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n479), .B1(new_n244), .B2(G33), .ZN(new_n609));
  AOI22_X1  g0409(.A1(new_n285), .A2(new_n609), .B1(new_n479), .B2(new_n282), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n597), .A2(new_n517), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(KEYINPUT85), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n265), .A2(G303), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n592), .ZN(new_n616));
  AOI22_X1  g0416(.A1(new_n614), .A2(new_n599), .B1(new_n616), .B2(new_n276), .ZN(new_n617));
  OAI211_X1 g0417(.A(new_n602), .B(new_n612), .C1(new_n617), .C2(new_n306), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n617), .A2(G179), .A3(new_n611), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n596), .B1(new_n600), .B2(new_n601), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n417), .B1(new_n608), .B2(new_n610), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT21), .ZN(new_n622));
  AND3_X1   g0422(.A1(new_n620), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n622), .B1(new_n620), .B2(new_n621), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n618), .B(new_n619), .C1(new_n623), .C2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  AND2_X1   g0426(.A1(G97), .A2(G107), .ZN(new_n627));
  NOR2_X1   g0427(.A1(G97), .A2(G107), .ZN(new_n628));
  OAI22_X1  g0428(.A1(new_n627), .A2(new_n628), .B1(KEYINPUT81), .B2(KEYINPUT6), .ZN(new_n629));
  NOR2_X1   g0429(.A1(KEYINPUT81), .A2(KEYINPUT6), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n630), .B1(KEYINPUT6), .B2(new_n552), .ZN(new_n631));
  XNOR2_X1  g0431(.A(G97), .B(G107), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n629), .B(G20), .C1(new_n631), .C2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n295), .A2(G77), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n636), .B1(new_n438), .B2(new_n270), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(new_n284), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n361), .A2(G97), .ZN(new_n639));
  AND3_X1   g0439(.A1(new_n499), .A2(new_n361), .A3(new_n500), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n639), .B1(new_n640), .B2(G97), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n521), .A2(new_n249), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n517), .B1(new_n642), .B2(new_n504), .ZN(new_n643));
  OAI211_X1 g0443(.A(G244), .B(new_n267), .C1(new_n257), .C2(new_n258), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT4), .ZN(new_n645));
  AOI22_X1  g0445(.A1(new_n644), .A2(new_n645), .B1(G33), .B2(G283), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n645), .A2(new_n218), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n259), .A2(new_n264), .A3(new_n267), .A4(new_n647), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n259), .A2(new_n264), .A3(G250), .A4(G1698), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n646), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n643), .B1(new_n650), .B2(new_n276), .ZN(new_n651));
  AOI22_X1  g0451(.A1(new_n638), .A2(new_n641), .B1(new_n278), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n650), .A2(new_n276), .ZN(new_n653));
  INV_X1    g0453(.A(new_n643), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(new_n417), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n651), .A2(new_n516), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n657), .B1(G200), .B2(new_n651), .ZN(new_n658));
  INV_X1    g0458(.A(new_n639), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n659), .B1(new_n501), .B2(new_n552), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n660), .B1(new_n637), .B2(new_n284), .ZN(new_n661));
  AOI22_X1  g0461(.A1(new_n652), .A2(new_n656), .B1(new_n658), .B2(new_n661), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n590), .A2(new_n626), .A3(new_n662), .ZN(new_n663));
  NOR3_X1   g0463(.A1(new_n471), .A2(new_n550), .A3(new_n663), .ZN(G372));
  INV_X1    g0464(.A(new_n328), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n455), .A2(new_n464), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n370), .A2(new_n385), .A3(new_n386), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(new_n302), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n394), .A2(new_n388), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n666), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n447), .A2(new_n468), .ZN(new_n671));
  OR2_X1    g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n337), .A2(new_n342), .A3(KEYINPUT92), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  AOI21_X1  g0474(.A(KEYINPUT92), .B1(new_n337), .B2(new_n342), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n665), .B1(new_n672), .B2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n471), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n581), .A2(new_n583), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT84), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n587), .A2(new_n585), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n681), .A2(new_n589), .A3(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n270), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n635), .B1(new_n459), .B2(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n641), .B1(new_n685), .B2(new_n299), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n651), .A2(new_n278), .ZN(new_n687));
  AND3_X1   g0487(.A1(new_n686), .A2(new_n656), .A3(new_n687), .ZN(new_n688));
  XNOR2_X1  g0488(.A(KEYINPUT91), .B(KEYINPUT26), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n683), .A2(new_n688), .A3(new_n578), .A4(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT26), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n682), .A2(new_n679), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(new_n578), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n686), .A2(new_n656), .A3(new_n687), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n692), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n691), .A2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(new_n694), .ZN(new_n698));
  INV_X1    g0498(.A(new_n537), .ZN(new_n699));
  AOI21_X1  g0499(.A(KEYINPUT90), .B1(new_n536), .B2(new_n532), .ZN(new_n700));
  OAI211_X1 g0500(.A(new_n662), .B(new_n698), .C1(new_n699), .C2(new_n700), .ZN(new_n701));
  AND2_X1   g0501(.A1(new_n543), .A2(new_n548), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n619), .B1(new_n623), .B2(new_n624), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  OAI211_X1 g0504(.A(new_n578), .B(new_n697), .C1(new_n701), .C2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n678), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n677), .A2(new_n706), .ZN(G369));
  NAND2_X1  g0507(.A1(new_n493), .A2(new_n212), .ZN(new_n708));
  OR2_X1    g0508(.A1(new_n708), .A2(KEYINPUT27), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(KEYINPUT27), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n709), .A2(G213), .A3(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(G343), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n611), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n626), .A2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n703), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n715), .B1(new_n716), .B2(new_n714), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(G330), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  AND2_X1   g0519(.A1(new_n544), .A2(new_n546), .ZN(new_n720));
  AND2_X1   g0520(.A1(new_n720), .A2(new_n713), .ZN(new_n721));
  INV_X1    g0521(.A(new_n713), .ZN(new_n722));
  OAI22_X1  g0522(.A1(new_n721), .A2(new_n550), .B1(new_n549), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n719), .A2(new_n723), .ZN(new_n724));
  XOR2_X1   g0524(.A(new_n713), .B(KEYINPUT93), .Z(new_n725));
  NAND2_X1  g0525(.A1(new_n702), .A2(new_n725), .ZN(new_n726));
  AND2_X1   g0526(.A1(new_n538), .A2(new_n549), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n716), .A2(new_n713), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n724), .A2(new_n726), .A3(new_n729), .ZN(G399));
  INV_X1    g0530(.A(new_n208), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n731), .A2(G41), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n270), .A2(new_n479), .A3(new_n555), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n733), .A2(G1), .A3(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n736), .B1(new_n216), .B2(new_n733), .ZN(new_n737));
  XNOR2_X1  g0537(.A(new_n737), .B(KEYINPUT28), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n701), .B1(new_n549), .B2(new_n716), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n690), .B1(new_n590), .B2(new_n688), .ZN(new_n740));
  NOR3_X1   g0540(.A1(new_n694), .A2(new_n695), .A3(new_n692), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n578), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  OAI211_X1 g0542(.A(KEYINPUT29), .B(new_n722), .C1(new_n739), .C2(new_n742), .ZN(new_n743));
  AND2_X1   g0543(.A1(new_n705), .A2(new_n725), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n743), .B1(new_n744), .B2(KEYINPUT29), .ZN(new_n745));
  OAI211_X1 g0545(.A(G179), .B(new_n522), .C1(new_n525), .C2(new_n528), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n574), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n617), .A2(new_n747), .A3(new_n651), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT30), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n617), .A2(new_n747), .A3(KEYINPUT30), .A4(new_n651), .ZN(new_n751));
  AOI21_X1  g0551(.A(G179), .B1(new_n514), .B2(new_n517), .ZN(new_n752));
  NAND4_X1  g0552(.A1(new_n655), .A2(new_n752), .A3(new_n620), .A4(new_n574), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n750), .A2(new_n751), .A3(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(new_n713), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT31), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n725), .A2(new_n756), .ZN(new_n757));
  AOI22_X1  g0557(.A1(new_n755), .A2(new_n756), .B1(new_n754), .B2(new_n757), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n538), .A2(new_n549), .A3(new_n725), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n758), .B1(new_n759), .B2(new_n663), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(G330), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n745), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n738), .B1(new_n763), .B2(G1), .ZN(G364));
  NOR2_X1   g0564(.A1(new_n717), .A2(G330), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n281), .A2(G20), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n244), .B1(new_n766), .B2(G45), .ZN(new_n767));
  AOI211_X1 g0567(.A(new_n765), .B(new_n719), .C1(new_n733), .C2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n767), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n732), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  OAI21_X1  g0571(.A(G20), .B1(KEYINPUT94), .B2(G169), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(KEYINPUT94), .A2(G169), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n211), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(G179), .A2(G200), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n212), .B1(new_n777), .B2(G190), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(new_n552), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n212), .A2(new_n278), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(G200), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(new_n516), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(new_n202), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n781), .A2(G190), .ZN(new_n785));
  AOI211_X1 g0585(.A(new_n779), .B(new_n784), .C1(G68), .C2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(KEYINPUT96), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n787), .B1(new_n212), .B2(G190), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n516), .A2(KEYINPUT96), .A3(G20), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n788), .A2(new_n789), .A3(new_n777), .ZN(new_n790));
  INV_X1    g0590(.A(G159), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  XNOR2_X1  g0592(.A(new_n792), .B(KEYINPUT32), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n780), .A2(new_n516), .A3(new_n306), .ZN(new_n794));
  AND2_X1   g0594(.A1(new_n794), .A2(KEYINPUT95), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n794), .A2(KEYINPUT95), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(G77), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n212), .A2(new_n516), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n800), .A2(G179), .A3(new_n306), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n306), .A2(G179), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  OAI22_X1  g0603(.A1(new_n801), .A2(new_n425), .B1(new_n803), .B2(new_n472), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n788), .A2(new_n789), .A3(new_n802), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n805), .A2(new_n219), .ZN(new_n806));
  NOR3_X1   g0606(.A1(new_n804), .A2(new_n806), .A3(new_n265), .ZN(new_n807));
  NAND4_X1  g0607(.A1(new_n786), .A2(new_n793), .A3(new_n799), .A4(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(G317), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(KEYINPUT33), .ZN(new_n810));
  OR2_X1    g0610(.A1(new_n809), .A2(KEYINPUT33), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n785), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n801), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n266), .B1(G322), .B2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n778), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n782), .A2(G326), .B1(G294), .B2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n805), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(G283), .ZN(new_n818));
  AND4_X1   g0618(.A1(new_n812), .A2(new_n814), .A3(new_n816), .A4(new_n818), .ZN(new_n819));
  XNOR2_X1  g0619(.A(new_n803), .B(KEYINPUT97), .ZN(new_n820));
  AOI22_X1  g0620(.A1(new_n798), .A2(G311), .B1(G303), .B2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n790), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n822), .A2(G329), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n819), .A2(new_n821), .A3(new_n823), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n776), .B1(new_n808), .B2(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(G13), .A2(G33), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n827), .A2(G20), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n775), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n266), .A2(G355), .A3(new_n208), .ZN(new_n830));
  AND2_X1   g0630(.A1(new_n242), .A2(G45), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n731), .A2(new_n402), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n832), .B1(G45), .B2(new_n216), .ZN(new_n833));
  OAI221_X1 g0633(.A(new_n830), .B1(G116), .B2(new_n208), .C1(new_n831), .C2(new_n833), .ZN(new_n834));
  AOI211_X1 g0634(.A(new_n771), .B(new_n825), .C1(new_n829), .C2(new_n834), .ZN(new_n835));
  XNOR2_X1  g0635(.A(new_n828), .B(KEYINPUT98), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n835), .B1(new_n717), .B2(new_n836), .ZN(new_n837));
  XNOR2_X1  g0637(.A(new_n837), .B(KEYINPUT99), .ZN(new_n838));
  OR2_X1    g0638(.A1(new_n768), .A2(new_n838), .ZN(G396));
  NOR2_X1   g0639(.A1(new_n775), .A2(new_n826), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n771), .B1(new_n840), .B2(new_n203), .ZN(new_n841));
  OAI22_X1  g0641(.A1(new_n783), .A2(new_n594), .B1(new_n778), .B2(new_n552), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n265), .B1(new_n507), .B2(new_n801), .ZN(new_n843));
  AND2_X1   g0643(.A1(new_n785), .A2(KEYINPUT100), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n785), .A2(KEYINPUT100), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(new_n847));
  AOI211_X1 g0647(.A(new_n842), .B(new_n843), .C1(new_n847), .C2(G283), .ZN(new_n848));
  INV_X1    g0648(.A(new_n820), .ZN(new_n849));
  OAI22_X1  g0649(.A1(new_n849), .A2(new_n219), .B1(new_n472), .B2(new_n805), .ZN(new_n850));
  INV_X1    g0650(.A(G311), .ZN(new_n851));
  OAI22_X1  g0651(.A1(new_n797), .A2(new_n479), .B1(new_n851), .B2(new_n790), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  AOI22_X1  g0653(.A1(G137), .A2(new_n782), .B1(new_n813), .B2(G143), .ZN(new_n854));
  INV_X1    g0654(.A(new_n785), .ZN(new_n855));
  OAI221_X1 g0655(.A(new_n854), .B1(new_n323), .B2(new_n855), .C1(new_n797), .C2(new_n791), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT34), .ZN(new_n857));
  OR2_X1    g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n431), .B1(new_n815), .B2(G58), .ZN(new_n859));
  AOI22_X1  g0659(.A1(G68), .A2(new_n817), .B1(new_n822), .B2(G132), .ZN(new_n860));
  OAI211_X1 g0660(.A(new_n859), .B(new_n860), .C1(new_n849), .C2(new_n202), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n861), .B1(new_n856), .B2(new_n857), .ZN(new_n862));
  AOI22_X1  g0662(.A1(new_n848), .A2(new_n853), .B1(new_n858), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n300), .A2(new_n713), .ZN(new_n864));
  INV_X1    g0664(.A(new_n301), .ZN(new_n865));
  AOI22_X1  g0665(.A1(new_n307), .A2(new_n864), .B1(new_n865), .B2(new_n279), .ZN(new_n866));
  NOR3_X1   g0666(.A1(new_n280), .A2(new_n301), .A3(new_n713), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  OAI221_X1 g0668(.A(new_n841), .B1(new_n776), .B2(new_n863), .C1(new_n868), .C2(new_n827), .ZN(new_n869));
  INV_X1    g0669(.A(new_n725), .ZN(new_n870));
  NOR3_X1   g0670(.A1(new_n866), .A2(new_n870), .A3(new_n867), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n705), .A2(new_n871), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n872), .B1(new_n744), .B2(new_n868), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n770), .B1(new_n873), .B2(new_n761), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n873), .A2(new_n761), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n869), .B1(new_n875), .B2(new_n876), .ZN(G384));
  OAI21_X1  g0677(.A(new_n629), .B1(new_n631), .B2(new_n632), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT35), .ZN(new_n879));
  OAI211_X1 g0679(.A(G116), .B(new_n213), .C1(new_n878), .C2(new_n879), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n880), .B1(new_n879), .B2(new_n878), .ZN(new_n881));
  XNOR2_X1  g0681(.A(new_n881), .B(KEYINPUT36), .ZN(new_n882));
  OR3_X1    g0682(.A1(new_n216), .A2(new_n203), .A3(new_n426), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n202), .A2(G68), .ZN(new_n884));
  AOI211_X1 g0684(.A(new_n244), .B(G13), .C1(new_n883), .C2(new_n884), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n882), .A2(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n440), .B1(new_n443), .B2(new_n429), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n457), .A2(new_n318), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(new_n462), .ZN(new_n889));
  INV_X1    g0689(.A(new_n711), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n469), .A2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(new_n889), .ZN(new_n894));
  OAI211_X1 g0694(.A(new_n463), .B(new_n891), .C1(new_n894), .C2(new_n419), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(KEYINPUT37), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n465), .A2(new_n466), .A3(new_n408), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT37), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n466), .A2(new_n890), .ZN(new_n899));
  NAND4_X1  g0699(.A1(new_n897), .A2(new_n898), .A3(new_n463), .A4(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n896), .A2(new_n900), .ZN(new_n901));
  AND3_X1   g0701(.A1(new_n893), .A2(KEYINPUT38), .A3(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(KEYINPUT38), .B1(new_n893), .B2(new_n901), .ZN(new_n903));
  OR2_X1    g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  OAI211_X1 g0704(.A(new_n388), .B(new_n713), .C1(new_n387), .C2(new_n394), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n388), .A2(new_n713), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n669), .A2(new_n667), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(new_n867), .ZN(new_n909));
  AOI21_X1  g0709(.A(KEYINPUT101), .B1(new_n872), .B2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT101), .ZN(new_n911));
  AOI211_X1 g0711(.A(new_n911), .B(new_n867), .C1(new_n705), .C2(new_n871), .ZN(new_n912));
  OAI211_X1 g0712(.A(new_n904), .B(new_n908), .C1(new_n910), .C2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n671), .A2(new_n711), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n913), .A2(KEYINPUT102), .A3(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT38), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n446), .A2(new_n711), .ZN(new_n917));
  AND2_X1   g0717(.A1(new_n469), .A2(new_n917), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n898), .B1(new_n899), .B2(KEYINPUT103), .ZN(new_n919));
  NAND4_X1  g0719(.A1(new_n919), .A2(new_n897), .A3(new_n463), .A4(new_n899), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT103), .ZN(new_n921));
  OAI21_X1  g0721(.A(KEYINPUT37), .B1(new_n917), .B2(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n897), .A2(new_n463), .A3(new_n899), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n920), .A2(new_n924), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n916), .B1(new_n918), .B2(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n893), .A2(KEYINPUT38), .A3(new_n901), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT39), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n902), .A2(new_n903), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(KEYINPUT39), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n669), .A2(new_n713), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n930), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n915), .A2(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(KEYINPUT102), .B1(new_n913), .B2(new_n914), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  OAI211_X1 g0739(.A(new_n743), .B(new_n678), .C1(new_n744), .C2(KEYINPUT29), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(new_n677), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n939), .B(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(G330), .ZN(new_n943));
  AND2_X1   g0743(.A1(new_n905), .A2(new_n907), .ZN(new_n944));
  INV_X1    g0744(.A(new_n868), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  AOI21_X1  g0746(.A(KEYINPUT31), .B1(new_n754), .B2(new_n713), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT104), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n754), .A2(KEYINPUT31), .A3(new_n713), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n947), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND4_X1  g0750(.A1(new_n754), .A2(KEYINPUT104), .A3(KEYINPUT31), .A4(new_n713), .ZN(new_n951));
  OAI211_X1 g0751(.A(new_n950), .B(new_n951), .C1(new_n663), .C2(new_n759), .ZN(new_n952));
  NAND4_X1  g0752(.A1(new_n928), .A2(new_n946), .A3(KEYINPUT40), .A4(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT40), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n759), .A2(new_n663), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n949), .A2(new_n948), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n755), .A2(new_n756), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n956), .A2(new_n957), .A3(new_n951), .ZN(new_n958));
  OAI211_X1 g0758(.A(new_n908), .B(new_n868), .C1(new_n955), .C2(new_n958), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n954), .B1(new_n931), .B2(new_n959), .ZN(new_n960));
  AND2_X1   g0760(.A1(new_n953), .A2(new_n960), .ZN(new_n961));
  AND4_X1   g0761(.A1(new_n626), .A2(new_n662), .A3(new_n578), .A4(new_n683), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n727), .A2(new_n962), .A3(new_n725), .ZN(new_n963));
  INV_X1    g0763(.A(new_n958), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n471), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n943), .B1(new_n961), .B2(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n966), .B1(new_n965), .B2(new_n961), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n942), .A2(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n244), .B2(new_n766), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n942), .A2(new_n967), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n886), .B1(new_n969), .B2(new_n970), .ZN(G367));
  NOR2_X1   g0771(.A1(new_n778), .A2(new_n346), .ZN(new_n972));
  OAI221_X1 g0772(.A(new_n266), .B1(new_n425), .B2(new_n803), .C1(new_n323), .C2(new_n801), .ZN(new_n973));
  AOI211_X1 g0773(.A(new_n972), .B(new_n973), .C1(G143), .C2(new_n782), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n974), .B1(new_n791), .B2(new_n846), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n817), .A2(G77), .ZN(new_n976));
  INV_X1    g0776(.A(G137), .ZN(new_n977));
  OAI221_X1 g0777(.A(new_n976), .B1(new_n977), .B2(new_n790), .C1(new_n797), .C2(new_n202), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n820), .A2(KEYINPUT46), .A3(G116), .ZN(new_n979));
  AOI22_X1  g0779(.A1(G97), .A2(new_n817), .B1(new_n822), .B2(G317), .ZN(new_n980));
  INV_X1    g0780(.A(G283), .ZN(new_n981));
  OAI211_X1 g0781(.A(new_n979), .B(new_n980), .C1(new_n981), .C2(new_n797), .ZN(new_n982));
  INV_X1    g0782(.A(new_n803), .ZN(new_n983));
  AOI21_X1  g0783(.A(KEYINPUT46), .B1(new_n983), .B2(G116), .ZN(new_n984));
  OAI221_X1 g0784(.A(new_n431), .B1(new_n778), .B2(new_n270), .C1(new_n801), .C2(new_n594), .ZN(new_n985));
  AOI211_X1 g0785(.A(new_n984), .B(new_n985), .C1(G311), .C2(new_n782), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n986), .B1(new_n507), .B2(new_n846), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n975), .A2(new_n978), .B1(new_n982), .B2(new_n987), .ZN(new_n988));
  XOR2_X1   g0788(.A(KEYINPUT106), .B(KEYINPUT47), .Z(new_n989));
  XNOR2_X1  g0789(.A(new_n988), .B(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(new_n775), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n587), .A2(new_n713), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n578), .A2(new_n992), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n993), .B1(new_n698), .B2(new_n992), .ZN(new_n994));
  INV_X1    g0794(.A(new_n836), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(new_n832), .ZN(new_n997));
  OAI221_X1 g0797(.A(new_n829), .B1(new_n291), .B2(new_n208), .C1(new_n235), .C2(new_n997), .ZN(new_n998));
  NAND4_X1  g0798(.A1(new_n991), .A2(new_n770), .A3(new_n996), .A4(new_n998), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(KEYINPUT107), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n658), .A2(new_n661), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1002), .A2(new_n695), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n725), .A2(new_n661), .ZN(new_n1004));
  OAI22_X1  g0804(.A1(new_n1003), .A2(new_n1004), .B1(new_n695), .B2(new_n725), .ZN(new_n1005));
  XOR2_X1   g0805(.A(new_n1005), .B(KEYINPUT105), .Z(new_n1006));
  NOR2_X1   g0806(.A1(new_n1006), .A2(new_n729), .ZN(new_n1007));
  XOR2_X1   g0807(.A(new_n1007), .B(KEYINPUT42), .Z(new_n1008));
  OR2_X1    g0808(.A1(new_n1006), .A2(new_n549), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n870), .B1(new_n1009), .B2(new_n695), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT43), .ZN(new_n1011));
  OAI22_X1  g0811(.A1(new_n1008), .A2(new_n1010), .B1(new_n1011), .B2(new_n994), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n994), .A2(new_n1011), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1012), .B(new_n1013), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n724), .A2(new_n1006), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1014), .B(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n729), .A2(new_n726), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1006), .A2(new_n1017), .ZN(new_n1018));
  XOR2_X1   g0818(.A(new_n1018), .B(KEYINPUT44), .Z(new_n1019));
  NOR2_X1   g0819(.A1(new_n1006), .A2(new_n1017), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(KEYINPUT45), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n724), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n729), .B1(new_n723), .B2(new_n728), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1025), .B(new_n718), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n1026), .A2(new_n762), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1019), .A2(new_n724), .A3(new_n1021), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1024), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1029), .A2(new_n763), .ZN(new_n1030));
  XOR2_X1   g0830(.A(new_n732), .B(KEYINPUT41), .Z(new_n1031));
  INV_X1    g0831(.A(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n769), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1001), .B1(new_n1016), .B2(new_n1033), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT108), .ZN(G387));
  OR2_X1    g0835(.A1(new_n723), .A2(new_n836), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n832), .B1(new_n232), .B2(new_n510), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n266), .A2(new_n208), .A3(new_n734), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n294), .A2(G50), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(KEYINPUT109), .B(KEYINPUT50), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1040), .B(new_n1041), .ZN(new_n1042));
  AOI21_X1  g0842(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1042), .A2(new_n735), .A3(new_n1043), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n1039), .A2(new_n1044), .B1(new_n219), .B2(new_n731), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n829), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n770), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n402), .B1(new_n803), .B2(new_n203), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n791), .A2(new_n783), .B1(new_n855), .B2(new_n294), .ZN(new_n1049));
  AOI211_X1 g0849(.A(new_n1048), .B(new_n1049), .C1(G50), .C2(new_n813), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(G97), .A2(new_n817), .B1(new_n822), .B2(G150), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n798), .A2(G68), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n291), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1053), .A2(new_n815), .ZN(new_n1054));
  NAND4_X1  g0854(.A1(new_n1050), .A2(new_n1051), .A3(new_n1052), .A4(new_n1054), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n402), .B1(new_n822), .B2(G326), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n803), .A2(new_n507), .B1(new_n778), .B2(new_n981), .ZN(new_n1057));
  XOR2_X1   g0857(.A(KEYINPUT110), .B(G322), .Z(new_n1058));
  AOI22_X1  g0858(.A1(new_n782), .A2(new_n1058), .B1(new_n813), .B2(G317), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n1059), .B1(new_n594), .B2(new_n797), .C1(new_n846), .C2(new_n851), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT48), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1057), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1062), .B1(new_n1061), .B2(new_n1060), .ZN(new_n1063));
  INV_X1    g0863(.A(KEYINPUT49), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n1056), .B1(new_n479), .B2(new_n805), .C1(new_n1063), .C2(new_n1064), .ZN(new_n1065));
  AND2_X1   g0865(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1055), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1047), .B1(new_n1067), .B2(new_n775), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1036), .A2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1069), .B1(new_n1026), .B2(new_n767), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n1027), .A2(new_n733), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1026), .A2(new_n762), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1070), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1073), .ZN(G393));
  INV_X1    g0874(.A(new_n1028), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n724), .B1(new_n1019), .B2(new_n1021), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n1075), .A2(new_n1076), .B1(new_n762), .B2(new_n1026), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1077), .A2(new_n1029), .A3(new_n732), .ZN(new_n1078));
  OAI21_X1  g0878(.A(KEYINPUT111), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1079));
  INV_X1    g0879(.A(KEYINPUT111), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1024), .A2(new_n1080), .A3(new_n1028), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1079), .A2(new_n1081), .A3(new_n769), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1006), .A2(new_n828), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n797), .A2(new_n507), .ZN(new_n1084));
  AOI211_X1 g0884(.A(new_n806), .B(new_n1084), .C1(new_n822), .C2(new_n1058), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n783), .A2(new_n809), .B1(new_n851), .B2(new_n801), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(new_n1086), .B(KEYINPUT52), .ZN(new_n1087));
  OAI221_X1 g0887(.A(new_n265), .B1(new_n479), .B2(new_n778), .C1(new_n981), .C2(new_n803), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1088), .B1(new_n847), .B2(G303), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1085), .A2(new_n1087), .A3(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(KEYINPUT51), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n783), .A2(new_n323), .B1(new_n791), .B2(new_n801), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n847), .A2(G50), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  OAI221_X1 g0893(.A(new_n402), .B1(new_n778), .B2(new_n203), .C1(new_n346), .C2(new_n803), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1094), .B1(G87), .B2(new_n817), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n294), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n798), .A2(new_n1096), .B1(G143), .B2(new_n822), .ZN(new_n1097));
  OR2_X1    g0897(.A1(new_n1092), .A2(new_n1091), .ZN(new_n1098));
  NAND4_X1  g0898(.A1(new_n1093), .A2(new_n1095), .A3(new_n1097), .A4(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n776), .B1(new_n1090), .B2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n239), .A2(new_n832), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1046), .B1(G97), .B2(new_n731), .ZN(new_n1102));
  AOI211_X1 g0902(.A(new_n771), .B(new_n1100), .C1(new_n1101), .C2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1083), .A2(new_n1103), .ZN(new_n1104));
  AND3_X1   g0904(.A1(new_n1082), .A2(KEYINPUT112), .A3(new_n1104), .ZN(new_n1105));
  AOI21_X1  g0905(.A(KEYINPUT112), .B1(new_n1082), .B2(new_n1104), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1078), .B1(new_n1105), .B2(new_n1106), .ZN(G390));
  NAND2_X1  g0907(.A1(new_n930), .A2(new_n932), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(new_n826), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n840), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n770), .B1(new_n1110), .B2(new_n1096), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(G68), .A2(new_n817), .B1(new_n822), .B2(G294), .ZN(new_n1112));
  OAI221_X1 g0912(.A(new_n1112), .B1(new_n797), .B2(new_n552), .C1(new_n472), .C2(new_n849), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n266), .B1(G116), .B2(new_n813), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n782), .A2(G283), .B1(G77), .B2(new_n815), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n1114), .B(new_n1115), .C1(new_n846), .C2(new_n270), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n265), .B1(G132), .B2(new_n813), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n782), .A2(G128), .B1(G159), .B2(new_n815), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n1117), .B(new_n1118), .C1(new_n846), .C2(new_n977), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n803), .A2(new_n323), .ZN(new_n1120));
  XNOR2_X1  g0920(.A(new_n1120), .B(KEYINPUT53), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(G50), .A2(new_n817), .B1(new_n822), .B2(G125), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(KEYINPUT54), .B(G143), .ZN(new_n1123));
  XOR2_X1   g0923(.A(new_n1123), .B(KEYINPUT116), .Z(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(new_n1125));
  OAI211_X1 g0925(.A(new_n1121), .B(new_n1122), .C1(new_n1125), .C2(new_n797), .ZN(new_n1126));
  OAI22_X1  g0926(.A1(new_n1113), .A2(new_n1116), .B1(new_n1119), .B2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1111), .B1(new_n1127), .B2(new_n775), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1109), .A2(new_n1128), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n908), .B1(new_n910), .B2(new_n912), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n933), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(new_n1108), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n928), .A2(new_n1131), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n866), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n722), .B(new_n1135), .C1(new_n739), .C2(new_n742), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(new_n909), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1134), .B1(new_n908), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  NAND4_X1  g0939(.A1(new_n908), .A2(G330), .A3(new_n760), .A4(new_n868), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1133), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n943), .B1(new_n964), .B2(new_n963), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1142), .A2(new_n868), .A3(new_n908), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n1130), .A2(new_n1131), .B1(new_n930), .B2(new_n932), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1144), .B1(new_n1145), .B2(new_n1138), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1141), .A2(new_n1146), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1129), .B1(new_n1147), .B2(new_n767), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT117), .ZN(new_n1149));
  OR2_X1    g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(KEYINPUT115), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n760), .A2(new_n868), .A3(G330), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1152), .A2(new_n944), .ZN(new_n1153));
  INV_X1    g0953(.A(KEYINPUT113), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1152), .A2(KEYINPUT113), .A3(new_n944), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1155), .A2(new_n1143), .A3(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n910), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n912), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT114), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n1161), .B(G330), .C1(new_n955), .C2(new_n958), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1162), .A2(new_n868), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1161), .B1(new_n952), .B2(G330), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n944), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  AND3_X1   g0965(.A1(new_n1136), .A2(new_n1140), .A3(new_n909), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n1157), .A2(new_n1160), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n678), .A2(new_n1142), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n940), .A2(new_n677), .A3(new_n1168), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1151), .B1(new_n1167), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1169), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(new_n1154), .A2(new_n1153), .B1(new_n946), .B2(new_n1142), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n1172), .A2(new_n1156), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1136), .A2(new_n1140), .A3(new_n909), .ZN(new_n1174));
  OAI21_X1  g0974(.A(G330), .B1(new_n955), .B2(new_n958), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1175), .A2(KEYINPUT114), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1176), .A2(new_n868), .A3(new_n1162), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1174), .B1(new_n1177), .B2(new_n944), .ZN(new_n1178));
  OAI211_X1 g0978(.A(KEYINPUT115), .B(new_n1171), .C1(new_n1173), .C2(new_n1178), .ZN(new_n1179));
  AND2_X1   g0979(.A1(new_n1170), .A2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1180), .A2(new_n1147), .ZN(new_n1181));
  AND2_X1   g0981(.A1(new_n1141), .A2(new_n1146), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1170), .A2(new_n1179), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1181), .A2(new_n732), .A3(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1150), .A2(new_n1185), .A3(new_n1186), .ZN(G378));
  NOR2_X1   g0987(.A1(new_n402), .A2(G41), .ZN(new_n1188));
  INV_X1    g0988(.A(G41), .ZN(new_n1189));
  AOI211_X1 g0989(.A(G50), .B(new_n1188), .C1(new_n261), .C2(new_n1189), .ZN(new_n1190));
  OAI221_X1 g0990(.A(new_n1188), .B1(new_n203), .B2(new_n803), .C1(new_n219), .C2(new_n801), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1191), .B1(new_n798), .B2(new_n1053), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n782), .A2(G116), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n972), .B1(new_n785), .B2(G97), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(G58), .A2(new_n817), .B1(new_n822), .B2(G283), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n1192), .A2(new_n1193), .A3(new_n1194), .A4(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT58), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1190), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(G132), .A2(new_n785), .B1(new_n813), .B2(G128), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1199), .B1(new_n1125), .B2(new_n803), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n782), .A2(G125), .B1(G150), .B2(new_n815), .ZN(new_n1201));
  XOR2_X1   g1001(.A(new_n1201), .B(KEYINPUT118), .Z(new_n1202));
  AOI211_X1 g1002(.A(new_n1200), .B(new_n1202), .C1(G137), .C2(new_n798), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1203), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n1204), .A2(KEYINPUT59), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n261), .B(new_n1189), .C1(new_n805), .C2(new_n791), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1206), .B1(G124), .B2(new_n822), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT59), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1207), .B1(new_n1203), .B2(new_n1208), .ZN(new_n1209));
  OAI221_X1 g1009(.A(new_n1198), .B1(new_n1197), .B2(new_n1196), .C1(new_n1205), .C2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1210), .A2(new_n775), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n771), .B1(new_n840), .B2(new_n202), .ZN(new_n1212));
  XNOR2_X1  g1012(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n327), .A2(new_n890), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1215), .B1(new_n676), .B2(new_n328), .ZN(new_n1216));
  INV_X1    g1016(.A(KEYINPUT92), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n343), .A2(new_n1217), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1218), .A2(new_n328), .A3(new_n673), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1215), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1214), .B1(new_n1216), .B2(new_n1221), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n676), .A2(new_n328), .A3(new_n1215), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1223), .A2(new_n1224), .A3(new_n1213), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1222), .A2(new_n1225), .ZN(new_n1226));
  OAI211_X1 g1026(.A(new_n1211), .B(new_n1212), .C1(new_n1226), .C2(new_n827), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1226), .A2(G330), .A3(new_n960), .A4(new_n953), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n953), .A2(new_n960), .A3(G330), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1225), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1213), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1229), .A2(new_n1232), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n936), .A2(new_n938), .B1(new_n1228), .B2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1233), .A2(new_n1228), .ZN(new_n1235));
  NOR3_X1   g1035(.A1(new_n1235), .A2(new_n935), .A3(new_n937), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n1234), .A2(new_n1236), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1227), .B1(new_n1237), .B2(new_n767), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT57), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1169), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1240), .B1(new_n1241), .B2(new_n1237), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1171), .B1(new_n1180), .B2(new_n1147), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n936), .A2(new_n938), .A3(new_n1228), .A4(new_n1233), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1235), .B1(new_n937), .B2(new_n935), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1240), .B1(new_n1244), .B2(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n733), .B1(new_n1243), .B2(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT119), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1242), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1249));
  OAI21_X1  g1049(.A(KEYINPUT57), .B1(new_n1234), .B2(new_n1236), .ZN(new_n1250));
  OAI211_X1 g1050(.A(new_n1248), .B(new_n732), .C1(new_n1250), .C2(new_n1241), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1251), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1239), .B1(new_n1249), .B2(new_n1252), .ZN(G375));
  OAI21_X1  g1053(.A(new_n770), .B1(new_n1110), .B2(G68), .ZN(new_n1254));
  OAI22_X1  g1054(.A1(new_n849), .A2(new_n791), .B1(new_n797), .B2(new_n323), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1255), .B1(G128), .B2(new_n822), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n782), .A2(G132), .ZN(new_n1257));
  OAI221_X1 g1057(.A(new_n1257), .B1(new_n202), .B2(new_n778), .C1(new_n977), .C2(new_n801), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1258), .B1(new_n847), .B2(new_n1124), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n402), .B1(new_n805), .B2(new_n425), .ZN(new_n1260));
  XOR2_X1   g1060(.A(new_n1260), .B(KEYINPUT121), .Z(new_n1261));
  NAND3_X1  g1061(.A1(new_n1256), .A2(new_n1259), .A3(new_n1261), .ZN(new_n1262));
  OAI221_X1 g1062(.A(new_n265), .B1(new_n981), .B2(new_n801), .C1(new_n783), .C2(new_n507), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1263), .B1(new_n847), .B2(G116), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n798), .A2(new_n684), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1264), .A2(new_n976), .A3(new_n1054), .A4(new_n1265), .ZN(new_n1266));
  AOI22_X1  g1066(.A1(new_n820), .A2(G97), .B1(G303), .B2(new_n822), .ZN(new_n1267));
  XOR2_X1   g1067(.A(new_n1267), .B(KEYINPUT120), .Z(new_n1268));
  OAI21_X1  g1068(.A(new_n1262), .B1(new_n1266), .B2(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1254), .B1(new_n1269), .B2(new_n775), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1270), .B1(new_n908), .B2(new_n827), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1271), .B1(new_n1167), .B2(new_n767), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1167), .A2(new_n1169), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1180), .A2(new_n1274), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1273), .B1(new_n1275), .B2(new_n1031), .ZN(G381));
  INV_X1    g1076(.A(new_n1078), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1082), .A2(new_n1104), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT112), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1082), .A2(KEYINPUT112), .A3(new_n1104), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1277), .B1(new_n1280), .B2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(G384), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(G393), .A2(G396), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1282), .A2(new_n1283), .A3(new_n1284), .ZN(new_n1285));
  NOR3_X1   g1085(.A1(G387), .A2(G381), .A3(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT122), .ZN(new_n1287));
  XNOR2_X1  g1087(.A(new_n1286), .B(new_n1287), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n732), .B1(new_n1250), .B2(new_n1241), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1289), .A2(KEYINPUT119), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1290), .A2(new_n1251), .A3(new_n1242), .ZN(new_n1291));
  INV_X1    g1091(.A(G378), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1291), .A2(new_n1292), .A3(new_n1239), .ZN(new_n1293));
  OR2_X1    g1093(.A1(new_n1288), .A2(new_n1293), .ZN(G407));
  NAND2_X1  g1094(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1243), .A2(new_n1295), .ZN(new_n1296));
  AOI22_X1  g1096(.A1(new_n1289), .A2(KEYINPUT119), .B1(new_n1296), .B2(new_n1240), .ZN(new_n1297));
  AOI211_X1 g1097(.A(G378), .B(new_n1238), .C1(new_n1297), .C2(new_n1251), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1298), .A2(G213), .A3(new_n712), .ZN(new_n1299));
  OAI211_X1 g1099(.A(G213), .B(new_n1299), .C1(new_n1288), .C2(new_n1293), .ZN(G409));
  NAND2_X1  g1100(.A1(G375), .A2(G378), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n712), .A2(G213), .ZN(new_n1302));
  NAND4_X1  g1102(.A1(new_n1243), .A2(KEYINPUT123), .A3(new_n1032), .A4(new_n1295), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT123), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1304), .B1(new_n1296), .B2(new_n1031), .ZN(new_n1305));
  NAND4_X1  g1105(.A1(new_n1292), .A2(new_n1303), .A3(new_n1305), .A4(new_n1239), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT60), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n733), .B1(new_n1274), .B2(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1308), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1309), .B1(new_n1275), .B2(KEYINPUT60), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1283), .B1(new_n1310), .B2(new_n1272), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1307), .B1(new_n1180), .B2(new_n1274), .ZN(new_n1312));
  OAI211_X1 g1112(.A(G384), .B(new_n1273), .C1(new_n1312), .C2(new_n1309), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1311), .A2(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1314), .ZN(new_n1315));
  NAND4_X1  g1115(.A1(new_n1301), .A2(new_n1302), .A3(new_n1306), .A4(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1316), .A2(KEYINPUT62), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1306), .A2(new_n1302), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1292), .B1(new_n1291), .B2(new_n1239), .ZN(new_n1319));
  NOR2_X1   g1119(.A1(new_n1318), .A2(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT62), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1320), .A2(new_n1321), .A3(new_n1315), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT61), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n712), .A2(G213), .A3(G2897), .ZN(new_n1324));
  AND3_X1   g1124(.A1(new_n1311), .A2(new_n1313), .A3(new_n1324), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1324), .B1(new_n1311), .B2(new_n1313), .ZN(new_n1326));
  NOR2_X1   g1126(.A1(new_n1325), .A2(new_n1326), .ZN(new_n1327));
  OAI21_X1  g1127(.A(new_n1327), .B1(new_n1318), .B2(new_n1319), .ZN(new_n1328));
  NAND4_X1  g1128(.A1(new_n1317), .A2(new_n1322), .A3(new_n1323), .A4(new_n1328), .ZN(new_n1329));
  INV_X1    g1129(.A(G396), .ZN(new_n1330));
  NOR2_X1   g1130(.A1(new_n1073), .A2(new_n1330), .ZN(new_n1331));
  OAI21_X1  g1131(.A(KEYINPUT108), .B1(new_n1284), .B2(new_n1331), .ZN(new_n1332));
  OAI211_X1 g1132(.A(new_n1332), .B(new_n1078), .C1(new_n1105), .C2(new_n1106), .ZN(new_n1333));
  NOR2_X1   g1133(.A1(new_n1284), .A2(new_n1331), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n1333), .B1(new_n1282), .B2(new_n1334), .ZN(new_n1335));
  INV_X1    g1135(.A(new_n1034), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1335), .A2(new_n1336), .ZN(new_n1337));
  OAI211_X1 g1137(.A(new_n1034), .B(new_n1333), .C1(new_n1282), .C2(new_n1334), .ZN(new_n1338));
  AND3_X1   g1138(.A1(new_n1337), .A2(KEYINPUT126), .A3(new_n1338), .ZN(new_n1339));
  AOI21_X1  g1139(.A(KEYINPUT126), .B1(new_n1337), .B2(new_n1338), .ZN(new_n1340));
  NOR2_X1   g1140(.A1(new_n1339), .A2(new_n1340), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1329), .A2(new_n1341), .ZN(new_n1342));
  INV_X1    g1142(.A(new_n1338), .ZN(new_n1343));
  OAI21_X1  g1143(.A(G390), .B1(new_n1284), .B2(new_n1331), .ZN(new_n1344));
  AOI21_X1  g1144(.A(new_n1034), .B1(new_n1344), .B2(new_n1333), .ZN(new_n1345));
  NOR2_X1   g1145(.A1(new_n1343), .A2(new_n1345), .ZN(new_n1346));
  AND3_X1   g1146(.A1(new_n1328), .A2(new_n1346), .A3(new_n1323), .ZN(new_n1347));
  XNOR2_X1  g1147(.A(KEYINPUT124), .B(KEYINPUT63), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1316), .A2(new_n1348), .ZN(new_n1349));
  INV_X1    g1149(.A(KEYINPUT63), .ZN(new_n1350));
  OAI21_X1  g1150(.A(KEYINPUT125), .B1(new_n1316), .B2(new_n1350), .ZN(new_n1351));
  INV_X1    g1151(.A(KEYINPUT125), .ZN(new_n1352));
  NAND4_X1  g1152(.A1(new_n1320), .A2(new_n1352), .A3(KEYINPUT63), .A4(new_n1315), .ZN(new_n1353));
  NAND4_X1  g1153(.A1(new_n1347), .A2(new_n1349), .A3(new_n1351), .A4(new_n1353), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1342), .A2(new_n1354), .ZN(G405));
  INV_X1    g1155(.A(KEYINPUT127), .ZN(new_n1356));
  OAI21_X1  g1156(.A(new_n1356), .B1(new_n1298), .B2(new_n1319), .ZN(new_n1357));
  NAND3_X1  g1157(.A1(new_n1301), .A2(KEYINPUT127), .A3(new_n1293), .ZN(new_n1358));
  AND3_X1   g1158(.A1(new_n1357), .A2(new_n1358), .A3(new_n1314), .ZN(new_n1359));
  AOI21_X1  g1159(.A(new_n1314), .B1(new_n1357), .B2(new_n1358), .ZN(new_n1360));
  INV_X1    g1160(.A(KEYINPUT126), .ZN(new_n1361));
  OAI21_X1  g1161(.A(new_n1361), .B1(new_n1343), .B2(new_n1345), .ZN(new_n1362));
  NAND3_X1  g1162(.A1(new_n1337), .A2(KEYINPUT126), .A3(new_n1338), .ZN(new_n1363));
  NAND2_X1  g1163(.A1(new_n1362), .A2(new_n1363), .ZN(new_n1364));
  NOR3_X1   g1164(.A1(new_n1359), .A2(new_n1360), .A3(new_n1364), .ZN(new_n1365));
  NOR3_X1   g1165(.A1(new_n1298), .A2(new_n1319), .A3(new_n1356), .ZN(new_n1366));
  AOI21_X1  g1166(.A(KEYINPUT127), .B1(new_n1301), .B2(new_n1293), .ZN(new_n1367));
  OAI21_X1  g1167(.A(new_n1315), .B1(new_n1366), .B2(new_n1367), .ZN(new_n1368));
  NAND3_X1  g1168(.A1(new_n1357), .A2(new_n1358), .A3(new_n1314), .ZN(new_n1369));
  AOI21_X1  g1169(.A(new_n1341), .B1(new_n1368), .B2(new_n1369), .ZN(new_n1370));
  NOR2_X1   g1170(.A1(new_n1365), .A2(new_n1370), .ZN(G402));
endmodule


