//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 0 0 0 1 1 1 0 1 1 0 0 1 0 1 1 0 0 0 0 1 0 1 1 1 1 0 0 1 1 0 1 0 1 0 0 1 0 1 0 1 0 0 0 0 1 1 1 0 0 0 1 0 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:40 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n594, new_n596,
    new_n597, new_n598, new_n599, new_n600, new_n601, new_n602, new_n603,
    new_n604, new_n605, new_n606, new_n607, new_n608, new_n609, new_n610,
    new_n611, new_n612, new_n613, new_n614, new_n615, new_n616, new_n617,
    new_n618, new_n619, new_n620, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n659, new_n660, new_n661, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n713, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT6), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT76), .ZN(new_n189));
  INV_X1    g003(.A(G104), .ZN(new_n190));
  AOI22_X1  g004(.A1(new_n189), .A2(KEYINPUT3), .B1(new_n190), .B2(G107), .ZN(new_n191));
  OAI22_X1  g005(.A1(new_n189), .A2(KEYINPUT3), .B1(new_n190), .B2(G107), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT3), .ZN(new_n193));
  INV_X1    g007(.A(G107), .ZN(new_n194));
  NAND4_X1  g008(.A1(new_n193), .A2(new_n194), .A3(KEYINPUT76), .A4(G104), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n191), .A2(new_n192), .A3(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G101), .ZN(new_n197));
  INV_X1    g011(.A(G101), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n191), .A2(new_n192), .A3(new_n198), .A4(new_n195), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n197), .A2(KEYINPUT4), .A3(new_n199), .ZN(new_n200));
  XNOR2_X1  g014(.A(G116), .B(G119), .ZN(new_n201));
  OR2_X1    g015(.A1(KEYINPUT2), .A2(G113), .ZN(new_n202));
  NAND2_X1  g016(.A1(KEYINPUT2), .A2(G113), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G119), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G116), .ZN(new_n206));
  INV_X1    g020(.A(G116), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G119), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  XNOR2_X1  g023(.A(KEYINPUT2), .B(G113), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n204), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT67), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n204), .A2(new_n211), .A3(KEYINPUT67), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT4), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n196), .A2(new_n216), .A3(G101), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n200), .A2(new_n214), .A3(new_n215), .A4(new_n217), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n209), .A2(new_n210), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT5), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n220), .A2(new_n205), .A3(G116), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT81), .ZN(new_n222));
  XNOR2_X1  g036(.A(new_n221), .B(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G113), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n224), .B1(new_n201), .B2(KEYINPUT5), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n219), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n190), .A2(G107), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n194), .A2(G104), .ZN(new_n228));
  OAI21_X1  g042(.A(G101), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  AND2_X1   g043(.A1(new_n199), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n226), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n218), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT82), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n218), .A2(KEYINPUT82), .A3(new_n231), .ZN(new_n235));
  XNOR2_X1  g049(.A(G110), .B(G122), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  AND4_X1   g051(.A1(new_n188), .A2(new_n234), .A3(new_n235), .A4(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n218), .A2(new_n231), .A3(new_n236), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(KEYINPUT6), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n236), .B1(new_n232), .B2(new_n233), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n240), .B1(new_n241), .B2(new_n235), .ZN(new_n242));
  OAI21_X1  g056(.A(KEYINPUT83), .B1(new_n238), .B2(new_n242), .ZN(new_n243));
  XNOR2_X1  g057(.A(G143), .B(G146), .ZN(new_n244));
  NAND2_X1  g058(.A1(KEYINPUT0), .A2(G128), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  XOR2_X1   g060(.A(KEYINPUT0), .B(G128), .Z(new_n247));
  OAI21_X1  g061(.A(new_n246), .B1(new_n247), .B2(new_n244), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(G125), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT66), .ZN(new_n250));
  INV_X1    g064(.A(G146), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G143), .ZN(new_n252));
  INV_X1    g066(.A(G143), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G146), .ZN(new_n254));
  AOI21_X1  g068(.A(G128), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  AND3_X1   g069(.A1(new_n253), .A2(KEYINPUT1), .A3(G146), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n250), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n251), .A2(G143), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(KEYINPUT1), .ZN(new_n259));
  OAI211_X1 g073(.A(new_n259), .B(KEYINPUT66), .C1(new_n244), .C2(G128), .ZN(new_n260));
  INV_X1    g074(.A(G128), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n261), .A2(KEYINPUT1), .ZN(new_n262));
  AOI22_X1  g076(.A1(new_n257), .A2(new_n260), .B1(new_n244), .B2(new_n262), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n249), .B1(new_n263), .B2(G125), .ZN(new_n264));
  INV_X1    g078(.A(G224), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n264), .B1(new_n265), .B2(G953), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n265), .A2(G953), .ZN(new_n267));
  OAI211_X1 g081(.A(new_n249), .B(new_n267), .C1(new_n263), .C2(G125), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n241), .A2(new_n235), .ZN(new_n270));
  INV_X1    g084(.A(new_n240), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT83), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n243), .A2(new_n269), .A3(new_n274), .ZN(new_n275));
  OAI21_X1  g089(.A(G210), .B1(G237), .B2(G902), .ZN(new_n276));
  INV_X1    g090(.A(G902), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n199), .A2(new_n229), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n226), .B1(KEYINPUT84), .B2(new_n278), .ZN(new_n279));
  XNOR2_X1  g093(.A(new_n236), .B(KEYINPUT8), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NOR3_X1   g095(.A1(new_n226), .A2(KEYINPUT84), .A3(new_n278), .ZN(new_n282));
  OAI221_X1 g096(.A(new_n268), .B1(new_n264), .B2(KEYINPUT7), .C1(new_n281), .C2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT7), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n239), .B1(new_n266), .B2(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n277), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(KEYINPUT85), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT85), .ZN(new_n288));
  OAI211_X1 g102(.A(new_n288), .B(new_n277), .C1(new_n283), .C2(new_n285), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  AND3_X1   g104(.A1(new_n275), .A2(new_n276), .A3(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n276), .B1(new_n275), .B2(new_n290), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n187), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(G221), .ZN(new_n294));
  XOR2_X1   g108(.A(KEYINPUT9), .B(G234), .Z(new_n295));
  AOI21_X1  g109(.A(new_n294), .B1(new_n295), .B2(new_n277), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(G469), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n262), .A2(new_n252), .A3(new_n254), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n253), .A2(G146), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n261), .B1(new_n300), .B2(new_n258), .ZN(new_n301));
  AOI21_X1  g115(.A(KEYINPUT66), .B1(new_n301), .B2(new_n259), .ZN(new_n302));
  NOR3_X1   g116(.A1(new_n255), .A2(new_n250), .A3(new_n256), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n299), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n304), .A2(KEYINPUT10), .A3(new_n230), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n301), .A2(new_n299), .A3(new_n259), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n230), .A2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT10), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT64), .ZN(new_n310));
  INV_X1    g124(.A(G134), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n310), .B1(new_n311), .B2(G137), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(KEYINPUT11), .ZN(new_n313));
  INV_X1    g127(.A(G131), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT11), .ZN(new_n315));
  OAI211_X1 g129(.A(new_n310), .B(new_n315), .C1(new_n311), .C2(G137), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n311), .A2(G137), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n313), .A2(new_n314), .A3(new_n316), .A4(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT65), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  AOI22_X1  g134(.A1(new_n312), .A2(KEYINPUT11), .B1(new_n311), .B2(G137), .ZN(new_n321));
  NAND4_X1  g135(.A1(new_n321), .A2(KEYINPUT65), .A3(new_n314), .A4(new_n316), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n316), .ZN(new_n323));
  AOI22_X1  g137(.A1(new_n320), .A2(new_n322), .B1(new_n323), .B2(G131), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n200), .A2(new_n248), .A3(new_n217), .ZN(new_n325));
  NAND4_X1  g139(.A1(new_n305), .A2(new_n309), .A3(new_n324), .A4(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  OAI211_X1 g141(.A(new_n299), .B(new_n278), .C1(new_n302), .C2(new_n303), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(new_n307), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n320), .A2(new_n322), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n323), .A2(G131), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n329), .A2(KEYINPUT77), .A3(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT78), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n324), .B1(new_n307), .B2(new_n328), .ZN(new_n336));
  AOI22_X1  g150(.A1(new_n335), .A2(KEYINPUT12), .B1(KEYINPUT78), .B2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT12), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n333), .A2(new_n334), .A3(new_n338), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n327), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(G953), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(G227), .ZN(new_n342));
  XNOR2_X1  g156(.A(new_n342), .B(KEYINPUT75), .ZN(new_n343));
  XNOR2_X1  g157(.A(G110), .B(G140), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n343), .B(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  AND3_X1   g160(.A1(new_n306), .A2(new_n199), .A3(new_n229), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n199), .A2(KEYINPUT10), .A3(new_n229), .ZN(new_n348));
  OAI22_X1  g162(.A1(new_n347), .A2(KEYINPUT10), .B1(new_n263), .B2(new_n348), .ZN(new_n349));
  AND3_X1   g163(.A1(new_n200), .A2(new_n248), .A3(new_n217), .ZN(new_n350));
  OAI21_X1  g164(.A(KEYINPUT79), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT79), .ZN(new_n352));
  NAND4_X1  g166(.A1(new_n305), .A2(new_n309), .A3(new_n352), .A4(new_n325), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n351), .A2(new_n332), .A3(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n326), .A2(new_n346), .ZN(new_n356));
  OAI22_X1  g170(.A1(new_n340), .A2(new_n346), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n298), .B1(new_n357), .B2(new_n277), .ZN(new_n358));
  XOR2_X1   g172(.A(KEYINPUT80), .B(G469), .Z(new_n359));
  AOI21_X1  g173(.A(new_n356), .B1(new_n337), .B2(new_n339), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n346), .B1(new_n354), .B2(new_n326), .ZN(new_n361));
  OAI211_X1 g175(.A(new_n277), .B(new_n359), .C1(new_n360), .C2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n297), .B1(new_n358), .B2(new_n363), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n293), .A2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(G234), .ZN(new_n366));
  OAI21_X1  g180(.A(G217), .B1(new_n366), .B2(G902), .ZN(new_n367));
  XNOR2_X1  g181(.A(new_n367), .B(KEYINPUT70), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT71), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n369), .A2(new_n261), .A3(G119), .ZN(new_n370));
  AOI21_X1  g184(.A(KEYINPUT71), .B1(new_n205), .B2(G128), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n205), .A2(G128), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n370), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  XNOR2_X1  g187(.A(KEYINPUT24), .B(G110), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT72), .ZN(new_n376));
  XNOR2_X1  g190(.A(new_n375), .B(new_n376), .ZN(new_n377));
  XNOR2_X1  g191(.A(G125), .B(G140), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(KEYINPUT16), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT16), .ZN(new_n380));
  INV_X1    g194(.A(G140), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n380), .A2(new_n381), .A3(G125), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n379), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(new_n251), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n379), .A2(G146), .A3(new_n382), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  OAI21_X1  g200(.A(KEYINPUT23), .B1(new_n261), .B2(G119), .ZN(new_n387));
  OAI21_X1  g201(.A(KEYINPUT73), .B1(new_n205), .B2(G128), .ZN(new_n388));
  XOR2_X1   g202(.A(new_n387), .B(new_n388), .Z(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(G110), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n377), .A2(new_n386), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n373), .A2(new_n374), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n392), .B1(new_n389), .B2(G110), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n378), .A2(new_n251), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n393), .A2(new_n385), .A3(new_n394), .ZN(new_n395));
  XNOR2_X1  g209(.A(KEYINPUT22), .B(G137), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n341), .A2(G221), .A3(G234), .ZN(new_n397));
  XNOR2_X1  g211(.A(new_n396), .B(new_n397), .ZN(new_n398));
  AND3_X1   g212(.A1(new_n391), .A2(new_n395), .A3(new_n398), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n398), .B1(new_n391), .B2(new_n395), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(KEYINPUT25), .B1(new_n401), .B2(new_n277), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT25), .ZN(new_n403));
  NOR4_X1   g217(.A1(new_n399), .A2(new_n400), .A3(new_n403), .A4(G902), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n368), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  OR3_X1    g219(.A1(new_n399), .A2(new_n400), .A3(KEYINPUT74), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n368), .A2(G902), .ZN(new_n407));
  OAI21_X1  g221(.A(KEYINPUT74), .B1(new_n399), .B2(new_n400), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n405), .A2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT30), .ZN(new_n412));
  INV_X1    g226(.A(new_n317), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n311), .A2(G137), .ZN(new_n414));
  OAI21_X1  g228(.A(G131), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  AND3_X1   g229(.A1(new_n304), .A2(new_n330), .A3(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n248), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n417), .B1(new_n330), .B2(new_n331), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n412), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n214), .A2(new_n215), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n304), .A2(new_n330), .A3(new_n415), .ZN(new_n422));
  OAI211_X1 g236(.A(new_n422), .B(KEYINPUT30), .C1(new_n324), .C2(new_n417), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n419), .A2(new_n421), .A3(new_n423), .ZN(new_n424));
  OAI211_X1 g238(.A(new_n422), .B(new_n420), .C1(new_n324), .C2(new_n417), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(G237), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n427), .A2(new_n341), .A3(G210), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n428), .B(new_n198), .ZN(new_n429));
  XNOR2_X1  g243(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n430));
  XOR2_X1   g244(.A(new_n429), .B(new_n430), .Z(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  AOI21_X1  g246(.A(KEYINPUT29), .B1(new_n426), .B2(new_n432), .ZN(new_n433));
  NOR3_X1   g247(.A1(new_n416), .A2(new_n418), .A3(new_n421), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n332), .A2(new_n248), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n420), .B1(new_n435), .B2(new_n422), .ZN(new_n436));
  OAI211_X1 g250(.A(KEYINPUT68), .B(KEYINPUT28), .C1(new_n434), .C2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT28), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n421), .B1(new_n416), .B2(new_n418), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n438), .B1(new_n439), .B2(new_n425), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT68), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n441), .B1(new_n425), .B2(new_n438), .ZN(new_n442));
  OAI211_X1 g256(.A(new_n437), .B(new_n431), .C1(new_n440), .C2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n433), .A2(new_n443), .ZN(new_n444));
  AOI21_X1  g258(.A(KEYINPUT69), .B1(new_n439), .B2(new_n425), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT69), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n436), .A2(new_n446), .ZN(new_n447));
  OAI21_X1  g261(.A(KEYINPUT28), .B1(new_n445), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n425), .A2(new_n438), .ZN(new_n449));
  NAND4_X1  g263(.A1(new_n448), .A2(KEYINPUT29), .A3(new_n431), .A4(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n444), .A2(new_n277), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(G472), .ZN(new_n452));
  NOR2_X1   g266(.A1(G472), .A2(G902), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n424), .A2(new_n431), .A3(new_n425), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(KEYINPUT31), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT31), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n424), .A2(new_n456), .A3(new_n431), .A4(new_n425), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  OAI21_X1  g272(.A(KEYINPUT28), .B1(new_n434), .B2(new_n436), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n449), .A2(KEYINPUT68), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n431), .B1(new_n461), .B2(new_n437), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n453), .B1(new_n458), .B2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT32), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  OAI211_X1 g279(.A(KEYINPUT32), .B(new_n453), .C1(new_n458), .C2(new_n462), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n452), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(G478), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n468), .A2(KEYINPUT15), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  XNOR2_X1  g284(.A(G128), .B(G143), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n471), .B(new_n311), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n472), .B(KEYINPUT91), .ZN(new_n473));
  XNOR2_X1  g287(.A(KEYINPUT88), .B(G122), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n474), .A2(new_n207), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT14), .ZN(new_n476));
  OAI21_X1  g290(.A(G107), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(G122), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n478), .A2(G116), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n475), .A2(new_n479), .ZN(new_n480));
  OR2_X1    g294(.A1(new_n477), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n477), .A2(new_n480), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n473), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n480), .A2(new_n194), .ZN(new_n484));
  OAI21_X1  g298(.A(G107), .B1(new_n475), .B2(new_n479), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  XOR2_X1   g300(.A(KEYINPUT89), .B(KEYINPUT13), .Z(new_n487));
  OR3_X1    g301(.A1(new_n487), .A2(new_n261), .A3(G143), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n311), .B1(new_n487), .B2(new_n471), .ZN(new_n489));
  AOI22_X1  g303(.A1(new_n488), .A2(new_n489), .B1(new_n311), .B2(new_n471), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n486), .A2(new_n490), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n491), .A2(KEYINPUT90), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT90), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n493), .B1(new_n486), .B2(new_n490), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n483), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n295), .A2(G217), .A3(new_n341), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n496), .ZN(new_n498));
  OAI211_X1 g312(.A(new_n483), .B(new_n498), .C1(new_n492), .C2(new_n494), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n470), .B1(new_n500), .B2(new_n277), .ZN(new_n501));
  AOI211_X1 g315(.A(G902), .B(new_n469), .C1(new_n497), .C2(new_n499), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(G952), .ZN(new_n504));
  AOI211_X1 g318(.A(G953), .B(new_n504), .C1(G234), .C2(G237), .ZN(new_n505));
  XOR2_X1   g319(.A(KEYINPUT21), .B(G898), .Z(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  AOI211_X1 g321(.A(new_n277), .B(new_n341), .C1(G234), .C2(G237), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n505), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  NOR2_X1   g324(.A1(G475), .A2(G902), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n427), .A2(new_n341), .A3(G214), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n512), .B(G143), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT18), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n513), .B1(new_n514), .B2(new_n314), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n512), .B(new_n253), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n516), .A2(KEYINPUT18), .A3(G131), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n378), .B(new_n251), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n515), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT86), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n515), .A2(new_n517), .A3(KEYINPUT86), .A4(new_n518), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(new_n386), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n516), .A2(KEYINPUT17), .A3(G131), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n516), .A2(G131), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n513), .A2(new_n314), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  OAI211_X1 g342(.A(new_n524), .B(new_n525), .C1(KEYINPUT17), .C2(new_n528), .ZN(new_n529));
  XNOR2_X1  g343(.A(G113), .B(G122), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n530), .B(new_n190), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n523), .A2(new_n529), .A3(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  XOR2_X1   g347(.A(new_n378), .B(KEYINPUT19), .Z(new_n534));
  OAI21_X1  g348(.A(new_n385), .B1(new_n534), .B2(G146), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT87), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  OAI211_X1 g351(.A(KEYINPUT87), .B(new_n385), .C1(new_n534), .C2(G146), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n537), .A2(new_n528), .A3(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n531), .B1(new_n539), .B2(new_n523), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n511), .B1(new_n533), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(KEYINPUT20), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT20), .ZN(new_n543));
  OAI211_X1 g357(.A(new_n543), .B(new_n511), .C1(new_n533), .C2(new_n540), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n531), .B1(new_n523), .B2(new_n529), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n277), .B1(new_n533), .B2(new_n545), .ZN(new_n546));
  AOI22_X1  g360(.A1(new_n542), .A2(new_n544), .B1(G475), .B2(new_n546), .ZN(new_n547));
  AND3_X1   g361(.A1(new_n503), .A2(new_n510), .A3(new_n547), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n365), .A2(new_n411), .A3(new_n467), .A4(new_n548), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n549), .B(G101), .ZN(G3));
  OAI211_X1 g364(.A(new_n510), .B(new_n187), .C1(new_n291), .C2(new_n292), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n355), .A2(new_n356), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n335), .A2(KEYINPUT12), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n336), .A2(KEYINPUT78), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n554), .A2(new_n339), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(new_n326), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n553), .B1(new_n557), .B2(new_n345), .ZN(new_n558));
  OAI21_X1  g372(.A(G469), .B1(new_n558), .B2(G902), .ZN(new_n559));
  AOI211_X1 g373(.A(new_n296), .B(new_n410), .C1(new_n559), .C2(new_n362), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n277), .B1(new_n458), .B2(new_n462), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(G472), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(new_n463), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(G902), .B1(new_n497), .B2(new_n499), .ZN(new_n565));
  XNOR2_X1  g379(.A(KEYINPUT93), .B(G478), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT33), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT92), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n568), .B1(new_n499), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n500), .A2(new_n570), .ZN(new_n571));
  OAI211_X1 g385(.A(new_n497), .B(new_n499), .C1(new_n569), .C2(new_n568), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n468), .A2(G902), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n567), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n575), .A2(new_n547), .ZN(new_n576));
  NAND4_X1  g390(.A1(new_n552), .A2(new_n560), .A3(new_n564), .A4(new_n576), .ZN(new_n577));
  XOR2_X1   g391(.A(KEYINPUT34), .B(G104), .Z(new_n578));
  XNOR2_X1  g392(.A(new_n577), .B(new_n578), .ZN(G6));
  INV_X1    g393(.A(new_n503), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(new_n547), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n551), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n582), .A2(new_n564), .A3(new_n560), .ZN(new_n583));
  XOR2_X1   g397(.A(KEYINPUT35), .B(G107), .Z(new_n584));
  XNOR2_X1  g398(.A(new_n583), .B(new_n584), .ZN(G9));
  NAND2_X1  g399(.A1(new_n391), .A2(new_n395), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT36), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n398), .A2(new_n587), .ZN(new_n588));
  XOR2_X1   g402(.A(new_n586), .B(new_n588), .Z(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(new_n407), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n405), .A2(new_n590), .ZN(new_n591));
  AND3_X1   g405(.A1(new_n562), .A2(new_n463), .A3(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n365), .A2(new_n548), .A3(new_n592), .ZN(new_n593));
  XOR2_X1   g407(.A(KEYINPUT37), .B(G110), .Z(new_n594));
  XNOR2_X1  g408(.A(new_n593), .B(new_n594), .ZN(G12));
  INV_X1    g409(.A(KEYINPUT94), .ZN(new_n596));
  INV_X1    g410(.A(new_n187), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n275), .A2(new_n290), .ZN(new_n598));
  INV_X1    g412(.A(new_n276), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n275), .A2(new_n276), .A3(new_n290), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n597), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n296), .B1(new_n559), .B2(new_n362), .ZN(new_n603));
  NAND4_X1  g417(.A1(new_n467), .A2(new_n602), .A3(new_n603), .A4(new_n591), .ZN(new_n604));
  INV_X1    g418(.A(G900), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n505), .B1(new_n508), .B2(new_n605), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n581), .A2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n596), .B1(new_n604), .B2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n591), .ZN(new_n610));
  INV_X1    g424(.A(new_n466), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n440), .A2(new_n442), .ZN(new_n612));
  AOI211_X1 g426(.A(new_n441), .B(new_n438), .C1(new_n439), .C2(new_n425), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n432), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n614), .A2(new_n455), .A3(new_n457), .ZN(new_n615));
  AOI21_X1  g429(.A(KEYINPUT32), .B1(new_n615), .B2(new_n453), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n611), .A2(new_n616), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n610), .B1(new_n617), .B2(new_n452), .ZN(new_n618));
  NAND4_X1  g432(.A1(new_n618), .A2(KEYINPUT94), .A3(new_n365), .A4(new_n607), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n609), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n620), .B(G128), .ZN(G30));
  NAND2_X1  g435(.A1(new_n600), .A2(new_n601), .ZN(new_n622));
  XNOR2_X1  g436(.A(KEYINPUT95), .B(KEYINPUT38), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n622), .B(new_n623), .ZN(new_n624));
  NOR4_X1   g438(.A1(new_n624), .A2(new_n503), .A3(new_n547), .A4(new_n597), .ZN(new_n625));
  XOR2_X1   g439(.A(new_n606), .B(KEYINPUT39), .Z(new_n626));
  NAND2_X1  g440(.A1(new_n603), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(KEYINPUT40), .ZN(new_n628));
  NAND2_X1  g442(.A1(G472), .A2(G902), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n445), .A2(new_n447), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n630), .A2(new_n431), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n454), .A2(G472), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n629), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  XOR2_X1   g447(.A(new_n633), .B(KEYINPUT96), .Z(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(new_n617), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n636), .A2(new_n591), .ZN(new_n637));
  OR2_X1    g451(.A1(new_n627), .A2(KEYINPUT40), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n625), .A2(new_n628), .A3(new_n637), .A4(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(G143), .ZN(G45));
  INV_X1    g454(.A(new_n547), .ZN(new_n641));
  INV_X1    g455(.A(new_n606), .ZN(new_n642));
  AOI211_X1 g456(.A(new_n468), .B(G902), .C1(new_n571), .C2(new_n572), .ZN(new_n643));
  OAI211_X1 g457(.A(new_n641), .B(new_n642), .C1(new_n643), .C2(new_n567), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n604), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(new_n251), .ZN(G48));
  INV_X1    g460(.A(new_n356), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n556), .A2(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(new_n361), .ZN(new_n649));
  AOI21_X1  g463(.A(G902), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  OAI211_X1 g464(.A(new_n362), .B(new_n297), .C1(new_n650), .C2(new_n298), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n467), .A2(new_n411), .A3(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n602), .A2(new_n510), .A3(new_n576), .ZN(new_n654));
  OR2_X1    g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(KEYINPUT41), .B(G113), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(KEYINPUT97), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n655), .B(new_n657), .ZN(G15));
  NOR2_X1   g472(.A1(new_n641), .A2(new_n503), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n602), .A2(new_n510), .A3(new_n659), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n653), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(new_n207), .ZN(G18));
  NOR2_X1   g476(.A1(new_n293), .A2(new_n651), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n618), .A2(new_n548), .A3(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(G119), .ZN(G21));
  NAND2_X1  g479(.A1(new_n354), .A2(new_n326), .ZN(new_n666));
  AOI22_X1  g480(.A1(new_n556), .A2(new_n647), .B1(new_n666), .B2(new_n345), .ZN(new_n667));
  OAI21_X1  g481(.A(G469), .B1(new_n667), .B2(G902), .ZN(new_n668));
  AND4_X1   g482(.A1(new_n510), .A2(new_n668), .A3(new_n297), .A4(new_n362), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n431), .B1(new_n448), .B2(new_n449), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n453), .B1(new_n458), .B2(new_n670), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n669), .A2(new_n411), .A3(new_n562), .A4(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT98), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n542), .A2(new_n544), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n546), .A2(G475), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n491), .B(KEYINPUT90), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n498), .B1(new_n676), .B2(new_n483), .ZN(new_n677));
  INV_X1    g491(.A(new_n499), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n277), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(new_n469), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n565), .A2(new_n470), .ZN(new_n681));
  AOI22_X1  g495(.A1(new_n674), .A2(new_n675), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n602), .A2(new_n673), .A3(new_n682), .ZN(new_n683));
  OAI211_X1 g497(.A(new_n682), .B(new_n187), .C1(new_n291), .C2(new_n292), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(KEYINPUT98), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n672), .B1(new_n683), .B2(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(new_n478), .ZN(G24));
  OR2_X1    g501(.A1(new_n458), .A2(new_n670), .ZN(new_n688));
  AOI22_X1  g502(.A1(new_n688), .A2(new_n453), .B1(new_n561), .B2(G472), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n689), .A2(KEYINPUT99), .A3(new_n591), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n562), .A2(new_n591), .A3(new_n671), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT99), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n644), .B1(new_n690), .B2(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(new_n663), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G125), .ZN(G27));
  NAND3_X1  g510(.A1(new_n600), .A2(new_n187), .A3(new_n601), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n697), .A2(new_n364), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n644), .A2(KEYINPUT42), .ZN(new_n699));
  AND4_X1   g513(.A1(new_n411), .A2(new_n698), .A3(new_n467), .A4(new_n699), .ZN(new_n700));
  NOR3_X1   g514(.A1(new_n644), .A2(new_n697), .A3(new_n364), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT101), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n466), .A2(new_n702), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n615), .A2(KEYINPUT101), .A3(KEYINPUT32), .A4(new_n453), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  AOI21_X1  g519(.A(KEYINPUT100), .B1(new_n463), .B2(new_n464), .ZN(new_n706));
  AND2_X1   g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n452), .B1(new_n705), .B2(new_n706), .ZN(new_n708));
  OAI211_X1 g522(.A(new_n411), .B(new_n701), .C1(new_n707), .C2(new_n708), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n700), .B1(new_n709), .B2(KEYINPUT42), .ZN(new_n710));
  XOR2_X1   g524(.A(KEYINPUT102), .B(G131), .Z(new_n711));
  XNOR2_X1  g525(.A(new_n710), .B(new_n711), .ZN(G33));
  NAND4_X1  g526(.A1(new_n698), .A2(new_n607), .A3(new_n411), .A4(new_n467), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G134), .ZN(G36));
  INV_X1    g528(.A(new_n697), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n563), .A2(new_n591), .ZN(new_n716));
  OR2_X1    g530(.A1(new_n716), .A2(KEYINPUT104), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n716), .A2(KEYINPUT104), .ZN(new_n718));
  INV_X1    g532(.A(new_n575), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n719), .A2(KEYINPUT43), .A3(new_n547), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT43), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n721), .B1(new_n575), .B2(new_n641), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n717), .A2(new_n718), .A3(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT44), .ZN(new_n725));
  OR2_X1    g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n724), .A2(new_n725), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT105), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  AOI21_X1  g543(.A(KEYINPUT105), .B1(new_n724), .B2(new_n725), .ZN(new_n730));
  OAI211_X1 g544(.A(new_n715), .B(new_n726), .C1(new_n729), .C2(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(G469), .A2(G902), .ZN(new_n732));
  AND2_X1   g546(.A1(new_n558), .A2(KEYINPUT45), .ZN(new_n733));
  OAI21_X1  g547(.A(G469), .B1(new_n558), .B2(KEYINPUT45), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n732), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT46), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n363), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n737), .B1(new_n736), .B2(new_n735), .ZN(new_n738));
  AND2_X1   g552(.A1(new_n738), .A2(new_n297), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(new_n626), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT103), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n739), .A2(KEYINPUT103), .A3(new_n626), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n731), .A2(new_n744), .ZN(new_n745));
  XOR2_X1   g559(.A(new_n745), .B(G137), .Z(G39));
  INV_X1    g560(.A(KEYINPUT47), .ZN(new_n747));
  AND3_X1   g561(.A1(new_n738), .A2(new_n747), .A3(new_n297), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n747), .B1(new_n738), .B2(new_n297), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NOR4_X1   g564(.A1(new_n467), .A2(new_n697), .A3(new_n644), .A4(new_n411), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(KEYINPUT106), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G140), .ZN(G42));
  INV_X1    g568(.A(new_n644), .ZN(new_n755));
  AOI21_X1  g569(.A(KEYINPUT99), .B1(new_n689), .B2(new_n591), .ZN(new_n756));
  AND4_X1   g570(.A1(KEYINPUT99), .A2(new_n562), .A3(new_n591), .A4(new_n671), .ZN(new_n757));
  OAI211_X1 g571(.A(new_n755), .B(new_n698), .C1(new_n756), .C2(new_n757), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n580), .A2(new_n641), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n610), .A2(new_n606), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n698), .A2(new_n467), .A3(new_n759), .A4(new_n760), .ZN(new_n761));
  AND3_X1   g575(.A1(new_n758), .A2(new_n713), .A3(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n467), .A2(new_n591), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n622), .A2(new_n652), .A3(new_n548), .A4(new_n187), .ZN(new_n764));
  OAI22_X1  g578(.A1(new_n653), .A2(new_n654), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NOR3_X1   g579(.A1(new_n765), .A2(new_n686), .A3(new_n661), .ZN(new_n766));
  AND4_X1   g580(.A1(new_n549), .A2(new_n583), .A3(new_n593), .A4(new_n577), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n710), .A2(new_n762), .A3(new_n766), .A4(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(new_n604), .ZN(new_n769));
  AOI22_X1  g583(.A1(new_n694), .A2(new_n663), .B1(new_n769), .B2(new_n755), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n683), .A2(new_n685), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n364), .A2(new_n606), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n771), .A2(new_n610), .A3(new_n635), .A4(new_n772), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n770), .A2(new_n620), .A3(new_n773), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n768), .B1(KEYINPUT52), .B2(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT110), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT52), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n770), .A2(new_n620), .A3(new_n773), .A4(new_n777), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n775), .A2(new_n776), .A3(KEYINPUT53), .A4(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT54), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n774), .A2(KEYINPUT52), .ZN(new_n781));
  INV_X1    g595(.A(new_n672), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n771), .A2(new_n782), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n410), .B1(new_n617), .B2(new_n452), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n784), .A2(new_n582), .A3(new_n652), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n783), .A2(new_n655), .A3(new_n785), .A4(new_n664), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n758), .A2(new_n713), .A3(new_n761), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n549), .A2(new_n583), .A3(new_n593), .A4(new_n577), .ZN(new_n788));
  NOR3_X1   g602(.A1(new_n786), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n781), .A2(new_n789), .A3(new_n710), .A4(new_n778), .ZN(new_n790));
  XOR2_X1   g604(.A(KEYINPUT109), .B(KEYINPUT53), .Z(new_n791));
  INV_X1    g605(.A(new_n791), .ZN(new_n792));
  AOI21_X1  g606(.A(KEYINPUT110), .B1(new_n790), .B2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT53), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n790), .A2(new_n794), .ZN(new_n795));
  OAI211_X1 g609(.A(new_n779), .B(new_n780), .C1(new_n793), .C2(new_n795), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n697), .A2(new_n651), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT111), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n723), .A2(new_n798), .A3(new_n505), .ZN(new_n799));
  INV_X1    g613(.A(new_n799), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n798), .B1(new_n723), .B2(new_n505), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n797), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  OR2_X1    g616(.A1(new_n707), .A2(new_n708), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n803), .A2(new_n411), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT114), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  OAI21_X1  g621(.A(KEYINPUT114), .B1(new_n802), .B2(new_n804), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT48), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n807), .A2(KEYINPUT48), .A3(new_n808), .ZN(new_n812));
  OAI211_X1 g626(.A(new_n411), .B(new_n689), .C1(new_n800), .C2(new_n801), .ZN(new_n813));
  INV_X1    g627(.A(new_n663), .ZN(new_n814));
  OAI211_X1 g628(.A(G952), .B(new_n341), .C1(new_n813), .C2(new_n814), .ZN(new_n815));
  AND4_X1   g629(.A1(new_n411), .A2(new_n636), .A3(new_n505), .A4(new_n797), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n815), .B1(new_n576), .B2(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n811), .A2(new_n812), .A3(new_n817), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n719), .A2(new_n641), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n816), .A2(new_n819), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n756), .A2(new_n757), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n820), .B1(new_n802), .B2(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n562), .A2(new_n411), .A3(new_n671), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n723), .A2(new_n505), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n824), .A2(KEYINPUT111), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n823), .B1(new_n825), .B2(new_n799), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n624), .A2(new_n597), .A3(new_n652), .ZN(new_n827));
  INV_X1    g641(.A(new_n827), .ZN(new_n828));
  OAI211_X1 g642(.A(new_n826), .B(new_n828), .C1(KEYINPUT112), .C2(KEYINPUT50), .ZN(new_n829));
  NOR2_X1   g643(.A1(KEYINPUT112), .A2(KEYINPUT50), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n830), .B1(new_n813), .B2(new_n827), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n822), .B1(new_n829), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n668), .A2(new_n362), .ZN(new_n833));
  OAI22_X1  g647(.A1(new_n748), .A2(new_n749), .B1(new_n297), .B2(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n834), .A2(new_n715), .A3(new_n826), .ZN(new_n835));
  AOI21_X1  g649(.A(KEYINPUT51), .B1(new_n832), .B2(new_n835), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n818), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n775), .A2(new_n778), .A3(new_n792), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n790), .A2(KEYINPUT53), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n838), .A2(KEYINPUT54), .A3(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT113), .ZN(new_n841));
  AOI211_X1 g655(.A(new_n697), .B(new_n813), .C1(new_n834), .C2(new_n841), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n842), .B1(new_n841), .B2(new_n834), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n843), .A2(KEYINPUT51), .A3(new_n832), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n796), .A2(new_n837), .A3(new_n840), .A4(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n504), .A2(new_n341), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  OR2_X1    g661(.A1(new_n833), .A2(KEYINPUT49), .ZN(new_n848));
  XOR2_X1   g662(.A(new_n848), .B(KEYINPUT107), .Z(new_n849));
  NAND3_X1  g663(.A1(new_n411), .A2(new_n187), .A3(new_n297), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n719), .A2(new_n547), .ZN(new_n851));
  AOI211_X1 g665(.A(new_n850), .B(new_n851), .C1(KEYINPUT49), .C2(new_n833), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n849), .A2(new_n624), .A3(new_n636), .A4(new_n852), .ZN(new_n853));
  XNOR2_X1  g667(.A(new_n853), .B(KEYINPUT108), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n847), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(KEYINPUT115), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT115), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n847), .A2(new_n857), .A3(new_n854), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n856), .A2(new_n858), .ZN(G75));
  OAI21_X1  g673(.A(new_n779), .B1(new_n793), .B2(new_n795), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n860), .A2(G210), .A3(G902), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT56), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n243), .A2(new_n274), .ZN(new_n863));
  XOR2_X1   g677(.A(new_n863), .B(new_n269), .Z(new_n864));
  XNOR2_X1  g678(.A(new_n864), .B(KEYINPUT55), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT116), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n865), .B1(new_n866), .B2(KEYINPUT56), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n861), .A2(new_n862), .A3(new_n867), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n867), .B1(new_n861), .B2(new_n862), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n341), .A2(G952), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n868), .A2(new_n869), .A3(new_n870), .ZN(G51));
  NAND2_X1  g685(.A1(new_n860), .A2(KEYINPUT54), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT118), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n872), .A2(new_n873), .A3(new_n796), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n860), .A2(KEYINPUT118), .A3(KEYINPUT54), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n732), .B(KEYINPUT117), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n876), .B(KEYINPUT57), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n874), .A2(new_n875), .A3(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n648), .A2(new_n649), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n790), .A2(KEYINPUT110), .A3(new_n794), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n790), .A2(new_n792), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(new_n776), .ZN(new_n883));
  INV_X1    g697(.A(new_n795), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n881), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n885), .A2(new_n277), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n733), .A2(new_n734), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n870), .B1(new_n880), .B2(new_n888), .ZN(G54));
  NAND3_X1  g703(.A1(new_n886), .A2(KEYINPUT58), .A3(G475), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n533), .A2(new_n540), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(new_n870), .ZN(new_n893));
  INV_X1    g707(.A(new_n891), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n886), .A2(KEYINPUT58), .A3(G475), .A4(new_n894), .ZN(new_n895));
  AND3_X1   g709(.A1(new_n892), .A2(new_n893), .A3(new_n895), .ZN(G60));
  NAND2_X1  g710(.A1(G478), .A2(G902), .ZN(new_n897));
  XOR2_X1   g711(.A(new_n897), .B(KEYINPUT59), .Z(new_n898));
  AOI21_X1  g712(.A(new_n898), .B1(new_n796), .B2(new_n840), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n893), .B1(new_n899), .B2(new_n573), .ZN(new_n900));
  AND2_X1   g714(.A1(new_n874), .A2(new_n875), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n898), .B1(new_n571), .B2(new_n572), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n900), .B1(new_n901), .B2(new_n902), .ZN(G63));
  NAND2_X1  g717(.A1(G217), .A2(G902), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(KEYINPUT60), .ZN(new_n905));
  INV_X1    g719(.A(new_n905), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n860), .A2(new_n589), .A3(new_n906), .ZN(new_n907));
  AND2_X1   g721(.A1(new_n907), .A2(new_n893), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT61), .ZN(new_n909));
  AND2_X1   g723(.A1(new_n406), .A2(new_n408), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n910), .B1(new_n860), .B2(new_n906), .ZN(new_n911));
  INV_X1    g725(.A(new_n911), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n908), .A2(KEYINPUT119), .A3(new_n909), .A4(new_n912), .ZN(new_n913));
  OR2_X1    g727(.A1(new_n909), .A2(KEYINPUT119), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n909), .A2(KEYINPUT119), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n907), .A2(new_n893), .ZN(new_n916));
  OAI211_X1 g730(.A(new_n914), .B(new_n915), .C1(new_n916), .C2(new_n911), .ZN(new_n917));
  AND2_X1   g731(.A1(new_n913), .A2(new_n917), .ZN(G66));
  OAI21_X1  g732(.A(G953), .B1(new_n507), .B2(new_n265), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n786), .A2(new_n788), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n919), .B1(new_n920), .B2(G953), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(KEYINPUT120), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n863), .B1(G898), .B2(new_n341), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n922), .B(new_n923), .Z(G69));
  AND2_X1   g738(.A1(new_n753), .A2(new_n713), .ZN(new_n925));
  AND2_X1   g739(.A1(new_n770), .A2(new_n620), .ZN(new_n926));
  AND2_X1   g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(new_n745), .ZN(new_n928));
  INV_X1    g742(.A(new_n804), .ZN(new_n929));
  NAND4_X1  g743(.A1(new_n742), .A2(new_n771), .A3(new_n929), .A4(new_n743), .ZN(new_n930));
  AND2_X1   g744(.A1(new_n930), .A2(new_n710), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n927), .A2(new_n928), .A3(KEYINPUT125), .A4(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT125), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n925), .A2(new_n710), .A3(new_n926), .A4(new_n930), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n933), .B1(new_n934), .B2(new_n745), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n932), .A2(new_n935), .A3(new_n341), .ZN(new_n936));
  NAND2_X1  g750(.A1(G900), .A2(G953), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n419), .A2(new_n423), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n534), .B(KEYINPUT121), .Z(new_n939));
  XNOR2_X1  g753(.A(new_n938), .B(new_n939), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n936), .A2(new_n937), .A3(new_n940), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n940), .B(KEYINPUT122), .ZN(new_n942));
  INV_X1    g756(.A(new_n627), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n581), .B1(new_n575), .B2(new_n547), .ZN(new_n944));
  NAND4_X1  g758(.A1(new_n784), .A2(new_n943), .A3(new_n715), .A4(new_n944), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n945), .B(KEYINPUT123), .Z(new_n946));
  NAND2_X1  g760(.A1(new_n753), .A2(new_n946), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n745), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n926), .A2(new_n639), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n949), .B(KEYINPUT62), .Z(new_n950));
  AND2_X1   g764(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n942), .B1(new_n951), .B2(G953), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n941), .A2(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(G227), .ZN(new_n954));
  OAI21_X1  g768(.A(G953), .B1(new_n954), .B2(new_n605), .ZN(new_n955));
  XOR2_X1   g769(.A(new_n955), .B(KEYINPUT124), .Z(new_n956));
  INV_X1    g770(.A(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n953), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n941), .A2(new_n952), .A3(new_n956), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n958), .A2(new_n959), .ZN(G72));
  XOR2_X1   g774(.A(new_n629), .B(KEYINPUT63), .Z(new_n961));
  INV_X1    g775(.A(new_n426), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n962), .A2(new_n431), .ZN(new_n963));
  INV_X1    g777(.A(new_n454), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n961), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n965), .B(KEYINPUT126), .Z(new_n966));
  NAND3_X1  g780(.A1(new_n838), .A2(new_n839), .A3(new_n966), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n967), .B(KEYINPUT127), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n948), .A2(new_n950), .A3(new_n920), .ZN(new_n969));
  AND2_X1   g783(.A1(new_n969), .A2(new_n961), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n426), .A2(new_n431), .ZN(new_n971));
  OAI211_X1 g785(.A(new_n968), .B(new_n893), .C1(new_n970), .C2(new_n971), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n932), .A2(new_n935), .A3(new_n920), .ZN(new_n973));
  AOI211_X1 g787(.A(new_n431), .B(new_n426), .C1(new_n973), .C2(new_n961), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n972), .A2(new_n974), .ZN(G57));
endmodule


