//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 1 1 0 1 0 0 0 1 0 1 1 1 1 0 0 0 1 1 1 1 1 0 0 1 1 1 1 1 0 0 0 0 0 1 1 1 0 1 1 0 1 0 0 1 0 0 1 1 1 0 1 0 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:01 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n560, new_n561, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n572, new_n573, new_n574, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n612, new_n613, new_n616, new_n618, new_n619,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n824, new_n825, new_n826, new_n827, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT65), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT66), .Z(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  AND2_X1   g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(G137), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  AND2_X1   g038(.A1(KEYINPUT67), .A2(G2105), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT67), .A2(G2105), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  AND2_X1   g042(.A1(new_n467), .A2(G2104), .ZN(new_n468));
  AOI22_X1  g043(.A1(new_n463), .A2(new_n466), .B1(G101), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  INV_X1    g045(.A(G125), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n470), .B1(new_n461), .B2(new_n471), .ZN(new_n472));
  XNOR2_X1  g047(.A(KEYINPUT67), .B(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n469), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(G160));
  NOR2_X1   g051(.A1(new_n461), .A2(new_n466), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  OAI221_X1 g053(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n466), .C2(G112), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n461), .A2(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G136), .ZN(new_n481));
  AND3_X1   g056(.A1(new_n478), .A2(new_n479), .A3(new_n481), .ZN(G162));
  AND2_X1   g057(.A1(G126), .A2(G2105), .ZN(new_n483));
  OAI21_X1  g058(.A(new_n483), .B1(new_n459), .B2(new_n460), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT68), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  OAI211_X1 g061(.A(KEYINPUT68), .B(new_n483), .C1(new_n459), .C2(new_n460), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(KEYINPUT69), .A2(KEYINPUT4), .ZN(new_n489));
  OR2_X1    g064(.A1(KEYINPUT69), .A2(KEYINPUT4), .ZN(new_n490));
  OAI21_X1  g065(.A(G138), .B1(new_n459), .B2(new_n460), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n489), .B(new_n490), .C1(new_n491), .C2(new_n473), .ZN(new_n492));
  INV_X1    g067(.A(G138), .ZN(new_n493));
  OR2_X1    g068(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n494));
  NAND2_X1  g069(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n496), .A2(KEYINPUT69), .A3(KEYINPUT4), .A4(new_n466), .ZN(new_n497));
  OAI21_X1  g072(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n498));
  INV_X1    g073(.A(G114), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n498), .B1(new_n499), .B2(G2105), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n488), .A2(new_n492), .A3(new_n497), .A4(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(G164));
  NAND2_X1  g078(.A1(G75), .A2(G543), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT5), .ZN(new_n505));
  INV_X1    g080(.A(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(KEYINPUT5), .A2(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AND2_X1   g084(.A1(new_n509), .A2(G62), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n504), .B1(new_n510), .B2(KEYINPUT70), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n509), .A2(KEYINPUT70), .A3(G62), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(new_n513));
  OAI21_X1  g088(.A(G651), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  OR2_X1    g089(.A1(KEYINPUT6), .A2(G651), .ZN(new_n515));
  NAND2_X1  g090(.A1(KEYINPUT6), .A2(G651), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n515), .A2(new_n516), .B1(new_n507), .B2(new_n508), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n506), .B1(new_n515), .B2(new_n516), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n517), .A2(G88), .B1(new_n518), .B2(G50), .ZN(new_n519));
  AND2_X1   g094(.A1(new_n514), .A2(new_n519), .ZN(G166));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n521), .B(KEYINPUT7), .ZN(new_n522));
  INV_X1    g097(.A(new_n518), .ZN(new_n523));
  INV_X1    g098(.A(G51), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  AND2_X1   g100(.A1(KEYINPUT5), .A2(G543), .ZN(new_n526));
  NOR2_X1   g101(.A1(KEYINPUT5), .A2(G543), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  AND2_X1   g103(.A1(KEYINPUT6), .A2(G651), .ZN(new_n529));
  NOR2_X1   g104(.A1(KEYINPUT6), .A2(G651), .ZN(new_n530));
  OAI21_X1  g105(.A(G89), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(G63), .A2(G651), .ZN(new_n532));
  AOI21_X1  g107(.A(new_n528), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n525), .A2(new_n533), .ZN(G168));
  INV_X1    g109(.A(G64), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n535), .B1(new_n507), .B2(new_n508), .ZN(new_n536));
  NAND2_X1  g111(.A1(G77), .A2(G543), .ZN(new_n537));
  INV_X1    g112(.A(new_n537), .ZN(new_n538));
  OAI21_X1  g113(.A(KEYINPUT71), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT71), .ZN(new_n540));
  OAI211_X1 g115(.A(new_n540), .B(new_n537), .C1(new_n528), .C2(new_n535), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n539), .A2(G651), .A3(new_n541), .ZN(new_n542));
  XNOR2_X1  g117(.A(KEYINPUT72), .B(G90), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n517), .A2(new_n543), .B1(new_n518), .B2(G52), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n542), .A2(new_n544), .ZN(G301));
  INV_X1    g120(.A(G301), .ZN(G171));
  INV_X1    g121(.A(G56), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n547), .B1(new_n507), .B2(new_n508), .ZN(new_n548));
  NAND2_X1  g123(.A1(G68), .A2(G543), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(new_n550));
  OAI21_X1  g125(.A(KEYINPUT73), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT73), .ZN(new_n552));
  OAI211_X1 g127(.A(new_n552), .B(new_n549), .C1(new_n528), .C2(new_n547), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n551), .A2(G651), .A3(new_n553), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n517), .A2(G81), .B1(new_n518), .B2(G43), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G860), .ZN(G153));
  NAND4_X1  g133(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND4_X1  g136(.A1(G319), .A2(G483), .A3(G661), .A4(new_n561), .ZN(G188));
  NAND2_X1  g137(.A1(new_n518), .A2(G53), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT9), .ZN(new_n564));
  NAND2_X1  g139(.A1(G78), .A2(G543), .ZN(new_n565));
  INV_X1    g140(.A(G65), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n565), .B1(new_n528), .B2(new_n566), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n567), .A2(G651), .B1(new_n517), .B2(G91), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n564), .A2(new_n568), .ZN(G299));
  INV_X1    g144(.A(G168), .ZN(G286));
  NAND2_X1  g145(.A1(new_n514), .A2(new_n519), .ZN(G303));
  NAND2_X1  g146(.A1(new_n517), .A2(G87), .ZN(new_n572));
  OAI21_X1  g147(.A(G651), .B1(new_n509), .B2(G74), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n518), .A2(G49), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(G288));
  OAI22_X1  g150(.A1(new_n527), .A2(new_n526), .B1(new_n529), .B2(new_n530), .ZN(new_n576));
  INV_X1    g151(.A(G86), .ZN(new_n577));
  OR3_X1    g152(.A1(new_n576), .A2(KEYINPUT74), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(G73), .A2(G543), .ZN(new_n579));
  INV_X1    g154(.A(G61), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n579), .B1(new_n528), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n581), .A2(G651), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n518), .A2(G48), .ZN(new_n583));
  OAI21_X1  g158(.A(KEYINPUT74), .B1(new_n576), .B2(new_n577), .ZN(new_n584));
  NAND4_X1  g159(.A1(new_n578), .A2(new_n582), .A3(new_n583), .A4(new_n584), .ZN(G305));
  XOR2_X1   g160(.A(KEYINPUT75), .B(G85), .Z(new_n586));
  NAND2_X1  g161(.A1(new_n517), .A2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(G47), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n588), .B2(new_n523), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n509), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n590));
  INV_X1    g165(.A(G651), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(G290));
  NAND2_X1  g169(.A1(G301), .A2(G868), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n517), .A2(KEYINPUT10), .A3(G92), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT10), .ZN(new_n597));
  INV_X1    g172(.A(G92), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n576), .B2(new_n598), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n596), .A2(new_n599), .B1(G54), .B2(new_n518), .ZN(new_n600));
  INV_X1    g175(.A(G66), .ZN(new_n601));
  INV_X1    g176(.A(G79), .ZN(new_n602));
  OAI22_X1  g177(.A1(new_n528), .A2(new_n601), .B1(new_n602), .B2(new_n506), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT76), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  OAI221_X1 g180(.A(KEYINPUT76), .B1(new_n602), .B2(new_n506), .C1(new_n528), .C2(new_n601), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n605), .A2(G651), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n600), .A2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n595), .B1(new_n609), .B2(G868), .ZN(G284));
  OAI21_X1  g185(.A(new_n595), .B1(new_n609), .B2(G868), .ZN(G321));
  INV_X1    g186(.A(G868), .ZN(new_n612));
  NAND2_X1  g187(.A1(G299), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n613), .B1(new_n612), .B2(G168), .ZN(G297));
  OAI21_X1  g189(.A(new_n613), .B1(new_n612), .B2(G168), .ZN(G280));
  INV_X1    g190(.A(G559), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n609), .B1(new_n616), .B2(G860), .ZN(G148));
  NAND2_X1  g192(.A1(new_n609), .A2(new_n616), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n618), .A2(G868), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n619), .B1(G868), .B2(new_n557), .ZN(G323));
  XNOR2_X1  g195(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g196(.A1(new_n494), .A2(new_n495), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n622), .A2(new_n468), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT12), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT13), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(G2100), .ZN(new_n626));
  AOI22_X1  g201(.A1(G123), .A2(new_n477), .B1(new_n480), .B2(G135), .ZN(new_n627));
  OAI221_X1 g202(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n466), .C2(G111), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(KEYINPUT77), .Z(new_n630));
  INV_X1    g205(.A(new_n630), .ZN(new_n631));
  AND2_X1   g206(.A1(new_n631), .A2(G2096), .ZN(new_n632));
  NOR2_X1   g207(.A1(new_n631), .A2(G2096), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n626), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT78), .ZN(G156));
  INV_X1    g210(.A(KEYINPUT14), .ZN(new_n636));
  XNOR2_X1  g211(.A(G2427), .B(G2438), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(G2430), .ZN(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT15), .B(G2435), .ZN(new_n639));
  AOI21_X1  g214(.A(new_n636), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n640), .B1(new_n639), .B2(new_n638), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2451), .B(G2454), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT16), .ZN(new_n643));
  XOR2_X1   g218(.A(G1341), .B(G1348), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n641), .B(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G2443), .B(G2446), .Z(new_n647));
  OAI21_X1  g222(.A(G14), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  AOI21_X1  g223(.A(new_n648), .B1(new_n647), .B2(new_n646), .ZN(G401));
  XNOR2_X1  g224(.A(G2072), .B(G2078), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT79), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT17), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2067), .B(G2678), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2084), .B(G2090), .ZN(new_n654));
  NOR3_X1   g229(.A1(new_n652), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n654), .B1(new_n651), .B2(new_n653), .ZN(new_n656));
  AOI21_X1  g231(.A(new_n656), .B1(new_n652), .B2(new_n653), .ZN(new_n657));
  INV_X1    g232(.A(new_n653), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n658), .A2(new_n654), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n651), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT18), .ZN(new_n661));
  NOR3_X1   g236(.A1(new_n655), .A2(new_n657), .A3(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2096), .B(G2100), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(G227));
  XOR2_X1   g239(.A(G1971), .B(G1976), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT19), .ZN(new_n666));
  XOR2_X1   g241(.A(G1956), .B(G2474), .Z(new_n667));
  XOR2_X1   g242(.A(G1961), .B(G1966), .Z(new_n668));
  NOR2_X1   g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  AND2_X1   g244(.A1(new_n666), .A2(new_n669), .ZN(new_n670));
  AND2_X1   g245(.A1(new_n667), .A2(new_n668), .ZN(new_n671));
  NOR3_X1   g246(.A1(new_n666), .A2(new_n671), .A3(new_n669), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n666), .A2(new_n671), .ZN(new_n673));
  XOR2_X1   g248(.A(KEYINPUT80), .B(KEYINPUT20), .Z(new_n674));
  AOI211_X1 g249(.A(new_n670), .B(new_n672), .C1(new_n673), .C2(new_n674), .ZN(new_n675));
  OAI21_X1  g250(.A(new_n675), .B1(new_n673), .B2(new_n674), .ZN(new_n676));
  XOR2_X1   g251(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT81), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n676), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1981), .B(G1986), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT82), .ZN(new_n681));
  OR2_X1    g256(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1991), .B(G1996), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n679), .A2(new_n681), .ZN(new_n684));
  AND3_X1   g259(.A1(new_n682), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n683), .B1(new_n682), .B2(new_n684), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n685), .A2(new_n686), .ZN(G229));
  INV_X1    g262(.A(G29), .ZN(new_n688));
  AND2_X1   g263(.A1(new_n688), .A2(G33), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n690));
  INV_X1    g265(.A(KEYINPUT25), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n480), .A2(G139), .ZN(new_n693));
  AOI22_X1  g268(.A1(new_n622), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n694));
  OAI211_X1 g269(.A(new_n692), .B(new_n693), .C1(new_n466), .C2(new_n694), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n695), .B(KEYINPUT90), .Z(new_n696));
  AOI21_X1  g271(.A(new_n689), .B1(new_n696), .B2(G29), .ZN(new_n697));
  INV_X1    g272(.A(G2072), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  XOR2_X1   g274(.A(new_n699), .B(KEYINPUT91), .Z(new_n700));
  INV_X1    g275(.A(G16), .ZN(new_n701));
  NOR2_X1   g276(.A1(G171), .A2(new_n701), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n702), .B1(G5), .B2(new_n701), .ZN(new_n703));
  INV_X1    g278(.A(G1961), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT98), .ZN(new_n706));
  XOR2_X1   g281(.A(KEYINPUT31), .B(G11), .Z(new_n707));
  XNOR2_X1  g282(.A(KEYINPUT30), .B(G28), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n707), .B1(new_n688), .B2(new_n708), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(new_n629), .B2(new_n688), .ZN(new_n710));
  INV_X1    g285(.A(G34), .ZN(new_n711));
  AND2_X1   g286(.A1(new_n711), .A2(KEYINPUT24), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n711), .A2(KEYINPUT24), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n688), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(G160), .B2(new_n688), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(G2084), .ZN(new_n716));
  INV_X1    g291(.A(G2078), .ZN(new_n717));
  NOR2_X1   g292(.A1(G164), .A2(new_n688), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n718), .B1(G27), .B2(new_n688), .ZN(new_n719));
  AOI211_X1 g294(.A(new_n710), .B(new_n716), .C1(new_n717), .C2(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(new_n719), .ZN(new_n721));
  AOI22_X1  g296(.A1(new_n703), .A2(new_n704), .B1(G2078), .B2(new_n721), .ZN(new_n722));
  NAND4_X1  g297(.A1(new_n700), .A2(new_n706), .A3(new_n720), .A4(new_n722), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n697), .A2(new_n698), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT92), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n688), .A2(G32), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n477), .A2(G129), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT93), .ZN(new_n729));
  AND2_X1   g304(.A1(new_n468), .A2(G105), .ZN(new_n730));
  NAND3_X1  g305(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(KEYINPUT26), .ZN(new_n732));
  AOI211_X1 g307(.A(new_n730), .B(new_n732), .C1(G141), .C2(new_n480), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n729), .A2(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(KEYINPUT94), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n734), .B(new_n735), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n727), .B1(new_n736), .B2(new_n688), .ZN(new_n737));
  XOR2_X1   g312(.A(KEYINPUT27), .B(G1996), .Z(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT95), .ZN(new_n739));
  OR2_X1    g314(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n737), .A2(new_n739), .ZN(new_n741));
  NOR2_X1   g316(.A1(G16), .A2(G21), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(G168), .B2(G16), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT96), .ZN(new_n744));
  XNOR2_X1  g319(.A(KEYINPUT97), .B(G1966), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n744), .B(new_n745), .ZN(new_n746));
  NAND4_X1  g321(.A1(new_n726), .A2(new_n740), .A3(new_n741), .A4(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(KEYINPUT99), .ZN(new_n748));
  OR3_X1    g323(.A1(new_n723), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n748), .B1(new_n723), .B2(new_n747), .ZN(new_n750));
  NOR2_X1   g325(.A1(G4), .A2(G16), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT87), .Z(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(new_n608), .B2(new_n701), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT88), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(G1348), .Z(new_n755));
  NOR2_X1   g330(.A1(G29), .A2(G35), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(G162), .B2(G29), .ZN(new_n757));
  XNOR2_X1  g332(.A(KEYINPUT29), .B(G2090), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n757), .B(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n688), .A2(G26), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT28), .ZN(new_n761));
  AOI22_X1  g336(.A1(G128), .A2(new_n477), .B1(new_n480), .B2(G140), .ZN(new_n762));
  OAI221_X1 g337(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n466), .C2(G116), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n764), .A2(G29), .ZN(new_n765));
  AND2_X1   g340(.A1(new_n765), .A2(KEYINPUT89), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n765), .A2(KEYINPUT89), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n761), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n759), .B1(G2067), .B2(new_n768), .ZN(new_n769));
  OR2_X1    g344(.A1(new_n701), .A2(KEYINPUT83), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n701), .A2(KEYINPUT83), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n773), .A2(G20), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(KEYINPUT23), .Z(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(G299), .B2(G16), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(G1956), .ZN(new_n777));
  OAI211_X1 g352(.A(new_n769), .B(new_n777), .C1(G2067), .C2(new_n768), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n772), .A2(G19), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(new_n557), .B2(new_n772), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(G1341), .ZN(new_n781));
  NOR3_X1   g356(.A1(new_n755), .A2(new_n778), .A3(new_n781), .ZN(new_n782));
  NAND3_X1  g357(.A1(new_n749), .A2(new_n750), .A3(new_n782), .ZN(new_n783));
  MUX2_X1   g358(.A(G6), .B(G305), .S(G16), .Z(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT84), .ZN(new_n785));
  XNOR2_X1  g360(.A(KEYINPUT32), .B(G1981), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n773), .A2(G22), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G166), .B2(new_n773), .ZN(new_n789));
  OR2_X1    g364(.A1(new_n789), .A2(G1971), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n701), .A2(G23), .ZN(new_n791));
  INV_X1    g366(.A(G288), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n791), .B1(new_n792), .B2(new_n701), .ZN(new_n793));
  XNOR2_X1  g368(.A(KEYINPUT33), .B(G1976), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT85), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n793), .B(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n789), .A2(G1971), .ZN(new_n797));
  AND3_X1   g372(.A1(new_n790), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n787), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n799), .A2(KEYINPUT34), .ZN(new_n800));
  OR2_X1    g375(.A1(new_n799), .A2(KEYINPUT34), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n688), .A2(G25), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n477), .A2(G119), .ZN(new_n803));
  OAI221_X1 g378(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n466), .C2(G107), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n480), .A2(G131), .ZN(new_n805));
  NAND3_X1  g380(.A1(new_n803), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  INV_X1    g381(.A(new_n806), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n802), .B1(new_n807), .B2(new_n688), .ZN(new_n808));
  XOR2_X1   g383(.A(KEYINPUT35), .B(G1991), .Z(new_n809));
  XOR2_X1   g384(.A(new_n808), .B(new_n809), .Z(new_n810));
  NOR2_X1   g385(.A1(new_n772), .A2(G24), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n811), .B1(new_n593), .B2(new_n772), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(G1986), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n810), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n801), .A2(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(KEYINPUT86), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  AOI21_X1  g392(.A(KEYINPUT86), .B1(new_n801), .B2(new_n814), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n800), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n819), .A2(KEYINPUT36), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT36), .ZN(new_n821));
  OAI211_X1 g396(.A(new_n821), .B(new_n800), .C1(new_n817), .C2(new_n818), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n783), .B1(new_n820), .B2(new_n822), .ZN(G311));
  AND3_X1   g398(.A1(new_n749), .A2(new_n750), .A3(new_n782), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n815), .B(new_n816), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n821), .B1(new_n825), .B2(new_n800), .ZN(new_n826));
  INV_X1    g401(.A(new_n822), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n824), .B1(new_n826), .B2(new_n827), .ZN(G150));
  OAI211_X1 g403(.A(G55), .B(G543), .C1(new_n529), .C2(new_n530), .ZN(new_n829));
  INV_X1    g404(.A(G93), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n829), .B1(new_n576), .B2(new_n830), .ZN(new_n831));
  OAI21_X1  g406(.A(G67), .B1(new_n526), .B2(new_n527), .ZN(new_n832));
  NAND2_X1  g407(.A1(G80), .A2(G543), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n591), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n831), .A2(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(G860), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT37), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n609), .A2(G559), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT38), .ZN(new_n840));
  OR2_X1    g415(.A1(new_n831), .A2(new_n834), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n556), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n835), .A2(new_n554), .A3(new_n555), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n840), .B(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT39), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT100), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n836), .B1(new_n845), .B2(new_n846), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n838), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n850), .B(KEYINPUT101), .Z(G145));
  AOI22_X1  g426(.A1(G130), .A2(new_n477), .B1(new_n480), .B2(G142), .ZN(new_n852));
  OAI221_X1 g427(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n466), .C2(G118), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(new_n624), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(new_n806), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(KEYINPUT103), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n492), .A2(new_n497), .ZN(new_n858));
  INV_X1    g433(.A(new_n858), .ZN(new_n859));
  AOI21_X1  g434(.A(KEYINPUT102), .B1(new_n488), .B2(new_n501), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT102), .ZN(new_n861));
  AOI211_X1 g436(.A(new_n861), .B(new_n500), .C1(new_n486), .C2(new_n487), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n859), .B1(new_n860), .B2(new_n862), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n736), .A2(new_n763), .A3(new_n762), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n734), .B(KEYINPUT94), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n865), .A2(new_n764), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n864), .A2(new_n696), .A3(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n696), .B1(new_n864), .B2(new_n866), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n863), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n869), .ZN(new_n871));
  AOI21_X1  g446(.A(KEYINPUT68), .B1(new_n622), .B2(new_n483), .ZN(new_n872));
  INV_X1    g447(.A(new_n487), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n501), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n874), .A2(new_n861), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n488), .A2(KEYINPUT102), .A3(new_n501), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n858), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n871), .A2(new_n867), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n857), .B1(new_n870), .B2(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n629), .B(new_n475), .ZN(new_n880));
  XOR2_X1   g455(.A(new_n880), .B(G162), .Z(new_n881));
  NOR2_X1   g456(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n870), .A2(new_n878), .A3(new_n856), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(G37), .ZN(new_n885));
  AND3_X1   g460(.A1(new_n870), .A2(new_n878), .A3(new_n857), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n881), .B1(new_n886), .B2(new_n879), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n884), .A2(new_n885), .A3(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n888), .B(new_n889), .ZN(G395));
  NAND2_X1  g465(.A1(new_n841), .A2(new_n612), .ZN(new_n891));
  NAND2_X1  g466(.A1(G303), .A2(new_n792), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n514), .A2(new_n519), .A3(G288), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  OR2_X1    g469(.A1(new_n593), .A2(G305), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n593), .A2(G305), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n894), .A2(new_n897), .ZN(new_n898));
  NAND4_X1  g473(.A1(new_n892), .A2(new_n895), .A3(new_n896), .A4(new_n893), .ZN(new_n899));
  AOI21_X1  g474(.A(KEYINPUT42), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  AND3_X1   g475(.A1(new_n898), .A2(KEYINPUT106), .A3(new_n899), .ZN(new_n901));
  AOI21_X1  g476(.A(KEYINPUT106), .B1(new_n898), .B2(new_n899), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n900), .B1(new_n904), .B2(KEYINPUT42), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n618), .B(new_n844), .ZN(new_n906));
  NAND4_X1  g481(.A1(new_n564), .A2(new_n600), .A3(new_n607), .A4(new_n568), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  AOI22_X1  g483(.A1(new_n564), .A2(new_n568), .B1(new_n600), .B2(new_n607), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n906), .A2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT105), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT41), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n913), .B1(new_n908), .B2(new_n909), .ZN(new_n914));
  NAND2_X1  g489(.A1(G299), .A2(new_n608), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n915), .A2(KEYINPUT41), .A3(new_n907), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  OAI211_X1 g492(.A(new_n911), .B(new_n912), .C1(new_n906), .C2(new_n917), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n918), .B1(new_n912), .B2(new_n911), .ZN(new_n919));
  XOR2_X1   g494(.A(new_n905), .B(new_n919), .Z(new_n920));
  OAI21_X1  g495(.A(new_n891), .B1(new_n920), .B2(new_n612), .ZN(G295));
  OAI21_X1  g496(.A(new_n891), .B1(new_n920), .B2(new_n612), .ZN(G331));
  INV_X1    g497(.A(KEYINPUT110), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT44), .ZN(new_n924));
  AOI21_X1  g499(.A(KEYINPUT107), .B1(new_n542), .B2(new_n544), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n542), .A2(new_n544), .A3(KEYINPUT107), .ZN(new_n927));
  INV_X1    g502(.A(new_n843), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n835), .B1(new_n554), .B2(new_n555), .ZN(new_n929));
  OAI211_X1 g504(.A(new_n926), .B(new_n927), .C1(new_n928), .C2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n927), .ZN(new_n931));
  OAI211_X1 g506(.A(new_n842), .B(new_n843), .C1(new_n931), .C2(new_n925), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(G286), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n930), .A2(new_n932), .A3(G168), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n934), .A2(new_n910), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n917), .B1(new_n934), .B2(new_n935), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT108), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n936), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  AND2_X1   g514(.A1(new_n914), .A2(new_n916), .ZN(new_n940));
  INV_X1    g515(.A(new_n935), .ZN(new_n941));
  AOI21_X1  g516(.A(G168), .B1(new_n930), .B2(new_n932), .ZN(new_n942));
  OAI211_X1 g517(.A(new_n940), .B(new_n938), .C1(new_n941), .C2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n904), .B1(new_n939), .B2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT109), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(new_n937), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n903), .A2(new_n948), .A3(new_n936), .ZN(new_n949));
  AND2_X1   g524(.A1(new_n949), .A2(new_n885), .ZN(new_n950));
  OAI211_X1 g525(.A(new_n904), .B(KEYINPUT109), .C1(new_n939), .C2(new_n944), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n947), .A2(new_n950), .A3(KEYINPUT43), .A4(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT43), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n949), .A2(new_n885), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n903), .B1(new_n948), .B2(new_n936), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n953), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n924), .B1(new_n952), .B2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(new_n957), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n947), .A2(new_n950), .A3(new_n953), .A4(new_n951), .ZN(new_n959));
  OAI21_X1  g534(.A(KEYINPUT43), .B1(new_n954), .B2(new_n955), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(new_n924), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n923), .B1(new_n958), .B2(new_n962), .ZN(new_n963));
  AOI21_X1  g538(.A(KEYINPUT44), .B1(new_n959), .B2(new_n960), .ZN(new_n964));
  NOR3_X1   g539(.A1(new_n957), .A2(new_n964), .A3(KEYINPUT110), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n963), .A2(new_n965), .ZN(G397));
  INV_X1    g541(.A(G1996), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n736), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n865), .A2(G1996), .ZN(new_n969));
  XOR2_X1   g544(.A(new_n764), .B(G2067), .Z(new_n970));
  NAND3_X1  g545(.A1(new_n968), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT45), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n972), .B1(new_n877), .B2(G1384), .ZN(new_n973));
  INV_X1    g548(.A(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n469), .A2(G40), .A3(new_n474), .ZN(new_n975));
  INV_X1    g550(.A(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n971), .A2(new_n978), .ZN(new_n979));
  XNOR2_X1  g554(.A(new_n979), .B(KEYINPUT111), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n807), .A2(new_n809), .ZN(new_n981));
  OAI22_X1  g556(.A1(new_n980), .A2(new_n981), .B1(G2067), .B2(new_n764), .ZN(new_n982));
  OR2_X1    g557(.A1(new_n807), .A2(new_n809), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n977), .B1(new_n983), .B2(new_n981), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n980), .A2(new_n984), .ZN(new_n985));
  OR2_X1    g560(.A1(G290), .A2(G1986), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n977), .A2(new_n986), .ZN(new_n987));
  XOR2_X1   g562(.A(new_n987), .B(KEYINPUT48), .Z(new_n988));
  AOI22_X1  g563(.A1(new_n982), .A2(new_n978), .B1(new_n985), .B2(new_n988), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n977), .B1(new_n736), .B2(new_n970), .ZN(new_n990));
  XNOR2_X1  g565(.A(new_n990), .B(KEYINPUT124), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT46), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n992), .B1(new_n977), .B2(G1996), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n978), .A2(KEYINPUT46), .A3(new_n967), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n991), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  XNOR2_X1  g570(.A(KEYINPUT125), .B(KEYINPUT47), .ZN(new_n996));
  INV_X1    g571(.A(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n991), .A2(new_n993), .A3(new_n994), .A4(new_n996), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(KEYINPUT126), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT126), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n998), .A2(new_n1002), .A3(new_n999), .ZN(new_n1003));
  AND3_X1   g578(.A1(new_n989), .A2(new_n1001), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT51), .ZN(new_n1005));
  INV_X1    g580(.A(G8), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT50), .ZN(new_n1007));
  INV_X1    g582(.A(G1384), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n863), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT112), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n502), .A2(new_n1008), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1010), .B1(new_n1011), .B2(KEYINPUT50), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1009), .A2(new_n1012), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n863), .A2(new_n1010), .A3(new_n1007), .A4(new_n1008), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(G2084), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n976), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT113), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n502), .A2(new_n1019), .A3(KEYINPUT45), .A4(new_n1008), .ZN(new_n1020));
  OAI21_X1  g595(.A(KEYINPUT113), .B1(new_n1011), .B2(new_n972), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n973), .A2(new_n976), .A3(new_n1020), .A4(new_n1021), .ZN(new_n1022));
  AOI22_X1  g597(.A1(new_n1015), .A2(new_n1018), .B1(new_n1022), .B2(new_n745), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1006), .B1(new_n1023), .B2(G168), .ZN(new_n1024));
  INV_X1    g599(.A(new_n745), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n863), .A2(new_n1008), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n975), .B1(new_n1026), .B2(new_n972), .ZN(new_n1027));
  AND2_X1   g602(.A1(new_n1021), .A2(new_n1020), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1025), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1017), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1030));
  OAI21_X1  g605(.A(G286), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1005), .B1(new_n1024), .B2(new_n1031), .ZN(new_n1032));
  AOI211_X1 g607(.A(KEYINPUT51), .B(new_n1006), .C1(new_n1023), .C2(G168), .ZN(new_n1033));
  OAI21_X1  g608(.A(KEYINPUT62), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1030), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1022), .A2(new_n745), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1035), .A2(new_n1036), .A3(G168), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1037), .A2(new_n1031), .A3(G8), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(KEYINPUT51), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT62), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1024), .A2(new_n1005), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1039), .A2(new_n1040), .A3(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n975), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1043), .A2(G1961), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT53), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n863), .A2(KEYINPUT45), .A3(new_n1008), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n975), .B1(new_n1011), .B2(new_n972), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1045), .B1(new_n1048), .B2(G2078), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1049), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1044), .A2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g626(.A(KEYINPUT119), .B1(new_n1022), .B2(G2078), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT119), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1027), .A2(new_n1028), .A3(new_n1053), .A4(new_n717), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1052), .A2(KEYINPUT53), .A3(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1051), .A2(new_n1055), .ZN(new_n1056));
  NOR2_X1   g631(.A1(G166), .A2(new_n1006), .ZN(new_n1057));
  XNOR2_X1  g632(.A(new_n1057), .B(KEYINPUT55), .ZN(new_n1058));
  AOI211_X1 g633(.A(G2090), .B(new_n975), .C1(new_n1013), .C2(new_n1014), .ZN(new_n1059));
  AOI21_X1  g634(.A(G1971), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1060));
  OAI211_X1 g635(.A(G8), .B(new_n1058), .C1(new_n1059), .C2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n863), .A2(new_n1008), .A3(new_n976), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n792), .A2(G1976), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1062), .A2(G8), .A3(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(KEYINPUT52), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n582), .A2(new_n583), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n576), .A2(new_n577), .ZN(new_n1067));
  OAI21_X1  g642(.A(G1981), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1068), .B1(G305), .B2(G1981), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT49), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  OAI211_X1 g646(.A(new_n1068), .B(KEYINPUT49), .C1(G305), .C2(G1981), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1071), .A2(G8), .A3(new_n1062), .A4(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(G1976), .ZN(new_n1074));
  AOI21_X1  g649(.A(KEYINPUT52), .B1(G288), .B2(new_n1074), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1062), .A2(G8), .A3(new_n1063), .A4(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1065), .A2(new_n1073), .A3(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1058), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1007), .B1(new_n863), .B2(new_n1008), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n976), .B1(new_n1011), .B2(KEYINPUT50), .ZN(new_n1080));
  NOR3_X1   g655(.A1(new_n1079), .A2(new_n1080), .A3(G2090), .ZN(new_n1081));
  OAI21_X1  g656(.A(G8), .B1(new_n1081), .B2(new_n1060), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1077), .B1(new_n1078), .B2(new_n1082), .ZN(new_n1083));
  AND4_X1   g658(.A1(G171), .A2(new_n1056), .A3(new_n1061), .A4(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1034), .A2(new_n1042), .A3(new_n1084), .ZN(new_n1085));
  AND3_X1   g660(.A1(new_n1073), .A2(new_n1074), .A3(new_n792), .ZN(new_n1086));
  NOR2_X1   g661(.A1(G305), .A2(G1981), .ZN(new_n1087));
  OAI211_X1 g662(.A(G8), .B(new_n1062), .C1(new_n1086), .C2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1088), .B1(new_n1061), .B2(new_n1077), .ZN(new_n1089));
  NOR3_X1   g664(.A1(new_n1023), .A2(new_n1006), .A3(G286), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1090), .A2(new_n1083), .A3(new_n1061), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT63), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  OAI221_X1 g668(.A(G8), .B1(new_n1058), .B2(KEYINPUT114), .C1(new_n1060), .C2(new_n1059), .ZN(new_n1094));
  OAI21_X1  g669(.A(G8), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT114), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1095), .A2(new_n1096), .A3(new_n1078), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1077), .A2(new_n1092), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1094), .A2(new_n1097), .A3(new_n1090), .A4(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1089), .B1(new_n1093), .B2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1083), .A2(new_n1061), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1101), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1045), .B1(KEYINPUT121), .B2(new_n717), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT120), .ZN(new_n1104));
  OAI221_X1 g679(.A(new_n1103), .B1(KEYINPUT121), .B2(new_n717), .C1(new_n975), .C2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1105), .B1(new_n1104), .B2(new_n975), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1106), .A2(new_n1046), .A3(new_n973), .ZN(new_n1107));
  OAI211_X1 g682(.A(new_n1107), .B(new_n1049), .C1(new_n1043), .C2(G1961), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(G171), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1109), .A2(KEYINPUT122), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1051), .A2(new_n1055), .A3(G301), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT122), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1108), .A2(new_n1112), .A3(G171), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1110), .A2(new_n1111), .A3(KEYINPUT54), .A4(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT54), .ZN(new_n1115));
  AOI21_X1  g690(.A(G301), .B1(new_n1051), .B2(new_n1055), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1108), .A2(G171), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1115), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1102), .A2(new_n1114), .A3(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT57), .ZN(new_n1120));
  XNOR2_X1  g695(.A(G299), .B(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(G1956), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1122), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1123));
  XNOR2_X1  g698(.A(KEYINPUT56), .B(G2072), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1046), .A2(new_n1047), .A3(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT115), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1121), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1128), .B1(new_n1127), .B2(new_n1126), .ZN(new_n1129));
  OR2_X1    g704(.A1(new_n1062), .A2(G2067), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1130), .B1(new_n1043), .B2(G1348), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1123), .A2(new_n1121), .A3(new_n1125), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1131), .A2(new_n609), .A3(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1129), .A2(new_n1133), .ZN(new_n1134));
  AND2_X1   g709(.A1(new_n1132), .A2(KEYINPUT118), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1132), .A2(KEYINPUT118), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT61), .ZN(new_n1137));
  NOR3_X1   g712(.A1(new_n1135), .A2(new_n1136), .A3(new_n1137), .ZN(new_n1138));
  XOR2_X1   g713(.A(KEYINPUT58), .B(G1341), .Z(new_n1139));
  NAND2_X1  g714(.A1(new_n1062), .A2(new_n1139), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1140), .B1(new_n1048), .B2(G1996), .ZN(new_n1141));
  NAND2_X1  g716(.A1(KEYINPUT116), .A2(KEYINPUT59), .ZN(new_n1142));
  AND3_X1   g717(.A1(new_n1141), .A2(new_n557), .A3(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1142), .B1(new_n1141), .B2(new_n557), .ZN(new_n1144));
  OAI211_X1 g719(.A(KEYINPUT60), .B(new_n1130), .C1(new_n1043), .C2(G1348), .ZN(new_n1145));
  OAI22_X1  g720(.A1(new_n1143), .A2(new_n1144), .B1(new_n1145), .B2(new_n609), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1138), .A2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1121), .B1(new_n1123), .B2(new_n1125), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT117), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  AOI211_X1 g725(.A(KEYINPUT117), .B(new_n1121), .C1(new_n1123), .C2(new_n1125), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1132), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT60), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n608), .B1(new_n1131), .B2(new_n1153), .ZN(new_n1154));
  AOI22_X1  g729(.A1(new_n1152), .A2(new_n1137), .B1(new_n1154), .B2(new_n1145), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1134), .B1(new_n1147), .B2(new_n1155), .ZN(new_n1156));
  OAI211_X1 g731(.A(new_n1085), .B(new_n1100), .C1(new_n1119), .C2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT123), .ZN(new_n1158));
  NAND2_X1  g733(.A1(G290), .A2(G1986), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n977), .B1(new_n986), .B2(new_n1159), .ZN(new_n1160));
  NOR3_X1   g735(.A1(new_n980), .A2(new_n1160), .A3(new_n984), .ZN(new_n1161));
  AND3_X1   g736(.A1(new_n1157), .A2(new_n1158), .A3(new_n1161), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1158), .B1(new_n1157), .B2(new_n1161), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1004), .B1(new_n1162), .B2(new_n1163), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g739(.A(G319), .ZN(new_n1166));
  NOR3_X1   g740(.A1(G227), .A2(G401), .A3(new_n1166), .ZN(new_n1167));
  OAI21_X1  g741(.A(new_n1167), .B1(new_n685), .B2(new_n686), .ZN(new_n1168));
  INV_X1    g742(.A(KEYINPUT127), .ZN(new_n1169));
  XNOR2_X1  g743(.A(new_n1168), .B(new_n1169), .ZN(new_n1170));
  NAND3_X1  g744(.A1(new_n1170), .A2(new_n888), .A3(new_n961), .ZN(G225));
  INV_X1    g745(.A(G225), .ZN(G308));
endmodule


