//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 0 0 1 1 0 1 0 1 0 0 1 0 0 0 0 1 0 0 0 0 0 1 1 1 0 1 0 1 0 1 0 1 0 1 1 1 1 1 1 1 1 0 0 1 1 0 0 0 0 0 1 1 0 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:29 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n691, new_n692, new_n693, new_n694, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n728, new_n729,
    new_n730, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n746, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n918, new_n919,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003;
  INV_X1    g000(.A(KEYINPUT84), .ZN(new_n187));
  INV_X1    g001(.A(G104), .ZN(new_n188));
  NOR3_X1   g002(.A1(new_n188), .A2(KEYINPUT3), .A3(G107), .ZN(new_n189));
  INV_X1    g003(.A(G107), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n190), .A2(G104), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n189), .A2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G101), .ZN(new_n193));
  OAI21_X1  g007(.A(KEYINPUT3), .B1(new_n188), .B2(G107), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(KEYINPUT82), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT82), .ZN(new_n196));
  OAI211_X1 g010(.A(new_n196), .B(KEYINPUT3), .C1(new_n188), .C2(G107), .ZN(new_n197));
  NAND4_X1  g011(.A1(new_n192), .A2(new_n193), .A3(new_n195), .A4(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n188), .A2(G107), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n190), .A2(G104), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT83), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n201), .A2(new_n202), .A3(G101), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n201), .A2(G101), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(KEYINPUT83), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n198), .A2(new_n203), .A3(new_n205), .ZN(new_n206));
  AND2_X1   g020(.A1(KEYINPUT65), .A2(G146), .ZN(new_n207));
  NOR2_X1   g021(.A1(KEYINPUT65), .A2(G146), .ZN(new_n208));
  OAI21_X1  g022(.A(G143), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT66), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G128), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n212), .A2(KEYINPUT1), .ZN(new_n213));
  OAI211_X1 g027(.A(KEYINPUT66), .B(G143), .C1(new_n207), .C2(new_n208), .ZN(new_n214));
  INV_X1    g028(.A(G146), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n215), .A2(G143), .ZN(new_n216));
  INV_X1    g030(.A(new_n216), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n211), .A2(new_n213), .A3(new_n214), .A4(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n215), .A2(G143), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n212), .B1(new_n219), .B2(KEYINPUT1), .ZN(new_n220));
  INV_X1    g034(.A(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(G143), .ZN(new_n222));
  OR2_X1    g036(.A1(KEYINPUT65), .A2(G146), .ZN(new_n223));
  NAND2_X1  g037(.A1(KEYINPUT65), .A2(G146), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n222), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n217), .B1(new_n225), .B2(KEYINPUT66), .ZN(new_n226));
  INV_X1    g040(.A(new_n214), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n221), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n206), .B1(new_n218), .B2(new_n228), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n187), .B1(new_n229), .B2(KEYINPUT10), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT0), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n231), .A2(new_n212), .ZN(new_n232));
  NAND4_X1  g046(.A1(new_n211), .A2(new_n214), .A3(new_n217), .A4(new_n232), .ZN(new_n233));
  XNOR2_X1  g047(.A(KEYINPUT65), .B(G146), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n219), .B1(new_n234), .B2(G143), .ZN(new_n235));
  INV_X1    g049(.A(new_n232), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n231), .A2(new_n212), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n235), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n233), .A2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  OR3_X1    g054(.A1(new_n188), .A2(KEYINPUT3), .A3(G107), .ZN(new_n241));
  NAND4_X1  g055(.A1(new_n195), .A2(new_n199), .A3(new_n241), .A4(new_n197), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT4), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n242), .A2(new_n243), .A3(G101), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n242), .A2(G101), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n245), .A2(KEYINPUT4), .A3(new_n198), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n240), .A2(new_n244), .A3(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT10), .ZN(new_n248));
  AND4_X1   g062(.A1(new_n213), .A2(new_n211), .A3(new_n214), .A4(new_n217), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n216), .B1(new_n209), .B2(new_n210), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n220), .B1(new_n250), .B2(new_n214), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  OAI211_X1 g066(.A(KEYINPUT84), .B(new_n248), .C1(new_n252), .C2(new_n206), .ZN(new_n253));
  AND3_X1   g067(.A1(new_n198), .A2(new_n203), .A3(new_n205), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT1), .ZN(new_n255));
  OAI21_X1  g069(.A(G128), .B1(new_n225), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(new_n235), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(new_n218), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n254), .A2(new_n258), .A3(KEYINPUT10), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n230), .A2(new_n247), .A3(new_n253), .A4(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(G137), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n261), .A2(G134), .ZN(new_n262));
  INV_X1    g076(.A(G134), .ZN(new_n263));
  OAI21_X1  g077(.A(KEYINPUT11), .B1(new_n263), .B2(G137), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT11), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n265), .A2(new_n261), .A3(G134), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n262), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(G131), .ZN(new_n268));
  XNOR2_X1  g082(.A(new_n267), .B(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT12), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n267), .A2(new_n268), .ZN(new_n271));
  AOI211_X1 g085(.A(G131), .B(new_n262), .C1(new_n264), .C2(new_n266), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n254), .B1(new_n249), .B2(new_n251), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n206), .A2(new_n257), .A3(new_n218), .ZN(new_n275));
  AOI211_X1 g089(.A(new_n270), .B(new_n273), .C1(new_n274), .C2(new_n275), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n275), .B1(new_n252), .B2(new_n206), .ZN(new_n277));
  AOI21_X1  g091(.A(KEYINPUT12), .B1(new_n277), .B2(new_n269), .ZN(new_n278));
  OAI22_X1  g092(.A1(new_n260), .A2(new_n269), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(KEYINPUT85), .ZN(new_n280));
  XNOR2_X1  g094(.A(G110), .B(G140), .ZN(new_n281));
  INV_X1    g095(.A(G953), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(G227), .ZN(new_n283));
  XNOR2_X1  g097(.A(new_n281), .B(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n277), .A2(new_n269), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(new_n270), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n277), .A2(KEYINPUT12), .A3(new_n269), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT85), .ZN(new_n290));
  AND2_X1   g104(.A1(new_n247), .A2(new_n259), .ZN(new_n291));
  NAND4_X1  g105(.A1(new_n291), .A2(new_n273), .A3(new_n230), .A4(new_n253), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n289), .A2(new_n290), .A3(new_n292), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n280), .A2(new_n285), .A3(new_n293), .ZN(new_n294));
  AND2_X1   g108(.A1(new_n292), .A2(new_n284), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n260), .A2(new_n269), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n294), .A2(G469), .A3(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(G469), .ZN(new_n299));
  XOR2_X1   g113(.A(KEYINPUT73), .B(G902), .Z(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  AND3_X1   g115(.A1(new_n289), .A2(new_n292), .A3(new_n284), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n284), .B1(new_n296), .B2(new_n292), .ZN(new_n303));
  OAI211_X1 g117(.A(new_n299), .B(new_n301), .C1(new_n302), .C2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(G469), .A2(G902), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n298), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  XOR2_X1   g120(.A(KEYINPUT9), .B(G234), .Z(new_n307));
  INV_X1    g121(.A(G902), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  AND2_X1   g123(.A1(new_n309), .A2(G221), .ZN(new_n310));
  XNOR2_X1  g124(.A(new_n310), .B(KEYINPUT81), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n306), .A2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT97), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n313), .B1(new_n212), .B2(G143), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n222), .A2(KEYINPUT97), .A3(G128), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n212), .A2(G143), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n316), .A2(new_n263), .A3(new_n317), .ZN(new_n318));
  XOR2_X1   g132(.A(new_n318), .B(KEYINPUT99), .Z(new_n319));
  XNOR2_X1  g133(.A(G116), .B(G122), .ZN(new_n320));
  XNOR2_X1  g134(.A(new_n320), .B(KEYINPUT96), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(new_n190), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT96), .ZN(new_n323));
  XNOR2_X1  g137(.A(new_n320), .B(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G107), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n322), .A2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT98), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT13), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n327), .B1(new_n316), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n316), .A2(new_n328), .ZN(new_n330));
  NAND4_X1  g144(.A1(new_n314), .A2(new_n315), .A3(KEYINPUT98), .A4(KEYINPUT13), .ZN(new_n331));
  NAND4_X1  g145(.A1(new_n329), .A2(new_n330), .A3(new_n317), .A4(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(G134), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n319), .A2(new_n326), .A3(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT14), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n320), .A2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(G116), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n337), .A2(KEYINPUT14), .A3(G122), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n336), .A2(G107), .A3(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT100), .ZN(new_n340));
  OR2_X1    g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n316), .A2(new_n317), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(G134), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(new_n318), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n339), .A2(new_n340), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n341), .A2(new_n344), .A3(new_n322), .A4(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n334), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n307), .A2(G217), .A3(new_n282), .ZN(new_n348));
  XOR2_X1   g162(.A(new_n348), .B(KEYINPUT101), .Z(new_n349));
  NAND2_X1  g163(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n349), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n334), .A2(new_n346), .A3(new_n351), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n350), .A2(KEYINPUT102), .A3(new_n352), .ZN(new_n353));
  OR3_X1    g167(.A1(new_n347), .A2(KEYINPUT102), .A3(new_n349), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n353), .A2(new_n354), .A3(new_n301), .ZN(new_n355));
  INV_X1    g169(.A(G478), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n356), .A2(KEYINPUT15), .ZN(new_n357));
  XNOR2_X1  g171(.A(new_n355), .B(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(G237), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n360), .A2(new_n282), .A3(G214), .ZN(new_n361));
  XNOR2_X1  g175(.A(new_n361), .B(G143), .ZN(new_n362));
  XNOR2_X1  g176(.A(new_n362), .B(new_n268), .ZN(new_n363));
  OR2_X1    g177(.A1(new_n363), .A2(KEYINPUT17), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n362), .A2(new_n268), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(KEYINPUT17), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT76), .ZN(new_n367));
  XNOR2_X1  g181(.A(KEYINPUT74), .B(G125), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT16), .ZN(new_n369));
  INV_X1    g183(.A(G140), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n368), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  NOR2_X1   g185(.A1(G125), .A2(G140), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n372), .B1(new_n368), .B2(G140), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n371), .B1(new_n373), .B2(new_n369), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n367), .B1(new_n374), .B2(new_n215), .ZN(new_n375));
  INV_X1    g189(.A(G125), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(KEYINPUT74), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT74), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(G125), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n377), .A2(new_n379), .A3(G140), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n376), .A2(new_n370), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n369), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  AND4_X1   g196(.A1(new_n369), .A2(new_n377), .A3(new_n379), .A4(new_n370), .ZN(new_n383));
  OAI211_X1 g197(.A(new_n367), .B(new_n215), .C1(new_n382), .C2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n375), .A2(new_n385), .ZN(new_n386));
  OAI211_X1 g200(.A(G146), .B(new_n371), .C1(new_n373), .C2(new_n369), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(KEYINPUT75), .ZN(new_n388));
  INV_X1    g202(.A(new_n382), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT75), .ZN(new_n390));
  NAND4_X1  g204(.A1(new_n389), .A2(new_n390), .A3(G146), .A4(new_n371), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n388), .A2(new_n391), .ZN(new_n392));
  NOR3_X1   g206(.A1(new_n386), .A2(KEYINPUT95), .A3(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT95), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n380), .A2(new_n381), .ZN(new_n395));
  AND3_X1   g209(.A1(new_n377), .A2(new_n379), .A3(new_n369), .ZN(new_n396));
  AOI22_X1  g210(.A1(new_n395), .A2(KEYINPUT16), .B1(new_n396), .B2(new_n370), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n390), .B1(new_n397), .B2(G146), .ZN(new_n398));
  NOR4_X1   g212(.A1(new_n382), .A2(new_n383), .A3(KEYINPUT75), .A4(new_n215), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  OAI21_X1  g214(.A(KEYINPUT76), .B1(new_n397), .B2(G146), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(new_n384), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n394), .B1(new_n400), .B2(new_n402), .ZN(new_n403));
  OAI211_X1 g217(.A(new_n364), .B(new_n366), .C1(new_n393), .C2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(KEYINPUT18), .A2(G131), .ZN(new_n405));
  XOR2_X1   g219(.A(new_n362), .B(new_n405), .Z(new_n406));
  INV_X1    g220(.A(KEYINPUT77), .ZN(new_n407));
  NAND2_X1  g221(.A1(G125), .A2(G140), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n407), .B1(new_n409), .B2(new_n372), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n381), .A2(KEYINPUT77), .A3(new_n408), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  AND3_X1   g226(.A1(new_n412), .A2(KEYINPUT78), .A3(new_n234), .ZN(new_n413));
  AOI21_X1  g227(.A(KEYINPUT78), .B1(new_n412), .B2(new_n234), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n395), .A2(new_n215), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n406), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  XNOR2_X1  g231(.A(G113), .B(G122), .ZN(new_n418));
  XNOR2_X1  g232(.A(new_n418), .B(new_n188), .ZN(new_n419));
  XNOR2_X1  g233(.A(new_n419), .B(KEYINPUT94), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n404), .A2(new_n417), .A3(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n419), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT19), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n412), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n373), .A2(KEYINPUT19), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n424), .A2(new_n425), .A3(new_n234), .ZN(new_n426));
  OR2_X1    g240(.A1(new_n426), .A2(KEYINPUT93), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(KEYINPUT93), .ZN(new_n428));
  AND4_X1   g242(.A1(new_n387), .A2(new_n427), .A3(new_n363), .A4(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(new_n417), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n422), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n421), .A2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT20), .ZN(new_n433));
  NOR2_X1   g247(.A1(G475), .A2(G902), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n432), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(new_n434), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n436), .B1(new_n421), .B2(new_n431), .ZN(new_n437));
  XNOR2_X1  g251(.A(KEYINPUT92), .B(KEYINPUT20), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n435), .B1(new_n437), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n282), .A2(G952), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n441), .B1(G234), .B2(G237), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(G234), .A2(G237), .ZN(new_n444));
  AND3_X1   g258(.A1(new_n300), .A2(G953), .A3(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  XOR2_X1   g260(.A(KEYINPUT21), .B(G898), .Z(new_n447));
  OAI21_X1  g261(.A(new_n443), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  XNOR2_X1  g262(.A(new_n448), .B(KEYINPUT103), .ZN(new_n449));
  INV_X1    g263(.A(new_n421), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n419), .B1(new_n404), .B2(new_n417), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n308), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(G475), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n359), .A2(new_n440), .A3(new_n449), .A4(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(G214), .B1(G237), .B2(G902), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT91), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n240), .A2(new_n368), .ZN(new_n457));
  INV_X1    g271(.A(new_n368), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n258), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n282), .A2(G224), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(new_n461), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n457), .A2(new_n459), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  XNOR2_X1  g279(.A(G110), .B(G122), .ZN(new_n466));
  INV_X1    g280(.A(G119), .ZN(new_n467));
  OAI21_X1  g281(.A(KEYINPUT71), .B1(new_n467), .B2(G116), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT71), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n469), .A2(new_n337), .A3(G119), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  OAI21_X1  g285(.A(KEYINPUT70), .B1(new_n337), .B2(G119), .ZN(new_n472));
  OR3_X1    g286(.A1(new_n337), .A2(KEYINPUT70), .A3(G119), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n471), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  XNOR2_X1  g288(.A(KEYINPUT2), .B(G113), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(new_n475), .ZN(new_n477));
  NAND4_X1  g291(.A1(new_n477), .A2(new_n471), .A3(new_n472), .A4(new_n473), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n246), .A2(new_n479), .A3(new_n244), .ZN(new_n480));
  AND2_X1   g294(.A1(new_n205), .A2(new_n203), .ZN(new_n481));
  INV_X1    g295(.A(G113), .ZN(new_n482));
  XNOR2_X1  g296(.A(KEYINPUT86), .B(KEYINPUT5), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n337), .A2(G119), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n485), .B1(new_n474), .B2(new_n483), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n481), .A2(new_n478), .A3(new_n486), .A4(new_n198), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n466), .B1(new_n480), .B2(new_n487), .ZN(new_n488));
  XNOR2_X1  g302(.A(KEYINPUT88), .B(KEYINPUT6), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n480), .A2(new_n487), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT87), .ZN(new_n492));
  INV_X1    g306(.A(new_n466), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n491), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(KEYINPUT6), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n480), .A2(new_n466), .A3(new_n487), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n496), .B1(new_n488), .B2(new_n492), .ZN(new_n497));
  OAI211_X1 g311(.A(new_n465), .B(new_n490), .C1(new_n495), .C2(new_n497), .ZN(new_n498));
  XNOR2_X1  g312(.A(new_n466), .B(KEYINPUT8), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n206), .A2(new_n478), .A3(new_n486), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT5), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n485), .B1(new_n474), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(new_n478), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n503), .B(KEYINPUT89), .ZN(new_n504));
  OAI211_X1 g318(.A(new_n499), .B(new_n500), .C1(new_n504), .C2(new_n206), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT7), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n506), .B1(new_n463), .B2(KEYINPUT90), .ZN(new_n507));
  OAI211_X1 g321(.A(new_n460), .B(new_n507), .C1(KEYINPUT90), .C2(new_n463), .ZN(new_n508));
  OAI211_X1 g322(.A(new_n457), .B(new_n459), .C1(new_n506), .C2(new_n463), .ZN(new_n509));
  NAND4_X1  g323(.A1(new_n505), .A2(new_n508), .A3(new_n509), .A4(new_n496), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n498), .A2(new_n308), .A3(new_n510), .ZN(new_n511));
  OAI21_X1  g325(.A(G210), .B1(G237), .B2(G902), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  NAND4_X1  g328(.A1(new_n498), .A2(new_n308), .A3(new_n512), .A4(new_n510), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n456), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  AND2_X1   g330(.A1(new_n515), .A2(new_n456), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n455), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NOR3_X1   g332(.A1(new_n312), .A2(new_n454), .A3(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT23), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n520), .B1(G119), .B2(new_n212), .ZN(new_n521));
  NOR3_X1   g335(.A1(new_n467), .A2(KEYINPUT23), .A3(G128), .ZN(new_n522));
  OAI22_X1  g336(.A1(new_n521), .A2(new_n522), .B1(G119), .B2(new_n212), .ZN(new_n523));
  XNOR2_X1  g337(.A(G119), .B(G128), .ZN(new_n524));
  XOR2_X1   g338(.A(KEYINPUT24), .B(G110), .Z(new_n525));
  OAI22_X1  g339(.A1(new_n523), .A2(G110), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  OAI211_X1 g340(.A(new_n387), .B(new_n526), .C1(new_n413), .C2(new_n414), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n527), .B(KEYINPUT79), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n525), .A2(new_n524), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n523), .A2(G110), .ZN(new_n530));
  OAI211_X1 g344(.A(new_n529), .B(new_n530), .C1(new_n386), .C2(new_n392), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n282), .A2(G221), .A3(G234), .ZN(new_n533));
  XNOR2_X1  g347(.A(new_n533), .B(KEYINPUT22), .ZN(new_n534));
  XNOR2_X1  g348(.A(new_n534), .B(new_n261), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n532), .A2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(new_n535), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n528), .A2(new_n531), .A3(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n536), .A2(new_n301), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(KEYINPUT25), .ZN(new_n540));
  INV_X1    g354(.A(G217), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n541), .B1(new_n301), .B2(G234), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT25), .ZN(new_n543));
  NAND4_X1  g357(.A1(new_n536), .A2(new_n543), .A3(new_n301), .A4(new_n538), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n540), .A2(new_n542), .A3(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT80), .ZN(new_n546));
  INV_X1    g360(.A(new_n538), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n537), .B1(new_n528), .B2(new_n531), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n542), .A2(G902), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n536), .A2(KEYINPUT80), .A3(new_n538), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  AND2_X1   g366(.A1(new_n545), .A2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  OR3_X1    g368(.A1(new_n261), .A2(KEYINPUT69), .A3(G134), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT68), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n556), .B1(new_n263), .B2(G137), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n261), .A2(KEYINPUT68), .A3(G134), .ZN(new_n558));
  OAI21_X1  g372(.A(KEYINPUT69), .B1(new_n261), .B2(G134), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n555), .A2(new_n557), .A3(new_n558), .A4(new_n559), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n272), .B1(G131), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n258), .A2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT72), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n258), .A2(new_n561), .A3(KEYINPUT72), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n240), .A2(new_n269), .ZN(new_n566));
  NAND4_X1  g380(.A1(new_n564), .A2(KEYINPUT30), .A3(new_n565), .A4(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT67), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n568), .B1(new_n239), .B2(new_n273), .ZN(new_n569));
  NAND4_X1  g383(.A1(new_n269), .A2(KEYINPUT67), .A3(new_n233), .A4(new_n238), .ZN(new_n570));
  AOI22_X1  g384(.A1(new_n569), .A2(new_n570), .B1(new_n258), .B2(new_n561), .ZN(new_n571));
  XOR2_X1   g385(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n572));
  OAI211_X1 g386(.A(new_n567), .B(new_n479), .C1(new_n571), .C2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(new_n479), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n564), .A2(new_n574), .A3(new_n565), .A4(new_n566), .ZN(new_n575));
  XNOR2_X1  g389(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n576), .B(G101), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n360), .A2(new_n282), .A3(G210), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n577), .B(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n573), .A2(new_n575), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(KEYINPUT31), .ZN(new_n581));
  INV_X1    g395(.A(new_n579), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT28), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n569), .A2(new_n570), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(new_n562), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(new_n479), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n583), .B1(new_n586), .B2(new_n575), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n566), .A2(new_n574), .A3(new_n562), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(new_n583), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n582), .B1(new_n587), .B2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT31), .ZN(new_n592));
  NAND4_X1  g406(.A1(new_n573), .A2(new_n592), .A3(new_n575), .A4(new_n579), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n581), .A2(new_n591), .A3(new_n593), .ZN(new_n594));
  NOR2_X1   g408(.A1(G472), .A2(G902), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(KEYINPUT32), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT32), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n594), .A2(new_n598), .A3(new_n595), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  NOR3_X1   g414(.A1(new_n587), .A2(new_n590), .A3(new_n582), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n579), .B1(new_n573), .B2(new_n575), .ZN(new_n602));
  NOR3_X1   g416(.A1(new_n601), .A2(KEYINPUT29), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n564), .A2(new_n566), .ZN(new_n604));
  INV_X1    g418(.A(new_n565), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n479), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n606), .A2(new_n575), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(KEYINPUT28), .ZN(new_n608));
  AND2_X1   g422(.A1(new_n579), .A2(KEYINPUT29), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n608), .A2(new_n589), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(new_n301), .ZN(new_n611));
  OAI21_X1  g425(.A(G472), .B1(new_n603), .B2(new_n611), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n554), .B1(new_n600), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n519), .A2(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n614), .B(G101), .ZN(G3));
  NAND2_X1  g429(.A1(new_n514), .A2(new_n515), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(new_n455), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(KEYINPUT104), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT33), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n353), .A2(new_n354), .A3(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n350), .A2(KEYINPUT33), .A3(new_n352), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n620), .A2(G478), .A3(new_n301), .A4(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n355), .A2(new_n356), .ZN(new_n623));
  AND2_X1   g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n624), .B1(new_n440), .B2(new_n453), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT104), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n616), .A2(new_n626), .A3(new_n455), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n618), .A2(new_n625), .A3(new_n449), .A4(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n594), .A2(new_n301), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(G472), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n553), .A2(new_n630), .A3(new_n596), .ZN(new_n631));
  NOR3_X1   g445(.A1(new_n628), .A2(new_n312), .A3(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(KEYINPUT34), .B(G104), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G6));
  AOI21_X1  g448(.A(new_n626), .B1(new_n616), .B2(new_n455), .ZN(new_n635));
  INV_X1    g449(.A(new_n455), .ZN(new_n636));
  AOI211_X1 g450(.A(KEYINPUT104), .B(new_n636), .C1(new_n514), .C2(new_n515), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n439), .B1(new_n432), .B2(new_n434), .ZN(new_n639));
  AOI211_X1 g453(.A(new_n436), .B(new_n438), .C1(new_n421), .C2(new_n431), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n404), .A2(new_n417), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n422), .ZN(new_n642));
  AOI21_X1  g456(.A(G902), .B1(new_n642), .B2(new_n421), .ZN(new_n643));
  INV_X1    g457(.A(G475), .ZN(new_n644));
  OAI22_X1  g458(.A1(new_n639), .A2(new_n640), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n645), .A2(new_n359), .ZN(new_n646));
  AND3_X1   g460(.A1(new_n638), .A2(new_n449), .A3(new_n646), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n631), .A2(new_n312), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  XOR2_X1   g463(.A(KEYINPUT35), .B(G107), .Z(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(G9));
  OAI21_X1  g465(.A(new_n532), .B1(KEYINPUT36), .B2(new_n535), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n535), .A2(KEYINPUT36), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n528), .A2(new_n531), .A3(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n652), .A2(new_n550), .A3(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(KEYINPUT105), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(new_n545), .ZN(new_n657));
  AND3_X1   g471(.A1(new_n657), .A2(new_n630), .A3(new_n596), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n519), .A2(new_n658), .ZN(new_n659));
  XOR2_X1   g473(.A(new_n659), .B(KEYINPUT37), .Z(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(G110), .ZN(G12));
  XNOR2_X1  g475(.A(new_n437), .B(new_n439), .ZN(new_n662));
  INV_X1    g476(.A(G900), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n442), .B1(new_n445), .B2(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n662), .A2(new_n358), .A3(new_n453), .A4(new_n665), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n666), .A2(new_n312), .ZN(new_n667));
  AND3_X1   g481(.A1(new_n594), .A2(new_n598), .A3(new_n595), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n598), .B1(new_n594), .B2(new_n595), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n612), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n667), .A2(new_n670), .A3(new_n638), .A4(new_n657), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G128), .ZN(G30));
  XNOR2_X1  g486(.A(new_n664), .B(KEYINPUT39), .ZN(new_n673));
  OR2_X1    g487(.A1(new_n312), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n674), .A2(KEYINPUT40), .ZN(new_n675));
  AOI211_X1 g489(.A(KEYINPUT20), .B(new_n436), .C1(new_n421), .C2(new_n431), .ZN(new_n676));
  OAI22_X1  g490(.A1(new_n639), .A2(new_n676), .B1(new_n643), .B2(new_n644), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(new_n358), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  AND2_X1   g493(.A1(new_n573), .A2(new_n575), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n680), .A2(new_n582), .ZN(new_n681));
  OAI21_X1  g495(.A(new_n308), .B1(new_n607), .B2(new_n579), .ZN(new_n682));
  OAI21_X1  g496(.A(G472), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n657), .B1(new_n600), .B2(new_n683), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n517), .B1(new_n616), .B2(KEYINPUT91), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT38), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n685), .B(new_n686), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n636), .B1(new_n674), .B2(KEYINPUT40), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n679), .A2(new_n684), .A3(new_n687), .A4(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G143), .ZN(G45));
  NAND2_X1  g504(.A1(new_n622), .A2(new_n623), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n677), .A2(new_n691), .A3(new_n665), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n692), .A2(new_n312), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n693), .A2(new_n670), .A3(new_n638), .A4(new_n657), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G146), .ZN(G48));
  OAI21_X1  g509(.A(new_n301), .B1(new_n302), .B2(new_n303), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(G469), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n697), .A2(KEYINPUT106), .A3(new_n304), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT106), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n696), .A2(new_n699), .A3(G469), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n310), .B1(new_n698), .B2(new_n700), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n701), .A2(new_n553), .A3(new_n670), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n702), .A2(new_n628), .ZN(new_n703));
  XOR2_X1   g517(.A(KEYINPUT41), .B(G113), .Z(new_n704));
  XNOR2_X1  g518(.A(new_n703), .B(new_n704), .ZN(G15));
  INV_X1    g519(.A(new_n702), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT107), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n706), .A2(new_n647), .A3(new_n707), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n638), .A2(new_n449), .A3(new_n646), .ZN(new_n709));
  OAI21_X1  g523(.A(KEYINPUT107), .B1(new_n709), .B2(new_n702), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G116), .ZN(G18));
  NAND4_X1  g526(.A1(new_n670), .A2(new_n627), .A3(new_n618), .A4(new_n657), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n698), .A2(new_n700), .ZN(new_n714));
  INV_X1    g528(.A(new_n310), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NOR3_X1   g530(.A1(new_n713), .A2(new_n454), .A3(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(new_n467), .ZN(G21));
  INV_X1    g532(.A(new_n678), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n638), .A2(new_n719), .A3(new_n701), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n583), .B1(new_n606), .B2(new_n575), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n582), .B1(new_n721), .B2(new_n590), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n722), .A2(new_n581), .A3(new_n593), .ZN(new_n723));
  AOI22_X1  g537(.A1(new_n629), .A2(G472), .B1(new_n595), .B2(new_n723), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n724), .A2(new_n553), .A3(new_n449), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n720), .A2(new_n725), .ZN(new_n726));
  XOR2_X1   g540(.A(new_n726), .B(G122), .Z(G24));
  AND2_X1   g541(.A1(new_n724), .A2(new_n657), .ZN(new_n728));
  INV_X1    g542(.A(new_n692), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n728), .A2(new_n729), .A3(new_n638), .A4(new_n701), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G125), .ZN(G27));
  AND2_X1   g545(.A1(new_n306), .A2(new_n715), .ZN(new_n732));
  NOR3_X1   g546(.A1(new_n516), .A2(new_n636), .A3(new_n517), .ZN(new_n733));
  AND2_X1   g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT109), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT42), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n735), .B1(KEYINPUT108), .B2(new_n736), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n737), .B1(new_n735), .B2(new_n736), .ZN(new_n738));
  INV_X1    g552(.A(new_n738), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n734), .A2(new_n613), .A3(new_n729), .A4(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(new_n737), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n732), .A2(new_n670), .A3(new_n553), .A4(new_n733), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n741), .B1(new_n742), .B2(new_n692), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n740), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G131), .ZN(G33));
  OR2_X1    g559(.A1(new_n742), .A2(new_n666), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G134), .ZN(G36));
  INV_X1    g561(.A(KEYINPUT46), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n284), .B1(new_n279), .B2(KEYINPUT85), .ZN(new_n749));
  AOI22_X1  g563(.A1(new_n749), .A2(new_n293), .B1(new_n296), .B2(new_n295), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT45), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n750), .B(new_n751), .ZN(new_n752));
  OAI211_X1 g566(.A(new_n748), .B(G469), .C1(new_n752), .C2(G902), .ZN(new_n753));
  OR2_X1    g567(.A1(new_n750), .A2(KEYINPUT45), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n750), .A2(KEYINPUT45), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n754), .A2(new_n755), .A3(G469), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n756), .A2(KEYINPUT46), .A3(new_n305), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n753), .A2(new_n757), .A3(new_n304), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(new_n715), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n759), .A2(new_n673), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT110), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n760), .B(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(new_n677), .ZN(new_n763));
  AOI21_X1  g577(.A(KEYINPUT43), .B1(new_n763), .B2(new_n691), .ZN(new_n764));
  INV_X1    g578(.A(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n763), .A2(KEYINPUT43), .A3(new_n691), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n630), .A2(new_n596), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n767), .A2(new_n768), .A3(new_n657), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT44), .ZN(new_n770));
  OAI21_X1  g584(.A(KEYINPUT111), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n733), .B(KEYINPUT112), .ZN(new_n772));
  INV_X1    g586(.A(new_n772), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n773), .B1(new_n769), .B2(new_n770), .ZN(new_n774));
  AOI22_X1  g588(.A1(new_n765), .A2(new_n766), .B1(new_n596), .B2(new_n630), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT111), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n775), .A2(new_n776), .A3(KEYINPUT44), .A4(new_n657), .ZN(new_n777));
  AND3_X1   g591(.A1(new_n771), .A2(new_n774), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n762), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G137), .ZN(G39));
  INV_X1    g594(.A(new_n733), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT47), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n759), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n758), .A2(KEYINPUT47), .A3(new_n715), .ZN(new_n784));
  AOI211_X1 g598(.A(new_n670), .B(new_n781), .C1(new_n783), .C2(new_n784), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n692), .A2(new_n553), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G140), .ZN(G42));
  INV_X1    g602(.A(new_n311), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n714), .A2(new_n789), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n783), .A2(new_n784), .A3(new_n790), .ZN(new_n791));
  AND2_X1   g605(.A1(new_n724), .A2(new_n553), .ZN(new_n792));
  INV_X1    g606(.A(new_n766), .ZN(new_n793));
  OAI211_X1 g607(.A(new_n442), .B(new_n792), .C1(new_n793), .C2(new_n764), .ZN(new_n794));
  OAI21_X1  g608(.A(KEYINPUT117), .B1(new_n773), .B2(new_n794), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n443), .B1(new_n765), .B2(new_n766), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT117), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n796), .A2(new_n772), .A3(new_n797), .A4(new_n792), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n795), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n791), .A2(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT50), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n796), .A2(new_n636), .A3(new_n792), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n687), .A2(new_n716), .ZN(new_n803));
  INV_X1    g617(.A(new_n803), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n801), .B1(new_n802), .B2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(new_n794), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n806), .A2(KEYINPUT50), .A3(new_n636), .A4(new_n803), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n716), .A2(new_n781), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n600), .A2(new_n683), .ZN(new_n810));
  AND4_X1   g624(.A1(new_n553), .A2(new_n809), .A3(new_n442), .A4(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n811), .A2(new_n763), .A3(new_n624), .ZN(new_n812));
  AND2_X1   g626(.A1(new_n796), .A2(new_n809), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n813), .A2(new_n728), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n800), .A2(new_n808), .A3(new_n812), .A4(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(KEYINPUT51), .ZN(new_n816));
  AOI22_X1  g630(.A1(new_n791), .A2(new_n799), .B1(new_n728), .B2(new_n813), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT51), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n817), .A2(new_n818), .A3(new_n812), .A4(new_n808), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n816), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n813), .A2(new_n613), .ZN(new_n821));
  XOR2_X1   g635(.A(KEYINPUT118), .B(KEYINPUT48), .Z(new_n822));
  XNOR2_X1  g636(.A(new_n821), .B(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n714), .A2(new_n618), .A3(new_n715), .A4(new_n627), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n794), .A2(new_n824), .ZN(new_n825));
  AOI211_X1 g639(.A(new_n441), .B(new_n825), .C1(new_n625), .C2(new_n811), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n820), .A2(new_n823), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n827), .A2(KEYINPUT119), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT119), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n820), .A2(new_n829), .A3(new_n823), .A4(new_n826), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT116), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n646), .A2(new_n311), .A3(new_n306), .A4(new_n665), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n713), .A2(new_n833), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n625), .A2(new_n724), .A3(new_n657), .A4(new_n665), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n824), .A2(new_n835), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT52), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n678), .A2(new_n635), .A3(new_n637), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n839), .A2(new_n684), .A3(new_n665), .A4(new_n732), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n837), .A2(new_n838), .A3(new_n694), .A4(new_n840), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n840), .A2(new_n671), .A3(new_n694), .A4(new_n730), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n842), .A2(KEYINPUT52), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(new_n518), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n454), .A2(new_n312), .ZN(new_n846));
  OAI211_X1 g660(.A(new_n845), .B(new_n846), .C1(new_n613), .C2(new_n658), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n312), .A2(new_n645), .A3(new_n664), .ZN(new_n848));
  AND3_X1   g662(.A1(new_n685), .A2(new_n455), .A3(new_n657), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n848), .A2(new_n670), .A3(new_n849), .A4(new_n359), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n677), .A2(new_n691), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n440), .A2(new_n358), .A3(new_n453), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n518), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n853), .A2(new_n648), .A3(new_n449), .ZN(new_n854));
  AND3_X1   g668(.A1(new_n847), .A2(new_n850), .A3(new_n854), .ZN(new_n855));
  OAI22_X1  g669(.A1(new_n720), .A2(new_n725), .B1(new_n702), .B2(new_n628), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n856), .A2(new_n717), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n855), .A2(new_n857), .A3(new_n711), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT113), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n734), .A2(new_n859), .A3(new_n729), .A4(new_n728), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n732), .A2(new_n733), .ZN(new_n861));
  OAI21_X1  g675(.A(KEYINPUT113), .B1(new_n861), .B2(new_n835), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n744), .A2(new_n863), .A3(new_n746), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n844), .A2(new_n858), .A3(new_n864), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n832), .B1(new_n865), .B2(KEYINPUT53), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n855), .A2(new_n857), .A3(new_n711), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n744), .A2(new_n863), .A3(new_n746), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n867), .A2(new_n843), .A3(new_n841), .A4(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT53), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n869), .A2(KEYINPUT116), .A3(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n866), .A2(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT54), .ZN(new_n873));
  AOI22_X1  g687(.A1(new_n841), .A2(new_n843), .B1(KEYINPUT115), .B2(new_n842), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n842), .A2(KEYINPUT115), .A3(new_n838), .ZN(new_n875));
  INV_X1    g689(.A(new_n875), .ZN(new_n876));
  NOR3_X1   g690(.A1(new_n874), .A2(new_n870), .A3(new_n876), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n858), .A2(new_n864), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n872), .A2(new_n873), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n869), .A2(KEYINPUT53), .ZN(new_n881));
  INV_X1    g695(.A(new_n874), .ZN(new_n882));
  OAI211_X1 g696(.A(new_n882), .B(new_n875), .C1(new_n878), .C2(KEYINPUT114), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n878), .A2(KEYINPUT114), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n884), .A2(new_n870), .ZN(new_n885));
  OAI211_X1 g699(.A(KEYINPUT54), .B(new_n881), .C1(new_n883), .C2(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n880), .A2(new_n886), .ZN(new_n887));
  OAI22_X1  g701(.A1(new_n831), .A2(new_n887), .B1(G952), .B2(G953), .ZN(new_n888));
  XOR2_X1   g702(.A(new_n714), .B(KEYINPUT49), .Z(new_n889));
  NOR4_X1   g703(.A1(new_n889), .A2(new_n554), .A3(new_n636), .A4(new_n789), .ZN(new_n890));
  INV_X1    g704(.A(new_n687), .ZN(new_n891));
  AND2_X1   g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n892), .A2(new_n763), .A3(new_n691), .A4(new_n810), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n888), .A2(new_n893), .ZN(G75));
  NOR3_X1   g708(.A1(new_n865), .A2(new_n832), .A3(KEYINPUT53), .ZN(new_n895));
  AOI21_X1  g709(.A(KEYINPUT116), .B1(new_n869), .B2(new_n870), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n879), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n897), .A2(new_n300), .A3(new_n513), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT56), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n490), .B1(new_n495), .B2(new_n497), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n900), .B(new_n465), .ZN(new_n901));
  XNOR2_X1  g715(.A(KEYINPUT120), .B(KEYINPUT55), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n901), .B(new_n902), .ZN(new_n903));
  AND3_X1   g717(.A1(new_n898), .A2(new_n899), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n903), .B1(new_n898), .B2(new_n899), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n282), .A2(G952), .ZN(new_n906));
  NOR3_X1   g720(.A1(new_n904), .A2(new_n905), .A3(new_n906), .ZN(G51));
  XOR2_X1   g721(.A(new_n305), .B(KEYINPUT57), .Z(new_n908));
  AOI221_X4 g722(.A(KEYINPUT54), .B1(new_n877), .B2(new_n878), .C1(new_n866), .C2(new_n871), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n873), .B1(new_n872), .B2(new_n879), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n908), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  OR2_X1    g725(.A1(new_n302), .A2(new_n303), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n897), .A2(G469), .A3(new_n300), .A4(new_n752), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n906), .B1(new_n913), .B2(new_n914), .ZN(G54));
  NAND4_X1  g729(.A1(new_n897), .A2(KEYINPUT58), .A3(G475), .A4(new_n300), .ZN(new_n916));
  INV_X1    g730(.A(new_n432), .ZN(new_n917));
  AND2_X1   g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n916), .A2(new_n917), .ZN(new_n919));
  NOR3_X1   g733(.A1(new_n918), .A2(new_n919), .A3(new_n906), .ZN(G60));
  INV_X1    g734(.A(new_n906), .ZN(new_n921));
  NAND2_X1  g735(.A1(G478), .A2(G902), .ZN(new_n922));
  XOR2_X1   g736(.A(new_n922), .B(KEYINPUT59), .Z(new_n923));
  AOI21_X1  g737(.A(new_n923), .B1(new_n880), .B2(new_n886), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n620), .A2(new_n621), .ZN(new_n925));
  INV_X1    g739(.A(new_n925), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n921), .B1(new_n924), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n897), .A2(KEYINPUT54), .ZN(new_n928));
  AOI211_X1 g742(.A(new_n925), .B(new_n923), .C1(new_n928), .C2(new_n880), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n927), .A2(new_n929), .ZN(G63));
  XNOR2_X1  g744(.A(KEYINPUT121), .B(KEYINPUT61), .ZN(new_n931));
  NAND2_X1  g745(.A1(G217), .A2(G902), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(KEYINPUT60), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n933), .B1(new_n872), .B2(new_n879), .ZN(new_n934));
  AND2_X1   g748(.A1(new_n652), .A2(new_n654), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n906), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n549), .A2(new_n551), .ZN(new_n937));
  AOI22_X1  g751(.A1(new_n866), .A2(new_n871), .B1(new_n878), .B2(new_n877), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n937), .B1(new_n938), .B2(new_n933), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n931), .B1(new_n936), .B2(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(new_n933), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n897), .A2(new_n935), .A3(new_n941), .ZN(new_n942));
  AND4_X1   g756(.A1(new_n921), .A2(new_n939), .A3(new_n931), .A4(new_n942), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n940), .A2(new_n943), .ZN(G66));
  AND2_X1   g758(.A1(new_n857), .A2(new_n711), .ZN(new_n945));
  AND2_X1   g759(.A1(new_n847), .A2(new_n854), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(new_n282), .ZN(new_n948));
  AND2_X1   g762(.A1(new_n447), .A2(G224), .ZN(new_n949));
  OAI211_X1 g763(.A(new_n948), .B(KEYINPUT122), .C1(new_n282), .C2(new_n949), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n950), .B1(KEYINPUT122), .B2(new_n948), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n900), .B1(G898), .B2(new_n282), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n951), .B(new_n952), .Z(G69));
  OR2_X1    g767(.A1(new_n571), .A2(new_n572), .ZN(new_n954));
  AND2_X1   g768(.A1(new_n954), .A2(new_n567), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n424), .A2(new_n425), .ZN(new_n956));
  XOR2_X1   g770(.A(new_n955), .B(new_n956), .Z(new_n957));
  OAI21_X1  g771(.A(new_n957), .B1(new_n663), .B2(new_n282), .ZN(new_n958));
  AND2_X1   g772(.A1(new_n839), .A2(new_n613), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n762), .B1(new_n778), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n671), .A2(new_n730), .ZN(new_n961));
  INV_X1    g775(.A(new_n694), .ZN(new_n962));
  OR3_X1    g776(.A1(new_n961), .A2(new_n962), .A3(KEYINPUT123), .ZN(new_n963));
  OAI21_X1  g777(.A(KEYINPUT123), .B1(new_n961), .B2(new_n962), .ZN(new_n964));
  AND2_X1   g778(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n744), .A2(new_n746), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n966), .B1(new_n785), .B2(new_n786), .ZN(new_n967));
  AND3_X1   g781(.A1(new_n960), .A2(new_n965), .A3(new_n967), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n958), .B1(new_n968), .B2(new_n282), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n963), .A2(new_n964), .A3(new_n689), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT62), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND4_X1  g786(.A1(new_n963), .A2(new_n964), .A3(KEYINPUT62), .A4(new_n689), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  AND2_X1   g788(.A1(new_n851), .A2(new_n852), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n670), .A2(new_n553), .ZN(new_n976));
  NOR4_X1   g790(.A1(new_n674), .A2(new_n975), .A3(new_n976), .A4(new_n781), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n977), .B1(new_n762), .B2(new_n778), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n974), .A2(new_n978), .A3(new_n787), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n957), .B1(new_n979), .B2(new_n282), .ZN(new_n980));
  OAI21_X1  g794(.A(KEYINPUT124), .B1(new_n969), .B2(new_n980), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n282), .B1(G227), .B2(G900), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n982), .B(KEYINPUT125), .ZN(new_n983));
  OAI211_X1 g797(.A(new_n981), .B(new_n983), .C1(KEYINPUT124), .C2(new_n980), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n982), .B1(new_n969), .B2(new_n980), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n984), .A2(new_n985), .ZN(G72));
  XNOR2_X1  g800(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n987));
  NAND2_X1  g801(.A1(G472), .A2(G902), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n987), .B(new_n988), .ZN(new_n989));
  INV_X1    g803(.A(new_n989), .ZN(new_n990));
  INV_X1    g804(.A(new_n602), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n990), .B1(new_n991), .B2(new_n580), .ZN(new_n992));
  OAI211_X1 g806(.A(new_n881), .B(new_n992), .C1(new_n883), .C2(new_n885), .ZN(new_n993));
  AND2_X1   g807(.A1(new_n993), .A2(new_n921), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n989), .B1(new_n979), .B2(new_n947), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n995), .A2(new_n681), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n960), .A2(new_n965), .A3(new_n967), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n989), .B1(new_n997), .B2(new_n947), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n998), .A2(new_n582), .A3(new_n680), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n994), .A2(new_n996), .A3(new_n999), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n1000), .A2(KEYINPUT127), .ZN(new_n1001));
  INV_X1    g815(.A(KEYINPUT127), .ZN(new_n1002));
  NAND4_X1  g816(.A1(new_n996), .A2(new_n994), .A3(new_n999), .A4(new_n1002), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1001), .A2(new_n1003), .ZN(G57));
endmodule


