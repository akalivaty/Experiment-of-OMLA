//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 0 1 1 0 1 1 0 1 0 1 0 1 0 0 1 0 0 1 1 0 1 1 1 0 1 1 0 0 1 1 1 1 0 0 1 0 0 0 1 0 0 1 0 1 1 1 1 1 1 0 0 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:46 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n712, new_n713, new_n714, new_n715, new_n716, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n747, new_n748, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n766,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n787, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n922, new_n923, new_n924, new_n925, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT73), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT70), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT2), .ZN(new_n190));
  INV_X1    g004(.A(G113), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n190), .A2(new_n191), .A3(KEYINPUT69), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT69), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n193), .B1(KEYINPUT2), .B2(G113), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(KEYINPUT2), .A2(G113), .ZN(new_n196));
  XNOR2_X1  g010(.A(G116), .B(G119), .ZN(new_n197));
  AND3_X1   g011(.A1(new_n195), .A2(new_n196), .A3(new_n197), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n197), .B1(new_n195), .B2(new_n196), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n189), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  NOR3_X1   g014(.A1(new_n193), .A2(KEYINPUT2), .A3(G113), .ZN(new_n201));
  AOI21_X1  g015(.A(KEYINPUT69), .B1(new_n190), .B2(new_n191), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n196), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(new_n197), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  AOI22_X1  g019(.A1(new_n192), .A2(new_n194), .B1(KEYINPUT2), .B2(G113), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(new_n197), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n205), .A2(KEYINPUT70), .A3(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n200), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(new_n209), .ZN(new_n210));
  AND2_X1   g024(.A1(KEYINPUT0), .A2(G128), .ZN(new_n211));
  INV_X1    g025(.A(G146), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G143), .ZN(new_n213));
  INV_X1    g027(.A(G143), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G146), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n211), .B1(new_n213), .B2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT64), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT0), .ZN(new_n218));
  INV_X1    g032(.A(G128), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n217), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  OAI21_X1  g034(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n216), .A2(new_n222), .A3(KEYINPUT65), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT66), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n224), .B1(new_n214), .B2(G146), .ZN(new_n225));
  NOR3_X1   g039(.A1(new_n212), .A2(KEYINPUT66), .A3(G143), .ZN(new_n226));
  OAI211_X1 g040(.A(new_n213), .B(new_n211), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  AND2_X1   g041(.A1(new_n223), .A2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT11), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n229), .A2(G137), .ZN(new_n230));
  AND2_X1   g044(.A1(KEYINPUT67), .A2(G134), .ZN(new_n231));
  NOR2_X1   g045(.A1(KEYINPUT67), .A2(G134), .ZN(new_n232));
  NOR3_X1   g046(.A1(new_n230), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(G137), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n234), .A2(KEYINPUT11), .A3(G134), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n229), .A2(G137), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  OAI21_X1  g051(.A(G131), .B1(new_n233), .B2(new_n237), .ZN(new_n238));
  OR2_X1    g052(.A1(KEYINPUT67), .A2(G134), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n234), .A2(KEYINPUT11), .ZN(new_n240));
  NAND2_X1  g054(.A1(KEYINPUT67), .A2(G134), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n239), .A2(new_n240), .A3(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(G131), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n242), .A2(new_n243), .A3(new_n235), .A4(new_n236), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n238), .A2(new_n244), .ZN(new_n245));
  AOI21_X1  g059(.A(KEYINPUT65), .B1(new_n216), .B2(new_n222), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n228), .A2(new_n245), .A3(new_n247), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n214), .A2(G146), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT1), .ZN(new_n250));
  OAI21_X1  g064(.A(G128), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n213), .A2(new_n215), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n219), .A2(KEYINPUT1), .ZN(new_n254));
  OAI211_X1 g068(.A(new_n213), .B(new_n254), .C1(new_n225), .C2(new_n226), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT68), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n243), .B1(G134), .B2(G137), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n239), .A2(new_n241), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n258), .B1(new_n259), .B2(G137), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n256), .A2(new_n257), .A3(new_n244), .A4(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n244), .A2(new_n260), .ZN(new_n262));
  OAI21_X1  g076(.A(KEYINPUT66), .B1(new_n212), .B2(G143), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n224), .A2(new_n214), .A3(G146), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n249), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  AOI22_X1  g079(.A1(new_n265), .A2(new_n254), .B1(new_n251), .B2(new_n252), .ZN(new_n266));
  OAI21_X1  g080(.A(KEYINPUT68), .B1(new_n262), .B2(new_n266), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n248), .A2(new_n261), .A3(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT71), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n269), .B1(new_n262), .B2(new_n266), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n256), .A2(KEYINPUT71), .A3(new_n244), .A4(new_n260), .ZN(new_n271));
  AND2_X1   g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n223), .A2(new_n227), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n273), .A2(new_n246), .ZN(new_n274));
  AOI22_X1  g088(.A1(new_n274), .A2(new_n245), .B1(new_n200), .B2(new_n208), .ZN(new_n275));
  AOI22_X1  g089(.A1(new_n210), .A2(new_n268), .B1(new_n272), .B2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT28), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n188), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  AND2_X1   g092(.A1(new_n268), .A2(new_n210), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n248), .A2(new_n209), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n270), .A2(new_n271), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  OAI211_X1 g096(.A(KEYINPUT73), .B(KEYINPUT28), .C1(new_n279), .C2(new_n282), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n262), .A2(new_n266), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n277), .B1(new_n280), .B2(new_n284), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n278), .A2(new_n283), .A3(new_n285), .ZN(new_n286));
  NOR2_X1   g100(.A1(G237), .A2(G953), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(G210), .ZN(new_n288));
  XNOR2_X1  g102(.A(new_n288), .B(KEYINPUT27), .ZN(new_n289));
  XNOR2_X1  g103(.A(KEYINPUT26), .B(G101), .ZN(new_n290));
  XNOR2_X1  g104(.A(new_n289), .B(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n291), .B1(new_n280), .B2(new_n281), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT72), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT30), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n268), .A2(new_n296), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n248), .A2(KEYINPUT30), .A3(new_n270), .A4(new_n271), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n297), .A2(new_n210), .A3(new_n298), .ZN(new_n299));
  OAI211_X1 g113(.A(KEYINPUT72), .B(new_n291), .C1(new_n280), .C2(new_n281), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n295), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT31), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND4_X1  g117(.A1(new_n295), .A2(new_n299), .A3(KEYINPUT31), .A4(new_n300), .ZN(new_n304));
  AOI22_X1  g118(.A1(new_n286), .A2(new_n292), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(G472), .ZN(new_n306));
  INV_X1    g120(.A(G902), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n306), .A2(new_n307), .A3(KEYINPUT74), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT74), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n309), .B1(G472), .B2(G902), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n187), .B1(new_n305), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n286), .A2(new_n292), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n303), .A2(new_n304), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NOR2_X1   g130(.A1(new_n312), .A2(new_n187), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(new_n285), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n319), .A2(new_n292), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n278), .A2(new_n283), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n272), .A2(new_n275), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n299), .A2(new_n322), .ZN(new_n323));
  AOI21_X1  g137(.A(KEYINPUT29), .B1(new_n323), .B2(new_n292), .ZN(new_n324));
  AND2_X1   g138(.A1(new_n321), .A2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(new_n248), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n210), .B1(new_n326), .B2(new_n281), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n277), .B1(new_n327), .B2(new_n322), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n285), .A2(KEYINPUT29), .A3(new_n291), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n307), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  OAI21_X1  g144(.A(G472), .B1(new_n325), .B2(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n313), .A2(new_n318), .A3(new_n331), .ZN(new_n332));
  XNOR2_X1  g146(.A(KEYINPUT9), .B(G234), .ZN(new_n333));
  OAI21_X1  g147(.A(G221), .B1(new_n333), .B2(G902), .ZN(new_n334));
  INV_X1    g148(.A(G469), .ZN(new_n335));
  INV_X1    g149(.A(new_n245), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n336), .A2(KEYINPUT82), .ZN(new_n337));
  INV_X1    g151(.A(G101), .ZN(new_n338));
  INV_X1    g152(.A(G107), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(G104), .ZN(new_n340));
  INV_X1    g154(.A(G104), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(G107), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n338), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT3), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n344), .A2(new_n339), .A3(G104), .ZN(new_n345));
  AND2_X1   g159(.A1(new_n345), .A2(new_n342), .ZN(new_n346));
  XOR2_X1   g160(.A(KEYINPUT80), .B(G101), .Z(new_n347));
  OAI21_X1  g161(.A(KEYINPUT3), .B1(new_n341), .B2(G107), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n346), .A2(KEYINPUT81), .A3(new_n347), .A4(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT81), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n348), .A2(new_n345), .A3(new_n342), .ZN(new_n351));
  XNOR2_X1  g165(.A(KEYINPUT80), .B(G101), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n350), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n343), .B1(new_n349), .B2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(new_n251), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n255), .B1(new_n355), .B2(new_n265), .ZN(new_n356));
  AND2_X1   g170(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n354), .A2(new_n256), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n337), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(KEYINPUT12), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n354), .A2(new_n356), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT10), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n266), .A2(new_n362), .ZN(new_n363));
  AOI22_X1  g177(.A1(new_n361), .A2(new_n362), .B1(new_n354), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n349), .A2(new_n353), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n351), .A2(KEYINPUT79), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT79), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n348), .A2(new_n345), .A3(new_n367), .A4(new_n342), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n366), .A2(G101), .A3(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n365), .A2(KEYINPUT4), .A3(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT4), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n366), .A2(new_n371), .A3(G101), .A4(new_n368), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n370), .A2(new_n274), .A3(new_n372), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n364), .A2(new_n336), .A3(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT12), .ZN(new_n375));
  OAI211_X1 g189(.A(new_n375), .B(new_n337), .C1(new_n357), .C2(new_n358), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n360), .A2(new_n374), .A3(new_n376), .ZN(new_n377));
  XNOR2_X1  g191(.A(G110), .B(G140), .ZN(new_n378));
  INV_X1    g192(.A(G227), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n379), .A2(G953), .ZN(new_n380));
  XNOR2_X1  g194(.A(new_n378), .B(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n377), .A2(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n336), .B1(new_n364), .B2(new_n373), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(new_n381), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n384), .A2(new_n374), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n382), .A2(new_n386), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n335), .B1(new_n387), .B2(new_n307), .ZN(new_n388));
  INV_X1    g202(.A(new_n374), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n381), .B1(new_n389), .B2(new_n383), .ZN(new_n390));
  NAND4_X1  g204(.A1(new_n360), .A2(new_n374), .A3(new_n385), .A4(new_n376), .ZN(new_n391));
  AOI211_X1 g205(.A(G469), .B(G902), .C1(new_n390), .C2(new_n391), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n334), .B1(new_n388), .B2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(G475), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT76), .ZN(new_n395));
  INV_X1    g209(.A(G140), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(G125), .ZN(new_n397));
  INV_X1    g211(.A(G125), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(G140), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n397), .A2(new_n399), .A3(KEYINPUT16), .ZN(new_n400));
  OR3_X1    g214(.A1(new_n398), .A2(KEYINPUT16), .A3(G140), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n395), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NOR3_X1   g216(.A1(new_n398), .A2(KEYINPUT16), .A3(G140), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n403), .A2(KEYINPUT76), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n212), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n401), .A2(new_n395), .ZN(new_n406));
  XNOR2_X1  g220(.A(G125), .B(G140), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n403), .B1(new_n407), .B2(KEYINPUT16), .ZN(new_n408));
  OAI211_X1 g222(.A(G146), .B(new_n406), .C1(new_n408), .C2(new_n395), .ZN(new_n409));
  INV_X1    g223(.A(G237), .ZN(new_n410));
  INV_X1    g224(.A(G953), .ZN(new_n411));
  AND4_X1   g225(.A1(G143), .A2(new_n410), .A3(new_n411), .A4(G214), .ZN(new_n412));
  AOI21_X1  g226(.A(G143), .B1(new_n287), .B2(G214), .ZN(new_n413));
  OAI21_X1  g227(.A(G131), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT17), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n410), .A2(new_n411), .A3(G214), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(new_n214), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n287), .A2(G143), .A3(G214), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n417), .A2(new_n243), .A3(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n414), .A2(new_n415), .A3(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n417), .A2(new_n418), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n421), .A2(KEYINPUT17), .A3(G131), .ZN(new_n422));
  NAND4_X1  g236(.A1(new_n405), .A2(new_n409), .A3(new_n420), .A4(new_n422), .ZN(new_n423));
  XNOR2_X1  g237(.A(G113), .B(G122), .ZN(new_n424));
  XNOR2_X1  g238(.A(new_n424), .B(new_n341), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n412), .A2(new_n413), .ZN(new_n426));
  NAND2_X1  g240(.A1(KEYINPUT18), .A2(G131), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n397), .A2(new_n399), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(G146), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n407), .A2(new_n212), .ZN(new_n430));
  AOI22_X1  g244(.A1(new_n426), .A2(new_n427), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(new_n427), .ZN(new_n432));
  AOI21_X1  g246(.A(KEYINPUT88), .B1(new_n421), .B2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT88), .ZN(new_n434));
  AOI211_X1 g248(.A(new_n434), .B(new_n427), .C1(new_n417), .C2(new_n418), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n431), .B1(new_n433), .B2(new_n435), .ZN(new_n436));
  AND3_X1   g250(.A1(new_n423), .A2(new_n425), .A3(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT89), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n423), .A2(new_n436), .ZN(new_n440));
  INV_X1    g254(.A(new_n425), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n439), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  AOI211_X1 g256(.A(KEYINPUT89), .B(new_n425), .C1(new_n423), .C2(new_n436), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n438), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n394), .B1(new_n444), .B2(new_n307), .ZN(new_n445));
  NOR2_X1   g259(.A1(G475), .A2(G902), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n414), .A2(new_n419), .ZN(new_n447));
  XNOR2_X1  g261(.A(new_n428), .B(KEYINPUT19), .ZN(new_n448));
  OAI211_X1 g262(.A(new_n409), .B(new_n447), .C1(G146), .C2(new_n448), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n425), .B1(new_n449), .B2(new_n436), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n446), .B1(new_n437), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(KEYINPUT20), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT20), .ZN(new_n453));
  OAI211_X1 g267(.A(new_n453), .B(new_n446), .C1(new_n437), .C2(new_n450), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n445), .B1(new_n452), .B2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(G478), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n456), .A2(KEYINPUT15), .ZN(new_n457));
  INV_X1    g271(.A(G122), .ZN(new_n458));
  OAI21_X1  g272(.A(KEYINPUT91), .B1(new_n458), .B2(G116), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT91), .ZN(new_n460));
  INV_X1    g274(.A(G116), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n460), .A2(new_n461), .A3(G122), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT14), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n459), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  OAI21_X1  g278(.A(KEYINPUT90), .B1(new_n461), .B2(G122), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT90), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n466), .A2(new_n458), .A3(G116), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n464), .A2(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n463), .B1(new_n459), .B2(new_n462), .ZN(new_n470));
  OAI21_X1  g284(.A(G107), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n231), .A2(new_n232), .ZN(new_n472));
  XNOR2_X1  g286(.A(G128), .B(G143), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n472), .B(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n459), .A2(new_n462), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT92), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n468), .A2(new_n475), .A3(new_n476), .A4(new_n339), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n468), .A2(new_n475), .A3(new_n339), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(KEYINPUT92), .ZN(new_n479));
  NAND4_X1  g293(.A1(new_n471), .A2(new_n474), .A3(new_n477), .A4(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n473), .A2(KEYINPUT13), .ZN(new_n481));
  NOR3_X1   g295(.A1(new_n219), .A2(KEYINPUT13), .A3(G143), .ZN(new_n482));
  INV_X1    g296(.A(G134), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  AOI22_X1  g298(.A1(new_n481), .A2(new_n484), .B1(new_n472), .B2(new_n473), .ZN(new_n485));
  INV_X1    g299(.A(new_n478), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n339), .B1(new_n468), .B2(new_n475), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n485), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(G217), .ZN(new_n489));
  NOR3_X1   g303(.A1(new_n333), .A2(new_n489), .A3(G953), .ZN(new_n490));
  AND3_X1   g304(.A1(new_n480), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n490), .B1(new_n480), .B2(new_n488), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n307), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n457), .B1(new_n493), .B2(KEYINPUT93), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n480), .A2(new_n488), .ZN(new_n495));
  INV_X1    g309(.A(new_n490), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n480), .A2(new_n488), .A3(new_n490), .ZN(new_n498));
  AOI21_X1  g312(.A(G902), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT93), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n493), .A2(KEYINPUT93), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n494), .B1(new_n503), .B2(new_n457), .ZN(new_n504));
  NAND2_X1  g318(.A1(G234), .A2(G237), .ZN(new_n505));
  AND3_X1   g319(.A1(new_n505), .A2(G952), .A3(new_n411), .ZN(new_n506));
  XOR2_X1   g320(.A(KEYINPUT21), .B(G898), .Z(new_n507));
  XNOR2_X1  g321(.A(new_n507), .B(KEYINPUT94), .ZN(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  AND3_X1   g323(.A1(new_n505), .A2(G902), .A3(G953), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n506), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n455), .A2(new_n504), .A3(new_n512), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n393), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n489), .B1(G234), .B2(new_n307), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT77), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n219), .A2(KEYINPUT23), .A3(G119), .ZN(new_n517));
  INV_X1    g331(.A(G119), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(G128), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n518), .A2(G128), .ZN(new_n520));
  OAI211_X1 g334(.A(new_n517), .B(new_n519), .C1(new_n520), .C2(KEYINPUT23), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(G110), .ZN(new_n522));
  XOR2_X1   g336(.A(KEYINPUT24), .B(G110), .Z(new_n523));
  XNOR2_X1  g337(.A(G119), .B(G128), .ZN(new_n524));
  AND3_X1   g338(.A1(new_n523), .A2(KEYINPUT75), .A3(new_n524), .ZN(new_n525));
  AOI21_X1  g339(.A(KEYINPUT75), .B1(new_n523), .B2(new_n524), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n522), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n527), .B1(new_n405), .B2(new_n409), .ZN(new_n528));
  OAI22_X1  g342(.A1(new_n521), .A2(G110), .B1(new_n523), .B2(new_n524), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n409), .A2(new_n529), .A3(new_n430), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n516), .B1(new_n528), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n405), .A2(new_n409), .ZN(new_n533));
  OR2_X1    g347(.A1(new_n525), .A2(new_n526), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n533), .A2(new_n522), .A3(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n535), .A2(KEYINPUT77), .A3(new_n530), .ZN(new_n536));
  XNOR2_X1  g350(.A(KEYINPUT22), .B(G137), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n411), .A2(G221), .A3(G234), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n537), .B(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n532), .A2(new_n536), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n535), .A2(new_n530), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n542), .A2(new_n516), .A3(new_n539), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(KEYINPUT25), .B1(new_n544), .B2(new_n307), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT25), .ZN(new_n546));
  AOI211_X1 g360(.A(new_n546), .B(G902), .C1(new_n541), .C2(new_n543), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n515), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT78), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  OAI211_X1 g364(.A(KEYINPUT78), .B(new_n515), .C1(new_n545), .C2(new_n547), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n515), .A2(G902), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n544), .A2(new_n552), .ZN(new_n553));
  AND3_X1   g367(.A1(new_n550), .A2(new_n551), .A3(new_n553), .ZN(new_n554));
  OAI21_X1  g368(.A(G214), .B1(G237), .B2(G902), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  OAI21_X1  g370(.A(G210), .B1(G237), .B2(G902), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT86), .ZN(new_n559));
  OAI21_X1  g373(.A(G125), .B1(new_n273), .B2(new_n246), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n266), .A2(new_n398), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n559), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n247), .A2(new_n227), .A3(new_n223), .ZN(new_n563));
  AOI21_X1  g377(.A(KEYINPUT86), .B1(new_n563), .B2(G125), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n411), .A2(G224), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  OAI211_X1 g381(.A(G224), .B(new_n411), .C1(new_n562), .C2(new_n564), .ZN(new_n568));
  AND2_X1   g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n197), .A2(KEYINPUT5), .ZN(new_n570));
  NOR3_X1   g384(.A1(new_n461), .A2(KEYINPUT5), .A3(G119), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n571), .A2(new_n191), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n198), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(new_n354), .ZN(new_n574));
  AND3_X1   g388(.A1(new_n365), .A2(KEYINPUT4), .A3(new_n369), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n200), .A2(new_n208), .A3(new_n372), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n574), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT83), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  OAI211_X1 g393(.A(KEYINPUT83), .B(new_n574), .C1(new_n575), .C2(new_n576), .ZN(new_n580));
  XOR2_X1   g394(.A(G110), .B(G122), .Z(new_n581));
  XNOR2_X1  g395(.A(new_n581), .B(KEYINPUT84), .ZN(new_n582));
  XOR2_X1   g396(.A(new_n582), .B(KEYINPUT85), .Z(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n579), .A2(new_n580), .A3(new_n584), .ZN(new_n585));
  OAI211_X1 g399(.A(new_n574), .B(new_n582), .C1(new_n575), .C2(new_n576), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(KEYINPUT6), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n583), .B1(new_n577), .B2(new_n578), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n589), .A2(KEYINPUT6), .A3(new_n580), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n569), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n582), .B(KEYINPUT8), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n573), .A2(new_n354), .A3(KEYINPUT87), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n593), .B1(new_n354), .B2(new_n573), .ZN(new_n594));
  AOI21_X1  g408(.A(KEYINPUT87), .B1(new_n573), .B2(new_n354), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n592), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n566), .A2(KEYINPUT7), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n598), .B1(new_n562), .B2(new_n564), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  NOR3_X1   g414(.A1(new_n562), .A2(new_n564), .A3(new_n598), .ZN(new_n601));
  OAI211_X1 g415(.A(new_n596), .B(new_n586), .C1(new_n600), .C2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(new_n307), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n558), .B1(new_n591), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n567), .A2(new_n568), .ZN(new_n605));
  AND3_X1   g419(.A1(new_n589), .A2(KEYINPUT6), .A3(new_n580), .ZN(new_n606));
  AOI22_X1  g420(.A1(new_n589), .A2(new_n580), .B1(KEYINPUT6), .B2(new_n586), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n605), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n586), .ZN(new_n609));
  INV_X1    g423(.A(new_n601), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n609), .B1(new_n610), .B2(new_n599), .ZN(new_n611));
  AOI21_X1  g425(.A(G902), .B1(new_n611), .B2(new_n596), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n608), .A2(new_n557), .A3(new_n612), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n556), .B1(new_n604), .B2(new_n613), .ZN(new_n614));
  NAND4_X1  g428(.A1(new_n332), .A2(new_n514), .A3(new_n554), .A4(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(new_n352), .ZN(G3));
  NAND2_X1  g430(.A1(new_n316), .A2(new_n307), .ZN(new_n617));
  AOI22_X1  g431(.A1(new_n617), .A2(G472), .B1(new_n311), .B2(new_n316), .ZN(new_n618));
  INV_X1    g432(.A(new_n334), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n335), .A2(new_n307), .ZN(new_n620));
  AND2_X1   g434(.A1(new_n382), .A2(new_n386), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n620), .B1(new_n621), .B2(G469), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n390), .A2(new_n391), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n623), .A2(new_n335), .A3(new_n307), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n619), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n618), .A2(new_n554), .A3(new_n625), .ZN(new_n626));
  AOI211_X1 g440(.A(new_n556), .B(new_n511), .C1(new_n604), .C2(new_n613), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n452), .A2(new_n454), .ZN(new_n628));
  AND2_X1   g442(.A1(new_n444), .A2(new_n307), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n628), .B1(new_n629), .B2(new_n394), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n456), .A2(new_n307), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n631), .B1(new_n499), .B2(new_n456), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT95), .ZN(new_n633));
  OAI21_X1  g447(.A(KEYINPUT33), .B1(new_n491), .B2(new_n492), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT33), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n497), .A2(new_n635), .A3(new_n498), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n634), .A2(new_n636), .A3(G478), .ZN(new_n637));
  AND3_X1   g451(.A1(new_n632), .A2(new_n633), .A3(new_n637), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n633), .B1(new_n632), .B2(new_n637), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n630), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n627), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n626), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(KEYINPUT34), .B(G104), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G6));
  INV_X1    g459(.A(new_n504), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT96), .ZN(new_n647));
  OR2_X1    g461(.A1(new_n454), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n452), .A2(new_n647), .A3(new_n454), .ZN(new_n649));
  OAI211_X1 g463(.A(new_n648), .B(new_n649), .C1(new_n445), .C2(KEYINPUT97), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT97), .ZN(new_n651));
  AOI211_X1 g465(.A(new_n651), .B(new_n394), .C1(new_n444), .C2(new_n307), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n627), .A2(new_n646), .A3(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n626), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(KEYINPUT35), .B(G107), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G9));
  INV_X1    g471(.A(KEYINPUT36), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n539), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(KEYINPUT99), .ZN(new_n660));
  XOR2_X1   g474(.A(new_n660), .B(KEYINPUT98), .Z(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(new_n542), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(new_n552), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n550), .A2(new_n551), .A3(new_n663), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n514), .A2(new_n618), .A3(new_n614), .A4(new_n664), .ZN(new_n665));
  XOR2_X1   g479(.A(KEYINPUT37), .B(G110), .Z(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(G12));
  INV_X1    g481(.A(KEYINPUT101), .ZN(new_n668));
  INV_X1    g482(.A(G900), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n510), .A2(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(new_n506), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  NOR4_X1   g487(.A1(new_n650), .A2(new_n504), .A3(new_n652), .A4(new_n673), .ZN(new_n674));
  AND3_X1   g488(.A1(new_n614), .A2(new_n674), .A3(KEYINPUT100), .ZN(new_n675));
  AOI21_X1  g489(.A(KEYINPUT100), .B1(new_n614), .B2(new_n674), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g491(.A(KEYINPUT32), .B1(new_n316), .B2(new_n311), .ZN(new_n678));
  INV_X1    g492(.A(new_n317), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n330), .B1(new_n321), .B2(new_n324), .ZN(new_n680));
  OAI22_X1  g494(.A1(new_n305), .A2(new_n679), .B1(new_n680), .B2(new_n306), .ZN(new_n681));
  OAI211_X1 g495(.A(new_n625), .B(new_n664), .C1(new_n678), .C2(new_n681), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n668), .B1(new_n677), .B2(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n614), .A2(new_n674), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT100), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n614), .A2(new_n674), .A3(KEYINPUT100), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(new_n682), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n688), .A2(new_n689), .A3(KEYINPUT101), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n683), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G128), .ZN(G30));
  NAND2_X1  g506(.A1(new_n604), .A2(new_n613), .ZN(new_n693));
  XOR2_X1   g507(.A(new_n693), .B(KEYINPUT38), .Z(new_n694));
  INV_X1    g508(.A(KEYINPUT40), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n672), .B(KEYINPUT39), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n625), .A2(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n694), .B1(new_n695), .B2(new_n698), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n305), .A2(new_n679), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n678), .A2(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(new_n301), .ZN(new_n702));
  AND2_X1   g516(.A1(new_n327), .A2(new_n322), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n703), .A2(new_n291), .ZN(new_n704));
  OAI21_X1  g518(.A(new_n307), .B1(new_n702), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(G472), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n664), .B1(new_n701), .B2(new_n706), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n646), .A2(new_n630), .A3(new_n555), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n708), .B1(new_n697), .B2(KEYINPUT40), .ZN(new_n709));
  AND3_X1   g523(.A1(new_n699), .A2(new_n707), .A3(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(new_n214), .ZN(G45));
  NOR2_X1   g525(.A1(new_n640), .A2(new_n673), .ZN(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n693), .A2(new_n555), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n689), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G146), .ZN(G48));
  NAND2_X1  g531(.A1(new_n623), .A2(new_n307), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(G469), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n719), .A2(new_n334), .A3(new_n624), .ZN(new_n720));
  INV_X1    g534(.A(new_n720), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n332), .A2(new_n554), .A3(new_n721), .ZN(new_n722));
  OR2_X1    g536(.A1(new_n722), .A2(new_n642), .ZN(new_n723));
  XNOR2_X1  g537(.A(KEYINPUT41), .B(G113), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n723), .B(new_n724), .ZN(G15));
  NOR2_X1   g539(.A1(new_n722), .A2(new_n654), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(new_n461), .ZN(G18));
  INV_X1    g541(.A(new_n513), .ZN(new_n728));
  OAI211_X1 g542(.A(new_n664), .B(new_n728), .C1(new_n681), .C2(new_n678), .ZN(new_n729));
  OAI21_X1  g543(.A(KEYINPUT102), .B1(new_n714), .B2(new_n720), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT102), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n721), .A2(new_n731), .A3(new_n614), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n729), .B1(new_n730), .B2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(new_n518), .ZN(G21));
  NOR2_X1   g548(.A1(new_n720), .A2(new_n511), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n708), .B1(new_n604), .B2(new_n613), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n311), .B(KEYINPUT103), .ZN(new_n737));
  INV_X1    g551(.A(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT104), .ZN(new_n739));
  OAI211_X1 g553(.A(new_n739), .B(new_n285), .C1(new_n703), .C2(new_n277), .ZN(new_n740));
  OAI21_X1  g554(.A(KEYINPUT104), .B1(new_n328), .B2(new_n319), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n740), .A2(new_n292), .A3(new_n741), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n738), .B1(new_n742), .B2(new_n315), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n743), .B1(new_n617), .B2(G472), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n735), .A2(new_n736), .A3(new_n554), .A4(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G122), .ZN(G24));
  NAND3_X1  g560(.A1(new_n744), .A2(new_n664), .A3(new_n712), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n747), .B1(new_n732), .B2(new_n730), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(new_n398), .ZN(G27));
  INV_X1    g563(.A(KEYINPUT106), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n750), .B1(new_n678), .B2(new_n700), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n313), .A2(KEYINPUT106), .A3(new_n318), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n751), .A2(new_n331), .A3(new_n752), .ZN(new_n753));
  OR2_X1    g567(.A1(new_n638), .A2(new_n639), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n754), .A2(KEYINPUT42), .A3(new_n630), .A4(new_n672), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n604), .A2(new_n613), .A3(new_n555), .ZN(new_n756));
  NOR3_X1   g570(.A1(new_n755), .A2(new_n393), .A3(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n753), .A2(new_n554), .A3(new_n757), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n756), .A2(new_n393), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n759), .A2(new_n332), .A3(new_n554), .A4(new_n712), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT42), .ZN(new_n761));
  AND3_X1   g575(.A1(new_n760), .A2(KEYINPUT105), .A3(new_n761), .ZN(new_n762));
  AOI21_X1  g576(.A(KEYINPUT105), .B1(new_n760), .B2(new_n761), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n758), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G131), .ZN(G33));
  NAND4_X1  g579(.A1(new_n759), .A2(new_n332), .A3(new_n554), .A4(new_n674), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G134), .ZN(G36));
  NAND2_X1  g581(.A1(new_n754), .A2(new_n455), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT43), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n768), .B(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(new_n618), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n770), .A2(new_n771), .A3(new_n664), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT44), .ZN(new_n773));
  OR2_X1    g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n621), .A2(KEYINPUT45), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT45), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n335), .B1(new_n387), .B2(new_n776), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n620), .B1(new_n775), .B2(new_n777), .ZN(new_n778));
  AND2_X1   g592(.A1(new_n778), .A2(KEYINPUT46), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n624), .B1(new_n778), .B2(KEYINPUT46), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n334), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(new_n696), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n756), .B1(new_n772), .B2(new_n773), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n774), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(G137), .ZN(G39));
  INV_X1    g600(.A(KEYINPUT47), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n781), .B(new_n787), .ZN(new_n788));
  NOR4_X1   g602(.A1(new_n713), .A2(new_n332), .A3(new_n554), .A4(new_n756), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G140), .ZN(G42));
  INV_X1    g605(.A(G952), .ZN(new_n792));
  AND2_X1   g606(.A1(new_n701), .A2(new_n706), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n720), .A2(new_n756), .ZN(new_n794));
  AND4_X1   g608(.A1(new_n554), .A2(new_n793), .A3(new_n506), .A4(new_n794), .ZN(new_n795));
  AOI211_X1 g609(.A(new_n792), .B(G953), .C1(new_n795), .C2(new_n641), .ZN(new_n796));
  AND3_X1   g610(.A1(new_n770), .A2(new_n506), .A3(new_n794), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n753), .A2(new_n554), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  XOR2_X1   g613(.A(KEYINPUT112), .B(KEYINPUT48), .Z(new_n800));
  OR2_X1    g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n799), .A2(new_n800), .ZN(new_n802));
  AND4_X1   g616(.A1(new_n554), .A2(new_n770), .A3(new_n506), .A4(new_n744), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n730), .A2(new_n732), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n796), .A2(new_n801), .A3(new_n802), .A4(new_n805), .ZN(new_n806));
  AND3_X1   g620(.A1(new_n694), .A2(new_n556), .A3(new_n721), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n803), .A2(new_n807), .ZN(new_n808));
  OR3_X1    g622(.A1(new_n808), .A2(KEYINPUT111), .A3(KEYINPUT50), .ZN(new_n809));
  INV_X1    g623(.A(new_n756), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n719), .A2(new_n624), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n811), .A2(new_n334), .ZN(new_n812));
  OAI211_X1 g626(.A(new_n810), .B(new_n803), .C1(new_n788), .C2(new_n812), .ZN(new_n813));
  XOR2_X1   g627(.A(KEYINPUT111), .B(KEYINPUT50), .Z(new_n814));
  NAND2_X1  g628(.A1(new_n744), .A2(new_n664), .ZN(new_n815));
  INV_X1    g629(.A(new_n815), .ZN(new_n816));
  AOI22_X1  g630(.A1(new_n808), .A2(new_n814), .B1(new_n816), .B2(new_n797), .ZN(new_n817));
  INV_X1    g631(.A(new_n754), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n795), .A2(new_n455), .A3(new_n818), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n809), .A2(new_n813), .A3(new_n817), .A4(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT51), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n806), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n822), .B1(new_n821), .B2(new_n820), .ZN(new_n823));
  OR2_X1    g637(.A1(new_n823), .A2(KEYINPUT113), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n745), .B1(new_n722), .B2(new_n642), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n825), .A2(new_n726), .A3(new_n733), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n759), .A2(new_n664), .A3(new_n712), .A4(new_n744), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n653), .A2(new_n504), .A3(new_n672), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT108), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n653), .A2(KEYINPUT108), .A3(new_n504), .A4(new_n672), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n830), .A2(new_n810), .A3(new_n831), .ZN(new_n832));
  OAI211_X1 g646(.A(new_n766), .B(new_n827), .C1(new_n832), .C2(new_n682), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT107), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n640), .A2(new_n834), .ZN(new_n835));
  OAI211_X1 g649(.A(new_n630), .B(KEYINPUT107), .C1(new_n638), .C2(new_n639), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n646), .A2(new_n455), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n835), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n838), .A2(new_n627), .ZN(new_n839));
  OAI211_X1 g653(.A(new_n615), .B(new_n665), .C1(new_n626), .C2(new_n839), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n833), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n764), .A2(new_n826), .A3(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(new_n748), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n455), .A2(new_n504), .A3(new_n556), .ZN(new_n844));
  XOR2_X1   g658(.A(new_n672), .B(KEYINPUT109), .Z(new_n845));
  AND4_X1   g659(.A1(new_n693), .A2(new_n625), .A3(new_n844), .A4(new_n845), .ZN(new_n846));
  AOI22_X1  g660(.A1(new_n715), .A2(new_n689), .B1(new_n707), .B2(new_n846), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n677), .A2(new_n668), .A3(new_n682), .ZN(new_n848));
  AOI21_X1  g662(.A(KEYINPUT101), .B1(new_n688), .B2(new_n689), .ZN(new_n849));
  OAI211_X1 g663(.A(new_n843), .B(new_n847), .C1(new_n848), .C2(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT52), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n748), .B1(new_n683), .B2(new_n690), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n853), .A2(KEYINPUT52), .A3(new_n847), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n842), .B1(new_n852), .B2(new_n854), .ZN(new_n855));
  XNOR2_X1  g669(.A(new_n855), .B(KEYINPUT53), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(KEYINPUT54), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n852), .A2(new_n854), .ZN(new_n858));
  INV_X1    g672(.A(new_n858), .ZN(new_n859));
  AND3_X1   g673(.A1(new_n753), .A2(new_n554), .A3(new_n757), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n760), .A2(new_n761), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT105), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n760), .A2(KEYINPUT105), .A3(new_n761), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n860), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  OR2_X1    g679(.A1(new_n722), .A2(new_n654), .ZN(new_n866));
  INV_X1    g680(.A(new_n729), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n804), .A2(new_n867), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n866), .A2(new_n723), .A3(new_n868), .A4(new_n745), .ZN(new_n869));
  OAI21_X1  g683(.A(KEYINPUT110), .B1(new_n865), .B2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT110), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n764), .A2(new_n826), .A3(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT53), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n833), .A2(new_n840), .A3(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n870), .A2(new_n872), .A3(new_n874), .ZN(new_n875));
  OAI22_X1  g689(.A1(new_n859), .A2(new_n875), .B1(new_n855), .B2(KEYINPUT53), .ZN(new_n876));
  OR2_X1    g690(.A1(new_n876), .A2(KEYINPUT54), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n823), .A2(KEYINPUT113), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n824), .A2(new_n857), .A3(new_n877), .A4(new_n878), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n879), .B1(G952), .B2(G953), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n811), .A2(KEYINPUT49), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n811), .A2(KEYINPUT49), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n334), .A2(new_n555), .ZN(new_n883));
  NOR4_X1   g697(.A1(new_n881), .A2(new_n882), .A3(new_n768), .A4(new_n883), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n884), .A2(new_n554), .A3(new_n793), .A4(new_n694), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n880), .A2(new_n885), .ZN(G75));
  NOR2_X1   g700(.A1(new_n411), .A2(G952), .ZN(new_n887));
  XOR2_X1   g701(.A(new_n887), .B(KEYINPUT115), .Z(new_n888));
  INV_X1    g702(.A(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(G210), .A2(G902), .ZN(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  AOI21_X1  g705(.A(KEYINPUT56), .B1(new_n876), .B2(new_n891), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n588), .A2(new_n590), .A3(new_n569), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n608), .A2(new_n893), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n894), .B(KEYINPUT55), .ZN(new_n895));
  INV_X1    g709(.A(new_n895), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n889), .B1(new_n892), .B2(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT114), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT56), .ZN(new_n899));
  AND3_X1   g713(.A1(new_n870), .A2(new_n872), .A3(new_n874), .ZN(new_n900));
  AND3_X1   g714(.A1(new_n764), .A2(new_n826), .A3(new_n841), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n850), .A2(new_n851), .ZN(new_n902));
  AOI21_X1  g716(.A(KEYINPUT52), .B1(new_n853), .B2(new_n847), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n901), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  AOI22_X1  g718(.A1(new_n858), .A2(new_n900), .B1(new_n904), .B2(new_n873), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n899), .B1(new_n905), .B2(new_n890), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n898), .B1(new_n906), .B2(new_n895), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n892), .A2(KEYINPUT114), .A3(new_n896), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n897), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT116), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  OAI211_X1 g725(.A(KEYINPUT116), .B(new_n897), .C1(new_n907), .C2(new_n908), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n911), .A2(new_n912), .ZN(G51));
  XNOR2_X1  g727(.A(new_n876), .B(KEYINPUT54), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n620), .B(KEYINPUT57), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n916), .A2(new_n623), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n905), .A2(new_n307), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n918), .A2(new_n775), .A3(new_n777), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n887), .B1(new_n917), .B2(new_n919), .ZN(G54));
  NAND3_X1  g734(.A1(new_n918), .A2(KEYINPUT58), .A3(G475), .ZN(new_n921));
  OR2_X1    g735(.A1(new_n437), .A2(new_n450), .ZN(new_n922));
  INV_X1    g736(.A(new_n922), .ZN(new_n923));
  AND2_X1   g737(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n921), .A2(new_n923), .ZN(new_n925));
  NOR3_X1   g739(.A1(new_n924), .A2(new_n925), .A3(new_n887), .ZN(G60));
  XOR2_X1   g740(.A(KEYINPUT118), .B(KEYINPUT59), .Z(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(new_n631), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n928), .B1(new_n877), .B2(new_n857), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n634), .A2(new_n636), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(KEYINPUT117), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n888), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(new_n931), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n933), .A2(new_n928), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n914), .A2(KEYINPUT119), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n914), .A2(new_n934), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT119), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n932), .B1(new_n935), .B2(new_n938), .ZN(G63));
  NAND2_X1  g753(.A1(G217), .A2(G902), .ZN(new_n940));
  XOR2_X1   g754(.A(new_n940), .B(KEYINPUT60), .Z(new_n941));
  NAND2_X1  g755(.A1(new_n876), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n942), .A2(KEYINPUT120), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT120), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n876), .A2(new_n944), .A3(new_n941), .ZN(new_n945));
  NAND4_X1  g759(.A1(new_n943), .A2(new_n543), .A3(new_n541), .A4(new_n945), .ZN(new_n946));
  AND3_X1   g760(.A1(new_n876), .A2(new_n944), .A3(new_n941), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n944), .B1(new_n876), .B2(new_n941), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n662), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n946), .A2(new_n949), .A3(new_n888), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT61), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n946), .A2(new_n949), .A3(KEYINPUT61), .A4(new_n888), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(G66));
  INV_X1    g768(.A(G224), .ZN(new_n955));
  OAI21_X1  g769(.A(G953), .B1(new_n509), .B2(new_n955), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n869), .A2(new_n840), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n956), .B1(new_n957), .B2(G953), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n958), .B(KEYINPUT121), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n959), .B(KEYINPUT122), .ZN(new_n960));
  OAI211_X1 g774(.A(new_n588), .B(new_n590), .C1(G898), .C2(new_n411), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n960), .B(new_n961), .Z(G69));
  NAND3_X1  g776(.A1(new_n783), .A2(new_n736), .A3(new_n798), .ZN(new_n963));
  AND4_X1   g777(.A1(new_n764), .A2(new_n790), .A3(new_n766), .A4(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT123), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n691), .A2(new_n716), .A3(new_n843), .ZN(new_n966));
  INV_X1    g780(.A(new_n966), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n965), .B1(new_n967), .B2(new_n785), .ZN(new_n968));
  AND4_X1   g782(.A1(new_n965), .A2(new_n785), .A3(new_n716), .A4(new_n853), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n964), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT124), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n970), .B(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n297), .A2(new_n298), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n973), .B(new_n448), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  OR3_X1    g789(.A1(new_n966), .A2(KEYINPUT62), .A3(new_n710), .ZN(new_n976));
  OAI21_X1  g790(.A(KEYINPUT62), .B1(new_n966), .B2(new_n710), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n697), .A2(new_n756), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n978), .A2(new_n332), .A3(new_n554), .A4(new_n838), .ZN(new_n979));
  AND3_X1   g793(.A1(new_n790), .A2(new_n785), .A3(new_n979), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n976), .A2(new_n977), .A3(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(new_n974), .ZN(new_n982));
  AOI21_X1  g796(.A(G953), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n982), .A2(new_n379), .ZN(new_n984));
  AOI211_X1 g798(.A(new_n669), .B(new_n411), .C1(new_n974), .C2(G227), .ZN(new_n985));
  AOI22_X1  g799(.A1(new_n975), .A2(new_n983), .B1(new_n984), .B2(new_n985), .ZN(G72));
  NAND2_X1  g800(.A1(G472), .A2(G902), .ZN(new_n987));
  XOR2_X1   g801(.A(new_n987), .B(KEYINPUT63), .Z(new_n988));
  AOI21_X1  g802(.A(new_n291), .B1(new_n299), .B2(new_n322), .ZN(new_n989));
  OAI211_X1 g803(.A(new_n856), .B(new_n988), .C1(new_n702), .C2(new_n989), .ZN(new_n990));
  INV_X1    g804(.A(new_n957), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n988), .B1(new_n981), .B2(new_n991), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n323), .B(KEYINPUT125), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n993), .A2(new_n292), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n992), .A2(new_n994), .ZN(new_n995));
  OAI211_X1 g809(.A(new_n990), .B(new_n995), .C1(G952), .C2(new_n411), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n993), .A2(new_n292), .ZN(new_n997));
  INV_X1    g811(.A(new_n988), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n998), .B1(new_n972), .B2(new_n957), .ZN(new_n999));
  INV_X1    g813(.A(KEYINPUT126), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n997), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  XNOR2_X1  g815(.A(new_n970), .B(KEYINPUT124), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n988), .B1(new_n1002), .B2(new_n991), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1003), .A2(KEYINPUT126), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n996), .B1(new_n1001), .B2(new_n1004), .ZN(G57));
endmodule


