

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755;

  NOR2_X1 U373 ( .A1(n582), .A2(n377), .ZN(n374) );
  OR2_X1 U374 ( .A1(n586), .A2(n579), .ZN(n618) );
  AND2_X1 U375 ( .A1(n611), .A2(G469), .ZN(n355) );
  XNOR2_X1 U376 ( .A(n393), .B(n733), .ZN(n455) );
  NAND2_X1 U377 ( .A1(n351), .A2(n535), .ZN(n540) );
  NAND2_X1 U378 ( .A1(n533), .A2(n532), .ZN(n351) );
  XNOR2_X2 U379 ( .A(n352), .B(n360), .ZN(n395) );
  NAND2_X1 U380 ( .A1(n397), .A2(n398), .ZN(n352) );
  NAND2_X2 U381 ( .A1(n399), .A2(n400), .ZN(n565) );
  XNOR2_X2 U382 ( .A(n429), .B(n428), .ZN(n431) );
  NOR2_X1 U383 ( .A1(G953), .A2(G237), .ZN(n476) );
  INV_X2 U384 ( .A(G953), .ZN(n446) );
  XNOR2_X2 U385 ( .A(G119), .B(G116), .ZN(n429) );
  NOR2_X2 U386 ( .A1(n560), .A2(n559), .ZN(n679) );
  XNOR2_X2 U387 ( .A(n445), .B(n444), .ZN(n735) );
  XNOR2_X2 U388 ( .A(n431), .B(n430), .ZN(n445) );
  XNOR2_X2 U389 ( .A(n745), .B(G146), .ZN(n437) );
  XNOR2_X2 U390 ( .A(n491), .B(n409), .ZN(n745) );
  NOR2_X1 U391 ( .A1(n622), .A2(n629), .ZN(n594) );
  OR2_X1 U392 ( .A1(n576), .A2(n575), .ZN(n586) );
  INV_X1 U393 ( .A(n542), .ZN(n550) );
  AND2_X1 U394 ( .A1(n615), .A2(n614), .ZN(n617) );
  OR2_X1 U395 ( .A1(n509), .A2(n508), .ZN(n511) );
  AND2_X1 U396 ( .A1(n565), .A2(n687), .ZN(n572) );
  XNOR2_X1 U397 ( .A(n424), .B(n423), .ZN(n542) );
  XNOR2_X1 U398 ( .A(n391), .B(n405), .ZN(n733) );
  XNOR2_X1 U399 ( .A(n451), .B(G134), .ZN(n491) );
  XNOR2_X1 U400 ( .A(n740), .B(n394), .ZN(n434) );
  XNOR2_X1 U401 ( .A(KEYINPUT66), .B(G101), .ZN(n394) );
  XNOR2_X1 U402 ( .A(KEYINPUT96), .B(KEYINPUT83), .ZN(n384) );
  XOR2_X1 U403 ( .A(n623), .B(KEYINPUT59), .Z(n624) );
  XNOR2_X2 U404 ( .A(n573), .B(n439), .ZN(n551) );
  XNOR2_X2 U405 ( .A(n353), .B(n354), .ZN(n500) );
  NOR2_X2 U406 ( .A1(n567), .A2(n467), .ZN(n353) );
  XOR2_X1 U407 ( .A(KEYINPUT87), .B(KEYINPUT0), .Z(n354) );
  XNOR2_X2 U408 ( .A(n554), .B(KEYINPUT19), .ZN(n567) );
  AND2_X2 U409 ( .A1(n649), .A2(G472), .ZN(n645) );
  XNOR2_X2 U410 ( .A(n388), .B(n387), .ZN(n640) );
  NOR2_X1 U411 ( .A1(n580), .A2(n703), .ZN(n378) );
  NAND2_X1 U412 ( .A1(n540), .A2(n539), .ZN(n541) );
  NAND2_X1 U413 ( .A1(n357), .A2(n378), .ZN(n371) );
  XNOR2_X1 U414 ( .A(n434), .B(KEYINPUT73), .ZN(n393) );
  NAND2_X1 U415 ( .A1(n586), .A2(n358), .ZN(n370) );
  INV_X1 U416 ( .A(n586), .ZN(n367) );
  INV_X1 U417 ( .A(G237), .ZN(n457) );
  NAND2_X1 U418 ( .A1(n402), .A2(n494), .ZN(n401) );
  XNOR2_X1 U419 ( .A(KEYINPUT69), .B(KEYINPUT8), .ZN(n412) );
  XOR2_X1 U420 ( .A(KEYINPUT103), .B(G122), .Z(n489) );
  XNOR2_X1 U421 ( .A(G116), .B(G107), .ZN(n488) );
  INV_X1 U422 ( .A(KEYINPUT65), .ZN(n403) );
  NAND2_X1 U423 ( .A1(n441), .A2(n440), .ZN(n443) );
  NAND2_X1 U424 ( .A1(n368), .A2(n365), .ZN(n601) );
  NAND2_X1 U425 ( .A1(n367), .A2(n366), .ZN(n365) );
  AND2_X1 U426 ( .A1(n370), .A2(n369), .ZN(n368) );
  NOR2_X1 U427 ( .A1(n702), .A2(n358), .ZN(n366) );
  INV_X1 U428 ( .A(KEYINPUT34), .ZN(n468) );
  BUF_X1 U429 ( .A(n517), .Z(n686) );
  AND2_X1 U430 ( .A1(n373), .A2(n375), .ZN(n372) );
  NAND2_X1 U431 ( .A1(n582), .A2(n377), .ZN(n375) );
  INV_X1 U432 ( .A(KEYINPUT67), .ZN(n385) );
  XNOR2_X1 U433 ( .A(G146), .B(G125), .ZN(n450) );
  NAND2_X1 U434 ( .A1(G234), .A2(G237), .ZN(n462) );
  NAND2_X1 U435 ( .A1(n702), .A2(n358), .ZN(n369) );
  XNOR2_X1 U436 ( .A(n565), .B(KEYINPUT1), .ZN(n517) );
  XNOR2_X1 U437 ( .A(n392), .B(KEYINPUT90), .ZN(n391) );
  XNOR2_X1 U438 ( .A(G110), .B(G107), .ZN(n392) );
  XNOR2_X1 U439 ( .A(n382), .B(n381), .ZN(n380) );
  XNOR2_X1 U440 ( .A(G119), .B(G137), .ZN(n382) );
  XNOR2_X1 U441 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(n381) );
  XNOR2_X1 U442 ( .A(G113), .B(G143), .ZN(n470) );
  XNOR2_X1 U443 ( .A(KEYINPUT12), .B(KEYINPUT11), .ZN(n472) );
  XNOR2_X1 U444 ( .A(n364), .B(n363), .ZN(n606) );
  INV_X1 U445 ( .A(KEYINPUT84), .ZN(n363) );
  XNOR2_X1 U446 ( .A(n591), .B(n590), .ZN(n718) );
  XNOR2_X1 U447 ( .A(KEYINPUT16), .B(G122), .ZN(n444) );
  XNOR2_X1 U448 ( .A(n493), .B(n492), .ZN(n657) );
  XNOR2_X1 U449 ( .A(n491), .B(n490), .ZN(n492) );
  NOR2_X1 U450 ( .A1(n446), .A2(G952), .ZN(n660) );
  INV_X1 U451 ( .A(G137), .ZN(n628) );
  NOR2_X1 U452 ( .A1(n556), .A2(n555), .ZN(n558) );
  INV_X1 U453 ( .A(KEYINPUT35), .ZN(n386) );
  INV_X1 U454 ( .A(KEYINPUT32), .ZN(n387) );
  NOR2_X1 U455 ( .A1(n530), .A2(n542), .ZN(n389) );
  XNOR2_X1 U456 ( .A(n390), .B(KEYINPUT107), .ZN(n641) );
  AND2_X1 U457 ( .A1(n604), .A2(KEYINPUT2), .ZN(n356) );
  AND2_X1 U458 ( .A1(n672), .A2(n377), .ZN(n357) );
  XNOR2_X1 U459 ( .A(KEYINPUT86), .B(KEYINPUT39), .ZN(n358) );
  INV_X1 U460 ( .A(KEYINPUT81), .ZN(n377) );
  AND2_X1 U461 ( .A1(G902), .A2(G469), .ZN(n359) );
  XNOR2_X1 U462 ( .A(KEYINPUT71), .B(KEYINPUT48), .ZN(n360) );
  XOR2_X1 U463 ( .A(n611), .B(n612), .Z(n361) );
  XNOR2_X1 U464 ( .A(KEYINPUT64), .B(KEYINPUT46), .ZN(n362) );
  INV_X1 U465 ( .A(G469), .ZN(n402) );
  NAND2_X1 U466 ( .A1(n395), .A2(n356), .ZN(n364) );
  NOR2_X1 U467 ( .A1(n623), .A2(G902), .ZN(n483) );
  XNOR2_X1 U468 ( .A(n481), .B(n743), .ZN(n623) );
  NOR2_X1 U469 ( .A1(n718), .A2(n592), .ZN(n593) );
  NOR2_X2 U470 ( .A1(n641), .A2(n640), .ZN(n537) );
  XNOR2_X2 U471 ( .A(G143), .B(G128), .ZN(n451) );
  NAND2_X1 U472 ( .A1(n601), .A2(n674), .ZN(n588) );
  NAND2_X1 U473 ( .A1(n395), .A2(n604), .ZN(n750) );
  NAND2_X1 U474 ( .A1(n372), .A2(n371), .ZN(n583) );
  NAND2_X1 U475 ( .A1(n374), .A2(n376), .ZN(n373) );
  NAND2_X1 U476 ( .A1(n378), .A2(n672), .ZN(n376) );
  XNOR2_X1 U477 ( .A(n404), .B(n379), .ZN(n416) );
  XNOR2_X1 U478 ( .A(n383), .B(n380), .ZN(n379) );
  XNOR2_X1 U479 ( .A(n411), .B(n384), .ZN(n383) );
  NOR2_X1 U480 ( .A1(n523), .A2(n385), .ZN(n521) );
  XNOR2_X2 U481 ( .A(n497), .B(n386), .ZN(n523) );
  AND2_X1 U482 ( .A1(n523), .A2(n385), .ZN(n536) );
  XNOR2_X1 U483 ( .A(n523), .B(G122), .ZN(n755) );
  NAND2_X1 U484 ( .A1(n500), .A2(n513), .ZN(n516) );
  NAND2_X1 U485 ( .A1(n528), .A2(n389), .ZN(n388) );
  NAND2_X1 U486 ( .A1(n528), .A2(n527), .ZN(n390) );
  XNOR2_X2 U487 ( .A(n516), .B(n515), .ZN(n528) );
  XNOR2_X2 U488 ( .A(KEYINPUT68), .B(KEYINPUT4), .ZN(n740) );
  AND2_X1 U489 ( .A1(n584), .A2(n583), .ZN(n397) );
  XNOR2_X1 U490 ( .A(n594), .B(n362), .ZN(n398) );
  NOR2_X1 U491 ( .A1(n355), .A2(n359), .ZN(n399) );
  OR2_X1 U492 ( .A1(n611), .A2(n401), .ZN(n400) );
  XNOR2_X1 U493 ( .A(n410), .B(n437), .ZN(n611) );
  NAND2_X1 U494 ( .A1(n649), .A2(G469), .ZN(n613) );
  AND2_X1 U495 ( .A1(n650), .A2(G478), .ZN(n659) );
  XNOR2_X2 U496 ( .A(n610), .B(n403), .ZN(n649) );
  AND2_X1 U497 ( .A1(G221), .A2(n485), .ZN(n404) );
  XNOR2_X1 U498 ( .A(G110), .B(G128), .ZN(n411) );
  INV_X1 U499 ( .A(n689), .ZN(n548) );
  AND2_X1 U500 ( .A1(n571), .A2(n548), .ZN(n549) );
  BUF_X1 U501 ( .A(n585), .Z(n577) );
  INV_X1 U502 ( .A(n660), .ZN(n614) );
  XNOR2_X1 U503 ( .A(G104), .B(KEYINPUT75), .ZN(n405) );
  XOR2_X1 U504 ( .A(G140), .B(KEYINPUT95), .Z(n407) );
  NAND2_X1 U505 ( .A1(G227), .A2(n446), .ZN(n406) );
  XNOR2_X1 U506 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U507 ( .A(n455), .B(n408), .ZN(n410) );
  XNOR2_X1 U508 ( .A(n628), .B(G131), .ZN(n409) );
  NAND2_X1 U509 ( .A1(n446), .A2(G234), .ZN(n413) );
  XNOR2_X1 U510 ( .A(n413), .B(n412), .ZN(n485) );
  XNOR2_X1 U511 ( .A(n450), .B(G140), .ZN(n415) );
  XOR2_X1 U512 ( .A(KEYINPUT70), .B(KEYINPUT10), .Z(n414) );
  XNOR2_X1 U513 ( .A(n415), .B(n414), .ZN(n743) );
  XNOR2_X1 U514 ( .A(n416), .B(n743), .ZN(n652) );
  INV_X1 U515 ( .A(G902), .ZN(n494) );
  NAND2_X1 U516 ( .A1(n652), .A2(n494), .ZN(n424) );
  XOR2_X1 U517 ( .A(KEYINPUT97), .B(KEYINPUT20), .Z(n420) );
  INV_X1 U518 ( .A(KEYINPUT15), .ZN(n417) );
  XNOR2_X1 U519 ( .A(n417), .B(G902), .ZN(n607) );
  INV_X1 U520 ( .A(n607), .ZN(n418) );
  NAND2_X1 U521 ( .A1(G234), .A2(n418), .ZN(n419) );
  XNOR2_X1 U522 ( .A(n420), .B(n419), .ZN(n425) );
  NAND2_X1 U523 ( .A1(G217), .A2(n425), .ZN(n422) );
  INV_X1 U524 ( .A(KEYINPUT25), .ZN(n421) );
  XNOR2_X1 U525 ( .A(n422), .B(n421), .ZN(n423) );
  NAND2_X1 U526 ( .A1(n425), .A2(G221), .ZN(n426) );
  XNOR2_X1 U527 ( .A(n426), .B(KEYINPUT21), .ZN(n689) );
  INV_X1 U528 ( .A(KEYINPUT98), .ZN(n427) );
  XNOR2_X1 U529 ( .A(n689), .B(n427), .ZN(n512) );
  AND2_X1 U530 ( .A1(n542), .A2(n512), .ZN(n687) );
  NAND2_X1 U531 ( .A1(n517), .A2(n687), .ZN(n498) );
  INV_X1 U532 ( .A(n498), .ZN(n441) );
  XNOR2_X2 U533 ( .A(G113), .B(KEYINPUT72), .ZN(n428) );
  XNOR2_X1 U534 ( .A(KEYINPUT91), .B(KEYINPUT3), .ZN(n430) );
  NAND2_X1 U535 ( .A1(n476), .A2(G210), .ZN(n432) );
  XNOR2_X1 U536 ( .A(n432), .B(KEYINPUT5), .ZN(n433) );
  XNOR2_X1 U537 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U538 ( .A(n445), .B(n435), .ZN(n436) );
  XNOR2_X1 U539 ( .A(n437), .B(n436), .ZN(n643) );
  OR2_X2 U540 ( .A1(n643), .A2(G902), .ZN(n438) );
  INV_X1 U541 ( .A(G472), .ZN(n642) );
  XNOR2_X2 U542 ( .A(n438), .B(n642), .ZN(n573) );
  XNOR2_X1 U543 ( .A(KEYINPUT105), .B(KEYINPUT6), .ZN(n439) );
  INV_X1 U544 ( .A(n551), .ZN(n440) );
  XNOR2_X1 U545 ( .A(KEYINPUT88), .B(KEYINPUT33), .ZN(n442) );
  XNOR2_X2 U546 ( .A(n443), .B(n442), .ZN(n719) );
  XOR2_X1 U547 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n449) );
  NAND2_X1 U548 ( .A1(G224), .A2(n446), .ZN(n447) );
  XNOR2_X1 U549 ( .A(n447), .B(KEYINPUT92), .ZN(n448) );
  XNOR2_X1 U550 ( .A(n449), .B(n448), .ZN(n453) );
  XNOR2_X1 U551 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U552 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U553 ( .A(n735), .B(n454), .ZN(n456) );
  XNOR2_X1 U554 ( .A(n456), .B(n455), .ZN(n630) );
  OR2_X2 U555 ( .A1(n630), .A2(n607), .ZN(n460) );
  NAND2_X1 U556 ( .A1(n494), .A2(n457), .ZN(n461) );
  NAND2_X1 U557 ( .A1(n461), .A2(G210), .ZN(n458) );
  XNOR2_X1 U558 ( .A(n458), .B(KEYINPUT93), .ZN(n459) );
  XNOR2_X2 U559 ( .A(n460), .B(n459), .ZN(n585) );
  NAND2_X1 U560 ( .A1(n461), .A2(G214), .ZN(n706) );
  AND2_X2 U561 ( .A1(n585), .A2(n706), .ZN(n554) );
  XNOR2_X1 U562 ( .A(n462), .B(KEYINPUT14), .ZN(n464) );
  NAND2_X1 U563 ( .A1(G952), .A2(n464), .ZN(n463) );
  XOR2_X1 U564 ( .A(KEYINPUT94), .B(n463), .Z(n716) );
  NAND2_X1 U565 ( .A1(n716), .A2(n446), .ZN(n546) );
  NAND2_X1 U566 ( .A1(G902), .A2(n464), .ZN(n543) );
  INV_X1 U567 ( .A(n543), .ZN(n465) );
  NOR2_X1 U568 ( .A1(G898), .A2(n446), .ZN(n736) );
  NAND2_X1 U569 ( .A1(n465), .A2(n736), .ZN(n466) );
  AND2_X1 U570 ( .A1(n546), .A2(n466), .ZN(n467) );
  NAND2_X1 U571 ( .A1(n719), .A2(n500), .ZN(n469) );
  XNOR2_X1 U572 ( .A(n469), .B(n468), .ZN(n496) );
  XOR2_X1 U573 ( .A(G104), .B(G122), .Z(n471) );
  XNOR2_X1 U574 ( .A(n471), .B(n470), .ZN(n475) );
  XOR2_X1 U575 ( .A(KEYINPUT101), .B(KEYINPUT100), .Z(n473) );
  XNOR2_X1 U576 ( .A(n473), .B(n472), .ZN(n474) );
  XNOR2_X1 U577 ( .A(n475), .B(n474), .ZN(n480) );
  XOR2_X1 U578 ( .A(KEYINPUT99), .B(G131), .Z(n478) );
  NAND2_X1 U579 ( .A1(G214), .A2(n476), .ZN(n477) );
  XNOR2_X1 U580 ( .A(n478), .B(n477), .ZN(n479) );
  XOR2_X1 U581 ( .A(n480), .B(n479), .Z(n481) );
  XNOR2_X1 U582 ( .A(KEYINPUT13), .B(KEYINPUT102), .ZN(n482) );
  XNOR2_X1 U583 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U584 ( .A(n484), .B(G475), .ZN(n509) );
  INV_X1 U585 ( .A(n509), .ZN(n503) );
  XOR2_X1 U586 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n487) );
  NAND2_X1 U587 ( .A1(G217), .A2(n485), .ZN(n486) );
  XNOR2_X1 U588 ( .A(n487), .B(n486), .ZN(n493) );
  XNOR2_X1 U589 ( .A(n489), .B(n488), .ZN(n490) );
  NAND2_X1 U590 ( .A1(n657), .A2(n494), .ZN(n495) );
  INV_X1 U591 ( .A(G478), .ZN(n656) );
  XNOR2_X1 U592 ( .A(n495), .B(n656), .ZN(n505) );
  NOR2_X1 U593 ( .A1(n503), .A2(n505), .ZN(n578) );
  NAND2_X1 U594 ( .A1(n496), .A2(n578), .ZN(n497) );
  NOR2_X1 U595 ( .A1(n498), .A2(n573), .ZN(n697) );
  NAND2_X1 U596 ( .A1(n500), .A2(n697), .ZN(n499) );
  XNOR2_X1 U597 ( .A(n499), .B(KEYINPUT31), .ZN(n677) );
  INV_X1 U598 ( .A(n500), .ZN(n502) );
  NAND2_X1 U599 ( .A1(n572), .A2(n573), .ZN(n501) );
  NOR2_X1 U600 ( .A1(n502), .A2(n501), .ZN(n665) );
  NOR2_X1 U601 ( .A1(n677), .A2(n665), .ZN(n507) );
  INV_X1 U602 ( .A(n505), .ZN(n508) );
  AND2_X1 U603 ( .A1(n503), .A2(n508), .ZN(n676) );
  INV_X1 U604 ( .A(KEYINPUT104), .ZN(n504) );
  XNOR2_X1 U605 ( .A(n676), .B(n504), .ZN(n602) );
  AND2_X1 U606 ( .A1(n505), .A2(n509), .ZN(n674) );
  INV_X1 U607 ( .A(n674), .ZN(n506) );
  AND2_X1 U608 ( .A1(n602), .A2(n506), .ZN(n703) );
  XNOR2_X1 U609 ( .A(n703), .B(KEYINPUT82), .ZN(n561) );
  OR2_X1 U610 ( .A1(n507), .A2(n561), .ZN(n520) );
  INV_X1 U611 ( .A(KEYINPUT106), .ZN(n510) );
  XNOR2_X2 U612 ( .A(n511), .B(n510), .ZN(n709) );
  AND2_X1 U613 ( .A1(n709), .A2(n512), .ZN(n513) );
  INV_X1 U614 ( .A(KEYINPUT74), .ZN(n514) );
  XNOR2_X1 U615 ( .A(n514), .B(KEYINPUT22), .ZN(n515) );
  NAND2_X1 U616 ( .A1(n551), .A2(n542), .ZN(n518) );
  NOR2_X1 U617 ( .A1(n686), .A2(n518), .ZN(n519) );
  NAND2_X1 U618 ( .A1(n528), .A2(n519), .ZN(n662) );
  NAND2_X1 U619 ( .A1(n520), .A2(n662), .ZN(n531) );
  NOR2_X1 U620 ( .A1(n521), .A2(n531), .ZN(n525) );
  NOR2_X1 U621 ( .A1(KEYINPUT67), .A2(KEYINPUT44), .ZN(n522) );
  NAND2_X1 U622 ( .A1(n523), .A2(n522), .ZN(n524) );
  NAND2_X1 U623 ( .A1(n525), .A2(n524), .ZN(n535) );
  INV_X1 U624 ( .A(n686), .ZN(n559) );
  AND2_X1 U625 ( .A1(n559), .A2(n573), .ZN(n526) );
  AND2_X1 U626 ( .A1(n550), .A2(n526), .ZN(n527) );
  XNOR2_X1 U627 ( .A(n551), .B(KEYINPUT76), .ZN(n529) );
  NAND2_X1 U628 ( .A1(n529), .A2(n686), .ZN(n530) );
  INV_X1 U629 ( .A(n537), .ZN(n533) );
  INV_X1 U630 ( .A(n531), .ZN(n532) );
  NAND2_X1 U631 ( .A1(n537), .A2(n536), .ZN(n538) );
  NAND2_X1 U632 ( .A1(n538), .A2(KEYINPUT44), .ZN(n539) );
  XNOR2_X2 U633 ( .A(n541), .B(KEYINPUT45), .ZN(n728) );
  NOR2_X1 U634 ( .A1(G900), .A2(n543), .ZN(n544) );
  NAND2_X1 U635 ( .A1(n544), .A2(G953), .ZN(n545) );
  NAND2_X1 U636 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U637 ( .A(n547), .B(KEYINPUT78), .ZN(n571) );
  NAND2_X1 U638 ( .A1(n550), .A2(n549), .ZN(n562) );
  NOR2_X1 U639 ( .A1(n551), .A2(n562), .ZN(n552) );
  XNOR2_X1 U640 ( .A(n552), .B(KEYINPUT108), .ZN(n553) );
  NAND2_X1 U641 ( .A1(n553), .A2(n674), .ZN(n595) );
  XNOR2_X1 U642 ( .A(n595), .B(KEYINPUT112), .ZN(n556) );
  INV_X1 U643 ( .A(n554), .ZN(n555) );
  INV_X1 U644 ( .A(KEYINPUT36), .ZN(n557) );
  XNOR2_X1 U645 ( .A(n558), .B(n557), .ZN(n560) );
  NOR2_X1 U646 ( .A1(n561), .A2(KEYINPUT47), .ZN(n569) );
  OR2_X1 U647 ( .A1(n573), .A2(n562), .ZN(n564) );
  INV_X1 U648 ( .A(KEYINPUT28), .ZN(n563) );
  XNOR2_X1 U649 ( .A(n564), .B(n563), .ZN(n566) );
  NAND2_X1 U650 ( .A1(n566), .A2(n565), .ZN(n592) );
  OR2_X1 U651 ( .A1(n592), .A2(n567), .ZN(n568) );
  XNOR2_X2 U652 ( .A(n568), .B(KEYINPUT77), .ZN(n672) );
  AND2_X1 U653 ( .A1(n569), .A2(n672), .ZN(n570) );
  NOR2_X1 U654 ( .A1(n679), .A2(n570), .ZN(n584) );
  NAND2_X1 U655 ( .A1(n572), .A2(n571), .ZN(n576) );
  INV_X1 U656 ( .A(n573), .ZN(n692) );
  NAND2_X1 U657 ( .A1(n692), .A2(n706), .ZN(n574) );
  XNOR2_X1 U658 ( .A(n574), .B(KEYINPUT30), .ZN(n575) );
  NAND2_X1 U659 ( .A1(n578), .A2(n577), .ZN(n579) );
  INV_X1 U660 ( .A(n618), .ZN(n580) );
  INV_X1 U661 ( .A(KEYINPUT47), .ZN(n581) );
  AND2_X1 U662 ( .A1(n618), .A2(n581), .ZN(n582) );
  INV_X1 U663 ( .A(n585), .ZN(n599) );
  XNOR2_X2 U664 ( .A(n599), .B(KEYINPUT38), .ZN(n708) );
  INV_X1 U665 ( .A(n708), .ZN(n702) );
  XOR2_X1 U666 ( .A(KEYINPUT110), .B(KEYINPUT40), .Z(n587) );
  XNOR2_X1 U667 ( .A(n588), .B(n587), .ZN(n622) );
  AND2_X1 U668 ( .A1(n706), .A2(n708), .ZN(n589) );
  NAND2_X1 U669 ( .A1(n709), .A2(n589), .ZN(n591) );
  XNOR2_X1 U670 ( .A(KEYINPUT111), .B(KEYINPUT41), .ZN(n590) );
  XNOR2_X1 U671 ( .A(n593), .B(KEYINPUT42), .ZN(n629) );
  XOR2_X1 U672 ( .A(KEYINPUT43), .B(KEYINPUT109), .Z(n598) );
  NOR2_X1 U673 ( .A1(n595), .A2(n686), .ZN(n596) );
  NAND2_X1 U674 ( .A1(n596), .A2(n706), .ZN(n597) );
  XNOR2_X1 U675 ( .A(n598), .B(n597), .ZN(n600) );
  AND2_X1 U676 ( .A1(n600), .A2(n599), .ZN(n620) );
  INV_X1 U677 ( .A(n601), .ZN(n603) );
  NOR2_X1 U678 ( .A1(n603), .A2(n602), .ZN(n619) );
  NOR2_X1 U679 ( .A1(n620), .A2(n619), .ZN(n604) );
  INV_X1 U680 ( .A(n750), .ZN(n605) );
  AND2_X2 U681 ( .A1(n728), .A2(n605), .ZN(n683) );
  NOR2_X1 U682 ( .A1(n683), .A2(KEYINPUT2), .ZN(n609) );
  NAND2_X1 U683 ( .A1(n606), .A2(n728), .ZN(n681) );
  NAND2_X1 U684 ( .A1(n681), .A2(n607), .ZN(n608) );
  NOR2_X2 U685 ( .A1(n609), .A2(n608), .ZN(n610) );
  XOR2_X1 U686 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n612) );
  XNOR2_X1 U687 ( .A(n613), .B(n361), .ZN(n615) );
  INV_X1 U688 ( .A(KEYINPUT119), .ZN(n616) );
  XNOR2_X1 U689 ( .A(n617), .B(n616), .ZN(G54) );
  XNOR2_X1 U690 ( .A(n618), .B(G143), .ZN(G45) );
  XOR2_X1 U691 ( .A(G134), .B(n619), .Z(G36) );
  XOR2_X1 U692 ( .A(G140), .B(KEYINPUT115), .Z(n621) );
  XOR2_X1 U693 ( .A(n621), .B(n620), .Z(G42) );
  XOR2_X1 U694 ( .A(G131), .B(n622), .Z(G33) );
  NAND2_X1 U695 ( .A1(n649), .A2(G475), .ZN(n625) );
  XNOR2_X1 U696 ( .A(n625), .B(n624), .ZN(n626) );
  NOR2_X2 U697 ( .A1(n626), .A2(n660), .ZN(n627) );
  XNOR2_X1 U698 ( .A(n627), .B(KEYINPUT60), .ZN(G60) );
  XNOR2_X1 U699 ( .A(n629), .B(n628), .ZN(G39) );
  NAND2_X1 U700 ( .A1(n649), .A2(G210), .ZN(n635) );
  BUF_X1 U701 ( .A(n630), .Z(n633) );
  XNOR2_X1 U702 ( .A(KEYINPUT79), .B(KEYINPUT54), .ZN(n631) );
  XNOR2_X1 U703 ( .A(n631), .B(KEYINPUT55), .ZN(n632) );
  XNOR2_X1 U704 ( .A(n633), .B(n632), .ZN(n634) );
  XNOR2_X1 U705 ( .A(n635), .B(n634), .ZN(n636) );
  NOR2_X2 U706 ( .A1(n636), .A2(n660), .ZN(n638) );
  XOR2_X1 U707 ( .A(KEYINPUT85), .B(KEYINPUT56), .Z(n637) );
  XNOR2_X1 U708 ( .A(n638), .B(n637), .ZN(G51) );
  XNOR2_X1 U709 ( .A(G119), .B(KEYINPUT127), .ZN(n639) );
  XNOR2_X1 U710 ( .A(n640), .B(n639), .ZN(G21) );
  XOR2_X1 U711 ( .A(G110), .B(n641), .Z(G12) );
  XOR2_X1 U712 ( .A(KEYINPUT62), .B(n643), .Z(n644) );
  XNOR2_X1 U713 ( .A(n645), .B(n644), .ZN(n646) );
  NOR2_X1 U714 ( .A1(n646), .A2(n660), .ZN(n648) );
  XNOR2_X1 U715 ( .A(KEYINPUT89), .B(KEYINPUT63), .ZN(n647) );
  XNOR2_X1 U716 ( .A(n648), .B(n647), .ZN(G57) );
  BUF_X1 U717 ( .A(n649), .Z(n650) );
  NAND2_X1 U718 ( .A1(n650), .A2(G217), .ZN(n654) );
  XNOR2_X1 U719 ( .A(KEYINPUT121), .B(KEYINPUT122), .ZN(n651) );
  XNOR2_X1 U720 ( .A(n652), .B(n651), .ZN(n653) );
  XNOR2_X1 U721 ( .A(n654), .B(n653), .ZN(n655) );
  NOR2_X1 U722 ( .A1(n655), .A2(n660), .ZN(G66) );
  XNOR2_X1 U723 ( .A(n657), .B(KEYINPUT120), .ZN(n658) );
  XNOR2_X1 U724 ( .A(n659), .B(n658), .ZN(n661) );
  NOR2_X1 U725 ( .A1(n661), .A2(n660), .ZN(G63) );
  XNOR2_X1 U726 ( .A(G101), .B(n662), .ZN(G3) );
  XOR2_X1 U727 ( .A(G104), .B(KEYINPUT113), .Z(n664) );
  NAND2_X1 U728 ( .A1(n665), .A2(n674), .ZN(n663) );
  XNOR2_X1 U729 ( .A(n664), .B(n663), .ZN(G6) );
  XOR2_X1 U730 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n667) );
  NAND2_X1 U731 ( .A1(n665), .A2(n676), .ZN(n666) );
  XNOR2_X1 U732 ( .A(n667), .B(n666), .ZN(n668) );
  XNOR2_X1 U733 ( .A(G107), .B(n668), .ZN(G9) );
  XOR2_X1 U734 ( .A(KEYINPUT29), .B(KEYINPUT114), .Z(n670) );
  NAND2_X1 U735 ( .A1(n672), .A2(n676), .ZN(n669) );
  XNOR2_X1 U736 ( .A(n670), .B(n669), .ZN(n671) );
  XNOR2_X1 U737 ( .A(G128), .B(n671), .ZN(G30) );
  NAND2_X1 U738 ( .A1(n672), .A2(n674), .ZN(n673) );
  XNOR2_X1 U739 ( .A(n673), .B(G146), .ZN(G48) );
  NAND2_X1 U740 ( .A1(n677), .A2(n674), .ZN(n675) );
  XNOR2_X1 U741 ( .A(n675), .B(G113), .ZN(G15) );
  NAND2_X1 U742 ( .A1(n677), .A2(n676), .ZN(n678) );
  XNOR2_X1 U743 ( .A(n678), .B(G116), .ZN(G18) );
  XNOR2_X1 U744 ( .A(n679), .B(G125), .ZN(n680) );
  XNOR2_X1 U745 ( .A(n680), .B(KEYINPUT37), .ZN(G27) );
  INV_X1 U746 ( .A(n681), .ZN(n685) );
  XNOR2_X1 U747 ( .A(KEYINPUT80), .B(KEYINPUT2), .ZN(n682) );
  NOR2_X1 U748 ( .A1(n683), .A2(n682), .ZN(n684) );
  NOR2_X1 U749 ( .A1(n685), .A2(n684), .ZN(n724) );
  NOR2_X1 U750 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U751 ( .A(KEYINPUT50), .B(n688), .ZN(n696) );
  NAND2_X1 U752 ( .A1(n689), .A2(n550), .ZN(n690) );
  XNOR2_X1 U753 ( .A(n690), .B(KEYINPUT49), .ZN(n691) );
  XNOR2_X1 U754 ( .A(n691), .B(KEYINPUT116), .ZN(n693) );
  NOR2_X1 U755 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U756 ( .A(n694), .B(KEYINPUT117), .ZN(n695) );
  OR2_X1 U757 ( .A1(n696), .A2(n695), .ZN(n699) );
  INV_X1 U758 ( .A(n697), .ZN(n698) );
  NAND2_X1 U759 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U760 ( .A(n700), .B(KEYINPUT51), .ZN(n701) );
  NOR2_X1 U761 ( .A1(n701), .A2(n718), .ZN(n714) );
  OR2_X1 U762 ( .A1(n703), .A2(n702), .ZN(n705) );
  INV_X1 U763 ( .A(n709), .ZN(n704) );
  NAND2_X1 U764 ( .A1(n705), .A2(n704), .ZN(n707) );
  NAND2_X1 U765 ( .A1(n707), .A2(n706), .ZN(n711) );
  NAND2_X1 U766 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U767 ( .A1(n711), .A2(n710), .ZN(n712) );
  AND2_X1 U768 ( .A1(n712), .A2(n719), .ZN(n713) );
  NOR2_X1 U769 ( .A1(n714), .A2(n713), .ZN(n715) );
  XOR2_X1 U770 ( .A(KEYINPUT52), .B(n715), .Z(n717) );
  NAND2_X1 U771 ( .A1(n717), .A2(n716), .ZN(n722) );
  INV_X1 U772 ( .A(n718), .ZN(n720) );
  NAND2_X1 U773 ( .A1(n720), .A2(n719), .ZN(n721) );
  NAND2_X1 U774 ( .A1(n722), .A2(n721), .ZN(n723) );
  NOR2_X1 U775 ( .A1(n724), .A2(n723), .ZN(n725) );
  XOR2_X1 U776 ( .A(KEYINPUT118), .B(n725), .Z(n726) );
  NOR2_X1 U777 ( .A1(G953), .A2(n726), .ZN(n727) );
  XNOR2_X1 U778 ( .A(KEYINPUT53), .B(n727), .ZN(G75) );
  NAND2_X1 U779 ( .A1(n728), .A2(n446), .ZN(n732) );
  NAND2_X1 U780 ( .A1(G953), .A2(G224), .ZN(n729) );
  XNOR2_X1 U781 ( .A(KEYINPUT61), .B(n729), .ZN(n730) );
  NAND2_X1 U782 ( .A1(n730), .A2(G898), .ZN(n731) );
  NAND2_X1 U783 ( .A1(n732), .A2(n731), .ZN(n739) );
  XNOR2_X1 U784 ( .A(n733), .B(G101), .ZN(n734) );
  XNOR2_X1 U785 ( .A(n735), .B(n734), .ZN(n737) );
  NOR2_X1 U786 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U787 ( .A(n739), .B(n738), .ZN(G69) );
  XNOR2_X1 U788 ( .A(KEYINPUT95), .B(KEYINPUT123), .ZN(n741) );
  XNOR2_X1 U789 ( .A(n740), .B(n741), .ZN(n742) );
  XNOR2_X1 U790 ( .A(n743), .B(n742), .ZN(n744) );
  XNOR2_X1 U791 ( .A(n745), .B(n744), .ZN(n748) );
  XNOR2_X1 U792 ( .A(n748), .B(G227), .ZN(n746) );
  NOR2_X1 U793 ( .A1(n446), .A2(n746), .ZN(n747) );
  NAND2_X1 U794 ( .A1(n747), .A2(G900), .ZN(n753) );
  XNOR2_X1 U795 ( .A(n748), .B(KEYINPUT124), .ZN(n749) );
  XNOR2_X1 U796 ( .A(n750), .B(n749), .ZN(n751) );
  NAND2_X1 U797 ( .A1(n751), .A2(n446), .ZN(n752) );
  NAND2_X1 U798 ( .A1(n753), .A2(n752), .ZN(n754) );
  XNOR2_X1 U799 ( .A(KEYINPUT125), .B(n754), .ZN(G72) );
  XNOR2_X1 U800 ( .A(KEYINPUT126), .B(n755), .ZN(G24) );
endmodule

