

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762;

  XNOR2_X2 U366 ( .A(n615), .B(n614), .ZN(n668) );
  NAND2_X2 U367 ( .A1(n449), .A2(n448), .ZN(n447) );
  NAND2_X2 U368 ( .A1(n367), .A2(n369), .ZN(n366) );
  INV_X1 U369 ( .A(n587), .ZN(n595) );
  XNOR2_X1 U370 ( .A(n411), .B(n734), .ZN(n408) );
  INV_X4 U371 ( .A(KEYINPUT4), .ZN(n409) );
  AND2_X1 U372 ( .A1(n405), .A2(n404), .ZN(n414) );
  XNOR2_X1 U373 ( .A(n586), .B(KEYINPUT32), .ZN(n755) );
  AND2_X1 U374 ( .A1(n592), .A2(n596), .ZN(n618) );
  XNOR2_X1 U375 ( .A(n584), .B(n583), .ZN(n592) );
  XNOR2_X1 U376 ( .A(n549), .B(n461), .ZN(n587) );
  XNOR2_X1 U377 ( .A(n520), .B(n519), .ZN(n540) );
  XNOR2_X1 U378 ( .A(n554), .B(n553), .ZN(n578) );
  OR2_X1 U379 ( .A1(n717), .A2(G902), .ZN(n365) );
  NOR2_X1 U380 ( .A1(n647), .A2(G902), .ZN(n520) );
  XNOR2_X1 U381 ( .A(n576), .B(KEYINPUT85), .ZN(n577) );
  XNOR2_X1 U382 ( .A(n742), .B(G146), .ZN(n516) );
  XNOR2_X1 U383 ( .A(n422), .B(G143), .ZN(n525) );
  NAND2_X1 U384 ( .A1(n595), .A2(n686), .ZN(n431) );
  XNOR2_X2 U385 ( .A(n378), .B(n353), .ZN(n413) );
  XNOR2_X1 U386 ( .A(n613), .B(n601), .ZN(n609) );
  AND2_X2 U387 ( .A1(n377), .A2(n368), .ZN(n354) );
  XNOR2_X2 U388 ( .A(n626), .B(KEYINPUT45), .ZN(n377) );
  XNOR2_X2 U389 ( .A(n409), .B(G101), .ZN(n509) );
  AND2_X1 U390 ( .A1(n444), .A2(n442), .ZN(n437) );
  NAND2_X1 U391 ( .A1(n440), .A2(KEYINPUT76), .ZN(n439) );
  NOR2_X1 U392 ( .A1(n447), .A2(n443), .ZN(n434) );
  NAND2_X1 U393 ( .A1(n755), .A2(n757), .ZN(n594) );
  NOR2_X1 U394 ( .A1(n588), .A2(n689), .ZN(n686) );
  NAND2_X1 U395 ( .A1(n373), .A2(n387), .ZN(n368) );
  BUF_X1 U396 ( .A(n540), .Z(n692) );
  NAND2_X1 U397 ( .A1(n549), .A2(n686), .ZN(n608) );
  INV_X1 U398 ( .A(KEYINPUT86), .ZN(n601) );
  XNOR2_X1 U399 ( .A(G146), .B(G125), .ZN(n524) );
  XOR2_X1 U400 ( .A(KEYINPUT90), .B(KEYINPUT5), .Z(n514) );
  XNOR2_X1 U401 ( .A(n393), .B(KEYINPUT46), .ZN(n392) );
  NAND2_X1 U402 ( .A1(n359), .A2(n394), .ZN(n393) );
  INV_X1 U403 ( .A(n762), .ZN(n394) );
  NOR2_X1 U404 ( .A1(n672), .A2(n349), .ZN(n423) );
  XNOR2_X1 U405 ( .A(n386), .B(G119), .ZN(n522) );
  XNOR2_X1 U406 ( .A(G113), .B(KEYINPUT3), .ZN(n386) );
  NAND2_X1 U407 ( .A1(n594), .A2(KEYINPUT44), .ZN(n404) );
  INV_X1 U408 ( .A(n594), .ZN(n622) );
  XNOR2_X1 U409 ( .A(n524), .B(n362), .ZN(n496) );
  XNOR2_X1 U410 ( .A(G140), .B(KEYINPUT10), .ZN(n362) );
  XNOR2_X1 U411 ( .A(n361), .B(KEYINPUT65), .ZN(n473) );
  INV_X1 U412 ( .A(G137), .ZN(n361) );
  INV_X1 U413 ( .A(n580), .ZN(n678) );
  XNOR2_X1 U414 ( .A(n546), .B(KEYINPUT38), .ZN(n676) );
  XNOR2_X1 U415 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X1 U416 ( .A(n410), .B(n457), .ZN(n734) );
  INV_X1 U417 ( .A(G104), .ZN(n457) );
  XNOR2_X1 U418 ( .A(KEYINPUT80), .B(G110), .ZN(n410) );
  XNOR2_X1 U419 ( .A(n397), .B(n523), .ZN(n736) );
  XNOR2_X1 U420 ( .A(n522), .B(KEYINPUT16), .ZN(n397) );
  XNOR2_X1 U421 ( .A(n474), .B(KEYINPUT88), .ZN(n376) );
  XNOR2_X1 U422 ( .A(G119), .B(G128), .ZN(n474) );
  XNOR2_X1 U423 ( .A(KEYINPUT23), .B(G110), .ZN(n375) );
  XNOR2_X1 U424 ( .A(n496), .B(n473), .ZN(n741) );
  XNOR2_X1 U425 ( .A(n509), .B(KEYINPUT66), .ZN(n411) );
  NAND2_X1 U426 ( .A1(n372), .A2(KEYINPUT2), .ZN(n371) );
  OR2_X1 U427 ( .A1(n665), .A2(n596), .ZN(n521) );
  NAND2_X1 U428 ( .A1(n413), .A2(n675), .ZN(n554) );
  OR2_X1 U429 ( .A1(n725), .A2(G902), .ZN(n364) );
  INV_X1 U430 ( .A(KEYINPUT25), .ZN(n481) );
  XNOR2_X1 U431 ( .A(G478), .B(n348), .ZN(n560) );
  INV_X1 U432 ( .A(KEYINPUT89), .ZN(n382) );
  NAND2_X1 U433 ( .A1(n608), .A2(n382), .ZN(n381) );
  OR2_X1 U434 ( .A1(n609), .A2(n384), .ZN(n383) );
  NAND2_X1 U435 ( .A1(n385), .A2(KEYINPUT89), .ZN(n384) );
  NAND2_X1 U436 ( .A1(n714), .A2(G475), .ZN(n403) );
  AND2_X1 U437 ( .A1(n443), .A2(KEYINPUT44), .ZN(n442) );
  INV_X1 U438 ( .A(KEYINPUT44), .ZN(n440) );
  INV_X1 U439 ( .A(KEYINPUT76), .ZN(n443) );
  NOR2_X1 U440 ( .A1(G953), .A2(G237), .ZN(n512) );
  XNOR2_X1 U441 ( .A(KEYINPUT64), .B(G131), .ZN(n499) );
  INV_X1 U442 ( .A(n627), .ZN(n373) );
  XNOR2_X1 U443 ( .A(KEYINPUT15), .B(G902), .ZN(n627) );
  INV_X1 U444 ( .A(G128), .ZN(n422) );
  XNOR2_X1 U445 ( .A(G104), .B(G122), .ZN(n500) );
  XNOR2_X1 U446 ( .A(G113), .B(G143), .ZN(n501) );
  XNOR2_X1 U447 ( .A(KEYINPUT93), .B(KEYINPUT12), .ZN(n493) );
  XOR2_X1 U448 ( .A(KEYINPUT94), .B(KEYINPUT11), .Z(n494) );
  NAND2_X1 U449 ( .A1(n373), .A2(KEYINPUT73), .ZN(n372) );
  NAND2_X1 U450 ( .A1(n627), .A2(n370), .ZN(n369) );
  INV_X1 U451 ( .A(KEYINPUT73), .ZN(n370) );
  NAND2_X1 U452 ( .A1(G234), .A2(G237), .ZN(n462) );
  NAND2_X1 U453 ( .A1(n676), .A2(n675), .ZN(n679) );
  INV_X1 U454 ( .A(n679), .ZN(n430) );
  AND2_X1 U455 ( .A1(n558), .A2(n547), .ZN(n580) );
  XNOR2_X1 U456 ( .A(n598), .B(n597), .ZN(n599) );
  INV_X1 U457 ( .A(KEYINPUT103), .ZN(n597) );
  INV_X1 U458 ( .A(G237), .ZN(n531) );
  NAND2_X1 U459 ( .A1(n446), .A2(n607), .ZN(n445) );
  INV_X1 U460 ( .A(n605), .ZN(n446) );
  INV_X1 U461 ( .A(KEYINPUT30), .ZN(n421) );
  XNOR2_X1 U462 ( .A(n516), .B(n419), .ZN(n647) );
  XNOR2_X1 U463 ( .A(n420), .B(n510), .ZN(n419) );
  XNOR2_X1 U464 ( .A(n511), .B(n515), .ZN(n420) );
  NOR2_X1 U465 ( .A1(n395), .A2(n392), .ZN(n564) );
  XNOR2_X1 U466 ( .A(n525), .B(n452), .ZN(n492) );
  INV_X1 U467 ( .A(G134), .ZN(n452) );
  XNOR2_X1 U468 ( .A(n487), .B(n486), .ZN(n523) );
  INV_X1 U469 ( .A(G122), .ZN(n486) );
  XNOR2_X1 U470 ( .A(n429), .B(n427), .ZN(n707) );
  XNOR2_X1 U471 ( .A(n428), .B(KEYINPUT41), .ZN(n427) );
  NAND2_X1 U472 ( .A1(n430), .A2(n580), .ZN(n429) );
  INV_X1 U473 ( .A(KEYINPUT106), .ZN(n428) );
  INV_X1 U474 ( .A(KEYINPUT39), .ZN(n551) );
  NAND2_X1 U475 ( .A1(n605), .A2(KEYINPUT35), .ZN(n448) );
  XNOR2_X1 U476 ( .A(n545), .B(KEYINPUT105), .ZN(n556) );
  NOR2_X1 U477 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U478 ( .A(n540), .B(n539), .ZN(n590) );
  XNOR2_X1 U479 ( .A(n376), .B(n375), .ZN(n477) );
  XNOR2_X1 U480 ( .A(n426), .B(n424), .ZN(n721) );
  XNOR2_X1 U481 ( .A(n523), .B(n425), .ZN(n424) );
  XNOR2_X1 U482 ( .A(n491), .B(n492), .ZN(n426) );
  XNOR2_X1 U483 ( .A(n489), .B(n488), .ZN(n425) );
  XNOR2_X1 U484 ( .A(n460), .B(n516), .ZN(n717) );
  XNOR2_X1 U485 ( .A(n537), .B(n416), .ZN(n538) );
  INV_X1 U486 ( .A(KEYINPUT36), .ZN(n416) );
  OR2_X1 U487 ( .A1(n560), .A2(n558), .ZN(n508) );
  AND2_X1 U488 ( .A1(n383), .A2(n356), .ZN(n380) );
  NAND2_X1 U489 ( .A1(n620), .A2(n619), .ZN(n641) );
  XNOR2_X1 U490 ( .A(n358), .B(KEYINPUT125), .ZN(G72) );
  INV_X1 U491 ( .A(KEYINPUT60), .ZN(n400) );
  AND2_X1 U492 ( .A1(n374), .A2(n371), .ZN(n347) );
  OR2_X1 U493 ( .A1(G902), .A2(n721), .ZN(n348) );
  XOR2_X1 U494 ( .A(n557), .B(KEYINPUT47), .Z(n349) );
  XOR2_X1 U495 ( .A(n458), .B(KEYINPUT87), .Z(n350) );
  XOR2_X1 U496 ( .A(n473), .B(G140), .Z(n351) );
  AND2_X1 U497 ( .A1(n732), .A2(n731), .ZN(n352) );
  XOR2_X1 U498 ( .A(n534), .B(n533), .Z(n353) );
  XOR2_X1 U499 ( .A(n482), .B(n481), .Z(n355) );
  AND2_X1 U500 ( .A1(n381), .A2(n610), .ZN(n356) );
  XOR2_X1 U501 ( .A(n646), .B(n645), .Z(n357) );
  INV_X1 U502 ( .A(KEYINPUT2), .ZN(n387) );
  INV_X1 U503 ( .A(G953), .ZN(n526) );
  AND2_X1 U504 ( .A1(n751), .A2(n752), .ZN(n358) );
  INV_X1 U505 ( .A(n759), .ZN(n359) );
  XNOR2_X1 U506 ( .A(n552), .B(KEYINPUT40), .ZN(n759) );
  NAND2_X1 U507 ( .A1(n456), .A2(n455), .ZN(n742) );
  XNOR2_X1 U508 ( .A(n388), .B(KEYINPUT69), .ZN(n562) );
  NAND2_X1 U509 ( .A1(n360), .A2(n414), .ZN(n621) );
  NAND2_X1 U510 ( .A1(n436), .A2(n433), .ZN(n360) );
  XNOR2_X1 U511 ( .A(n417), .B(n459), .ZN(n460) );
  NOR2_X1 U512 ( .A1(n565), .A2(n665), .ZN(n552) );
  XNOR2_X1 U513 ( .A(n363), .B(n551), .ZN(n565) );
  NAND2_X1 U514 ( .A1(n562), .A2(n676), .ZN(n363) );
  XNOR2_X2 U515 ( .A(n364), .B(n355), .ZN(n588) );
  XNOR2_X2 U516 ( .A(n365), .B(G469), .ZN(n549) );
  NOR2_X4 U517 ( .A1(n347), .A2(n366), .ZN(n714) );
  NAND2_X1 U518 ( .A1(n354), .A2(n412), .ZN(n367) );
  NAND2_X1 U519 ( .A1(n412), .A2(n377), .ZN(n374) );
  XNOR2_X1 U520 ( .A(n374), .B(n387), .ZN(n711) );
  NAND2_X1 U521 ( .A1(n377), .A2(n526), .ZN(n732) );
  INV_X1 U522 ( .A(n413), .ZN(n546) );
  NAND2_X1 U523 ( .A1(n630), .A2(n627), .ZN(n378) );
  XNOR2_X1 U524 ( .A(n398), .B(n736), .ZN(n630) );
  NAND2_X2 U525 ( .A1(n380), .A2(n379), .ZN(n657) );
  NAND2_X1 U526 ( .A1(n609), .A2(n382), .ZN(n379) );
  INV_X1 U527 ( .A(n608), .ZN(n385) );
  NAND2_X1 U528 ( .A1(n390), .A2(n389), .ZN(n388) );
  NOR2_X1 U529 ( .A1(n608), .A2(n550), .ZN(n389) );
  XNOR2_X1 U530 ( .A(n391), .B(n421), .ZN(n390) );
  NAND2_X1 U531 ( .A1(n590), .A2(n675), .ZN(n391) );
  NAND2_X1 U532 ( .A1(n423), .A2(n396), .ZN(n395) );
  INV_X1 U533 ( .A(n644), .ZN(n396) );
  XNOR2_X1 U534 ( .A(n408), .B(n399), .ZN(n398) );
  XNOR2_X1 U535 ( .A(n530), .B(n529), .ZN(n399) );
  XNOR2_X1 U536 ( .A(n401), .B(n400), .ZN(G60) );
  NAND2_X1 U537 ( .A1(n402), .A2(n651), .ZN(n401) );
  XNOR2_X1 U538 ( .A(n403), .B(n357), .ZN(n402) );
  XNOR2_X1 U539 ( .A(n406), .B(KEYINPUT99), .ZN(n405) );
  NAND2_X1 U540 ( .A1(n407), .A2(n641), .ZN(n406) );
  NAND2_X1 U541 ( .A1(n617), .A2(n616), .ZN(n407) );
  XNOR2_X1 U542 ( .A(n408), .B(n350), .ZN(n417) );
  INV_X1 U543 ( .A(n747), .ZN(n412) );
  NAND2_X1 U544 ( .A1(n415), .A2(n570), .ZN(n747) );
  XNOR2_X1 U545 ( .A(n564), .B(KEYINPUT48), .ZN(n415) );
  NAND2_X1 U546 ( .A1(n447), .A2(n442), .ZN(n441) );
  NAND2_X1 U547 ( .A1(n441), .A2(n439), .ZN(n438) );
  XNOR2_X2 U548 ( .A(n418), .B(KEYINPUT0), .ZN(n613) );
  NOR2_X2 U549 ( .A1(n578), .A2(n577), .ZN(n418) );
  XOR2_X1 U550 ( .A(KEYINPUT42), .B(n548), .Z(n762) );
  INV_X1 U551 ( .A(n431), .ZN(n611) );
  NOR2_X1 U552 ( .A1(n431), .A2(n596), .ZN(n600) );
  NAND2_X1 U553 ( .A1(n435), .A2(n432), .ZN(n753) );
  INV_X1 U554 ( .A(n447), .ZN(n432) );
  NAND2_X1 U555 ( .A1(n435), .A2(n434), .ZN(n433) );
  INV_X1 U556 ( .A(n444), .ZN(n435) );
  NOR2_X1 U557 ( .A1(n438), .A2(n437), .ZN(n436) );
  NOR2_X1 U558 ( .A1(n606), .A2(n445), .ZN(n444) );
  NAND2_X1 U559 ( .A1(n606), .A2(KEYINPUT35), .ZN(n449) );
  XNOR2_X1 U560 ( .A(n719), .B(n718), .ZN(n720) );
  BUF_X1 U561 ( .A(n595), .Z(n685) );
  XOR2_X1 U562 ( .A(n716), .B(n715), .Z(n450) );
  XOR2_X1 U563 ( .A(n569), .B(KEYINPUT43), .Z(n451) );
  INV_X1 U564 ( .A(KEYINPUT91), .ZN(n517) );
  INV_X1 U565 ( .A(KEYINPUT101), .ZN(n539) );
  XNOR2_X1 U566 ( .A(n477), .B(n476), .ZN(n478) );
  BUF_X1 U567 ( .A(n630), .Z(n631) );
  XNOR2_X1 U568 ( .A(n648), .B(KEYINPUT62), .ZN(n649) );
  XNOR2_X1 U569 ( .A(n479), .B(n478), .ZN(n725) );
  INV_X1 U570 ( .A(KEYINPUT35), .ZN(n607) );
  XNOR2_X1 U571 ( .A(n717), .B(n450), .ZN(n718) );
  INV_X1 U572 ( .A(n492), .ZN(n454) );
  INV_X1 U573 ( .A(n499), .ZN(n453) );
  NAND2_X1 U574 ( .A1(n454), .A2(n499), .ZN(n456) );
  NAND2_X1 U575 ( .A1(n453), .A2(n492), .ZN(n455) );
  AND2_X1 U576 ( .A1(G227), .A2(n526), .ZN(n458) );
  XNOR2_X1 U577 ( .A(n351), .B(G107), .ZN(n459) );
  INV_X1 U578 ( .A(KEYINPUT1), .ZN(n461) );
  XNOR2_X1 U579 ( .A(n462), .B(KEYINPUT82), .ZN(n463) );
  XNOR2_X1 U580 ( .A(KEYINPUT14), .B(n463), .ZN(n465) );
  NAND2_X1 U581 ( .A1(G952), .A2(n465), .ZN(n705) );
  NOR2_X1 U582 ( .A1(G953), .A2(n705), .ZN(n464) );
  XNOR2_X1 U583 ( .A(KEYINPUT83), .B(n464), .ZN(n575) );
  INV_X1 U584 ( .A(n575), .ZN(n468) );
  AND2_X1 U585 ( .A1(n465), .A2(G953), .ZN(n466) );
  NAND2_X1 U586 ( .A1(G902), .A2(n466), .ZN(n572) );
  NOR2_X1 U587 ( .A1(G900), .A2(n572), .ZN(n467) );
  NOR2_X1 U588 ( .A1(n468), .A2(n467), .ZN(n469) );
  XNOR2_X1 U589 ( .A(KEYINPUT72), .B(n469), .ZN(n550) );
  INV_X1 U590 ( .A(n550), .ZN(n485) );
  NAND2_X1 U591 ( .A1(G234), .A2(n627), .ZN(n470) );
  XNOR2_X1 U592 ( .A(KEYINPUT20), .B(n470), .ZN(n480) );
  AND2_X1 U593 ( .A1(n480), .A2(G221), .ZN(n472) );
  INV_X1 U594 ( .A(KEYINPUT21), .ZN(n471) );
  XNOR2_X1 U595 ( .A(n472), .B(n471), .ZN(n689) );
  XNOR2_X1 U596 ( .A(n741), .B(KEYINPUT24), .ZN(n479) );
  NAND2_X1 U597 ( .A1(G234), .A2(n526), .ZN(n475) );
  XOR2_X1 U598 ( .A(KEYINPUT8), .B(n475), .Z(n490) );
  NAND2_X1 U599 ( .A1(n490), .A2(G221), .ZN(n476) );
  NAND2_X1 U600 ( .A1(n480), .A2(G217), .ZN(n482) );
  INV_X1 U601 ( .A(n588), .ZN(n483) );
  NOR2_X1 U602 ( .A1(n689), .A2(n483), .ZN(n484) );
  NAND2_X1 U603 ( .A1(n485), .A2(n484), .ZN(n541) );
  XOR2_X1 U604 ( .A(G116), .B(G107), .Z(n487) );
  XOR2_X1 U605 ( .A(KEYINPUT95), .B(KEYINPUT96), .Z(n489) );
  XNOR2_X1 U606 ( .A(KEYINPUT9), .B(KEYINPUT7), .ZN(n488) );
  NAND2_X1 U607 ( .A1(G217), .A2(n490), .ZN(n491) );
  XNOR2_X1 U608 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U609 ( .A(n496), .B(n495), .ZN(n498) );
  NAND2_X1 U610 ( .A1(G214), .A2(n512), .ZN(n497) );
  XNOR2_X1 U611 ( .A(n498), .B(n497), .ZN(n505) );
  XNOR2_X1 U612 ( .A(KEYINPUT92), .B(n499), .ZN(n503) );
  INV_X1 U613 ( .A(G143), .ZN(n643) );
  XNOR2_X1 U614 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U615 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U616 ( .A(n505), .B(n504), .ZN(n646) );
  INV_X1 U617 ( .A(G902), .ZN(n532) );
  NAND2_X1 U618 ( .A1(n646), .A2(n532), .ZN(n507) );
  XNOR2_X1 U619 ( .A(KEYINPUT13), .B(G475), .ZN(n506) );
  XNOR2_X1 U620 ( .A(n507), .B(n506), .ZN(n558) );
  XOR2_X1 U621 ( .A(n508), .B(KEYINPUT97), .Z(n665) );
  XOR2_X1 U622 ( .A(n509), .B(G116), .Z(n511) );
  XNOR2_X1 U623 ( .A(n522), .B(G137), .ZN(n510) );
  NAND2_X1 U624 ( .A1(n512), .A2(G210), .ZN(n513) );
  XNOR2_X1 U625 ( .A(n514), .B(n513), .ZN(n515) );
  INV_X1 U626 ( .A(G472), .ZN(n518) );
  XNOR2_X1 U627 ( .A(n692), .B(KEYINPUT6), .ZN(n596) );
  NOR2_X1 U628 ( .A1(n541), .A2(n521), .ZN(n567) );
  XNOR2_X1 U629 ( .A(KEYINPUT107), .B(n567), .ZN(n536) );
  XNOR2_X1 U630 ( .A(n525), .B(n524), .ZN(n530) );
  XNOR2_X1 U631 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n528) );
  NAND2_X1 U632 ( .A1(n526), .A2(G224), .ZN(n527) );
  XNOR2_X1 U633 ( .A(n528), .B(n527), .ZN(n529) );
  NAND2_X1 U634 ( .A1(n532), .A2(n531), .ZN(n535) );
  NAND2_X1 U635 ( .A1(n535), .A2(G210), .ZN(n534) );
  XNOR2_X1 U636 ( .A(KEYINPUT71), .B(KEYINPUT81), .ZN(n533) );
  NAND2_X1 U637 ( .A1(n535), .A2(G214), .ZN(n675) );
  NOR2_X1 U638 ( .A1(n536), .A2(n554), .ZN(n537) );
  NOR2_X1 U639 ( .A1(n587), .A2(n538), .ZN(n672) );
  INV_X1 U640 ( .A(n590), .ZN(n542) );
  XNOR2_X1 U641 ( .A(KEYINPUT28), .B(n543), .ZN(n544) );
  NAND2_X1 U642 ( .A1(n544), .A2(n549), .ZN(n545) );
  INV_X1 U643 ( .A(n560), .ZN(n547) );
  INV_X1 U644 ( .A(n707), .ZN(n699) );
  NAND2_X1 U645 ( .A1(n556), .A2(n699), .ZN(n548) );
  INV_X1 U646 ( .A(KEYINPUT19), .ZN(n553) );
  INV_X1 U647 ( .A(n578), .ZN(n555) );
  NAND2_X1 U648 ( .A1(n556), .A2(n555), .ZN(n663) );
  NAND2_X1 U649 ( .A1(n558), .A2(n560), .ZN(n669) );
  AND2_X1 U650 ( .A1(n665), .A2(n669), .ZN(n680) );
  NOR2_X1 U651 ( .A1(n663), .A2(n680), .ZN(n557) );
  INV_X1 U652 ( .A(n558), .ZN(n559) );
  NAND2_X1 U653 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U654 ( .A(KEYINPUT104), .B(n561), .Z(n604) );
  NAND2_X1 U655 ( .A1(n562), .A2(n604), .ZN(n563) );
  NOR2_X1 U656 ( .A1(n563), .A2(n546), .ZN(n644) );
  OR2_X1 U657 ( .A1(n669), .A2(n565), .ZN(n566) );
  XNOR2_X1 U658 ( .A(n566), .B(KEYINPUT108), .ZN(n760) );
  NAND2_X1 U659 ( .A1(n567), .A2(n675), .ZN(n568) );
  NOR2_X1 U660 ( .A1(n685), .A2(n568), .ZN(n569) );
  NAND2_X1 U661 ( .A1(n451), .A2(n546), .ZN(n642) );
  AND2_X1 U662 ( .A1(n760), .A2(n642), .ZN(n570) );
  XNOR2_X1 U663 ( .A(n588), .B(KEYINPUT98), .ZN(n688) );
  AND2_X1 U664 ( .A1(n685), .A2(n688), .ZN(n571) );
  XNOR2_X1 U665 ( .A(KEYINPUT100), .B(n571), .ZN(n585) );
  INV_X1 U666 ( .A(n572), .ZN(n573) );
  XOR2_X1 U667 ( .A(G898), .B(KEYINPUT84), .Z(n733) );
  NAND2_X1 U668 ( .A1(n573), .A2(n733), .ZN(n574) );
  NAND2_X1 U669 ( .A1(n575), .A2(n574), .ZN(n576) );
  INV_X1 U670 ( .A(n689), .ZN(n579) );
  AND2_X1 U671 ( .A1(n580), .A2(n579), .ZN(n581) );
  NAND2_X1 U672 ( .A1(n613), .A2(n581), .ZN(n584) );
  INV_X1 U673 ( .A(KEYINPUT68), .ZN(n582) );
  XNOR2_X1 U674 ( .A(n582), .B(KEYINPUT22), .ZN(n583) );
  NAND2_X1 U675 ( .A1(n585), .A2(n618), .ZN(n586) );
  NAND2_X1 U676 ( .A1(n588), .A2(n587), .ZN(n589) );
  NOR2_X1 U677 ( .A1(n590), .A2(n589), .ZN(n591) );
  NAND2_X1 U678 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U679 ( .A(n593), .B(KEYINPUT102), .ZN(n757) );
  XNOR2_X1 U680 ( .A(KEYINPUT33), .B(KEYINPUT78), .ZN(n598) );
  XNOR2_X1 U681 ( .A(n600), .B(n599), .ZN(n674) );
  NOR2_X1 U682 ( .A1(n674), .A2(n609), .ZN(n603) );
  XNOR2_X1 U683 ( .A(KEYINPUT67), .B(KEYINPUT34), .ZN(n602) );
  XNOR2_X1 U684 ( .A(n603), .B(n602), .ZN(n606) );
  XOR2_X1 U685 ( .A(n604), .B(KEYINPUT70), .Z(n605) );
  INV_X1 U686 ( .A(n692), .ZN(n610) );
  NAND2_X1 U687 ( .A1(n692), .A2(n611), .ZN(n697) );
  INV_X1 U688 ( .A(n697), .ZN(n612) );
  NAND2_X1 U689 ( .A1(n613), .A2(n612), .ZN(n615) );
  INV_X1 U690 ( .A(KEYINPUT31), .ZN(n614) );
  NAND2_X1 U691 ( .A1(n657), .A2(n668), .ZN(n617) );
  INV_X1 U692 ( .A(n680), .ZN(n616) );
  XNOR2_X1 U693 ( .A(n618), .B(KEYINPUT74), .ZN(n620) );
  NOR2_X1 U694 ( .A1(n688), .A2(n685), .ZN(n619) );
  XNOR2_X1 U695 ( .A(n621), .B(KEYINPUT75), .ZN(n625) );
  NOR2_X1 U696 ( .A1(n753), .A2(KEYINPUT44), .ZN(n623) );
  NAND2_X1 U697 ( .A1(n623), .A2(n622), .ZN(n624) );
  NAND2_X1 U698 ( .A1(n625), .A2(n624), .ZN(n626) );
  NAND2_X1 U699 ( .A1(n714), .A2(G210), .ZN(n634) );
  XOR2_X1 U700 ( .A(KEYINPUT55), .B(KEYINPUT77), .Z(n629) );
  XNOR2_X1 U701 ( .A(KEYINPUT54), .B(KEYINPUT118), .ZN(n628) );
  XNOR2_X1 U702 ( .A(n629), .B(n628), .ZN(n632) );
  XOR2_X1 U703 ( .A(n632), .B(n631), .Z(n633) );
  XNOR2_X1 U704 ( .A(n634), .B(n633), .ZN(n638) );
  INV_X1 U705 ( .A(G952), .ZN(n635) );
  NAND2_X1 U706 ( .A1(n635), .A2(G953), .ZN(n637) );
  INV_X1 U707 ( .A(KEYINPUT79), .ZN(n636) );
  XNOR2_X1 U708 ( .A(n637), .B(n636), .ZN(n651) );
  NAND2_X1 U709 ( .A1(n638), .A2(n651), .ZN(n640) );
  INV_X1 U710 ( .A(KEYINPUT56), .ZN(n639) );
  XNOR2_X1 U711 ( .A(n640), .B(n639), .ZN(G51) );
  XNOR2_X1 U712 ( .A(n641), .B(G101), .ZN(G3) );
  XNOR2_X1 U713 ( .A(n642), .B(G140), .ZN(G42) );
  XNOR2_X1 U714 ( .A(n644), .B(n643), .ZN(G45) );
  XOR2_X1 U715 ( .A(KEYINPUT121), .B(KEYINPUT59), .Z(n645) );
  INV_X1 U716 ( .A(n651), .ZN(n728) );
  NAND2_X1 U717 ( .A1(n714), .A2(G472), .ZN(n650) );
  XNOR2_X1 U718 ( .A(KEYINPUT109), .B(n647), .ZN(n648) );
  XNOR2_X1 U719 ( .A(n650), .B(n649), .ZN(n652) );
  NAND2_X1 U720 ( .A1(n652), .A2(n651), .ZN(n653) );
  XNOR2_X1 U721 ( .A(n653), .B(KEYINPUT63), .ZN(G57) );
  NOR2_X1 U722 ( .A1(n665), .A2(n657), .ZN(n654) );
  XOR2_X1 U723 ( .A(G104), .B(n654), .Z(G6) );
  XOR2_X1 U724 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n656) );
  XNOR2_X1 U725 ( .A(G107), .B(KEYINPUT110), .ZN(n655) );
  XNOR2_X1 U726 ( .A(n656), .B(n655), .ZN(n659) );
  NOR2_X1 U727 ( .A1(n669), .A2(n657), .ZN(n658) );
  XOR2_X1 U728 ( .A(n659), .B(n658), .Z(G9) );
  NOR2_X1 U729 ( .A1(n663), .A2(n669), .ZN(n661) );
  XNOR2_X1 U730 ( .A(KEYINPUT29), .B(KEYINPUT112), .ZN(n660) );
  XNOR2_X1 U731 ( .A(n661), .B(n660), .ZN(n662) );
  XNOR2_X1 U732 ( .A(G128), .B(n662), .ZN(G30) );
  NOR2_X1 U733 ( .A1(n663), .A2(n665), .ZN(n664) );
  XOR2_X1 U734 ( .A(G146), .B(n664), .Z(G48) );
  NOR2_X1 U735 ( .A1(n665), .A2(n668), .ZN(n667) );
  XNOR2_X1 U736 ( .A(G113), .B(KEYINPUT113), .ZN(n666) );
  XNOR2_X1 U737 ( .A(n667), .B(n666), .ZN(G15) );
  NOR2_X1 U738 ( .A1(n669), .A2(n668), .ZN(n670) );
  XOR2_X1 U739 ( .A(KEYINPUT114), .B(n670), .Z(n671) );
  XNOR2_X1 U740 ( .A(G116), .B(n671), .ZN(G18) );
  XNOR2_X1 U741 ( .A(G125), .B(n672), .ZN(n673) );
  XNOR2_X1 U742 ( .A(n673), .B(KEYINPUT37), .ZN(G27) );
  BUF_X1 U743 ( .A(n674), .Z(n706) );
  NOR2_X1 U744 ( .A1(n676), .A2(n675), .ZN(n677) );
  NOR2_X1 U745 ( .A1(n678), .A2(n677), .ZN(n682) );
  NOR2_X1 U746 ( .A1(n680), .A2(n679), .ZN(n681) );
  NOR2_X1 U747 ( .A1(n682), .A2(n681), .ZN(n683) );
  NOR2_X1 U748 ( .A1(n706), .A2(n683), .ZN(n684) );
  XNOR2_X1 U749 ( .A(n684), .B(KEYINPUT117), .ZN(n702) );
  NOR2_X1 U750 ( .A1(n686), .A2(n685), .ZN(n687) );
  XOR2_X1 U751 ( .A(KEYINPUT50), .B(n687), .Z(n695) );
  NAND2_X1 U752 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U753 ( .A(KEYINPUT49), .B(n690), .ZN(n691) );
  NOR2_X1 U754 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U755 ( .A(KEYINPUT116), .B(n693), .ZN(n694) );
  NAND2_X1 U756 ( .A1(n695), .A2(n694), .ZN(n696) );
  NAND2_X1 U757 ( .A1(n697), .A2(n696), .ZN(n698) );
  XOR2_X1 U758 ( .A(KEYINPUT51), .B(n698), .Z(n700) );
  NAND2_X1 U759 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U760 ( .A1(n702), .A2(n701), .ZN(n703) );
  XOR2_X1 U761 ( .A(KEYINPUT52), .B(n703), .Z(n704) );
  NOR2_X1 U762 ( .A1(n705), .A2(n704), .ZN(n709) );
  NOR2_X1 U763 ( .A1(n707), .A2(n706), .ZN(n708) );
  NOR2_X1 U764 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U765 ( .A1(n711), .A2(n710), .ZN(n712) );
  NOR2_X1 U766 ( .A1(n712), .A2(G953), .ZN(n713) );
  XNOR2_X1 U767 ( .A(n713), .B(KEYINPUT53), .ZN(G75) );
  BUF_X2 U768 ( .A(n714), .Z(n724) );
  NAND2_X1 U769 ( .A1(n724), .A2(G469), .ZN(n719) );
  XOR2_X1 U770 ( .A(KEYINPUT119), .B(KEYINPUT120), .Z(n716) );
  XNOR2_X1 U771 ( .A(KEYINPUT58), .B(KEYINPUT57), .ZN(n715) );
  NOR2_X1 U772 ( .A1(n728), .A2(n720), .ZN(G54) );
  NAND2_X1 U773 ( .A1(n724), .A2(G478), .ZN(n722) );
  XNOR2_X1 U774 ( .A(n722), .B(n721), .ZN(n723) );
  NOR2_X1 U775 ( .A1(n728), .A2(n723), .ZN(G63) );
  NAND2_X1 U776 ( .A1(n724), .A2(G217), .ZN(n726) );
  XNOR2_X1 U777 ( .A(n726), .B(n725), .ZN(n727) );
  NOR2_X1 U778 ( .A1(n728), .A2(n727), .ZN(G66) );
  NAND2_X1 U779 ( .A1(G953), .A2(G224), .ZN(n729) );
  XOR2_X1 U780 ( .A(KEYINPUT61), .B(n729), .Z(n730) );
  OR2_X1 U781 ( .A1(n733), .A2(n730), .ZN(n731) );
  NAND2_X1 U782 ( .A1(n733), .A2(G953), .ZN(n738) );
  XNOR2_X1 U783 ( .A(n734), .B(G101), .ZN(n735) );
  XNOR2_X1 U784 ( .A(n736), .B(n735), .ZN(n737) );
  NAND2_X1 U785 ( .A1(n738), .A2(n737), .ZN(n739) );
  XNOR2_X1 U786 ( .A(n739), .B(KEYINPUT122), .ZN(n740) );
  XNOR2_X1 U787 ( .A(n352), .B(n740), .ZN(G69) );
  XNOR2_X1 U788 ( .A(n741), .B(KEYINPUT123), .ZN(n744) );
  XNOR2_X1 U789 ( .A(n742), .B(KEYINPUT4), .ZN(n743) );
  XNOR2_X1 U790 ( .A(n744), .B(n743), .ZN(n748) );
  XOR2_X1 U791 ( .A(G227), .B(n748), .Z(n745) );
  NAND2_X1 U792 ( .A1(n745), .A2(G900), .ZN(n746) );
  NAND2_X1 U793 ( .A1(n746), .A2(G953), .ZN(n752) );
  XNOR2_X1 U794 ( .A(n748), .B(n747), .ZN(n749) );
  NOR2_X1 U795 ( .A1(G953), .A2(n749), .ZN(n750) );
  XOR2_X1 U796 ( .A(KEYINPUT124), .B(n750), .Z(n751) );
  XOR2_X1 U797 ( .A(n753), .B(G122), .Z(n754) );
  XNOR2_X1 U798 ( .A(KEYINPUT126), .B(n754), .ZN(G24) );
  XOR2_X1 U799 ( .A(G119), .B(n755), .Z(n756) );
  XNOR2_X1 U800 ( .A(KEYINPUT127), .B(n756), .ZN(G21) );
  XOR2_X1 U801 ( .A(G110), .B(n757), .Z(n758) );
  XNOR2_X1 U802 ( .A(KEYINPUT111), .B(n758), .ZN(G12) );
  XOR2_X1 U803 ( .A(G131), .B(n759), .Z(G33) );
  XOR2_X1 U804 ( .A(G134), .B(n760), .Z(n761) );
  XNOR2_X1 U805 ( .A(KEYINPUT115), .B(n761), .ZN(G36) );
  XOR2_X1 U806 ( .A(G137), .B(n762), .Z(G39) );
endmodule

