//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 0 0 1 0 1 1 1 0 1 1 0 0 1 1 1 0 0 1 1 0 1 0 1 0 0 0 0 1 1 1 1 0 1 0 1 0 0 0 1 1 1 1 0 0 0 1 0 0 1 1 1 0 0 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:42 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n564,
    new_n566, new_n567, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n582, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n619, new_n622, new_n624, new_n625, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1226,
    new_n1227, new_n1228, new_n1229;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(G261));
  INV_X1    g028(.A(G261), .ZN(G325));
  INV_X1    g029(.A(G2106), .ZN(new_n455));
  INV_X1    g030(.A(G567), .ZN(new_n456));
  OAI22_X1  g031(.A1(new_n451), .A2(new_n455), .B1(new_n456), .B2(new_n452), .ZN(new_n457));
  XNOR2_X1  g032(.A(new_n457), .B(KEYINPUT64), .ZN(G319));
  INV_X1    g033(.A(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n459), .A2(G2105), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G101), .ZN(new_n461));
  OR2_X1    g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G137), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n461), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n464), .A2(G125), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n465), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n468), .A2(new_n471), .ZN(G160));
  OR2_X1    g047(.A1(G100), .A2(G2105), .ZN(new_n473));
  OAI211_X1 g048(.A(new_n473), .B(G2104), .C1(G112), .C2(new_n465), .ZN(new_n474));
  XNOR2_X1  g049(.A(new_n474), .B(KEYINPUT66), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT65), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n466), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n464), .A2(KEYINPUT65), .A3(new_n465), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  AND2_X1   g055(.A1(new_n480), .A2(G136), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n465), .B1(new_n462), .B2(new_n463), .ZN(new_n482));
  AOI211_X1 g057(.A(new_n475), .B(new_n481), .C1(G124), .C2(new_n482), .ZN(G162));
  AND2_X1   g058(.A1(KEYINPUT68), .A2(G138), .ZN(new_n484));
  AND2_X1   g059(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n485));
  NOR2_X1   g060(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n465), .B(new_n484), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(KEYINPUT4), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n464), .A2(new_n489), .A3(new_n465), .A4(new_n484), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  OAI21_X1  g066(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(G114), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G2105), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n493), .A2(KEYINPUT67), .A3(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT67), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n465), .A2(G114), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n497), .B1(new_n498), .B2(new_n492), .ZN(new_n499));
  AOI22_X1  g074(.A1(new_n496), .A2(new_n499), .B1(new_n482), .B2(G126), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n491), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(G164));
  INV_X1    g077(.A(G543), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT5), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n503), .B1(new_n504), .B2(KEYINPUT69), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT69), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n506), .A2(KEYINPUT5), .A3(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  AOI22_X1  g083(.A1(new_n508), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n509));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  OR2_X1    g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  XOR2_X1   g086(.A(KEYINPUT70), .B(G88), .Z(new_n512));
  XNOR2_X1  g087(.A(KEYINPUT6), .B(G651), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n512), .A2(new_n508), .A3(new_n513), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n513), .A2(G50), .A3(G543), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n514), .A2(KEYINPUT71), .A3(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(new_n516), .ZN(new_n517));
  AOI21_X1  g092(.A(KEYINPUT71), .B1(new_n514), .B2(new_n515), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n511), .B1(new_n517), .B2(new_n518), .ZN(G303));
  INV_X1    g094(.A(G303), .ZN(G166));
  INV_X1    g095(.A(KEYINPUT74), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n508), .A2(G89), .A3(new_n513), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT73), .ZN(new_n523));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  INV_X1    g099(.A(new_n524), .ZN(new_n525));
  NOR2_X1   g100(.A1(KEYINPUT72), .A2(KEYINPUT7), .ZN(new_n526));
  INV_X1    g101(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(KEYINPUT72), .A2(KEYINPUT7), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n525), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(new_n528), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n524), .B1(new_n530), .B2(new_n526), .ZN(new_n531));
  NAND4_X1  g106(.A1(new_n522), .A2(new_n523), .A3(new_n529), .A4(new_n531), .ZN(new_n532));
  AND2_X1   g107(.A1(KEYINPUT6), .A2(G651), .ZN(new_n533));
  NOR2_X1   g108(.A1(KEYINPUT6), .A2(G651), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n535), .A2(new_n503), .ZN(new_n536));
  AND2_X1   g111(.A1(G63), .A2(G651), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n536), .A2(G51), .B1(new_n508), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n532), .A2(new_n538), .ZN(new_n539));
  AND2_X1   g114(.A1(new_n529), .A2(new_n531), .ZN(new_n540));
  AOI21_X1  g115(.A(new_n523), .B1(new_n540), .B2(new_n522), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n521), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n522), .A2(new_n529), .A3(new_n531), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(KEYINPUT73), .ZN(new_n544));
  NAND4_X1  g119(.A1(new_n544), .A2(KEYINPUT74), .A3(new_n532), .A4(new_n538), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n542), .A2(new_n545), .ZN(G168));
  AOI22_X1  g121(.A1(new_n508), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n547), .A2(new_n510), .ZN(new_n548));
  AND3_X1   g123(.A1(new_n506), .A2(KEYINPUT5), .A3(G543), .ZN(new_n549));
  AOI21_X1  g124(.A(G543), .B1(new_n506), .B2(KEYINPUT5), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n513), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(G90), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n513), .A2(G543), .ZN(new_n553));
  INV_X1    g128(.A(G52), .ZN(new_n554));
  OAI22_X1  g129(.A1(new_n551), .A2(new_n552), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n548), .A2(new_n555), .ZN(G171));
  AOI22_X1  g131(.A1(new_n508), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n557), .A2(new_n510), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n508), .A2(G81), .A3(new_n513), .ZN(new_n559));
  INV_X1    g134(.A(G43), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n559), .B1(new_n560), .B2(new_n553), .ZN(new_n561));
  NOR2_X1   g136(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G860), .ZN(G153));
  NAND4_X1  g138(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT75), .ZN(G176));
  NAND2_X1  g140(.A1(G1), .A2(G3), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT8), .ZN(new_n567));
  NAND4_X1  g142(.A1(G319), .A2(G483), .A3(G661), .A4(new_n567), .ZN(G188));
  INV_X1    g143(.A(KEYINPUT76), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n551), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n508), .A2(KEYINPUT76), .A3(new_n513), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n570), .A2(G91), .A3(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(G65), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n573), .B1(new_n505), .B2(new_n507), .ZN(new_n574));
  AND2_X1   g149(.A1(G78), .A2(G543), .ZN(new_n575));
  OAI21_X1  g150(.A(G651), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  OAI211_X1 g151(.A(G53), .B(G543), .C1(new_n533), .C2(new_n534), .ZN(new_n577));
  XNOR2_X1  g152(.A(new_n577), .B(KEYINPUT9), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n572), .A2(new_n576), .A3(new_n578), .ZN(G299));
  INV_X1    g154(.A(G171), .ZN(G301));
  INV_X1    g155(.A(G168), .ZN(G286));
  NAND3_X1  g156(.A1(new_n570), .A2(G87), .A3(new_n571), .ZN(new_n582));
  INV_X1    g157(.A(G74), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n505), .A2(new_n583), .A3(new_n507), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n536), .A2(G49), .B1(G651), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n582), .A2(new_n585), .ZN(G288));
  NAND3_X1  g161(.A1(new_n570), .A2(G86), .A3(new_n571), .ZN(new_n587));
  INV_X1    g162(.A(G61), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n588), .B1(new_n505), .B2(new_n507), .ZN(new_n589));
  AND2_X1   g164(.A1(G73), .A2(G543), .ZN(new_n590));
  OAI21_X1  g165(.A(G651), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT77), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  OAI211_X1 g168(.A(KEYINPUT77), .B(G651), .C1(new_n589), .C2(new_n590), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n513), .A2(G48), .A3(G543), .ZN(new_n595));
  NAND4_X1  g170(.A1(new_n587), .A2(new_n593), .A3(new_n594), .A4(new_n595), .ZN(G305));
  NAND2_X1  g171(.A1(new_n508), .A2(G60), .ZN(new_n597));
  INV_X1    g172(.A(G72), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n598), .B2(new_n503), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n599), .A2(G651), .ZN(new_n600));
  XNOR2_X1  g175(.A(KEYINPUT78), .B(G85), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n508), .A2(new_n513), .A3(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT79), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n513), .A2(G47), .A3(G543), .ZN(new_n604));
  AND3_X1   g179(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n603), .B1(new_n602), .B2(new_n604), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n600), .B1(new_n605), .B2(new_n606), .ZN(G290));
  NAND2_X1  g182(.A1(G301), .A2(G868), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n536), .A2(G54), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n508), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n610), .B2(new_n510), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n570), .A2(G92), .A3(new_n571), .ZN(new_n612));
  INV_X1    g187(.A(KEYINPUT10), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND4_X1  g189(.A1(new_n570), .A2(KEYINPUT10), .A3(G92), .A4(new_n571), .ZN(new_n615));
  AOI21_X1  g190(.A(new_n611), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n608), .B1(new_n616), .B2(G868), .ZN(G284));
  OAI21_X1  g192(.A(new_n608), .B1(new_n616), .B2(G868), .ZN(G321));
  NOR2_X1   g193(.A1(G299), .A2(G868), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n619), .B1(G168), .B2(G868), .ZN(G297));
  AOI21_X1  g195(.A(new_n619), .B1(G168), .B2(G868), .ZN(G280));
  INV_X1    g196(.A(G559), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n616), .B1(new_n622), .B2(G860), .ZN(G148));
  INV_X1    g198(.A(new_n616), .ZN(new_n624));
  OAI21_X1  g199(.A(G868), .B1(new_n624), .B2(G559), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n625), .B1(G868), .B2(new_n562), .ZN(G323));
  XNOR2_X1  g201(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g202(.A1(new_n464), .A2(new_n460), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT12), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT13), .ZN(new_n630));
  INV_X1    g205(.A(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n482), .A2(G123), .ZN(new_n632));
  NOR2_X1   g207(.A1(new_n465), .A2(G111), .ZN(new_n633));
  OAI21_X1  g208(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n634));
  INV_X1    g209(.A(G135), .ZN(new_n635));
  OAI221_X1 g210(.A(new_n632), .B1(new_n633), .B2(new_n634), .C1(new_n479), .C2(new_n635), .ZN(new_n636));
  AOI22_X1  g211(.A1(new_n631), .A2(G2100), .B1(G2096), .B2(new_n636), .ZN(new_n637));
  OR2_X1    g212(.A1(new_n636), .A2(G2096), .ZN(new_n638));
  OAI211_X1 g213(.A(new_n637), .B(new_n638), .C1(G2100), .C2(new_n631), .ZN(G156));
  XOR2_X1   g214(.A(G1341), .B(G1348), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT80), .ZN(new_n641));
  XOR2_X1   g216(.A(G2451), .B(G2454), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT16), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n641), .B(new_n643), .Z(new_n644));
  INV_X1    g219(.A(KEYINPUT14), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2427), .B(G2438), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(G2430), .ZN(new_n647));
  XNOR2_X1  g222(.A(KEYINPUT15), .B(G2435), .ZN(new_n648));
  AOI21_X1  g223(.A(new_n645), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n649), .B1(new_n648), .B2(new_n647), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n644), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2443), .B(G2446), .ZN(new_n652));
  OR2_X1    g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n651), .A2(new_n652), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n653), .A2(G14), .A3(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(new_n655), .B(KEYINPUT81), .Z(G401));
  XNOR2_X1  g231(.A(G2072), .B(G2078), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n657), .B(KEYINPUT17), .Z(new_n658));
  XNOR2_X1  g233(.A(G2067), .B(G2678), .ZN(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(G2084), .B(G2090), .Z(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  OAI21_X1  g238(.A(new_n663), .B1(new_n659), .B2(new_n657), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n665), .B(KEYINPUT82), .Z(new_n666));
  NAND3_X1  g241(.A1(new_n662), .A2(new_n659), .A3(new_n657), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT18), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n663), .A2(new_n659), .ZN(new_n669));
  AOI21_X1  g244(.A(new_n668), .B1(new_n658), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n666), .A2(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(G2096), .B(G2100), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(G227));
  XNOR2_X1  g248(.A(G1971), .B(G1976), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT84), .ZN(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT83), .B(KEYINPUT19), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1956), .B(G2474), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1961), .B(G1966), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT20), .ZN(new_n682));
  AND2_X1   g257(.A1(new_n678), .A2(new_n679), .ZN(new_n683));
  NOR3_X1   g258(.A1(new_n677), .A2(new_n680), .A3(new_n683), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n684), .B1(new_n677), .B2(new_n683), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XOR2_X1   g263(.A(G1991), .B(G1996), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1981), .B(G1986), .ZN(new_n691));
  OR2_X1    g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n690), .A2(new_n691), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(G229));
  NAND2_X1  g270(.A1(G166), .A2(G16), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n696), .B1(G16), .B2(G22), .ZN(new_n697));
  INV_X1    g272(.A(G1971), .ZN(new_n698));
  XOR2_X1   g273(.A(KEYINPUT32), .B(G1981), .Z(new_n699));
  INV_X1    g274(.A(G16), .ZN(new_n700));
  AND2_X1   g275(.A1(new_n700), .A2(G6), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n701), .B1(G305), .B2(G16), .ZN(new_n702));
  AOI22_X1  g277(.A1(new_n697), .A2(new_n698), .B1(new_n699), .B2(new_n702), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n703), .B1(new_n698), .B2(new_n697), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n700), .A2(G23), .ZN(new_n705));
  AND2_X1   g280(.A1(new_n582), .A2(new_n585), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n705), .B1(new_n706), .B2(new_n700), .ZN(new_n707));
  XNOR2_X1  g282(.A(KEYINPUT33), .B(G1976), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(new_n702), .B2(new_n699), .ZN(new_n710));
  NOR3_X1   g285(.A1(new_n704), .A2(KEYINPUT34), .A3(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(G29), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(G25), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n480), .A2(G131), .ZN(new_n714));
  NOR2_X1   g289(.A1(G95), .A2(G2105), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT85), .ZN(new_n716));
  INV_X1    g291(.A(G107), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n459), .B1(new_n717), .B2(G2105), .ZN(new_n718));
  AOI22_X1  g293(.A1(new_n716), .A2(new_n718), .B1(G119), .B2(new_n482), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n714), .A2(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n713), .B1(new_n721), .B2(new_n712), .ZN(new_n722));
  XOR2_X1   g297(.A(KEYINPUT35), .B(G1991), .Z(new_n723));
  XOR2_X1   g298(.A(new_n722), .B(new_n723), .Z(new_n724));
  NAND2_X1  g299(.A1(new_n700), .A2(G24), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n602), .A2(new_n604), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n726), .A2(KEYINPUT79), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(new_n728));
  AOI22_X1  g303(.A1(new_n727), .A2(new_n728), .B1(G651), .B2(new_n599), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n725), .B1(new_n729), .B2(new_n700), .ZN(new_n730));
  XNOR2_X1  g305(.A(KEYINPUT86), .B(G1986), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  NOR3_X1   g307(.A1(new_n711), .A2(new_n724), .A3(new_n732), .ZN(new_n733));
  OAI21_X1  g308(.A(KEYINPUT34), .B1(new_n704), .B2(new_n710), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g310(.A(KEYINPUT36), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n712), .A2(G35), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(G162), .B2(new_n712), .ZN(new_n739));
  XOR2_X1   g314(.A(KEYINPUT29), .B(G2090), .Z(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  XOR2_X1   g316(.A(KEYINPUT31), .B(G11), .Z(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT90), .ZN(new_n743));
  INV_X1    g318(.A(KEYINPUT30), .ZN(new_n744));
  AND2_X1   g319(.A1(new_n744), .A2(G28), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n712), .B1(new_n744), .B2(G28), .ZN(new_n746));
  OAI221_X1 g321(.A(new_n743), .B1(new_n745), .B2(new_n746), .C1(new_n636), .C2(new_n712), .ZN(new_n747));
  NAND2_X1  g322(.A1(G160), .A2(G29), .ZN(new_n748));
  XNOR2_X1  g323(.A(KEYINPUT24), .B(G34), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n749), .A2(new_n712), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT87), .ZN(new_n751));
  AOI21_X1  g326(.A(G2084), .B1(new_n748), .B2(new_n751), .ZN(new_n752));
  AND3_X1   g327(.A1(new_n748), .A2(G2084), .A3(new_n751), .ZN(new_n753));
  NOR3_X1   g328(.A1(new_n747), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n700), .A2(G19), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(new_n562), .B2(new_n700), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(G1341), .Z(new_n757));
  NAND2_X1  g332(.A1(new_n712), .A2(G26), .ZN(new_n758));
  XOR2_X1   g333(.A(new_n758), .B(KEYINPUT28), .Z(new_n759));
  NAND2_X1  g334(.A1(new_n480), .A2(G140), .ZN(new_n760));
  OAI21_X1  g335(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n761));
  INV_X1    g336(.A(G116), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n761), .B1(new_n762), .B2(G2105), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(G128), .B2(new_n482), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n760), .A2(new_n764), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n759), .B1(new_n765), .B2(G29), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(G2067), .ZN(new_n767));
  AND4_X1   g342(.A1(new_n741), .A2(new_n754), .A3(new_n757), .A4(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n712), .A2(G32), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n480), .A2(G141), .ZN(new_n770));
  AND2_X1   g345(.A1(new_n460), .A2(G105), .ZN(new_n771));
  NAND3_X1  g346(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT26), .ZN(new_n773));
  AOI211_X1 g348(.A(new_n771), .B(new_n773), .C1(G129), .C2(new_n482), .ZN(new_n774));
  AND2_X1   g349(.A1(new_n770), .A2(new_n774), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n769), .B1(new_n775), .B2(new_n712), .ZN(new_n776));
  XNOR2_X1  g351(.A(KEYINPUT27), .B(G1996), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n712), .A2(G27), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G164), .B2(new_n712), .ZN(new_n780));
  XOR2_X1   g355(.A(new_n780), .B(G2078), .Z(new_n781));
  NAND2_X1  g356(.A1(new_n778), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n712), .A2(G33), .ZN(new_n783));
  NAND3_X1  g358(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n784), .B(KEYINPUT25), .Z(new_n785));
  AOI22_X1  g360(.A1(new_n464), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n785), .B1(new_n786), .B2(new_n465), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(new_n480), .B2(G139), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n783), .B1(new_n788), .B2(new_n712), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(G2072), .ZN(new_n790));
  NOR2_X1   g365(.A1(G5), .A2(G16), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(G171), .B2(G16), .ZN(new_n792));
  XNOR2_X1  g367(.A(KEYINPUT91), .B(G1961), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NOR3_X1   g369(.A1(new_n782), .A2(new_n790), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n700), .A2(G20), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT23), .ZN(new_n797));
  INV_X1    g372(.A(G299), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n797), .B1(new_n798), .B2(new_n700), .ZN(new_n799));
  INV_X1    g374(.A(G1956), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  NOR2_X1   g376(.A1(G4), .A2(G16), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(new_n616), .B2(G16), .ZN(new_n803));
  INV_X1    g378(.A(G1348), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  NAND4_X1  g380(.A1(new_n768), .A2(new_n795), .A3(new_n801), .A4(new_n805), .ZN(new_n806));
  NOR2_X1   g381(.A1(G16), .A2(G21), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n807), .B1(G168), .B2(G16), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT88), .ZN(new_n809));
  XOR2_X1   g384(.A(KEYINPUT89), .B(G1966), .Z(new_n810));
  AND2_X1   g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n809), .A2(new_n810), .ZN(new_n812));
  OR3_X1    g387(.A1(new_n806), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n737), .A2(new_n813), .ZN(G311));
  INV_X1    g389(.A(G311), .ZN(G150));
  NAND2_X1  g390(.A1(new_n536), .A2(G55), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n508), .A2(G93), .A3(new_n513), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n508), .A2(G67), .ZN(new_n819));
  NAND2_X1  g394(.A1(G80), .A2(G543), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n510), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  OAI21_X1  g396(.A(KEYINPUT92), .B1(new_n818), .B2(new_n821), .ZN(new_n822));
  OAI221_X1 g397(.A(new_n559), .B1(new_n560), .B2(new_n553), .C1(new_n557), .C2(new_n510), .ZN(new_n823));
  INV_X1    g398(.A(G67), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n824), .B1(new_n505), .B2(new_n507), .ZN(new_n825));
  INV_X1    g400(.A(new_n820), .ZN(new_n826));
  OAI21_X1  g401(.A(G651), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT92), .ZN(new_n828));
  NAND4_X1  g403(.A1(new_n827), .A2(new_n816), .A3(new_n828), .A4(new_n817), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n822), .A2(new_n823), .A3(new_n829), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n818), .A2(new_n821), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n562), .A2(new_n831), .A3(new_n828), .ZN(new_n832));
  AND2_X1   g407(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT38), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n616), .A2(G559), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n834), .B(new_n835), .ZN(new_n836));
  OR2_X1    g411(.A1(new_n836), .A2(KEYINPUT39), .ZN(new_n837));
  INV_X1    g412(.A(G860), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n836), .A2(KEYINPUT39), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n837), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n831), .A2(new_n838), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT37), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n840), .A2(new_n842), .ZN(G145));
  NAND2_X1  g418(.A1(new_n482), .A2(G130), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n465), .A2(G118), .ZN(new_n845));
  OAI21_X1  g420(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n844), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n847), .B1(new_n480), .B2(G142), .ZN(new_n848));
  XOR2_X1   g423(.A(new_n848), .B(new_n629), .Z(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(new_n720), .ZN(new_n850));
  INV_X1    g425(.A(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(new_n765), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n852), .A2(new_n775), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n770), .A2(new_n774), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n765), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n856), .A2(G164), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(new_n788), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n856), .A2(G164), .ZN(new_n860));
  NOR3_X1   g435(.A1(new_n858), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  AND2_X1   g436(.A1(new_n853), .A2(new_n855), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n862), .A2(new_n501), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n788), .B1(new_n863), .B2(new_n857), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n851), .B1(new_n861), .B2(new_n864), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n859), .B1(new_n858), .B2(new_n860), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n863), .A2(new_n788), .A3(new_n857), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n866), .A2(new_n850), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n865), .A2(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n636), .B(G160), .ZN(new_n870));
  XNOR2_X1  g445(.A(G162), .B(new_n870), .ZN(new_n871));
  AOI21_X1  g446(.A(G37), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n868), .A2(KEYINPUT93), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT93), .ZN(new_n874));
  NAND4_X1  g449(.A1(new_n866), .A2(new_n874), .A3(new_n850), .A4(new_n867), .ZN(new_n875));
  INV_X1    g450(.A(new_n871), .ZN(new_n876));
  NAND4_X1  g451(.A1(new_n873), .A2(new_n875), .A3(new_n865), .A4(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n872), .A2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT94), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n872), .A2(KEYINPUT94), .A3(new_n877), .ZN(new_n881));
  AND3_X1   g456(.A1(new_n880), .A2(KEYINPUT40), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(KEYINPUT40), .B1(new_n880), .B2(new_n881), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n882), .A2(new_n883), .ZN(G395));
  INV_X1    g459(.A(KEYINPUT97), .ZN(new_n885));
  OAI211_X1 g460(.A(G288), .B(new_n511), .C1(new_n518), .C2(new_n517), .ZN(new_n886));
  AND2_X1   g461(.A1(new_n593), .A2(new_n594), .ZN(new_n887));
  INV_X1    g462(.A(new_n595), .ZN(new_n888));
  AND3_X1   g463(.A1(new_n508), .A2(KEYINPUT76), .A3(new_n513), .ZN(new_n889));
  AOI21_X1  g464(.A(KEYINPUT76), .B1(new_n508), .B2(new_n513), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n888), .B1(new_n891), .B2(G86), .ZN(new_n892));
  NAND3_X1  g467(.A1(G290), .A2(new_n887), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(G303), .A2(new_n706), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n729), .A2(G305), .ZN(new_n895));
  AND4_X1   g470(.A1(new_n886), .A2(new_n893), .A3(new_n894), .A4(new_n895), .ZN(new_n896));
  AOI22_X1  g471(.A1(new_n895), .A2(new_n893), .B1(new_n894), .B2(new_n886), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n885), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n893), .A2(new_n895), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n894), .A2(new_n886), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND4_X1  g476(.A1(new_n893), .A2(new_n894), .A3(new_n895), .A4(new_n886), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n901), .A2(KEYINPUT98), .A3(new_n902), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n898), .B1(new_n885), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(KEYINPUT42), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT42), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n903), .A2(new_n906), .ZN(new_n907));
  AND2_X1   g482(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  OR2_X1    g483(.A1(new_n908), .A2(KEYINPUT99), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n572), .A2(KEYINPUT95), .A3(new_n576), .A4(new_n578), .ZN(new_n910));
  INV_X1    g485(.A(new_n611), .ZN(new_n911));
  AOI21_X1  g486(.A(KEYINPUT10), .B1(new_n891), .B2(G92), .ZN(new_n912));
  INV_X1    g487(.A(new_n615), .ZN(new_n913));
  OAI211_X1 g488(.A(new_n910), .B(new_n911), .C1(new_n912), .C2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT95), .ZN(new_n915));
  NAND2_X1  g490(.A1(G299), .A2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n914), .A2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT41), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n616), .A2(new_n916), .A3(new_n910), .ZN(new_n920));
  AND3_X1   g495(.A1(new_n918), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n919), .B1(new_n918), .B2(new_n920), .ZN(new_n922));
  OAI21_X1  g497(.A(KEYINPUT96), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT96), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n918), .A2(new_n919), .A3(new_n920), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n924), .B1(new_n925), .B2(KEYINPUT41), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n923), .A2(new_n926), .ZN(new_n927));
  AND3_X1   g502(.A1(new_n616), .A2(new_n916), .A3(new_n910), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n916), .B1(new_n616), .B2(new_n910), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n616), .A2(new_n622), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n830), .A2(new_n832), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n931), .B(new_n932), .ZN(new_n933));
  MUX2_X1   g508(.A(new_n927), .B(new_n930), .S(new_n933), .Z(new_n934));
  NAND2_X1  g509(.A1(new_n908), .A2(KEYINPUT99), .ZN(new_n935));
  AND3_X1   g510(.A1(new_n909), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n934), .B1(new_n909), .B2(new_n935), .ZN(new_n937));
  OAI21_X1  g512(.A(G868), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n938), .B1(G868), .B2(new_n831), .ZN(G295));
  OAI21_X1  g514(.A(new_n938), .B1(G868), .B2(new_n831), .ZN(G331));
  INV_X1    g515(.A(KEYINPUT101), .ZN(new_n941));
  NAND2_X1  g516(.A1(G168), .A2(G171), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n542), .A2(new_n545), .A3(G301), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n942), .A2(new_n833), .A3(new_n943), .ZN(new_n944));
  AND3_X1   g519(.A1(new_n542), .A2(new_n545), .A3(G301), .ZN(new_n945));
  AOI21_X1  g520(.A(G301), .B1(new_n542), .B2(new_n545), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n932), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n944), .A2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n949), .B1(new_n923), .B2(new_n926), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n930), .A2(new_n944), .A3(new_n947), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n901), .A2(KEYINPUT97), .A3(new_n902), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n951), .A2(new_n952), .A3(new_n898), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n941), .B1(new_n950), .B2(new_n953), .ZN(new_n954));
  OAI21_X1  g529(.A(KEYINPUT41), .B1(new_n928), .B2(new_n929), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n924), .B1(new_n955), .B2(new_n925), .ZN(new_n956));
  AOI21_X1  g531(.A(KEYINPUT96), .B1(new_n930), .B2(new_n919), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n948), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n898), .A2(new_n952), .ZN(new_n959));
  INV_X1    g534(.A(new_n959), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n958), .A2(KEYINPUT101), .A3(new_n960), .A4(new_n951), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n949), .A2(KEYINPUT102), .A3(new_n930), .ZN(new_n962));
  AOI22_X1  g537(.A1(new_n925), .A2(new_n955), .B1(new_n944), .B2(new_n947), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT102), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n951), .A2(new_n964), .ZN(new_n965));
  OAI211_X1 g540(.A(new_n962), .B(new_n959), .C1(new_n963), .C2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(G37), .ZN(new_n967));
  NAND4_X1  g542(.A1(new_n954), .A2(new_n961), .A3(new_n966), .A4(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT103), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n953), .B1(new_n927), .B2(new_n948), .ZN(new_n971));
  AOI21_X1  g546(.A(G37), .B1(new_n971), .B2(KEYINPUT101), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n972), .A2(KEYINPUT103), .A3(new_n954), .A4(new_n966), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n970), .A2(new_n973), .A3(KEYINPUT43), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(KEYINPUT104), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT104), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n970), .A2(new_n973), .A3(new_n976), .A4(KEYINPUT43), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n954), .A2(new_n961), .A3(new_n967), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n960), .B1(new_n958), .B2(new_n951), .ZN(new_n979));
  NOR3_X1   g554(.A1(new_n978), .A2(KEYINPUT43), .A3(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT44), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n975), .A2(new_n977), .A3(new_n982), .ZN(new_n983));
  OAI21_X1  g558(.A(KEYINPUT43), .B1(new_n978), .B2(new_n979), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n984), .B1(KEYINPUT43), .B2(new_n968), .ZN(new_n985));
  XNOR2_X1  g560(.A(KEYINPUT100), .B(KEYINPUT44), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n983), .A2(new_n987), .ZN(G397));
  INV_X1    g563(.A(G1384), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n501), .A2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(G40), .ZN(new_n991));
  NOR3_X1   g566(.A1(new_n468), .A2(new_n471), .A3(new_n991), .ZN(new_n992));
  XNOR2_X1  g567(.A(KEYINPUT105), .B(KEYINPUT45), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n990), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  XNOR2_X1  g569(.A(new_n994), .B(KEYINPUT106), .ZN(new_n995));
  INV_X1    g570(.A(new_n995), .ZN(new_n996));
  OR2_X1    g571(.A1(new_n996), .A2(KEYINPUT107), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(KEYINPUT107), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  XNOR2_X1  g574(.A(new_n765), .B(G2067), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n1000), .A2(new_n854), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT46), .ZN(new_n1002));
  INV_X1    g577(.A(G1996), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n995), .A2(new_n1003), .ZN(new_n1004));
  OAI22_X1  g579(.A1(new_n999), .A2(new_n1001), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1002), .ZN(new_n1006));
  XNOR2_X1  g581(.A(new_n1006), .B(KEYINPUT125), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT126), .ZN(new_n1008));
  OR3_X1    g583(.A1(new_n1005), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1008), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT47), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n775), .A2(new_n1003), .ZN(new_n1014));
  OAI211_X1 g589(.A(new_n997), .B(new_n998), .C1(new_n1000), .C2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1015), .B1(new_n854), .B2(new_n1004), .ZN(new_n1016));
  AND2_X1   g591(.A1(new_n997), .A2(new_n998), .ZN(new_n1017));
  XOR2_X1   g592(.A(new_n720), .B(new_n723), .Z(new_n1018));
  AOI21_X1  g593(.A(new_n1016), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  NOR3_X1   g594(.A1(new_n996), .A2(G1986), .A3(G290), .ZN(new_n1020));
  XNOR2_X1  g595(.A(KEYINPUT127), .B(KEYINPUT48), .ZN(new_n1021));
  XNOR2_X1  g596(.A(new_n1020), .B(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n721), .A2(new_n723), .ZN(new_n1023));
  OAI22_X1  g598(.A1(new_n1016), .A2(new_n1023), .B1(G2067), .B2(new_n765), .ZN(new_n1024));
  AOI22_X1  g599(.A1(new_n1019), .A2(new_n1022), .B1(new_n1024), .B2(new_n1017), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1009), .A2(KEYINPUT47), .A3(new_n1010), .ZN(new_n1026));
  AND3_X1   g601(.A1(new_n1013), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(G1981), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n887), .A2(new_n892), .A3(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1029), .ZN(new_n1030));
  XNOR2_X1  g605(.A(KEYINPUT109), .B(G86), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n508), .A2(new_n513), .A3(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(new_n595), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(KEYINPUT110), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT110), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1032), .A2(new_n1035), .A3(new_n595), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n1034), .A2(new_n593), .A3(new_n594), .A4(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(G1981), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1029), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT49), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(G8), .ZN(new_n1042));
  AOI21_X1  g617(.A(G1384), .B1(new_n491), .B2(new_n500), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT108), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  AOI211_X1 g620(.A(KEYINPUT108), .B(G1384), .C1(new_n491), .C2(new_n500), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1042), .B1(new_n1047), .B2(new_n992), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1029), .A2(new_n1038), .A3(KEYINPUT49), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1041), .A2(new_n1048), .A3(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT111), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1041), .A2(new_n1048), .A3(KEYINPUT111), .A4(new_n1049), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NOR2_X1   g629(.A1(G288), .A2(G1976), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1030), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1048), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n990), .A2(KEYINPUT108), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1058), .A2(new_n992), .A3(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n706), .A2(G1976), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1060), .A2(G8), .A3(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(KEYINPUT52), .ZN(new_n1063));
  INV_X1    g638(.A(G1976), .ZN(new_n1064));
  AOI21_X1  g639(.A(KEYINPUT52), .B1(G288), .B2(new_n1064), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1060), .A2(G8), .A3(new_n1061), .A4(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1063), .A2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1067), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(G303), .A2(G8), .ZN(new_n1070));
  XNOR2_X1  g645(.A(new_n1070), .B(KEYINPUT55), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT50), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1058), .A2(new_n1073), .A3(new_n1059), .ZN(new_n1074));
  INV_X1    g649(.A(G2090), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n992), .B1(new_n1043), .B2(new_n1073), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1074), .A2(new_n1075), .A3(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n990), .A2(new_n993), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1043), .A2(KEYINPUT45), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1079), .A2(new_n992), .A3(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(new_n698), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1078), .A2(new_n1082), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1072), .A2(new_n1083), .A3(G8), .ZN(new_n1084));
  OAI22_X1  g659(.A1(new_n1056), .A2(new_n1057), .B1(new_n1069), .B2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(KEYINPUT63), .ZN(new_n1086));
  INV_X1    g661(.A(G2084), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1074), .A2(new_n1087), .A3(new_n1077), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(KEYINPUT113), .ZN(new_n1089));
  AOI21_X1  g664(.A(KEYINPUT45), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n992), .B1(new_n990), .B2(new_n993), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n810), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT113), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1074), .A2(new_n1077), .A3(new_n1093), .A4(new_n1087), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1089), .A2(new_n1092), .A3(new_n1094), .ZN(new_n1095));
  NOR2_X1   g670(.A1(G286), .A2(new_n1042), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT114), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1095), .A2(KEYINPUT114), .A3(new_n1096), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1086), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT115), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1083), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1071), .B1(new_n1103), .B2(new_n1042), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1067), .ZN(new_n1105));
  AND4_X1   g680(.A1(new_n1102), .A2(new_n1054), .A3(new_n1104), .A4(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1102), .B1(new_n1068), .B2(new_n1104), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1101), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT63), .ZN(new_n1109));
  AND3_X1   g684(.A1(new_n1095), .A2(KEYINPUT114), .A3(new_n1096), .ZN(new_n1110));
  AOI21_X1  g685(.A(KEYINPUT114), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT112), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1113), .B1(new_n990), .B2(KEYINPUT50), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1043), .A2(KEYINPUT112), .A3(new_n1073), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  OAI21_X1  g691(.A(KEYINPUT50), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1116), .A2(new_n992), .A3(new_n1117), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1082), .B1(new_n1118), .B2(G2090), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(G8), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(new_n1071), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1068), .A2(new_n1121), .A3(new_n1084), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1109), .B1(new_n1112), .B2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1085), .B1(new_n1108), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT51), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1089), .A2(G168), .A3(new_n1092), .A4(new_n1094), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1126), .A2(G8), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1095), .A2(G286), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1125), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1127), .A2(KEYINPUT51), .ZN(new_n1131));
  OAI21_X1  g706(.A(KEYINPUT62), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1129), .ZN(new_n1133));
  OAI21_X1  g708(.A(KEYINPUT51), .B1(new_n1133), .B2(new_n1127), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1131), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT62), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1134), .A2(new_n1135), .A3(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT118), .ZN(new_n1138));
  NOR3_X1   g713(.A1(new_n1045), .A2(new_n1046), .A3(KEYINPUT50), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1138), .B1(new_n1139), .B2(new_n1076), .ZN(new_n1140));
  INV_X1    g715(.A(G1961), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1074), .A2(KEYINPUT118), .A3(new_n1077), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1140), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT53), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1145), .A2(G2078), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1144), .A2(new_n1146), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1145), .B1(new_n1081), .B2(G2078), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1143), .A2(new_n1147), .A3(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1149), .A2(G171), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1122), .A2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1132), .A2(new_n1137), .A3(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1124), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1079), .A2(new_n992), .ZN(new_n1155));
  OR2_X1    g730(.A1(new_n1155), .A2(KEYINPUT124), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1155), .A2(KEYINPUT124), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1156), .A2(new_n1080), .A3(new_n1146), .A4(new_n1157), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1143), .A2(new_n1158), .A3(new_n1148), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1150), .B1(G171), .B2(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT54), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(new_n1122), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1161), .B1(new_n1159), .B2(G171), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1164), .B1(G171), .B2(new_n1149), .ZN(new_n1165));
  NAND4_X1  g740(.A1(new_n1154), .A2(new_n1162), .A3(new_n1163), .A4(new_n1165), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n572), .A2(KEYINPUT116), .A3(new_n576), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT57), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  XNOR2_X1  g744(.A(new_n1169), .B(G299), .ZN(new_n1170));
  XNOR2_X1  g745(.A(KEYINPUT117), .B(KEYINPUT56), .ZN(new_n1171));
  XNOR2_X1  g746(.A(new_n1171), .B(G2072), .ZN(new_n1172));
  INV_X1    g747(.A(new_n1172), .ZN(new_n1173));
  NOR2_X1   g748(.A1(new_n1081), .A2(new_n1173), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1174), .B1(new_n1118), .B2(new_n800), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1170), .B1(new_n1175), .B2(KEYINPUT119), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT119), .ZN(new_n1177));
  AOI211_X1 g752(.A(new_n1177), .B(new_n1174), .C1(new_n800), .C2(new_n1118), .ZN(new_n1178));
  NOR2_X1   g753(.A1(new_n1176), .A2(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(new_n1170), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1175), .A2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1140), .A2(new_n804), .A3(new_n1142), .ZN(new_n1182));
  INV_X1    g757(.A(G2067), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1047), .A2(new_n1183), .A3(new_n992), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n624), .B1(new_n1182), .B2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g760(.A(new_n1179), .B1(new_n1181), .B2(new_n1185), .ZN(new_n1186));
  INV_X1    g761(.A(KEYINPUT61), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1187), .B1(new_n1175), .B2(new_n1180), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n1188), .B1(new_n1176), .B2(new_n1178), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT122), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  OAI211_X1 g766(.A(KEYINPUT122), .B(new_n1188), .C1(new_n1176), .C2(new_n1178), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  INV_X1    g768(.A(new_n1181), .ZN(new_n1194));
  NOR2_X1   g769(.A1(new_n1175), .A2(new_n1180), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n1187), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1182), .A2(new_n1184), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1197), .A2(new_n624), .ZN(new_n1198));
  NAND3_X1  g773(.A1(new_n1182), .A2(new_n616), .A3(new_n1184), .ZN(new_n1199));
  NAND3_X1  g774(.A1(new_n1198), .A2(KEYINPUT60), .A3(new_n1199), .ZN(new_n1200));
  OR2_X1    g775(.A1(new_n1199), .A2(KEYINPUT60), .ZN(new_n1201));
  XOR2_X1   g776(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n1202));
  OAI21_X1  g777(.A(KEYINPUT120), .B1(new_n1081), .B2(G1996), .ZN(new_n1203));
  NAND2_X1  g778(.A1(G160), .A2(G40), .ZN(new_n1204));
  AOI21_X1  g779(.A(new_n1204), .B1(new_n990), .B2(new_n993), .ZN(new_n1205));
  INV_X1    g780(.A(KEYINPUT120), .ZN(new_n1206));
  NAND4_X1  g781(.A1(new_n1205), .A2(new_n1206), .A3(new_n1003), .A4(new_n1080), .ZN(new_n1207));
  XOR2_X1   g782(.A(KEYINPUT58), .B(G1341), .Z(new_n1208));
  NAND2_X1  g783(.A1(new_n1060), .A2(new_n1208), .ZN(new_n1209));
  NAND3_X1  g784(.A1(new_n1203), .A2(new_n1207), .A3(new_n1209), .ZN(new_n1210));
  AOI21_X1  g785(.A(new_n1202), .B1(new_n1210), .B2(new_n562), .ZN(new_n1211));
  INV_X1    g786(.A(KEYINPUT59), .ZN(new_n1212));
  NOR2_X1   g787(.A1(new_n1212), .A2(KEYINPUT121), .ZN(new_n1213));
  AND2_X1   g788(.A1(new_n1210), .A2(new_n562), .ZN(new_n1214));
  AOI21_X1  g789(.A(new_n1211), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  NAND4_X1  g790(.A1(new_n1196), .A2(new_n1200), .A3(new_n1201), .A4(new_n1215), .ZN(new_n1216));
  OAI21_X1  g791(.A(new_n1186), .B1(new_n1193), .B2(new_n1216), .ZN(new_n1217));
  INV_X1    g792(.A(KEYINPUT123), .ZN(new_n1218));
  AOI21_X1  g793(.A(new_n1166), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  OAI211_X1 g794(.A(KEYINPUT123), .B(new_n1186), .C1(new_n1193), .C2(new_n1216), .ZN(new_n1220));
  AOI21_X1  g795(.A(new_n1153), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1221));
  XNOR2_X1  g796(.A(new_n729), .B(G1986), .ZN(new_n1222));
  OAI21_X1  g797(.A(new_n1019), .B1(new_n996), .B2(new_n1222), .ZN(new_n1223));
  OAI21_X1  g798(.A(new_n1027), .B1(new_n1221), .B2(new_n1223), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g799(.A1(new_n880), .A2(new_n881), .ZN(new_n1226));
  NOR2_X1   g800(.A1(G227), .A2(new_n457), .ZN(new_n1227));
  NAND2_X1  g801(.A1(new_n1227), .A2(new_n655), .ZN(new_n1228));
  AOI21_X1  g802(.A(new_n1228), .B1(new_n692), .B2(new_n693), .ZN(new_n1229));
  NAND3_X1  g803(.A1(new_n1226), .A2(new_n985), .A3(new_n1229), .ZN(G225));
  INV_X1    g804(.A(G225), .ZN(G308));
endmodule


