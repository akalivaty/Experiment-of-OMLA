//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 1 1 0 1 0 0 1 0 0 0 1 1 0 0 0 0 1 1 1 0 1 0 1 1 1 0 0 0 1 1 1 0 0 1 0 1 0 1 0 0 1 0 0 0 1 1 1 1 0 1 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:09 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n720, new_n721, new_n722, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n752, new_n753, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012;
  INV_X1    g000(.A(KEYINPUT73), .ZN(new_n187));
  INV_X1    g001(.A(G116), .ZN(new_n188));
  OAI21_X1  g002(.A(KEYINPUT66), .B1(new_n188), .B2(G119), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT66), .ZN(new_n190));
  INV_X1    g004(.A(G119), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n190), .A2(new_n191), .A3(G116), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n188), .A2(G119), .ZN(new_n193));
  AND3_X1   g007(.A1(new_n189), .A2(new_n192), .A3(new_n193), .ZN(new_n194));
  NOR2_X1   g008(.A1(KEYINPUT2), .A2(G113), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT65), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT2), .ZN(new_n197));
  INV_X1    g011(.A(G113), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n196), .B1(new_n197), .B2(new_n198), .ZN(new_n199));
  NAND3_X1  g013(.A1(KEYINPUT65), .A2(KEYINPUT2), .A3(G113), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n195), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n194), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(new_n200), .ZN(new_n203));
  AOI21_X1  g017(.A(KEYINPUT65), .B1(KEYINPUT2), .B2(G113), .ZN(new_n204));
  OAI22_X1  g018(.A1(new_n203), .A2(new_n204), .B1(KEYINPUT2), .B2(G113), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n189), .A2(new_n192), .A3(new_n193), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n202), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT70), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G146), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G143), .ZN(new_n212));
  INV_X1    g026(.A(G143), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G146), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n212), .A2(new_n214), .A3(KEYINPUT0), .A4(G128), .ZN(new_n215));
  XNOR2_X1  g029(.A(G143), .B(G146), .ZN(new_n216));
  XNOR2_X1  g030(.A(KEYINPUT0), .B(G128), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n215), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT11), .ZN(new_n220));
  INV_X1    g034(.A(G134), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n220), .B1(new_n221), .B2(G137), .ZN(new_n222));
  INV_X1    g036(.A(G137), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n223), .A2(KEYINPUT11), .A3(G134), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n221), .A2(G137), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n222), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(G131), .ZN(new_n227));
  INV_X1    g041(.A(G131), .ZN(new_n228));
  NAND4_X1  g042(.A1(new_n222), .A2(new_n224), .A3(new_n228), .A4(new_n225), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n219), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n202), .A2(new_n207), .A3(KEYINPUT70), .ZN(new_n232));
  AND3_X1   g046(.A1(new_n210), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n221), .A2(G137), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n223), .A2(G134), .ZN(new_n235));
  OAI21_X1  g049(.A(G131), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  AND3_X1   g050(.A1(new_n229), .A2(new_n236), .A3(KEYINPUT67), .ZN(new_n237));
  AOI21_X1  g051(.A(KEYINPUT67), .B1(new_n229), .B2(new_n236), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT1), .ZN(new_n240));
  AND4_X1   g054(.A1(new_n240), .A2(new_n212), .A3(new_n214), .A4(G128), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(G128), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n213), .A2(G146), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n211), .A2(G143), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n243), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(KEYINPUT1), .ZN(new_n247));
  AOI21_X1  g061(.A(KEYINPUT64), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  AOI21_X1  g062(.A(G128), .B1(new_n212), .B2(new_n214), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT64), .ZN(new_n250));
  NOR3_X1   g064(.A1(new_n240), .A2(new_n211), .A3(G143), .ZN(new_n251));
  NOR3_X1   g065(.A1(new_n249), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n242), .B1(new_n248), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n239), .A2(new_n253), .ZN(new_n254));
  AOI21_X1  g068(.A(KEYINPUT28), .B1(new_n233), .B2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  XOR2_X1   g070(.A(KEYINPUT71), .B(KEYINPUT27), .Z(new_n257));
  INV_X1    g071(.A(G237), .ZN(new_n258));
  INV_X1    g072(.A(G953), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n258), .A2(new_n259), .A3(G210), .ZN(new_n260));
  XNOR2_X1  g074(.A(new_n257), .B(new_n260), .ZN(new_n261));
  XNOR2_X1  g075(.A(KEYINPUT26), .B(G101), .ZN(new_n262));
  XOR2_X1   g076(.A(new_n261), .B(new_n262), .Z(new_n263));
  INV_X1    g077(.A(KEYINPUT29), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n229), .A2(new_n236), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT67), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n229), .A2(new_n236), .A3(KEYINPUT67), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n250), .B1(new_n249), .B2(new_n251), .ZN(new_n271));
  OAI211_X1 g085(.A(new_n247), .B(KEYINPUT64), .C1(new_n216), .C2(G128), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n241), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  OAI21_X1  g087(.A(KEYINPUT68), .B1(new_n270), .B2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT68), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n239), .A2(new_n253), .A3(new_n275), .ZN(new_n276));
  AND2_X1   g090(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n274), .A2(new_n276), .A3(new_n231), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n210), .A2(new_n232), .ZN(new_n279));
  AOI22_X1  g093(.A1(new_n277), .A2(new_n233), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT28), .ZN(new_n281));
  OAI211_X1 g095(.A(new_n256), .B(new_n265), .C1(new_n280), .C2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(G902), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n274), .A2(new_n276), .A3(KEYINPUT30), .A4(new_n231), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n231), .B1(new_n273), .B2(new_n266), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT30), .ZN(new_n287));
  AOI22_X1  g101(.A1(new_n286), .A2(new_n287), .B1(new_n207), .B2(new_n202), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n285), .A2(KEYINPUT69), .A3(new_n288), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n233), .A2(new_n274), .A3(new_n276), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(KEYINPUT69), .B1(new_n285), .B2(new_n288), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n263), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n286), .A2(new_n208), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT72), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n286), .A2(KEYINPUT72), .A3(new_n208), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n290), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n255), .B1(new_n298), .B2(KEYINPUT28), .ZN(new_n299));
  INV_X1    g113(.A(new_n263), .ZN(new_n300));
  AOI21_X1  g114(.A(KEYINPUT29), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n284), .B1(new_n293), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(G472), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n187), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n285), .A2(new_n288), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT69), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND4_X1  g121(.A1(new_n307), .A2(new_n290), .A3(new_n300), .A4(new_n289), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT31), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  AND2_X1   g124(.A1(new_n289), .A2(new_n290), .ZN(new_n311));
  NAND4_X1  g125(.A1(new_n311), .A2(KEYINPUT31), .A3(new_n300), .A4(new_n307), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n299), .A2(new_n300), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  NOR2_X1   g130(.A1(G472), .A2(G902), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n316), .A2(KEYINPUT32), .A3(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT32), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n314), .B1(new_n310), .B2(new_n312), .ZN(new_n320));
  INV_X1    g134(.A(new_n317), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n319), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n299), .A2(new_n300), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n323), .A2(new_n293), .A3(new_n264), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n278), .A2(new_n279), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(new_n290), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n255), .B1(new_n326), .B2(KEYINPUT28), .ZN(new_n327));
  AOI21_X1  g141(.A(G902), .B1(new_n327), .B2(new_n265), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n324), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n329), .A2(KEYINPUT73), .A3(G472), .ZN(new_n330));
  NAND4_X1  g144(.A1(new_n304), .A2(new_n318), .A3(new_n322), .A4(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(G217), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n332), .B1(G234), .B2(new_n283), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT25), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n243), .A2(G119), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n191), .A2(G128), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  XNOR2_X1  g152(.A(new_n338), .B(KEYINPUT74), .ZN(new_n339));
  XOR2_X1   g153(.A(KEYINPUT24), .B(G110), .Z(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  XNOR2_X1  g155(.A(new_n341), .B(KEYINPUT75), .ZN(new_n342));
  INV_X1    g156(.A(G140), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(G125), .ZN(new_n344));
  INV_X1    g158(.A(G125), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(G140), .ZN(new_n346));
  AND2_X1   g160(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(KEYINPUT16), .ZN(new_n348));
  OR2_X1    g162(.A1(new_n344), .A2(KEYINPUT16), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(new_n211), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n348), .A2(G146), .A3(new_n349), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n243), .A2(KEYINPUT23), .A3(G119), .ZN(new_n353));
  INV_X1    g167(.A(new_n336), .ZN(new_n354));
  OAI211_X1 g168(.A(new_n337), .B(new_n353), .C1(new_n354), .C2(KEYINPUT23), .ZN(new_n355));
  AOI22_X1  g169(.A1(new_n351), .A2(new_n352), .B1(G110), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n342), .A2(new_n356), .ZN(new_n357));
  OAI22_X1  g171(.A1(new_n339), .A2(new_n340), .B1(G110), .B2(new_n355), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n347), .A2(new_n211), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n358), .A2(new_n352), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n357), .A2(new_n360), .ZN(new_n361));
  XNOR2_X1  g175(.A(KEYINPUT22), .B(G137), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n259), .A2(G221), .A3(G234), .ZN(new_n363));
  XNOR2_X1  g177(.A(new_n362), .B(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n361), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n357), .A2(new_n360), .A3(new_n364), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n335), .B1(new_n368), .B2(G902), .ZN(new_n369));
  NAND4_X1  g183(.A1(new_n366), .A2(KEYINPUT25), .A3(new_n283), .A4(new_n367), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n334), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NOR3_X1   g185(.A1(new_n368), .A2(G902), .A3(new_n333), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  AND2_X1   g187(.A1(new_n331), .A2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT98), .ZN(new_n375));
  INV_X1    g189(.A(G104), .ZN(new_n376));
  OAI21_X1  g190(.A(KEYINPUT3), .B1(new_n376), .B2(G107), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT3), .ZN(new_n378));
  INV_X1    g192(.A(G107), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n378), .A2(new_n379), .A3(G104), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n376), .A2(G107), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n377), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(G101), .ZN(new_n383));
  INV_X1    g197(.A(G101), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n377), .A2(new_n380), .A3(new_n384), .A4(new_n381), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n383), .A2(KEYINPUT4), .A3(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT4), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n382), .A2(new_n387), .A3(G101), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n386), .A2(new_n219), .A3(new_n388), .ZN(new_n389));
  OAI21_X1  g203(.A(KEYINPUT77), .B1(new_n379), .B2(G104), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT77), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n391), .A2(new_n376), .A3(G107), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n379), .A2(G104), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n390), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(G101), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n395), .A2(KEYINPUT10), .A3(new_n385), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n389), .B1(new_n273), .B2(new_n396), .ZN(new_n397));
  XOR2_X1   g211(.A(KEYINPUT79), .B(KEYINPUT10), .Z(new_n398));
  OAI21_X1  g212(.A(KEYINPUT78), .B1(new_n249), .B2(new_n251), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT78), .ZN(new_n400));
  OAI211_X1 g214(.A(new_n247), .B(new_n400), .C1(new_n216), .C2(G128), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n399), .A2(new_n242), .A3(new_n401), .ZN(new_n402));
  AND2_X1   g216(.A1(new_n395), .A2(new_n385), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n398), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n230), .B1(new_n397), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n402), .A2(new_n403), .ZN(new_n406));
  INV_X1    g220(.A(new_n398), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n396), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n253), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n230), .A2(KEYINPUT80), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT80), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n227), .A2(new_n412), .A3(new_n229), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  NAND4_X1  g228(.A1(new_n408), .A2(new_n389), .A3(new_n410), .A4(new_n414), .ZN(new_n415));
  XNOR2_X1  g229(.A(G110), .B(G140), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n259), .A2(G227), .ZN(new_n417));
  XNOR2_X1  g231(.A(new_n416), .B(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n405), .A2(new_n415), .A3(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  XNOR2_X1  g234(.A(new_n418), .B(KEYINPUT76), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n271), .A2(new_n272), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n395), .A2(new_n385), .ZN(new_n424));
  AND3_X1   g238(.A1(new_n423), .A2(new_n242), .A3(new_n424), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n247), .B1(new_n216), .B2(G128), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n241), .B1(new_n426), .B2(KEYINPUT78), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n424), .B1(new_n427), .B2(new_n401), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n230), .B1(new_n425), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(KEYINPUT12), .ZN(new_n430));
  INV_X1    g244(.A(new_n230), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n423), .A2(new_n242), .A3(new_n424), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n431), .B1(new_n406), .B2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT12), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n430), .A2(new_n415), .A3(new_n435), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n422), .B1(new_n436), .B2(KEYINPUT81), .ZN(new_n437));
  XNOR2_X1  g251(.A(new_n433), .B(KEYINPUT12), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT81), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n438), .A2(new_n439), .A3(new_n415), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n420), .B1(new_n437), .B2(new_n440), .ZN(new_n441));
  OAI21_X1  g255(.A(G469), .B1(new_n441), .B2(G902), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT83), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n418), .B1(new_n405), .B2(new_n415), .ZN(new_n444));
  NAND4_X1  g258(.A1(new_n430), .A2(new_n415), .A3(new_n418), .A4(new_n435), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT82), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n444), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND4_X1  g261(.A1(new_n438), .A2(KEYINPUT82), .A3(new_n415), .A4(new_n418), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(G469), .ZN(new_n450));
  AND4_X1   g264(.A1(new_n443), .A2(new_n449), .A3(new_n450), .A4(new_n283), .ZN(new_n451));
  AOI21_X1  g265(.A(G902), .B1(new_n447), .B2(new_n448), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n443), .B1(new_n452), .B2(new_n450), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n442), .B1(new_n451), .B2(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(G214), .B1(G237), .B2(G902), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  OAI21_X1  g270(.A(G210), .B1(G237), .B2(G902), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n219), .A2(G125), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n459), .B1(new_n273), .B2(G125), .ZN(new_n460));
  INV_X1    g274(.A(G224), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n461), .A2(G953), .ZN(new_n462));
  XNOR2_X1  g276(.A(new_n460), .B(new_n462), .ZN(new_n463));
  NAND4_X1  g277(.A1(new_n189), .A2(new_n192), .A3(KEYINPUT5), .A4(new_n193), .ZN(new_n464));
  NOR3_X1   g278(.A1(new_n188), .A2(KEYINPUT5), .A3(G119), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n465), .A2(new_n198), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  NAND4_X1  g281(.A1(new_n202), .A2(new_n467), .A3(new_n385), .A4(new_n395), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(KEYINPUT84), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT84), .ZN(new_n470));
  AOI22_X1  g284(.A1(new_n194), .A2(new_n201), .B1(new_n464), .B2(new_n466), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n403), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n208), .A2(new_n388), .A3(new_n386), .ZN(new_n473));
  XNOR2_X1  g287(.A(G110), .B(G122), .ZN(new_n474));
  NAND4_X1  g288(.A1(new_n469), .A2(new_n472), .A3(new_n473), .A4(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT86), .ZN(new_n476));
  AND2_X1   g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n475), .A2(new_n476), .ZN(new_n478));
  OAI21_X1  g292(.A(KEYINPUT6), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n469), .A2(new_n472), .A3(new_n473), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n474), .B(KEYINPUT85), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n479), .A2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n482), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(KEYINPUT6), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n463), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT7), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n462), .A2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n460), .A2(new_n489), .ZN(new_n490));
  OAI211_X1 g304(.A(new_n459), .B(new_n488), .C1(new_n273), .C2(G125), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  OR2_X1    g306(.A1(new_n403), .A2(new_n471), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(new_n468), .ZN(new_n494));
  XNOR2_X1  g308(.A(new_n474), .B(KEYINPUT8), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n492), .A2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT87), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n492), .A2(new_n496), .A3(KEYINPUT87), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  OR2_X1    g315(.A1(new_n475), .A2(new_n476), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n475), .A2(new_n476), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n283), .B1(new_n501), .B2(new_n505), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n458), .B1(new_n486), .B2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT6), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n508), .B1(new_n502), .B2(new_n503), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n485), .B1(new_n509), .B2(new_n484), .ZN(new_n510));
  INV_X1    g324(.A(new_n463), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AND3_X1   g326(.A1(new_n492), .A2(new_n496), .A3(KEYINPUT87), .ZN(new_n513));
  AOI21_X1  g327(.A(KEYINPUT87), .B1(new_n492), .B2(new_n496), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g329(.A(G902), .B1(new_n515), .B2(new_n504), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n512), .A2(new_n457), .A3(new_n516), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n456), .B1(new_n507), .B2(new_n517), .ZN(new_n518));
  XNOR2_X1  g332(.A(KEYINPUT9), .B(G234), .ZN(new_n519));
  OAI21_X1  g333(.A(G221), .B1(new_n519), .B2(G902), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n454), .A2(new_n518), .A3(new_n520), .ZN(new_n521));
  XNOR2_X1  g335(.A(KEYINPUT88), .B(G143), .ZN(new_n522));
  AND3_X1   g336(.A1(new_n258), .A2(new_n259), .A3(G214), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n258), .A2(new_n259), .A3(G214), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n525), .B1(KEYINPUT88), .B2(new_n213), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT18), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n527), .B1(new_n528), .B2(new_n228), .ZN(new_n529));
  XNOR2_X1  g343(.A(new_n529), .B(KEYINPUT90), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT89), .ZN(new_n531));
  XNOR2_X1  g345(.A(new_n347), .B(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(G146), .ZN(new_n533));
  OAI21_X1  g347(.A(G131), .B1(new_n524), .B2(new_n526), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  AOI22_X1  g349(.A1(new_n533), .A2(new_n359), .B1(new_n535), .B2(KEYINPUT18), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n530), .A2(new_n536), .ZN(new_n537));
  XNOR2_X1  g351(.A(G113), .B(G122), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n538), .B(new_n376), .ZN(new_n539));
  AND2_X1   g353(.A1(new_n351), .A2(new_n352), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n535), .A2(KEYINPUT17), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n527), .A2(new_n228), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(new_n534), .ZN(new_n543));
  OAI211_X1 g357(.A(new_n540), .B(new_n541), .C1(KEYINPUT17), .C2(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n537), .A2(new_n539), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n532), .A2(KEYINPUT19), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(KEYINPUT91), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT91), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n532), .A2(new_n548), .A3(KEYINPUT19), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT19), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n347), .A2(new_n550), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n547), .A2(new_n211), .A3(new_n549), .A4(new_n551), .ZN(new_n552));
  AND2_X1   g366(.A1(new_n543), .A2(new_n352), .ZN(new_n553));
  AOI22_X1  g367(.A1(new_n552), .A2(new_n553), .B1(new_n530), .B2(new_n536), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n545), .B1(new_n554), .B2(new_n539), .ZN(new_n555));
  NOR2_X1   g369(.A1(G475), .A2(G902), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(KEYINPUT20), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT20), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n555), .A2(new_n559), .A3(new_n556), .ZN(new_n560));
  INV_X1    g374(.A(new_n545), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n539), .B1(new_n537), .B2(new_n544), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n283), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  AOI22_X1  g377(.A1(new_n558), .A2(new_n560), .B1(G475), .B2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(G122), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(G116), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n188), .A2(G122), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n566), .A2(new_n567), .A3(new_n379), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n566), .A2(new_n567), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n569), .A2(KEYINPUT14), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT14), .ZN(new_n571));
  OAI21_X1  g385(.A(G107), .B1(new_n567), .B2(new_n571), .ZN(new_n572));
  OAI21_X1  g386(.A(KEYINPUT92), .B1(new_n243), .B2(G143), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT92), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n574), .A2(new_n213), .A3(G128), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n576), .B1(G128), .B2(new_n213), .ZN(new_n577));
  AND2_X1   g391(.A1(new_n577), .A2(G134), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n577), .A2(G134), .ZN(new_n579));
  OAI221_X1 g393(.A(new_n568), .B1(new_n570), .B2(new_n572), .C1(new_n578), .C2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n569), .A2(G107), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(new_n568), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n582), .B1(new_n577), .B2(G134), .ZN(new_n583));
  AND2_X1   g397(.A1(new_n573), .A2(new_n575), .ZN(new_n584));
  OAI21_X1  g398(.A(KEYINPUT93), .B1(new_n584), .B2(KEYINPUT13), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n584), .A2(KEYINPUT94), .A3(KEYINPUT13), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n213), .A2(G128), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n573), .A2(new_n575), .A3(KEYINPUT13), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT94), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n587), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT93), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT13), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n576), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n585), .A2(new_n586), .A3(new_n590), .A4(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n583), .B1(new_n594), .B2(G134), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT95), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  AOI211_X1 g411(.A(KEYINPUT95), .B(new_n583), .C1(new_n594), .C2(G134), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n580), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NOR3_X1   g413(.A1(new_n519), .A2(new_n332), .A3(G953), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  OAI211_X1 g416(.A(new_n580), .B(new_n600), .C1(new_n597), .C2(new_n598), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(new_n283), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT96), .ZN(new_n606));
  INV_X1    g420(.A(G478), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n607), .A2(KEYINPUT15), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n605), .A2(new_n606), .A3(new_n608), .ZN(new_n609));
  AOI21_X1  g423(.A(G902), .B1(new_n602), .B2(new_n603), .ZN(new_n610));
  INV_X1    g424(.A(new_n608), .ZN(new_n611));
  OAI21_X1  g425(.A(KEYINPUT96), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n609), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n604), .A2(new_n283), .A3(new_n611), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT97), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n610), .A2(KEYINPUT97), .A3(new_n611), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(G952), .ZN(new_n619));
  AOI211_X1 g433(.A(G953), .B(new_n619), .C1(G234), .C2(G237), .ZN(new_n620));
  AOI211_X1 g434(.A(new_n283), .B(new_n259), .C1(G234), .C2(G237), .ZN(new_n621));
  XNOR2_X1  g435(.A(KEYINPUT21), .B(G898), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n620), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n564), .A2(new_n613), .A3(new_n618), .A4(new_n624), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n375), .B1(new_n521), .B2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n520), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n449), .A2(new_n450), .A3(new_n283), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(KEYINPUT83), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n452), .A2(new_n443), .A3(new_n450), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n627), .B1(new_n631), .B2(new_n442), .ZN(new_n632));
  INV_X1    g446(.A(new_n625), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n632), .A2(new_n633), .A3(KEYINPUT98), .A4(new_n518), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n374), .A2(new_n626), .A3(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(G101), .ZN(G3));
  NAND2_X1  g450(.A1(new_n437), .A2(new_n440), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(new_n419), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n450), .B1(new_n638), .B2(new_n283), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n639), .B1(new_n630), .B2(new_n629), .ZN(new_n640));
  INV_X1    g454(.A(new_n373), .ZN(new_n641));
  NOR3_X1   g455(.A1(new_n640), .A2(new_n641), .A3(new_n627), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n605), .A2(new_n607), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n604), .A2(KEYINPUT33), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT99), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n599), .A2(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT100), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n601), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n603), .A2(new_n647), .ZN(new_n650));
  OAI211_X1 g464(.A(new_n599), .B(new_n645), .C1(new_n647), .C2(new_n601), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n649), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n644), .B1(KEYINPUT33), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n283), .A2(G478), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n643), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n558), .A2(new_n560), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n563), .A2(G475), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n507), .A2(new_n517), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n660), .A2(new_n624), .A3(new_n455), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  OAI21_X1  g476(.A(G472), .B1(new_n320), .B2(G902), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n316), .A2(new_n317), .ZN(new_n664));
  AND2_X1   g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n642), .A2(new_n662), .A3(new_n665), .ZN(new_n666));
  XOR2_X1   g480(.A(KEYINPUT34), .B(G104), .Z(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G6));
  INV_X1    g482(.A(new_n612), .ZN(new_n669));
  NOR3_X1   g483(.A1(new_n610), .A2(KEYINPUT96), .A3(new_n611), .ZN(new_n670));
  AND3_X1   g484(.A1(new_n610), .A2(KEYINPUT97), .A3(new_n611), .ZN(new_n671));
  AOI21_X1  g485(.A(KEYINPUT97), .B1(new_n610), .B2(new_n611), .ZN(new_n672));
  OAI22_X1  g486(.A1(new_n669), .A2(new_n670), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(new_n564), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n661), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n642), .A2(new_n675), .A3(new_n665), .ZN(new_n676));
  XOR2_X1   g490(.A(KEYINPUT35), .B(G107), .Z(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G9));
  NOR2_X1   g492(.A1(new_n365), .A2(KEYINPUT36), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(KEYINPUT101), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n361), .B(new_n680), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n333), .A2(G902), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  OR2_X1    g498(.A1(new_n371), .A2(new_n684), .ZN(new_n685));
  AND3_X1   g499(.A1(new_n685), .A2(new_n664), .A3(new_n663), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n626), .A2(new_n634), .A3(new_n686), .ZN(new_n687));
  XOR2_X1   g501(.A(KEYINPUT37), .B(G110), .Z(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(G12));
  INV_X1    g503(.A(new_n521), .ZN(new_n690));
  INV_X1    g504(.A(G900), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n621), .A2(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(new_n620), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n674), .A2(new_n695), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n690), .A2(new_n331), .A3(new_n696), .A4(new_n685), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G128), .ZN(G30));
  XNOR2_X1  g512(.A(KEYINPUT103), .B(KEYINPUT39), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n694), .B(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n632), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(KEYINPUT40), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT40), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n632), .A2(new_n704), .A3(new_n701), .ZN(new_n705));
  AND3_X1   g519(.A1(new_n507), .A2(new_n517), .A3(KEYINPUT38), .ZN(new_n706));
  AOI21_X1  g520(.A(KEYINPUT38), .B1(new_n507), .B2(new_n517), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n673), .A2(new_n658), .ZN(new_n709));
  NOR3_X1   g523(.A1(new_n709), .A2(new_n456), .A3(new_n685), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n703), .A2(new_n705), .A3(new_n708), .A4(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n311), .A2(new_n307), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(new_n300), .ZN(new_n713));
  OAI211_X1 g527(.A(new_n713), .B(new_n283), .C1(new_n300), .C2(new_n326), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(G472), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n318), .A2(new_n322), .A3(new_n715), .ZN(new_n716));
  XOR2_X1   g530(.A(new_n716), .B(KEYINPUT102), .Z(new_n717));
  NOR2_X1   g531(.A1(new_n711), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(new_n213), .ZN(G45));
  NAND3_X1  g533(.A1(new_n655), .A2(new_n658), .A3(new_n694), .ZN(new_n720));
  INV_X1    g534(.A(new_n720), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n690), .A2(new_n331), .A3(new_n685), .A4(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G146), .ZN(G48));
  OR2_X1    g537(.A1(new_n452), .A2(new_n450), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n631), .A2(new_n520), .A3(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(new_n725), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n662), .A2(new_n331), .A3(new_n373), .A4(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(KEYINPUT41), .B(G113), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n727), .B(new_n728), .ZN(G15));
  NAND4_X1  g543(.A1(new_n675), .A2(new_n331), .A3(new_n373), .A4(new_n726), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G116), .ZN(G18));
  NAND2_X1  g545(.A1(new_n660), .A2(new_n455), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n725), .A2(new_n732), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n371), .A2(new_n684), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n625), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n733), .A2(new_n331), .A3(new_n735), .ZN(new_n736));
  XOR2_X1   g550(.A(KEYINPUT104), .B(G119), .Z(new_n737));
  XNOR2_X1  g551(.A(new_n736), .B(new_n737), .ZN(G21));
  NOR2_X1   g552(.A1(new_n725), .A2(new_n623), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n256), .B1(new_n280), .B2(new_n281), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT105), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n327), .A2(KEYINPUT105), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n742), .A2(new_n743), .A3(new_n263), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(new_n313), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n745), .A2(new_n317), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(new_n663), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n747), .A2(new_n641), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n709), .A2(new_n732), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n739), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G122), .ZN(G24));
  NOR2_X1   g565(.A1(new_n747), .A2(new_n734), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n733), .A2(new_n752), .A3(new_n721), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G125), .ZN(G27));
  NAND3_X1  g568(.A1(new_n507), .A2(new_n517), .A3(new_n455), .ZN(new_n755));
  NOR3_X1   g569(.A1(new_n640), .A2(new_n627), .A3(new_n755), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n756), .A2(new_n331), .A3(new_n721), .A4(new_n373), .ZN(new_n757));
  XOR2_X1   g571(.A(KEYINPUT106), .B(KEYINPUT42), .Z(new_n758));
  INV_X1    g572(.A(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  AOI21_X1  g574(.A(KEYINPUT73), .B1(new_n329), .B2(G472), .ZN(new_n761));
  AOI211_X1 g575(.A(new_n187), .B(new_n303), .C1(new_n324), .C2(new_n328), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT107), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n318), .A2(new_n764), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n316), .A2(KEYINPUT107), .A3(KEYINPUT32), .A4(new_n317), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n763), .A2(new_n765), .A3(new_n322), .A4(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT42), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n720), .A2(new_n768), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n767), .A2(new_n769), .A3(new_n373), .A4(new_n756), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n760), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G131), .ZN(G33));
  NAND4_X1  g586(.A1(new_n374), .A2(KEYINPUT108), .A3(new_n696), .A4(new_n756), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n756), .A2(new_n696), .A3(new_n331), .A4(new_n373), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT108), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n773), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G134), .ZN(G36));
  NOR2_X1   g592(.A1(new_n665), .A2(new_n734), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n655), .A2(new_n564), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(KEYINPUT43), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT43), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n655), .A2(new_n782), .A3(new_n564), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n779), .A2(new_n781), .A3(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT44), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  AND2_X1   g600(.A1(new_n781), .A2(new_n783), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n787), .A2(KEYINPUT44), .A3(new_n779), .ZN(new_n788));
  INV_X1    g602(.A(new_n755), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n786), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT110), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n786), .A2(new_n788), .A3(KEYINPUT110), .A4(new_n789), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n450), .A2(new_n283), .ZN(new_n794));
  INV_X1    g608(.A(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT45), .ZN(new_n796));
  OAI21_X1  g610(.A(KEYINPUT109), .B1(new_n638), .B2(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT109), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n441), .A2(new_n798), .A3(KEYINPUT45), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  OAI21_X1  g614(.A(G469), .B1(new_n441), .B2(KEYINPUT45), .ZN(new_n801));
  OAI211_X1 g615(.A(KEYINPUT46), .B(new_n795), .C1(new_n800), .C2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT46), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n801), .B1(new_n797), .B2(new_n799), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n803), .B1(new_n804), .B2(new_n794), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n802), .A2(new_n805), .A3(new_n631), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n806), .A2(new_n520), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n807), .A2(new_n700), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n792), .A2(new_n793), .A3(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(G137), .ZN(G39));
  INV_X1    g624(.A(KEYINPUT47), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n807), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n806), .A2(KEYINPUT47), .A3(new_n520), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT111), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n721), .A2(new_n641), .A3(new_n789), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n815), .B1(new_n816), .B2(new_n331), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n720), .A2(new_n373), .A3(new_n755), .ZN(new_n818));
  INV_X1    g632(.A(new_n331), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n818), .A2(KEYINPUT111), .A3(new_n819), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n817), .A2(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT112), .ZN(new_n822));
  AND3_X1   g636(.A1(new_n814), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n822), .B1(new_n814), .B2(new_n821), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  XNOR2_X1  g639(.A(new_n825), .B(new_n343), .ZN(G42));
  NAND3_X1  g640(.A1(new_n373), .A2(new_n520), .A3(new_n455), .ZN(new_n827));
  NOR3_X1   g641(.A1(new_n708), .A2(new_n780), .A3(new_n827), .ZN(new_n828));
  AND2_X1   g642(.A1(new_n631), .A2(new_n724), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n829), .B(KEYINPUT49), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n717), .A2(new_n828), .A3(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT54), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n635), .A2(new_n666), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT113), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n635), .A2(KEYINPUT113), .A3(new_n666), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT114), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n837), .B1(new_n661), .B2(new_n674), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n658), .B1(new_n613), .B2(new_n618), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n839), .A2(KEYINPUT114), .A3(new_n624), .A4(new_n518), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n838), .A2(new_n840), .A3(new_n642), .A4(new_n665), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n687), .A2(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n835), .A2(new_n836), .A3(new_n843), .ZN(new_n844));
  AND4_X1   g658(.A1(new_n727), .A2(new_n730), .A3(new_n736), .A4(new_n750), .ZN(new_n845));
  INV_X1    g659(.A(new_n673), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n331), .A2(new_n564), .A3(new_n846), .ZN(new_n847));
  OR2_X1    g661(.A1(new_n659), .A2(new_n747), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n849), .A2(new_n685), .A3(new_n694), .A4(new_n756), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n845), .A2(new_n777), .A3(new_n771), .A4(new_n850), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n844), .A2(new_n851), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n685), .A2(new_n695), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n749), .A2(new_n632), .A3(new_n716), .A4(new_n853), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n697), .A2(new_n722), .A3(new_n753), .A4(new_n854), .ZN(new_n855));
  XOR2_X1   g669(.A(new_n855), .B(KEYINPUT52), .Z(new_n856));
  AOI21_X1  g670(.A(KEYINPUT53), .B1(new_n852), .B2(new_n856), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n842), .B1(new_n833), .B2(new_n834), .ZN(new_n858));
  AOI22_X1  g672(.A1(new_n776), .A2(new_n773), .B1(new_n760), .B2(new_n770), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n727), .A2(new_n730), .A3(new_n736), .A4(new_n750), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n756), .A2(new_n685), .A3(new_n694), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n861), .B1(new_n847), .B2(new_n848), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n858), .A2(new_n836), .A3(new_n859), .A4(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT53), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n855), .B(KEYINPUT52), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n832), .B1(new_n857), .B2(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n852), .A2(KEYINPUT53), .A3(new_n856), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n865), .B1(new_n864), .B2(new_n866), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n869), .A2(new_n870), .A3(KEYINPUT54), .ZN(new_n871));
  AND2_X1   g685(.A1(new_n868), .A2(new_n871), .ZN(new_n872));
  AND3_X1   g686(.A1(new_n787), .A2(new_n620), .A3(new_n748), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n708), .A2(new_n455), .A3(new_n725), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT50), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n875), .B(new_n876), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n725), .A2(new_n755), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n717), .A2(new_n373), .A3(new_n620), .A4(new_n878), .ZN(new_n879));
  OR3_X1    g693(.A1(new_n879), .A2(new_n658), .A3(new_n655), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n787), .A2(new_n620), .A3(new_n878), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(new_n752), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n877), .A2(new_n880), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n829), .A2(new_n627), .ZN(new_n884));
  INV_X1    g698(.A(new_n884), .ZN(new_n885));
  OAI211_X1 g699(.A(new_n789), .B(new_n873), .C1(new_n814), .C2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(new_n886), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n883), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n888), .A2(KEYINPUT51), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n873), .A2(new_n733), .ZN(new_n890));
  AOI211_X1 g704(.A(new_n619), .B(G953), .C1(new_n890), .C2(KEYINPUT115), .ZN(new_n891));
  OAI221_X1 g705(.A(new_n891), .B1(KEYINPUT115), .B2(new_n890), .C1(new_n659), .C2(new_n879), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n881), .A2(new_n373), .A3(new_n767), .ZN(new_n893));
  XOR2_X1   g707(.A(new_n893), .B(KEYINPUT48), .Z(new_n894));
  OR2_X1    g708(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT51), .ZN(new_n896));
  NOR3_X1   g710(.A1(new_n883), .A2(new_n896), .A3(new_n887), .ZN(new_n897));
  NOR4_X1   g711(.A1(new_n872), .A2(new_n889), .A3(new_n895), .A4(new_n897), .ZN(new_n898));
  NOR2_X1   g712(.A1(G952), .A2(G953), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n831), .B1(new_n898), .B2(new_n899), .ZN(G75));
  INV_X1    g714(.A(KEYINPUT117), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n283), .B1(new_n869), .B2(new_n870), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(G210), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT56), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n510), .A2(new_n511), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n905), .A2(new_n486), .ZN(new_n906));
  XOR2_X1   g720(.A(new_n906), .B(KEYINPUT55), .Z(new_n907));
  INV_X1    g721(.A(KEYINPUT116), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n907), .B1(new_n908), .B2(new_n904), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n903), .A2(new_n904), .A3(new_n909), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n259), .A2(G952), .ZN(new_n911));
  INV_X1    g725(.A(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n909), .B1(new_n903), .B2(new_n904), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n901), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n903), .A2(new_n904), .ZN(new_n916));
  INV_X1    g730(.A(new_n909), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n918), .A2(KEYINPUT117), .A3(new_n910), .A4(new_n912), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n915), .A2(new_n919), .ZN(G51));
  XNOR2_X1  g734(.A(KEYINPUT118), .B(KEYINPUT57), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(new_n794), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n872), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(new_n449), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n902), .A2(new_n804), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n911), .B1(new_n924), .B2(new_n925), .ZN(G54));
  AND2_X1   g740(.A1(KEYINPUT58), .A2(G475), .ZN(new_n927));
  AND3_X1   g741(.A1(new_n902), .A2(new_n555), .A3(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n555), .B1(new_n902), .B2(new_n927), .ZN(new_n929));
  NOR3_X1   g743(.A1(new_n928), .A2(new_n929), .A3(new_n911), .ZN(G60));
  NAND2_X1  g744(.A1(G478), .A2(G902), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(KEYINPUT59), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n868), .A2(new_n871), .A3(new_n932), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n653), .B(KEYINPUT119), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(new_n934), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n868), .A2(new_n871), .A3(new_n932), .A4(new_n936), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n935), .A2(new_n912), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(KEYINPUT120), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT120), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n935), .A2(new_n940), .A3(new_n912), .A4(new_n937), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n939), .A2(new_n941), .ZN(G63));
  NAND2_X1  g756(.A1(G217), .A2(G902), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(KEYINPUT60), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n944), .B1(new_n869), .B2(new_n870), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(new_n681), .ZN(new_n946));
  INV_X1    g760(.A(new_n368), .ZN(new_n947));
  OAI211_X1 g761(.A(new_n946), .B(new_n912), .C1(new_n947), .C2(new_n945), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT61), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n948), .B(new_n949), .ZN(G66));
  OAI21_X1  g764(.A(new_n259), .B1(new_n844), .B2(new_n860), .ZN(new_n951));
  OAI21_X1  g765(.A(G953), .B1(new_n622), .B2(new_n461), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n951), .A2(KEYINPUT121), .A3(new_n952), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n953), .B1(KEYINPUT121), .B2(new_n951), .ZN(new_n954));
  OAI211_X1 g768(.A(new_n483), .B(new_n485), .C1(G898), .C2(new_n259), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n955), .B(KEYINPUT122), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n954), .B(new_n956), .ZN(G69));
  AND4_X1   g771(.A1(new_n373), .A2(new_n808), .A3(new_n749), .A4(new_n767), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n825), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n697), .A2(new_n722), .A3(new_n753), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n960), .A2(KEYINPUT124), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT124), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n697), .A2(new_n722), .A3(new_n753), .A4(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  AND2_X1   g778(.A1(new_n964), .A2(new_n859), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n959), .A2(new_n259), .A3(new_n809), .A4(new_n965), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n547), .A2(new_n549), .A3(new_n551), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n967), .B(KEYINPUT123), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n286), .A2(new_n287), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n285), .A2(new_n969), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n968), .B(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(G900), .A2(G953), .ZN(new_n972));
  AND2_X1   g786(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n966), .A2(new_n973), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n718), .B1(new_n961), .B2(new_n963), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT62), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n975), .B(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(new_n702), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n755), .B1(new_n659), .B2(new_n674), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n374), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  OAI211_X1 g794(.A(new_n809), .B(new_n980), .C1(new_n823), .C2(new_n824), .ZN(new_n981));
  OAI21_X1  g795(.A(KEYINPUT125), .B1(new_n977), .B2(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(new_n718), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n964), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n984), .A2(new_n976), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n964), .A2(KEYINPUT62), .A3(new_n983), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g801(.A(new_n980), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n814), .A2(new_n821), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n989), .A2(KEYINPUT112), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n814), .A2(new_n821), .A3(new_n822), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n988), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  INV_X1    g806(.A(KEYINPUT125), .ZN(new_n993));
  NAND4_X1  g807(.A1(new_n987), .A2(new_n992), .A3(new_n993), .A4(new_n809), .ZN(new_n994));
  AOI21_X1  g808(.A(G953), .B1(new_n982), .B2(new_n994), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n974), .B1(new_n995), .B2(new_n971), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n259), .B1(G227), .B2(G900), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n997), .B1(new_n974), .B2(KEYINPUT126), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  OAI221_X1 g813(.A(new_n974), .B1(KEYINPUT126), .B2(new_n997), .C1(new_n995), .C2(new_n971), .ZN(new_n1000));
  AND2_X1   g814(.A1(new_n999), .A2(new_n1000), .ZN(G72));
  NOR2_X1   g815(.A1(new_n844), .A2(new_n860), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n982), .A2(new_n994), .A3(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g817(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n1004));
  NOR2_X1   g818(.A1(new_n303), .A2(new_n283), .ZN(new_n1005));
  XOR2_X1   g819(.A(new_n1004), .B(new_n1005), .Z(new_n1006));
  AOI21_X1  g820(.A(new_n713), .B1(new_n1003), .B2(new_n1006), .ZN(new_n1007));
  NAND4_X1  g821(.A1(new_n959), .A2(new_n809), .A3(new_n1002), .A4(new_n965), .ZN(new_n1008));
  AOI211_X1 g822(.A(new_n300), .B(new_n712), .C1(new_n1008), .C2(new_n1006), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n293), .A2(new_n308), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1010), .A2(new_n1006), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n1011), .B1(new_n869), .B2(new_n870), .ZN(new_n1012));
  NOR4_X1   g826(.A1(new_n1007), .A2(new_n1009), .A3(new_n911), .A4(new_n1012), .ZN(G57));
endmodule


