

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585;

  XNOR2_X1 U321 ( .A(n332), .B(n331), .ZN(n333) );
  NOR2_X1 U322 ( .A1(n533), .A2(n416), .ZN(n418) );
  XNOR2_X1 U323 ( .A(n479), .B(n478), .ZN(n520) );
  XNOR2_X1 U324 ( .A(KEYINPUT108), .B(KEYINPUT37), .ZN(n478) );
  AND2_X1 U325 ( .A1(G232GAT), .A2(G233GAT), .ZN(n289) );
  XOR2_X1 U326 ( .A(G64GAT), .B(G92GAT), .Z(n290) );
  XNOR2_X1 U327 ( .A(n388), .B(KEYINPUT45), .ZN(n389) );
  NOR2_X1 U328 ( .A1(n570), .A2(n390), .ZN(n391) );
  XNOR2_X1 U329 ( .A(n334), .B(n333), .ZN(n336) );
  INV_X1 U330 ( .A(KEYINPUT54), .ZN(n417) );
  XNOR2_X1 U331 ( .A(n405), .B(n289), .ZN(n352) );
  INV_X1 U332 ( .A(KEYINPUT99), .ZN(n410) );
  NOR2_X1 U333 ( .A1(n475), .A2(n474), .ZN(n486) );
  XNOR2_X1 U334 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U335 ( .A(n353), .B(n352), .ZN(n360) );
  XNOR2_X1 U336 ( .A(n411), .B(n410), .ZN(n412) );
  NOR2_X1 U337 ( .A1(n521), .A2(n419), .ZN(n568) );
  XNOR2_X1 U338 ( .A(n345), .B(n344), .ZN(n573) );
  XNOR2_X1 U339 ( .A(n350), .B(KEYINPUT64), .ZN(n554) );
  XNOR2_X1 U340 ( .A(n413), .B(n412), .ZN(n414) );
  XOR2_X1 U341 ( .A(KEYINPUT120), .B(n457), .Z(n563) );
  XNOR2_X1 U342 ( .A(n480), .B(KEYINPUT38), .ZN(n505) );
  XNOR2_X1 U343 ( .A(G183GAT), .B(KEYINPUT122), .ZN(n458) );
  XNOR2_X1 U344 ( .A(n481), .B(KEYINPUT106), .ZN(n482) );
  XNOR2_X1 U345 ( .A(n459), .B(n458), .ZN(G1350GAT) );
  XNOR2_X1 U346 ( .A(n483), .B(n482), .ZN(G1328GAT) );
  XOR2_X1 U347 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n292) );
  XNOR2_X1 U348 ( .A(G155GAT), .B(KEYINPUT97), .ZN(n291) );
  XNOR2_X1 U349 ( .A(n292), .B(n291), .ZN(n299) );
  XOR2_X1 U350 ( .A(G85GAT), .B(G162GAT), .Z(n294) );
  XNOR2_X1 U351 ( .A(G127GAT), .B(G148GAT), .ZN(n293) );
  XNOR2_X1 U352 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U353 ( .A(n295), .B(G120GAT), .Z(n297) );
  XOR2_X1 U354 ( .A(G113GAT), .B(G1GAT), .Z(n318) );
  XNOR2_X1 U355 ( .A(G29GAT), .B(n318), .ZN(n296) );
  XNOR2_X1 U356 ( .A(n297), .B(n296), .ZN(n298) );
  XNOR2_X1 U357 ( .A(n299), .B(n298), .ZN(n308) );
  XOR2_X1 U358 ( .A(KEYINPUT1), .B(G57GAT), .Z(n301) );
  NAND2_X1 U359 ( .A1(G225GAT), .A2(G233GAT), .ZN(n300) );
  XNOR2_X1 U360 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U361 ( .A(n302), .B(KEYINPUT6), .Z(n306) );
  XNOR2_X1 U362 ( .A(G134GAT), .B(KEYINPUT85), .ZN(n303) );
  XNOR2_X1 U363 ( .A(n303), .B(KEYINPUT0), .ZN(n444) );
  XNOR2_X1 U364 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n304) );
  XNOR2_X1 U365 ( .A(n304), .B(KEYINPUT2), .ZN(n423) );
  XNOR2_X1 U366 ( .A(n444), .B(n423), .ZN(n305) );
  XNOR2_X1 U367 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U368 ( .A(n308), .B(n307), .ZN(n521) );
  XOR2_X1 U369 ( .A(G8GAT), .B(G141GAT), .Z(n310) );
  XNOR2_X1 U370 ( .A(G197GAT), .B(G22GAT), .ZN(n309) );
  XNOR2_X1 U371 ( .A(n310), .B(n309), .ZN(n314) );
  XOR2_X1 U372 ( .A(KEYINPUT29), .B(KEYINPUT67), .Z(n312) );
  XNOR2_X1 U373 ( .A(KEYINPUT30), .B(KEYINPUT66), .ZN(n311) );
  XNOR2_X1 U374 ( .A(n312), .B(n311), .ZN(n313) );
  XNOR2_X1 U375 ( .A(n314), .B(n313), .ZN(n327) );
  XOR2_X1 U376 ( .A(G15GAT), .B(G50GAT), .Z(n316) );
  XNOR2_X1 U377 ( .A(G169GAT), .B(G36GAT), .ZN(n315) );
  XNOR2_X1 U378 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U379 ( .A(n318), .B(n317), .Z(n320) );
  NAND2_X1 U380 ( .A1(G229GAT), .A2(G233GAT), .ZN(n319) );
  XNOR2_X1 U381 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U382 ( .A(n321), .B(KEYINPUT68), .Z(n325) );
  XOR2_X1 U383 ( .A(G29GAT), .B(G43GAT), .Z(n323) );
  XNOR2_X1 U384 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n322) );
  XNOR2_X1 U385 ( .A(n323), .B(n322), .ZN(n353) );
  XNOR2_X1 U386 ( .A(n353), .B(KEYINPUT69), .ZN(n324) );
  XNOR2_X1 U387 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U388 ( .A(n327), .B(n326), .ZN(n570) );
  XNOR2_X1 U389 ( .A(G99GAT), .B(G85GAT), .ZN(n328) );
  XNOR2_X1 U390 ( .A(n328), .B(KEYINPUT74), .ZN(n361) );
  XNOR2_X1 U391 ( .A(n361), .B(KEYINPUT77), .ZN(n334) );
  XOR2_X1 U392 ( .A(KEYINPUT72), .B(KEYINPUT31), .Z(n330) );
  XNOR2_X1 U393 ( .A(KEYINPUT76), .B(KEYINPUT71), .ZN(n329) );
  XNOR2_X1 U394 ( .A(n330), .B(n329), .ZN(n332) );
  AND2_X1 U395 ( .A1(G230GAT), .A2(G233GAT), .ZN(n331) );
  XOR2_X1 U396 ( .A(G120GAT), .B(G71GAT), .Z(n445) );
  XOR2_X1 U397 ( .A(G57GAT), .B(KEYINPUT13), .Z(n371) );
  XOR2_X1 U398 ( .A(n445), .B(n371), .Z(n335) );
  XNOR2_X1 U399 ( .A(n336), .B(n335), .ZN(n340) );
  XOR2_X1 U400 ( .A(KEYINPUT33), .B(KEYINPUT75), .Z(n338) );
  XNOR2_X1 U401 ( .A(KEYINPUT32), .B(KEYINPUT70), .ZN(n337) );
  XNOR2_X1 U402 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U403 ( .A(n340), .B(n339), .ZN(n345) );
  XOR2_X1 U404 ( .A(G78GAT), .B(G148GAT), .Z(n342) );
  XNOR2_X1 U405 ( .A(G106GAT), .B(KEYINPUT73), .ZN(n341) );
  XNOR2_X1 U406 ( .A(n342), .B(n341), .ZN(n424) );
  XNOR2_X1 U407 ( .A(G176GAT), .B(G204GAT), .ZN(n343) );
  XNOR2_X1 U408 ( .A(n290), .B(n343), .ZN(n406) );
  XOR2_X1 U409 ( .A(n424), .B(n406), .Z(n344) );
  INV_X1 U410 ( .A(n573), .ZN(n347) );
  INV_X1 U411 ( .A(KEYINPUT41), .ZN(n346) );
  NAND2_X1 U412 ( .A1(n347), .A2(n346), .ZN(n349) );
  NAND2_X1 U413 ( .A1(n573), .A2(KEYINPUT41), .ZN(n348) );
  NAND2_X1 U414 ( .A1(n349), .A2(n348), .ZN(n350) );
  NAND2_X1 U415 ( .A1(n570), .A2(n554), .ZN(n351) );
  XNOR2_X1 U416 ( .A(n351), .B(KEYINPUT46), .ZN(n386) );
  XOR2_X1 U417 ( .A(G36GAT), .B(G190GAT), .Z(n405) );
  XOR2_X1 U418 ( .A(KEYINPUT81), .B(KEYINPUT9), .Z(n355) );
  XNOR2_X1 U419 ( .A(G106GAT), .B(G92GAT), .ZN(n354) );
  XNOR2_X1 U420 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U421 ( .A(n356), .B(KEYINPUT80), .Z(n358) );
  XOR2_X1 U422 ( .A(G50GAT), .B(G162GAT), .Z(n432) );
  XNOR2_X1 U423 ( .A(G218GAT), .B(n432), .ZN(n357) );
  XNOR2_X1 U424 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U425 ( .A(n360), .B(n359), .ZN(n368) );
  XOR2_X1 U426 ( .A(n361), .B(KEYINPUT10), .Z(n366) );
  XOR2_X1 U427 ( .A(KEYINPUT78), .B(KEYINPUT65), .Z(n363) );
  XNOR2_X1 U428 ( .A(G134GAT), .B(KEYINPUT79), .ZN(n362) );
  XNOR2_X1 U429 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U430 ( .A(n364), .B(KEYINPUT11), .ZN(n365) );
  XNOR2_X1 U431 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X2 U432 ( .A(n368), .B(n367), .Z(n562) );
  XOR2_X1 U433 ( .A(G78GAT), .B(G211GAT), .Z(n370) );
  XNOR2_X1 U434 ( .A(G183GAT), .B(G71GAT), .ZN(n369) );
  XNOR2_X1 U435 ( .A(n370), .B(n369), .ZN(n384) );
  XOR2_X1 U436 ( .A(G8GAT), .B(KEYINPUT82), .Z(n409) );
  XOR2_X1 U437 ( .A(n371), .B(n409), .Z(n373) );
  XOR2_X1 U438 ( .A(G15GAT), .B(G127GAT), .Z(n440) );
  XOR2_X1 U439 ( .A(G22GAT), .B(G155GAT), .Z(n431) );
  XNOR2_X1 U440 ( .A(n440), .B(n431), .ZN(n372) );
  XNOR2_X1 U441 ( .A(n373), .B(n372), .ZN(n377) );
  XOR2_X1 U442 ( .A(KEYINPUT84), .B(KEYINPUT14), .Z(n375) );
  NAND2_X1 U443 ( .A1(G231GAT), .A2(G233GAT), .ZN(n374) );
  XNOR2_X1 U444 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U445 ( .A(n377), .B(n376), .Z(n382) );
  XOR2_X1 U446 ( .A(KEYINPUT15), .B(KEYINPUT12), .Z(n379) );
  XNOR2_X1 U447 ( .A(G1GAT), .B(G64GAT), .ZN(n378) );
  XNOR2_X1 U448 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U449 ( .A(n380), .B(KEYINPUT83), .ZN(n381) );
  XNOR2_X1 U450 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U451 ( .A(n384), .B(n383), .ZN(n484) );
  INV_X1 U452 ( .A(n484), .ZN(n577) );
  NOR2_X1 U453 ( .A1(n562), .A2(n577), .ZN(n385) );
  AND2_X1 U454 ( .A1(n386), .A2(n385), .ZN(n387) );
  XNOR2_X1 U455 ( .A(n387), .B(KEYINPUT47), .ZN(n393) );
  XOR2_X1 U456 ( .A(n562), .B(KEYINPUT36), .Z(n583) );
  NOR2_X1 U457 ( .A1(n484), .A2(n583), .ZN(n388) );
  NAND2_X1 U458 ( .A1(n389), .A2(n573), .ZN(n390) );
  XNOR2_X1 U459 ( .A(KEYINPUT117), .B(n391), .ZN(n392) );
  NAND2_X1 U460 ( .A1(n393), .A2(n392), .ZN(n395) );
  INV_X1 U461 ( .A(KEYINPUT48), .ZN(n394) );
  XNOR2_X1 U462 ( .A(n395), .B(n394), .ZN(n533) );
  XOR2_X1 U463 ( .A(KEYINPUT88), .B(KEYINPUT19), .Z(n397) );
  XNOR2_X1 U464 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n396) );
  XNOR2_X1 U465 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U466 ( .A(n398), .B(KEYINPUT89), .Z(n400) );
  XNOR2_X1 U467 ( .A(G169GAT), .B(G183GAT), .ZN(n399) );
  XNOR2_X1 U468 ( .A(n400), .B(n399), .ZN(n453) );
  XNOR2_X1 U469 ( .A(G211GAT), .B(KEYINPUT95), .ZN(n401) );
  XNOR2_X1 U470 ( .A(n401), .B(KEYINPUT94), .ZN(n402) );
  XOR2_X1 U471 ( .A(n402), .B(KEYINPUT21), .Z(n404) );
  XNOR2_X1 U472 ( .A(G197GAT), .B(G218GAT), .ZN(n403) );
  XNOR2_X1 U473 ( .A(n404), .B(n403), .ZN(n436) );
  XNOR2_X1 U474 ( .A(n453), .B(n436), .ZN(n415) );
  XOR2_X1 U475 ( .A(n406), .B(n405), .Z(n408) );
  NAND2_X1 U476 ( .A1(G226GAT), .A2(G233GAT), .ZN(n407) );
  XNOR2_X1 U477 ( .A(n408), .B(n407), .ZN(n413) );
  XNOR2_X1 U478 ( .A(n409), .B(KEYINPUT98), .ZN(n411) );
  XOR2_X1 U479 ( .A(n415), .B(n414), .Z(n525) );
  XNOR2_X1 U480 ( .A(KEYINPUT119), .B(n525), .ZN(n416) );
  XOR2_X1 U481 ( .A(KEYINPUT23), .B(G204GAT), .Z(n421) );
  NAND2_X1 U482 ( .A1(G228GAT), .A2(G233GAT), .ZN(n420) );
  XNOR2_X1 U483 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U484 ( .A(n422), .B(KEYINPUT93), .Z(n426) );
  XNOR2_X1 U485 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U486 ( .A(n426), .B(n425), .ZN(n430) );
  XOR2_X1 U487 ( .A(KEYINPUT92), .B(KEYINPUT22), .Z(n428) );
  XNOR2_X1 U488 ( .A(KEYINPUT96), .B(KEYINPUT24), .ZN(n427) );
  XNOR2_X1 U489 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U490 ( .A(n430), .B(n429), .Z(n434) );
  XNOR2_X1 U491 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U492 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U493 ( .A(n436), .B(n435), .ZN(n471) );
  NAND2_X1 U494 ( .A1(n568), .A2(n471), .ZN(n437) );
  XNOR2_X1 U495 ( .A(n437), .B(KEYINPUT55), .ZN(n456) );
  XOR2_X1 U496 ( .A(KEYINPUT90), .B(KEYINPUT20), .Z(n439) );
  XNOR2_X1 U497 ( .A(G190GAT), .B(G99GAT), .ZN(n438) );
  XNOR2_X1 U498 ( .A(n439), .B(n438), .ZN(n441) );
  XOR2_X1 U499 ( .A(n441), .B(n440), .Z(n443) );
  XNOR2_X1 U500 ( .A(G43GAT), .B(G113GAT), .ZN(n442) );
  XNOR2_X1 U501 ( .A(n443), .B(n442), .ZN(n449) );
  XOR2_X1 U502 ( .A(n445), .B(n444), .Z(n447) );
  NAND2_X1 U503 ( .A1(G227GAT), .A2(G233GAT), .ZN(n446) );
  XNOR2_X1 U504 ( .A(n447), .B(n446), .ZN(n448) );
  XOR2_X1 U505 ( .A(n449), .B(n448), .Z(n455) );
  XOR2_X1 U506 ( .A(KEYINPUT87), .B(KEYINPUT91), .Z(n451) );
  XNOR2_X1 U507 ( .A(G176GAT), .B(KEYINPUT86), .ZN(n450) );
  XNOR2_X1 U508 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U509 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U510 ( .A(n455), .B(n454), .ZN(n536) );
  NAND2_X1 U511 ( .A1(n456), .A2(n536), .ZN(n457) );
  NAND2_X1 U512 ( .A1(n563), .A2(n577), .ZN(n459) );
  XOR2_X1 U513 ( .A(n554), .B(KEYINPUT111), .Z(n539) );
  NAND2_X1 U514 ( .A1(n539), .A2(n563), .ZN(n463) );
  XOR2_X1 U515 ( .A(G176GAT), .B(KEYINPUT121), .Z(n461) );
  XOR2_X1 U516 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n460) );
  XNOR2_X1 U517 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U518 ( .A(n463), .B(n462), .ZN(G1349GAT) );
  NAND2_X1 U519 ( .A1(n525), .A2(n536), .ZN(n464) );
  NAND2_X1 U520 ( .A1(n464), .A2(n471), .ZN(n465) );
  XNOR2_X1 U521 ( .A(n465), .B(KEYINPUT101), .ZN(n466) );
  XOR2_X1 U522 ( .A(KEYINPUT25), .B(n466), .Z(n469) );
  XNOR2_X1 U523 ( .A(n525), .B(KEYINPUT27), .ZN(n472) );
  NOR2_X1 U524 ( .A1(n536), .A2(n471), .ZN(n467) );
  XNOR2_X1 U525 ( .A(KEYINPUT26), .B(n467), .ZN(n569) );
  AND2_X1 U526 ( .A1(n472), .A2(n569), .ZN(n468) );
  NOR2_X1 U527 ( .A1(n469), .A2(n468), .ZN(n470) );
  NOR2_X1 U528 ( .A1(n521), .A2(n470), .ZN(n475) );
  XNOR2_X1 U529 ( .A(KEYINPUT28), .B(n471), .ZN(n498) );
  NAND2_X1 U530 ( .A1(n472), .A2(n521), .ZN(n473) );
  XOR2_X1 U531 ( .A(KEYINPUT100), .B(n473), .Z(n549) );
  NAND2_X1 U532 ( .A1(n498), .A2(n549), .ZN(n534) );
  NOR2_X1 U533 ( .A1(n536), .A2(n534), .ZN(n474) );
  NOR2_X1 U534 ( .A1(n577), .A2(n486), .ZN(n476) );
  XNOR2_X1 U535 ( .A(n476), .B(KEYINPUT107), .ZN(n477) );
  NOR2_X1 U536 ( .A1(n583), .A2(n477), .ZN(n479) );
  NAND2_X1 U537 ( .A1(n570), .A2(n573), .ZN(n489) );
  NOR2_X1 U538 ( .A1(n520), .A2(n489), .ZN(n480) );
  NAND2_X1 U539 ( .A1(n521), .A2(n505), .ZN(n483) );
  XOR2_X1 U540 ( .A(G29GAT), .B(KEYINPUT39), .Z(n481) );
  NOR2_X1 U541 ( .A1(n562), .A2(n484), .ZN(n485) );
  XNOR2_X1 U542 ( .A(n485), .B(KEYINPUT16), .ZN(n488) );
  INV_X1 U543 ( .A(n486), .ZN(n487) );
  NAND2_X1 U544 ( .A1(n488), .A2(n487), .ZN(n509) );
  NOR2_X1 U545 ( .A1(n489), .A2(n509), .ZN(n499) );
  NAND2_X1 U546 ( .A1(n499), .A2(n521), .ZN(n493) );
  XOR2_X1 U547 ( .A(KEYINPUT103), .B(KEYINPUT102), .Z(n491) );
  XNOR2_X1 U548 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n490) );
  XNOR2_X1 U549 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U550 ( .A(n493), .B(n492), .ZN(G1324GAT) );
  NAND2_X1 U551 ( .A1(n525), .A2(n499), .ZN(n494) );
  XNOR2_X1 U552 ( .A(n494), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U553 ( .A(KEYINPUT104), .B(KEYINPUT35), .Z(n496) );
  NAND2_X1 U554 ( .A1(n499), .A2(n536), .ZN(n495) );
  XNOR2_X1 U555 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U556 ( .A(G15GAT), .B(n497), .ZN(G1326GAT) );
  XOR2_X1 U557 ( .A(G22GAT), .B(KEYINPUT105), .Z(n501) );
  INV_X1 U558 ( .A(n498), .ZN(n530) );
  NAND2_X1 U559 ( .A1(n499), .A2(n530), .ZN(n500) );
  XNOR2_X1 U560 ( .A(n501), .B(n500), .ZN(G1327GAT) );
  NAND2_X1 U561 ( .A1(n505), .A2(n525), .ZN(n502) );
  XNOR2_X1 U562 ( .A(n502), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U563 ( .A1(n505), .A2(n536), .ZN(n503) );
  XNOR2_X1 U564 ( .A(n503), .B(KEYINPUT40), .ZN(n504) );
  XNOR2_X1 U565 ( .A(G43GAT), .B(n504), .ZN(G1330GAT) );
  XOR2_X1 U566 ( .A(KEYINPUT109), .B(KEYINPUT110), .Z(n507) );
  NAND2_X1 U567 ( .A1(n505), .A2(n530), .ZN(n506) );
  XNOR2_X1 U568 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U569 ( .A(G50GAT), .B(n508), .ZN(G1331GAT) );
  XNOR2_X1 U570 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n511) );
  INV_X1 U571 ( .A(n570), .ZN(n551) );
  NAND2_X1 U572 ( .A1(n539), .A2(n551), .ZN(n519) );
  NOR2_X1 U573 ( .A1(n519), .A2(n509), .ZN(n515) );
  NAND2_X1 U574 ( .A1(n521), .A2(n515), .ZN(n510) );
  XNOR2_X1 U575 ( .A(n511), .B(n510), .ZN(G1332GAT) );
  NAND2_X1 U576 ( .A1(n525), .A2(n515), .ZN(n512) );
  XNOR2_X1 U577 ( .A(n512), .B(KEYINPUT112), .ZN(n513) );
  XNOR2_X1 U578 ( .A(G64GAT), .B(n513), .ZN(G1333GAT) );
  NAND2_X1 U579 ( .A1(n515), .A2(n536), .ZN(n514) );
  XNOR2_X1 U580 ( .A(n514), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U581 ( .A(KEYINPUT43), .B(KEYINPUT113), .Z(n517) );
  NAND2_X1 U582 ( .A1(n515), .A2(n530), .ZN(n516) );
  XNOR2_X1 U583 ( .A(n517), .B(n516), .ZN(n518) );
  XOR2_X1 U584 ( .A(G78GAT), .B(n518), .Z(G1335GAT) );
  XOR2_X1 U585 ( .A(KEYINPUT114), .B(KEYINPUT115), .Z(n523) );
  NOR2_X1 U586 ( .A1(n520), .A2(n519), .ZN(n529) );
  NAND2_X1 U587 ( .A1(n529), .A2(n521), .ZN(n522) );
  XNOR2_X1 U588 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X1 U589 ( .A(G85GAT), .B(n524), .ZN(G1336GAT) );
  NAND2_X1 U590 ( .A1(n525), .A2(n529), .ZN(n526) );
  XNOR2_X1 U591 ( .A(n526), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U592 ( .A1(n529), .A2(n536), .ZN(n527) );
  XNOR2_X1 U593 ( .A(n527), .B(KEYINPUT116), .ZN(n528) );
  XNOR2_X1 U594 ( .A(G99GAT), .B(n528), .ZN(G1338GAT) );
  NAND2_X1 U595 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U596 ( .A(n531), .B(KEYINPUT44), .ZN(n532) );
  XNOR2_X1 U597 ( .A(G106GAT), .B(n532), .ZN(G1339GAT) );
  NOR2_X1 U598 ( .A1(n533), .A2(n534), .ZN(n535) );
  NAND2_X1 U599 ( .A1(n536), .A2(n535), .ZN(n538) );
  NOR2_X1 U600 ( .A1(n551), .A2(n538), .ZN(n537) );
  XOR2_X1 U601 ( .A(G113GAT), .B(n537), .Z(G1340GAT) );
  XOR2_X1 U602 ( .A(G120GAT), .B(KEYINPUT49), .Z(n541) );
  INV_X1 U603 ( .A(n538), .ZN(n544) );
  NAND2_X1 U604 ( .A1(n544), .A2(n539), .ZN(n540) );
  XNOR2_X1 U605 ( .A(n541), .B(n540), .ZN(G1341GAT) );
  NAND2_X1 U606 ( .A1(n544), .A2(n577), .ZN(n542) );
  XNOR2_X1 U607 ( .A(n542), .B(KEYINPUT50), .ZN(n543) );
  XNOR2_X1 U608 ( .A(G127GAT), .B(n543), .ZN(G1342GAT) );
  XOR2_X1 U609 ( .A(KEYINPUT118), .B(KEYINPUT51), .Z(n546) );
  NAND2_X1 U610 ( .A1(n544), .A2(n562), .ZN(n545) );
  XNOR2_X1 U611 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U612 ( .A(G134GAT), .B(n547), .ZN(G1343GAT) );
  INV_X1 U613 ( .A(n569), .ZN(n548) );
  NOR2_X1 U614 ( .A1(n548), .A2(n533), .ZN(n550) );
  NAND2_X1 U615 ( .A1(n550), .A2(n549), .ZN(n553) );
  NOR2_X1 U616 ( .A1(n551), .A2(n553), .ZN(n552) );
  XOR2_X1 U617 ( .A(G141GAT), .B(n552), .Z(G1344GAT) );
  XOR2_X1 U618 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n556) );
  INV_X1 U619 ( .A(n553), .ZN(n559) );
  NAND2_X1 U620 ( .A1(n559), .A2(n554), .ZN(n555) );
  XNOR2_X1 U621 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U622 ( .A(G148GAT), .B(n557), .ZN(G1345GAT) );
  NAND2_X1 U623 ( .A1(n559), .A2(n577), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n558), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U625 ( .A1(n562), .A2(n559), .ZN(n560) );
  XNOR2_X1 U626 ( .A(n560), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U627 ( .A1(n570), .A2(n563), .ZN(n561) );
  XNOR2_X1 U628 ( .A(G169GAT), .B(n561), .ZN(G1348GAT) );
  NAND2_X1 U629 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n564), .B(KEYINPUT58), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n565), .B(G190GAT), .ZN(G1351GAT) );
  XOR2_X1 U632 ( .A(KEYINPUT123), .B(KEYINPUT59), .Z(n567) );
  XNOR2_X1 U633 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n566) );
  XNOR2_X1 U634 ( .A(n567), .B(n566), .ZN(n572) );
  NAND2_X1 U635 ( .A1(n569), .A2(n568), .ZN(n582) );
  INV_X1 U636 ( .A(n582), .ZN(n578) );
  NAND2_X1 U637 ( .A1(n578), .A2(n570), .ZN(n571) );
  XOR2_X1 U638 ( .A(n572), .B(n571), .Z(G1352GAT) );
  XOR2_X1 U639 ( .A(KEYINPUT61), .B(KEYINPUT124), .Z(n575) );
  OR2_X1 U640 ( .A1(n582), .A2(n573), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U642 ( .A(G204GAT), .B(n576), .ZN(G1353GAT) );
  NAND2_X1 U643 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n579), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U645 ( .A(KEYINPUT125), .B(KEYINPUT126), .Z(n581) );
  XNOR2_X1 U646 ( .A(G218GAT), .B(KEYINPUT62), .ZN(n580) );
  XNOR2_X1 U647 ( .A(n581), .B(n580), .ZN(n585) );
  NOR2_X1 U648 ( .A1(n583), .A2(n582), .ZN(n584) );
  XOR2_X1 U649 ( .A(n585), .B(n584), .Z(G1355GAT) );
endmodule

