//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 0 0 1 0 0 1 0 0 0 0 0 0 1 1 1 0 1 1 0 1 1 1 0 1 1 0 1 1 1 0 1 1 1 1 0 0 0 0 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:50 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n257, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1077, new_n1078,
    new_n1079, new_n1080, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1134, new_n1135, new_n1136, new_n1137, new_n1138, new_n1139,
    new_n1140, new_n1141, new_n1142, new_n1143, new_n1144, new_n1145,
    new_n1146, new_n1147, new_n1148, new_n1149, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1167, new_n1168, new_n1169, new_n1170, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  AOI22_X1  g0008(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n209));
  INV_X1    g0009(.A(G116), .ZN(new_n210));
  INV_X1    g0010(.A(G270), .ZN(new_n211));
  OAI21_X1  g0011(.A(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n213));
  INV_X1    g0013(.A(G68), .ZN(new_n214));
  INV_X1    g0014(.A(G238), .ZN(new_n215));
  INV_X1    g0015(.A(G257), .ZN(new_n216));
  OAI221_X1 g0016(.A(new_n213), .B1(new_n214), .B2(new_n215), .C1(new_n205), .C2(new_n216), .ZN(new_n217));
  AOI211_X1 g0017(.A(new_n212), .B(new_n217), .C1(G58), .C2(G232), .ZN(new_n218));
  INV_X1    g0018(.A(G1), .ZN(new_n219));
  INV_X1    g0019(.A(G20), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n218), .A2(new_n221), .ZN(new_n222));
  XOR2_X1   g0022(.A(new_n222), .B(KEYINPUT65), .Z(new_n223));
  NAND2_X1  g0023(.A1(new_n223), .A2(KEYINPUT1), .ZN(new_n224));
  XOR2_X1   g0024(.A(new_n224), .B(KEYINPUT66), .Z(new_n225));
  INV_X1    g0025(.A(G13), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n221), .A2(new_n226), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n228), .B(G250), .C1(G257), .C2(G264), .ZN(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT64), .B(KEYINPUT0), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  INV_X1    g0031(.A(new_n201), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n232), .A2(G50), .ZN(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(new_n234));
  NAND2_X1  g0034(.A1(G1), .A2(G13), .ZN(new_n235));
  INV_X1    g0035(.A(new_n235), .ZN(new_n236));
  NAND3_X1  g0036(.A1(new_n234), .A2(G20), .A3(new_n236), .ZN(new_n237));
  OAI21_X1  g0037(.A(new_n237), .B1(new_n223), .B2(KEYINPUT1), .ZN(new_n238));
  NOR3_X1   g0038(.A1(new_n225), .A2(new_n231), .A3(new_n238), .ZN(G361));
  XOR2_X1   g0039(.A(G238), .B(G244), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G232), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT2), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(G226), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G250), .B(G257), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT67), .ZN(new_n245));
  INV_X1    g0045(.A(G264), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(new_n211), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n243), .B(new_n248), .Z(G358));
  XNOR2_X1  g0049(.A(G87), .B(G97), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n250), .B(G107), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n251), .B(new_n210), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n252), .B(KEYINPUT68), .ZN(new_n253));
  XNOR2_X1  g0053(.A(G50), .B(G68), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n254), .B(G58), .ZN(new_n255));
  INV_X1    g0055(.A(G77), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n255), .B(new_n256), .ZN(new_n257));
  XNOR2_X1  g0057(.A(new_n253), .B(new_n257), .ZN(G351));
  INV_X1    g0058(.A(G58), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(KEYINPUT71), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT71), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G58), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT72), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n259), .A2(KEYINPUT8), .ZN(new_n265));
  AOI22_X1  g0065(.A1(new_n263), .A2(KEYINPUT8), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n266), .B1(new_n264), .B2(new_n265), .ZN(new_n267));
  INV_X1    g0067(.A(G33), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n268), .A2(G20), .ZN(new_n269));
  AOI22_X1  g0069(.A1(new_n267), .A2(new_n269), .B1(G20), .B2(new_n203), .ZN(new_n270));
  INV_X1    g0070(.A(G150), .ZN(new_n271));
  NOR2_X1   g0071(.A1(G20), .A2(G33), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n270), .B1(new_n271), .B2(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n236), .B1(new_n221), .B2(G33), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n219), .A2(G13), .A3(G20), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n279), .A2(G50), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n275), .B1(G1), .B2(new_n220), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n280), .B1(new_n281), .B2(G50), .ZN(new_n282));
  XNOR2_X1  g0082(.A(new_n282), .B(KEYINPUT73), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n277), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT3), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(new_n268), .ZN(new_n287));
  NAND2_X1  g0087(.A1(KEYINPUT3), .A2(G33), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G1698), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G222), .ZN(new_n292));
  OAI22_X1  g0092(.A1(new_n291), .A2(new_n292), .B1(new_n256), .B2(new_n289), .ZN(new_n293));
  AND2_X1   g0093(.A1(KEYINPUT3), .A2(G33), .ZN(new_n294));
  NOR2_X1   g0094(.A1(KEYINPUT3), .A2(G33), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n296), .A2(new_n290), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n293), .B1(G223), .B2(new_n297), .ZN(new_n298));
  XNOR2_X1  g0098(.A(new_n298), .B(KEYINPUT70), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n235), .B1(G33), .B2(G41), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G179), .ZN(new_n302));
  XNOR2_X1  g0102(.A(KEYINPUT69), .B(G45), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  OAI211_X1 g0104(.A(new_n219), .B(G274), .C1(new_n304), .C2(G41), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(new_n300), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n219), .B1(G41), .B2(G45), .ZN(new_n308));
  AND2_X1   g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n306), .B1(G226), .B2(new_n309), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n301), .A2(new_n302), .A3(new_n310), .ZN(new_n311));
  OR2_X1    g0111(.A1(new_n311), .A2(KEYINPUT74), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(KEYINPUT74), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n285), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n301), .A2(new_n310), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n314), .B1(G169), .B2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT9), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n284), .B1(KEYINPUT77), .B2(new_n319), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n319), .A2(KEYINPUT77), .ZN(new_n321));
  OR2_X1    g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n320), .A2(new_n321), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n316), .A2(G190), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n315), .A2(G200), .ZN(new_n325));
  NAND4_X1  g0125(.A1(new_n322), .A2(new_n323), .A3(new_n324), .A4(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(KEYINPUT10), .ZN(new_n327));
  AND2_X1   g0127(.A1(new_n324), .A2(new_n325), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT10), .ZN(new_n329));
  NAND4_X1  g0129(.A1(new_n328), .A2(new_n329), .A3(new_n322), .A4(new_n323), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n318), .B1(new_n327), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(G20), .A2(G77), .ZN(new_n332));
  XNOR2_X1  g0132(.A(KEYINPUT8), .B(G58), .ZN(new_n333));
  INV_X1    g0133(.A(new_n269), .ZN(new_n334));
  XNOR2_X1  g0134(.A(KEYINPUT15), .B(G87), .ZN(new_n335));
  OAI221_X1 g0135(.A(new_n332), .B1(new_n333), .B2(new_n273), .C1(new_n334), .C2(new_n335), .ZN(new_n336));
  AOI22_X1  g0136(.A1(new_n336), .A2(new_n276), .B1(new_n256), .B2(new_n279), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n337), .B1(new_n256), .B2(new_n281), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n289), .A2(G232), .A3(new_n290), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n289), .A2(G1698), .ZN(new_n340));
  OAI221_X1 g0140(.A(new_n339), .B1(new_n206), .B2(new_n289), .C1(new_n340), .C2(new_n215), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n306), .B1(new_n341), .B2(new_n300), .ZN(new_n342));
  INV_X1    g0142(.A(G244), .ZN(new_n343));
  INV_X1    g0143(.A(new_n309), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n342), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n338), .B1(new_n345), .B2(G200), .ZN(new_n346));
  XOR2_X1   g0146(.A(new_n346), .B(KEYINPUT76), .Z(new_n347));
  INV_X1    g0147(.A(G190), .ZN(new_n348));
  OR2_X1    g0148(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT75), .ZN(new_n350));
  XNOR2_X1  g0150(.A(new_n349), .B(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n347), .A2(new_n351), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n296), .A2(G1698), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(G226), .ZN(new_n354));
  NAND2_X1  g0154(.A1(G33), .A2(G97), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n289), .A2(G232), .A3(G1698), .ZN(new_n356));
  AND3_X1   g0156(.A1(new_n354), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  OAI221_X1 g0157(.A(new_n305), .B1(new_n215), .B2(new_n344), .C1(new_n357), .C2(new_n307), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT13), .ZN(new_n359));
  XNOR2_X1  g0159(.A(new_n358), .B(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(G169), .ZN(new_n361));
  OAI21_X1  g0161(.A(KEYINPUT14), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  XNOR2_X1  g0162(.A(new_n358), .B(KEYINPUT13), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT14), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n363), .A2(new_n364), .A3(G169), .ZN(new_n365));
  OAI211_X1 g0165(.A(new_n362), .B(new_n365), .C1(new_n302), .C2(new_n363), .ZN(new_n366));
  AOI22_X1  g0166(.A1(new_n269), .A2(G77), .B1(new_n272), .B2(G50), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n367), .B1(new_n220), .B2(G68), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n368), .A2(KEYINPUT11), .A3(new_n276), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n369), .B1(new_n214), .B2(new_n281), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n278), .A2(G68), .ZN(new_n371));
  XNOR2_X1  g0171(.A(new_n371), .B(KEYINPUT12), .ZN(new_n372));
  AOI21_X1  g0172(.A(KEYINPUT11), .B1(new_n368), .B2(new_n276), .ZN(new_n373));
  NOR3_X1   g0173(.A1(new_n370), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n366), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n360), .A2(G190), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n363), .A2(G200), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n377), .A2(new_n378), .A3(new_n374), .ZN(new_n379));
  AND2_X1   g0179(.A1(new_n345), .A2(new_n361), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n338), .B1(new_n345), .B2(G179), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n376), .A2(new_n379), .A3(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT7), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n385), .A2(G20), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n386), .A2(new_n287), .A3(new_n288), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(KEYINPUT78), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n287), .A2(new_n220), .A3(new_n288), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(new_n385), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT78), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n386), .A2(new_n287), .A3(new_n391), .A4(new_n288), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n388), .A2(new_n390), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(G68), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n260), .A2(new_n262), .A3(G68), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(new_n232), .ZN(new_n396));
  AOI22_X1  g0196(.A1(new_n396), .A2(G20), .B1(G159), .B2(new_n272), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n394), .A2(KEYINPUT16), .A3(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT16), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n272), .A2(G159), .ZN(new_n400));
  XNOR2_X1  g0200(.A(KEYINPUT71), .B(G58), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n201), .B1(new_n401), .B2(G68), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n400), .B1(new_n402), .B2(new_n220), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n214), .B1(new_n390), .B2(new_n387), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n399), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n398), .A2(new_n276), .A3(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(KEYINPUT79), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n267), .A2(new_n278), .ZN(new_n408));
  INV_X1    g0208(.A(new_n281), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n408), .B1(new_n267), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n396), .A2(G20), .ZN(new_n411));
  AOI22_X1  g0211(.A1(new_n389), .A2(new_n385), .B1(new_n296), .B2(new_n386), .ZN(new_n412));
  OAI211_X1 g0212(.A(new_n411), .B(new_n400), .C1(new_n412), .C2(new_n214), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n275), .B1(new_n413), .B2(new_n399), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT79), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n414), .A2(new_n415), .A3(new_n398), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n407), .A2(new_n410), .A3(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT80), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n407), .A2(KEYINPUT80), .A3(new_n410), .A4(new_n416), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n289), .A2(G226), .A3(G1698), .ZN(new_n422));
  NAND2_X1  g0222(.A1(G33), .A2(G87), .ZN(new_n423));
  OAI211_X1 g0223(.A(G223), .B(new_n290), .C1(new_n294), .C2(new_n295), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n422), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(new_n300), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n309), .A2(G232), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n426), .A2(new_n427), .A3(new_n305), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n428), .A2(new_n302), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n429), .B1(G169), .B2(new_n428), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  AOI21_X1  g0231(.A(KEYINPUT18), .B1(new_n421), .B2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT18), .ZN(new_n433));
  AOI211_X1 g0233(.A(new_n433), .B(new_n430), .C1(new_n419), .C2(new_n420), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT17), .ZN(new_n435));
  AND4_X1   g0235(.A1(new_n415), .A2(new_n398), .A3(new_n276), .A4(new_n405), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n415), .B1(new_n414), .B2(new_n398), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT81), .ZN(new_n439));
  INV_X1    g0239(.A(G200), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n428), .A2(new_n440), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n426), .A2(new_n427), .A3(new_n348), .A4(new_n305), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n438), .A2(new_n439), .A3(new_n410), .A4(new_n443), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n407), .A2(new_n410), .A3(new_n443), .A4(new_n416), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(KEYINPUT81), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n435), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n445), .A2(KEYINPUT17), .ZN(new_n448));
  OAI22_X1  g0248(.A1(new_n432), .A2(new_n434), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n384), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n331), .A2(new_n352), .A3(new_n450), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n289), .A2(G238), .A3(new_n290), .ZN(new_n452));
  NAND2_X1  g0252(.A1(G33), .A2(G116), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n452), .B(new_n453), .C1(new_n340), .C2(new_n343), .ZN(new_n454));
  INV_X1    g0254(.A(G45), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n455), .A2(G1), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n300), .A2(new_n456), .ZN(new_n457));
  AOI22_X1  g0257(.A1(new_n454), .A2(new_n300), .B1(G250), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n456), .A2(G274), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n458), .A2(G179), .A3(new_n459), .ZN(new_n460));
  AND2_X1   g0260(.A1(new_n458), .A2(new_n459), .ZN(new_n461));
  OAI211_X1 g0261(.A(KEYINPUT85), .B(new_n460), .C1(new_n461), .C2(new_n361), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT85), .ZN(new_n463));
  AND3_X1   g0263(.A1(new_n458), .A2(G179), .A3(new_n459), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n361), .B1(new_n458), .B2(new_n459), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n463), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n289), .A2(new_n220), .A3(G68), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT19), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n220), .B1(new_n355), .B2(new_n468), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n469), .B1(G87), .B2(new_n207), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n468), .B1(new_n355), .B2(G20), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n467), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  AOI22_X1  g0272(.A1(new_n472), .A2(new_n276), .B1(new_n279), .B2(new_n335), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n221), .A2(G33), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n268), .A2(G1), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(KEYINPUT83), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n474), .A2(new_n476), .A3(new_n235), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n278), .B1(new_n475), .B2(KEYINPUT83), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  XNOR2_X1  g0280(.A(new_n335), .B(KEYINPUT86), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n473), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n462), .A2(new_n466), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n458), .A2(new_n459), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(G200), .ZN(new_n485));
  AOI21_X1  g0285(.A(KEYINPUT87), .B1(new_n479), .B2(G87), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT87), .ZN(new_n487));
  INV_X1    g0287(.A(G87), .ZN(new_n488));
  NOR4_X1   g0288(.A1(new_n477), .A2(new_n487), .A3(new_n478), .A4(new_n488), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n473), .B1(new_n486), .B2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT88), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n485), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n461), .A2(G190), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n440), .B1(new_n458), .B2(new_n459), .ZN(new_n495));
  OAI21_X1  g0295(.A(KEYINPUT88), .B1(new_n495), .B2(new_n490), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n493), .A2(new_n494), .A3(new_n496), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n453), .A2(G20), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n289), .A2(new_n220), .A3(G87), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(KEYINPUT22), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT22), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n289), .A2(new_n501), .A3(new_n220), .A4(G87), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n498), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT24), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n220), .A2(G107), .ZN(new_n505));
  XNOR2_X1  g0305(.A(new_n505), .B(KEYINPUT23), .ZN(new_n506));
  AND3_X1   g0306(.A1(new_n503), .A2(new_n504), .A3(new_n506), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n504), .B1(new_n503), .B2(new_n506), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n276), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n479), .A2(G107), .ZN(new_n510));
  NAND2_X1  g0310(.A1(G33), .A2(G294), .ZN(new_n511));
  INV_X1    g0311(.A(G250), .ZN(new_n512));
  OAI221_X1 g0312(.A(new_n511), .B1(new_n340), .B2(new_n216), .C1(new_n512), .C2(new_n291), .ZN(new_n513));
  AND2_X1   g0313(.A1(KEYINPUT5), .A2(G41), .ZN(new_n514));
  NOR2_X1   g0314(.A1(KEYINPUT5), .A2(G41), .ZN(new_n515));
  OR2_X1    g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n300), .B1(new_n516), .B2(new_n456), .ZN(new_n517));
  AOI22_X1  g0317(.A1(new_n513), .A2(new_n300), .B1(G264), .B2(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n516), .A2(G274), .A3(new_n456), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n518), .A2(G190), .A3(new_n519), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n278), .A2(G107), .ZN(new_n521));
  XNOR2_X1  g0321(.A(new_n521), .B(KEYINPUT25), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n509), .A2(new_n510), .A3(new_n520), .A4(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n518), .A2(new_n519), .ZN(new_n524));
  INV_X1    g0324(.A(new_n524), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n525), .A2(new_n440), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n483), .B(new_n497), .C1(new_n523), .C2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n296), .A2(G303), .ZN(new_n528));
  OAI221_X1 g0328(.A(new_n528), .B1(new_n340), .B2(new_n246), .C1(new_n216), .C2(new_n291), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(new_n300), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n517), .A2(G270), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n530), .A2(new_n519), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(G200), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n279), .A2(new_n210), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n479), .A2(G116), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n275), .B1(G20), .B2(new_n210), .ZN(new_n536));
  NAND2_X1  g0336(.A1(G33), .A2(G283), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n537), .B(new_n220), .C1(G33), .C2(new_n205), .ZN(new_n538));
  AND3_X1   g0338(.A1(new_n536), .A2(KEYINPUT20), .A3(new_n538), .ZN(new_n539));
  AOI21_X1  g0339(.A(KEYINPUT20), .B1(new_n536), .B2(new_n538), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n534), .B(new_n535), .C1(new_n539), .C2(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(new_n541), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n533), .B(new_n542), .C1(new_n348), .C2(new_n532), .ZN(new_n543));
  AOI22_X1  g0343(.A1(new_n529), .A2(new_n300), .B1(G270), .B2(new_n517), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n541), .A2(new_n544), .A3(G179), .A4(new_n519), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n361), .B1(new_n544), .B2(new_n519), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT21), .ZN(new_n547));
  AND3_X1   g0347(.A1(new_n546), .A2(new_n547), .A3(new_n541), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n547), .B1(new_n546), .B2(new_n541), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n543), .B(new_n545), .C1(new_n548), .C2(new_n549), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n527), .A2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT4), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n552), .B1(new_n291), .B2(new_n343), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n353), .A2(KEYINPUT4), .A3(G244), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n297), .A2(G250), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n553), .A2(new_n554), .A3(new_n555), .A4(new_n537), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(new_n300), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n517), .A2(G257), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n557), .A2(new_n519), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(G169), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n560), .B1(new_n302), .B2(new_n559), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n279), .A2(new_n205), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n479), .A2(G97), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n272), .A2(G77), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT6), .ZN(new_n565));
  NOR3_X1   g0365(.A1(new_n565), .A2(new_n205), .A3(G107), .ZN(new_n566));
  XNOR2_X1  g0366(.A(G97), .B(G107), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n566), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  OAI221_X1 g0368(.A(new_n564), .B1(new_n568), .B2(new_n220), .C1(new_n412), .C2(new_n206), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT82), .ZN(new_n570));
  AND3_X1   g0370(.A1(new_n569), .A2(new_n570), .A3(new_n276), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n570), .B1(new_n569), .B2(new_n276), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n562), .B(new_n563), .C1(new_n571), .C2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n561), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n559), .A2(G200), .ZN(new_n575));
  AOI22_X1  g0375(.A1(new_n556), .A2(new_n300), .B1(G257), .B2(new_n517), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n576), .A2(G190), .A3(new_n519), .ZN(new_n577));
  AND2_X1   g0377(.A1(new_n573), .A2(KEYINPUT84), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n573), .A2(KEYINPUT84), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n575), .B(new_n577), .C1(new_n578), .C2(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n509), .A2(new_n510), .A3(new_n522), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n525), .A2(new_n302), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n581), .B(new_n582), .C1(G169), .C2(new_n525), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n551), .A2(new_n574), .A3(new_n580), .A4(new_n583), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n451), .A2(new_n584), .ZN(G372));
  NAND2_X1  g0385(.A1(new_n431), .A2(new_n417), .ZN(new_n586));
  XNOR2_X1  g0386(.A(new_n586), .B(KEYINPUT18), .ZN(new_n587));
  INV_X1    g0387(.A(new_n587), .ZN(new_n588));
  OR2_X1    g0388(.A1(new_n447), .A2(new_n448), .ZN(new_n589));
  INV_X1    g0389(.A(new_n589), .ZN(new_n590));
  AOI22_X1  g0390(.A1(new_n366), .A2(new_n375), .B1(new_n379), .B2(new_n382), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n588), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n327), .A2(new_n330), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n318), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n460), .B1(new_n461), .B2(new_n361), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n495), .A2(new_n490), .ZN(new_n596));
  AOI22_X1  g0396(.A1(new_n595), .A2(new_n482), .B1(new_n596), .B2(new_n494), .ZN(new_n597));
  INV_X1    g0397(.A(new_n572), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n569), .A2(new_n570), .A3(new_n276), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT84), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n600), .A2(new_n601), .A3(new_n562), .A4(new_n563), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n573), .A2(KEYINPUT84), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n597), .A2(new_n602), .A3(new_n603), .A4(new_n561), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n604), .A2(KEYINPUT26), .ZN(new_n605));
  AND2_X1   g0405(.A1(new_n595), .A2(new_n482), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n483), .A2(new_n497), .ZN(new_n608));
  OAI21_X1  g0408(.A(KEYINPUT26), .B1(new_n608), .B2(new_n574), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n545), .B1(new_n548), .B2(new_n549), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(KEYINPUT89), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT89), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n612), .B(new_n545), .C1(new_n548), .C2(new_n549), .ZN(new_n613));
  AND3_X1   g0413(.A1(new_n611), .A2(new_n583), .A3(new_n613), .ZN(new_n614));
  OR2_X1    g0414(.A1(new_n523), .A2(new_n526), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n580), .A2(new_n574), .A3(new_n615), .A4(new_n597), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n607), .B(new_n609), .C1(new_n614), .C2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(new_n617), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n594), .B1(new_n451), .B2(new_n618), .ZN(G369));
  NAND2_X1  g0419(.A1(new_n611), .A2(new_n613), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n226), .A2(G20), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(new_n219), .ZN(new_n622));
  OR2_X1    g0422(.A1(new_n622), .A2(KEYINPUT27), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(KEYINPUT27), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n623), .A2(G213), .A3(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(G343), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n542), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n620), .A2(new_n629), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n630), .B1(new_n550), .B2(new_n629), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(G330), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n583), .A2(new_n627), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n581), .A2(new_n627), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n615), .A2(new_n634), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n633), .B1(new_n635), .B2(new_n583), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n632), .A2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n610), .A2(new_n628), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n637), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n641), .A2(new_n633), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n639), .A2(new_n642), .ZN(G399));
  NOR2_X1   g0443(.A1(new_n227), .A2(G41), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  NOR3_X1   g0445(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n645), .A2(G1), .A3(new_n646), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n647), .B1(new_n233), .B2(new_n645), .ZN(new_n648));
  XNOR2_X1  g0448(.A(new_n648), .B(KEYINPUT28), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT91), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n559), .A2(new_n302), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n532), .A2(new_n484), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n651), .A2(KEYINPUT30), .A3(new_n652), .A4(new_n518), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n519), .B1(new_n576), .B2(new_n544), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n654), .A2(new_n302), .A3(new_n524), .A4(new_n484), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT30), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n576), .A2(G179), .A3(new_n518), .A4(new_n519), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n544), .A2(new_n519), .A3(new_n459), .A4(new_n458), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n656), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n653), .A2(new_n655), .A3(new_n659), .ZN(new_n660));
  XOR2_X1   g0460(.A(KEYINPUT90), .B(KEYINPUT31), .Z(new_n661));
  NAND3_X1  g0461(.A1(new_n660), .A2(new_n627), .A3(new_n661), .ZN(new_n662));
  AND2_X1   g0462(.A1(new_n660), .A2(new_n627), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT31), .ZN(new_n664));
  OAI211_X1 g0464(.A(new_n650), .B(new_n662), .C1(new_n663), .C2(new_n664), .ZN(new_n665));
  AND3_X1   g0465(.A1(new_n660), .A2(new_n627), .A3(new_n661), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n664), .B1(new_n660), .B2(new_n627), .ZN(new_n667));
  OAI21_X1  g0467(.A(KEYINPUT91), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  OAI211_X1 g0468(.A(new_n665), .B(new_n668), .C1(new_n584), .C2(new_n627), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(G330), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT92), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n669), .A2(KEYINPUT92), .A3(G330), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  NOR3_X1   g0475(.A1(new_n618), .A2(KEYINPUT29), .A3(new_n627), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT29), .ZN(new_n677));
  OR3_X1    g0477(.A1(new_n608), .A2(KEYINPUT26), .A3(new_n574), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n606), .B1(new_n604), .B2(KEYINPUT26), .ZN(new_n679));
  INV_X1    g0479(.A(new_n610), .ZN(new_n680));
  AND2_X1   g0480(.A1(new_n680), .A2(new_n583), .ZN(new_n681));
  OAI211_X1 g0481(.A(new_n678), .B(new_n679), .C1(new_n616), .C2(new_n681), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n677), .B1(new_n682), .B2(new_n628), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n676), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n675), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n649), .B1(new_n686), .B2(G1), .ZN(G364));
  AOI21_X1  g0487(.A(new_n219), .B1(new_n621), .B2(G45), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n644), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n220), .A2(G190), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n440), .A2(G179), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  XOR2_X1   g0494(.A(new_n694), .B(KEYINPUT97), .Z(new_n695));
  NOR2_X1   g0495(.A1(G179), .A2(G200), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n692), .A2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  AOI22_X1  g0498(.A1(new_n695), .A2(G283), .B1(G329), .B2(new_n698), .ZN(new_n699));
  XOR2_X1   g0499(.A(new_n699), .B(KEYINPUT98), .Z(new_n700));
  NAND3_X1  g0500(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n701), .A2(new_n348), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(G326), .ZN(new_n703));
  INV_X1    g0503(.A(G294), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n220), .B1(new_n696), .B2(G190), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n703), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n220), .A2(new_n348), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n302), .A2(G200), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(G322), .ZN(new_n710));
  INV_X1    g0510(.A(G303), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n707), .A2(new_n693), .ZN(new_n712));
  OAI221_X1 g0512(.A(new_n296), .B1(new_n709), .B2(new_n710), .C1(new_n711), .C2(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n701), .A2(G190), .ZN(new_n714));
  XNOR2_X1  g0514(.A(KEYINPUT99), .B(KEYINPUT33), .ZN(new_n715));
  XNOR2_X1  g0515(.A(new_n715), .B(G317), .ZN(new_n716));
  AOI211_X1 g0516(.A(new_n706), .B(new_n713), .C1(new_n714), .C2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(G311), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n692), .A2(new_n708), .ZN(new_n719));
  OAI211_X1 g0519(.A(new_n700), .B(new_n717), .C1(new_n718), .C2(new_n719), .ZN(new_n720));
  XNOR2_X1  g0520(.A(new_n720), .B(KEYINPUT100), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n719), .A2(new_n256), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n698), .A2(G159), .ZN(new_n723));
  XNOR2_X1  g0523(.A(new_n723), .B(KEYINPUT32), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n724), .B1(G68), .B2(new_n714), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n705), .A2(new_n205), .ZN(new_n726));
  OAI221_X1 g0526(.A(new_n289), .B1(new_n709), .B2(new_n263), .C1(new_n488), .C2(new_n712), .ZN(new_n727));
  AOI211_X1 g0527(.A(new_n726), .B(new_n727), .C1(G50), .C2(new_n702), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n695), .A2(G107), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n725), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n721), .B1(new_n722), .B2(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n235), .B1(G20), .B2(new_n361), .ZN(new_n732));
  OR2_X1    g0532(.A1(new_n732), .A2(KEYINPUT95), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(KEYINPUT95), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n691), .B1(new_n731), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n228), .A2(new_n296), .ZN(new_n737));
  XOR2_X1   g0537(.A(new_n737), .B(KEYINPUT93), .Z(new_n738));
  OAI221_X1 g0538(.A(new_n738), .B1(new_n233), .B2(new_n304), .C1(new_n257), .C2(new_n455), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n228), .A2(G355), .A3(new_n289), .ZN(new_n740));
  OAI211_X1 g0540(.A(new_n739), .B(new_n740), .C1(G116), .C2(new_n228), .ZN(new_n741));
  INV_X1    g0541(.A(new_n735), .ZN(new_n742));
  NOR2_X1   g0542(.A1(G13), .A2(G33), .ZN(new_n743));
  XOR2_X1   g0543(.A(new_n743), .B(KEYINPUT94), .Z(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(new_n220), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n742), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g0546(.A(new_n746), .B(KEYINPUT96), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n741), .A2(new_n748), .ZN(new_n749));
  OAI211_X1 g0549(.A(new_n736), .B(new_n749), .C1(new_n631), .C2(new_n745), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n632), .A2(new_n691), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n631), .A2(G330), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n750), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  XNOR2_X1  g0553(.A(new_n753), .B(KEYINPUT101), .ZN(G396));
  NOR2_X1   g0554(.A1(new_n383), .A2(new_n627), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n338), .A2(new_n627), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n352), .A2(new_n756), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n755), .B1(new_n757), .B2(new_n383), .ZN(new_n758));
  XNOR2_X1  g0558(.A(new_n674), .B(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n618), .A2(new_n627), .ZN(new_n760));
  XNOR2_X1  g0560(.A(new_n759), .B(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(new_n691), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n296), .B1(new_n712), .B2(new_n206), .ZN(new_n763));
  XOR2_X1   g0563(.A(new_n763), .B(KEYINPUT102), .Z(new_n764));
  NAND2_X1  g0564(.A1(new_n695), .A2(G87), .ZN(new_n765));
  INV_X1    g0565(.A(new_n709), .ZN(new_n766));
  AOI22_X1  g0566(.A1(G294), .A2(new_n766), .B1(new_n698), .B2(G311), .ZN(new_n767));
  AND3_X1   g0567(.A1(new_n764), .A2(new_n765), .A3(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n702), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(new_n711), .ZN(new_n770));
  AOI211_X1 g0570(.A(new_n726), .B(new_n770), .C1(G283), .C2(new_n714), .ZN(new_n771));
  OAI211_X1 g0571(.A(new_n768), .B(new_n771), .C1(new_n210), .C2(new_n719), .ZN(new_n772));
  XOR2_X1   g0572(.A(new_n772), .B(KEYINPUT103), .Z(new_n773));
  INV_X1    g0573(.A(G132), .ZN(new_n774));
  OAI221_X1 g0574(.A(new_n289), .B1(new_n697), .B2(new_n774), .C1(new_n263), .C2(new_n705), .ZN(new_n775));
  AND2_X1   g0575(.A1(new_n695), .A2(G68), .ZN(new_n776));
  INV_X1    g0576(.A(new_n719), .ZN(new_n777));
  AOI22_X1  g0577(.A1(new_n777), .A2(G159), .B1(G137), .B2(new_n702), .ZN(new_n778));
  INV_X1    g0578(.A(G143), .ZN(new_n779));
  INV_X1    g0579(.A(new_n714), .ZN(new_n780));
  OAI221_X1 g0580(.A(new_n778), .B1(new_n779), .B2(new_n709), .C1(new_n271), .C2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(KEYINPUT34), .ZN(new_n782));
  AOI211_X1 g0582(.A(new_n775), .B(new_n776), .C1(new_n781), .C2(new_n782), .ZN(new_n783));
  OAI221_X1 g0583(.A(new_n783), .B1(new_n782), .B2(new_n781), .C1(new_n202), .C2(new_n712), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n773), .A2(new_n784), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n691), .B1(new_n785), .B2(new_n735), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n735), .A2(new_n743), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n744), .ZN(new_n789));
  OAI221_X1 g0589(.A(new_n786), .B1(G77), .B2(new_n788), .C1(new_n758), .C2(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n762), .A2(new_n790), .ZN(G384));
  NAND2_X1  g0591(.A1(new_n394), .A2(new_n397), .ZN(new_n792));
  NOR2_X1   g0592(.A1(KEYINPUT104), .A2(KEYINPUT16), .ZN(new_n793));
  XNOR2_X1  g0593(.A(new_n792), .B(new_n793), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n410), .B1(new_n794), .B2(new_n275), .ZN(new_n795));
  INV_X1    g0595(.A(new_n625), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n795), .A2(new_n431), .ZN(new_n799));
  AND2_X1   g0599(.A1(new_n445), .A2(KEYINPUT81), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n445), .A2(KEYINPUT81), .ZN(new_n801));
  OAI211_X1 g0601(.A(new_n797), .B(new_n799), .C1(new_n800), .C2(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(KEYINPUT37), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n625), .B1(new_n419), .B2(new_n420), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(KEYINPUT80), .B1(new_n438), .B2(new_n410), .ZN(new_n806));
  INV_X1    g0606(.A(new_n420), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n431), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(KEYINPUT37), .B1(new_n444), .B2(new_n446), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n805), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  AOI22_X1  g0610(.A1(new_n449), .A2(new_n798), .B1(new_n803), .B2(new_n810), .ZN(new_n811));
  OAI21_X1  g0611(.A(KEYINPUT105), .B1(new_n811), .B2(KEYINPUT38), .ZN(new_n812));
  INV_X1    g0612(.A(KEYINPUT105), .ZN(new_n813));
  INV_X1    g0613(.A(KEYINPUT38), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n808), .A2(new_n433), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n421), .A2(KEYINPUT18), .A3(new_n431), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n797), .B1(new_n817), .B2(new_n589), .ZN(new_n818));
  AND2_X1   g0618(.A1(new_n803), .A2(new_n810), .ZN(new_n819));
  OAI211_X1 g0619(.A(new_n813), .B(new_n814), .C1(new_n818), .C2(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n811), .A2(KEYINPUT38), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n812), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n375), .A2(new_n627), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n376), .A2(new_n379), .A3(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n379), .ZN(new_n825));
  OAI211_X1 g0625(.A(new_n375), .B(new_n627), .C1(new_n825), .C2(new_n366), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n663), .A2(new_n661), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n828), .B1(new_n584), .B2(new_n627), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n663), .A2(new_n664), .ZN(new_n830));
  AND4_X1   g0630(.A1(new_n758), .A2(new_n827), .A3(new_n829), .A4(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n822), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT40), .ZN(new_n833));
  AOI21_X1  g0633(.A(KEYINPUT106), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT106), .ZN(new_n835));
  AOI211_X1 g0635(.A(new_n835), .B(KEYINPUT40), .C1(new_n822), .C2(new_n831), .ZN(new_n836));
  OR2_X1    g0636(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n805), .B1(new_n589), .B2(new_n588), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n586), .A2(new_n445), .ZN(new_n839));
  OAI21_X1  g0639(.A(KEYINPUT37), .B1(new_n804), .B2(new_n839), .ZN(new_n840));
  AND2_X1   g0640(.A1(new_n810), .A2(new_n840), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n814), .B1(new_n838), .B2(new_n841), .ZN(new_n842));
  AND3_X1   g0642(.A1(new_n821), .A2(new_n842), .A3(KEYINPUT107), .ZN(new_n843));
  AOI21_X1  g0643(.A(KEYINPUT107), .B1(new_n821), .B2(new_n842), .ZN(new_n844));
  OAI211_X1 g0644(.A(KEYINPUT40), .B(new_n831), .C1(new_n843), .C2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n837), .A2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n451), .ZN(new_n847));
  AND2_X1   g0647(.A1(new_n829), .A2(new_n830), .ZN(new_n848));
  AND2_X1   g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  XOR2_X1   g0649(.A(new_n849), .B(KEYINPUT108), .Z(new_n850));
  XNOR2_X1  g0650(.A(new_n846), .B(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n851), .A2(G330), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n757), .A2(new_n383), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n617), .A2(new_n628), .A3(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n755), .ZN(new_n855));
  AND2_X1   g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n857), .A2(new_n827), .A3(new_n822), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n587), .A2(new_n625), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n821), .A2(new_n842), .ZN(new_n860));
  OR2_X1    g0660(.A1(new_n860), .A2(KEYINPUT39), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n822), .A2(KEYINPUT39), .ZN(new_n862));
  AND2_X1   g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n376), .A2(new_n627), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(new_n865));
  OAI211_X1 g0665(.A(new_n858), .B(new_n859), .C1(new_n863), .C2(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n847), .B1(new_n683), .B2(new_n676), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n594), .ZN(new_n868));
  XOR2_X1   g0668(.A(new_n866), .B(new_n868), .Z(new_n869));
  XNOR2_X1  g0669(.A(new_n852), .B(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n870), .B1(new_n219), .B2(new_n621), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT35), .ZN(new_n872));
  AOI211_X1 g0672(.A(new_n220), .B(new_n235), .C1(new_n568), .C2(new_n872), .ZN(new_n873));
  OAI211_X1 g0673(.A(new_n873), .B(G116), .C1(new_n872), .C2(new_n568), .ZN(new_n874));
  XNOR2_X1  g0674(.A(new_n874), .B(KEYINPUT36), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n234), .A2(G77), .A3(new_n395), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n876), .B1(G50), .B2(new_n214), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n877), .A2(G1), .A3(new_n226), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n871), .A2(new_n875), .A3(new_n878), .ZN(G367));
  INV_X1    g0679(.A(KEYINPUT109), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n578), .A2(new_n579), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(new_n627), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n882), .A2(new_n574), .A3(new_n580), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n881), .A2(new_n561), .A3(new_n627), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n641), .A2(new_n880), .A3(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT42), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n880), .B1(new_n641), .B2(new_n885), .ZN(new_n889));
  OR3_X1    g0689(.A1(new_n887), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n885), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n574), .B1(new_n891), .B2(new_n583), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(new_n628), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n888), .B1(new_n887), .B2(new_n889), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n890), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n639), .A2(new_n891), .ZN(new_n896));
  INV_X1    g0696(.A(new_n896), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n491), .A2(new_n628), .ZN(new_n898));
  MUX2_X1   g0698(.A(new_n597), .B(new_n606), .S(new_n898), .Z(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(KEYINPUT43), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n895), .A2(new_n897), .A3(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n899), .A2(KEYINPUT43), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n897), .B1(new_n895), .B2(new_n900), .ZN(new_n905));
  OR3_X1    g0705(.A1(new_n902), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n904), .B1(new_n902), .B2(new_n905), .ZN(new_n907));
  XNOR2_X1  g0707(.A(new_n644), .B(KEYINPUT41), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n642), .A2(new_n885), .ZN(new_n910));
  OR2_X1    g0710(.A1(new_n910), .A2(KEYINPUT110), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(KEYINPUT110), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT45), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n642), .A2(new_n885), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n916), .B(KEYINPUT44), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n911), .A2(KEYINPUT45), .A3(new_n912), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n915), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(new_n638), .ZN(new_n920));
  NAND4_X1  g0720(.A1(new_n915), .A2(new_n917), .A3(new_n639), .A4(new_n918), .ZN(new_n921));
  XOR2_X1   g0721(.A(new_n636), .B(new_n640), .Z(new_n922));
  XNOR2_X1  g0722(.A(new_n922), .B(new_n632), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n685), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n920), .A2(new_n921), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n909), .B1(new_n925), .B2(new_n686), .ZN(new_n926));
  OAI211_X1 g0726(.A(new_n906), .B(new_n907), .C1(new_n926), .C2(new_n689), .ZN(new_n927));
  INV_X1    g0727(.A(new_n705), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(G68), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n296), .B1(new_n714), .B2(G159), .ZN(new_n930));
  OAI211_X1 g0730(.A(new_n929), .B(new_n930), .C1(new_n779), .C2(new_n769), .ZN(new_n931));
  AOI22_X1  g0731(.A1(G150), .A2(new_n766), .B1(new_n777), .B2(G50), .ZN(new_n932));
  INV_X1    g0732(.A(G137), .ZN(new_n933));
  OAI221_X1 g0733(.A(new_n932), .B1(new_n256), .B2(new_n694), .C1(new_n933), .C2(new_n697), .ZN(new_n934));
  INV_X1    g0734(.A(new_n712), .ZN(new_n935));
  AOI211_X1 g0735(.A(new_n931), .B(new_n934), .C1(new_n401), .C2(new_n935), .ZN(new_n936));
  XOR2_X1   g0736(.A(new_n936), .B(KEYINPUT111), .Z(new_n937));
  OAI21_X1  g0737(.A(new_n296), .B1(new_n780), .B2(new_n704), .ZN(new_n938));
  INV_X1    g0738(.A(G283), .ZN(new_n939));
  OAI22_X1  g0739(.A1(new_n205), .A2(new_n694), .B1(new_n719), .B2(new_n939), .ZN(new_n940));
  AOI211_X1 g0740(.A(new_n938), .B(new_n940), .C1(G317), .C2(new_n698), .ZN(new_n941));
  OAI22_X1  g0741(.A1(new_n769), .A2(new_n718), .B1(new_n705), .B2(new_n206), .ZN(new_n942));
  OR3_X1    g0742(.A1(new_n712), .A2(KEYINPUT46), .A3(new_n210), .ZN(new_n943));
  OAI21_X1  g0743(.A(KEYINPUT46), .B1(new_n712), .B2(new_n210), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n942), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  OAI211_X1 g0745(.A(new_n941), .B(new_n945), .C1(new_n711), .C2(new_n709), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n937), .A2(new_n946), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n947), .B(KEYINPUT47), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(new_n735), .ZN(new_n949));
  OR2_X1    g0749(.A1(new_n899), .A2(new_n745), .ZN(new_n950));
  INV_X1    g0750(.A(new_n738), .ZN(new_n951));
  OAI221_X1 g0751(.A(new_n748), .B1(new_n228), .B2(new_n335), .C1(new_n248), .C2(new_n951), .ZN(new_n952));
  NAND4_X1  g0752(.A1(new_n949), .A2(new_n690), .A3(new_n950), .A4(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n927), .A2(new_n953), .ZN(G387));
  INV_X1    g0754(.A(new_n924), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n645), .B1(new_n685), .B2(new_n923), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n333), .A2(G50), .ZN(new_n958));
  INV_X1    g0758(.A(new_n958), .ZN(new_n959));
  OAI221_X1 g0759(.A(new_n646), .B1(new_n214), .B2(new_n256), .C1(new_n959), .C2(KEYINPUT50), .ZN(new_n960));
  AOI211_X1 g0760(.A(G45), .B(new_n960), .C1(KEYINPUT50), .C2(new_n959), .ZN(new_n961));
  INV_X1    g0761(.A(new_n243), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n738), .B1(new_n962), .B2(new_n303), .ZN(new_n963));
  OR3_X1    g0763(.A1(new_n646), .A2(new_n227), .A3(new_n296), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n961), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n965), .B1(new_n206), .B2(new_n227), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n690), .B1(new_n966), .B2(new_n747), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n967), .B(KEYINPUT112), .ZN(new_n968));
  AOI22_X1  g0768(.A1(new_n777), .A2(G303), .B1(G322), .B2(new_n702), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n969), .B1(new_n718), .B2(new_n780), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n970), .B1(G317), .B2(new_n766), .ZN(new_n971));
  XOR2_X1   g0771(.A(new_n971), .B(KEYINPUT48), .Z(new_n972));
  OAI221_X1 g0772(.A(new_n972), .B1(new_n939), .B2(new_n705), .C1(new_n704), .C2(new_n712), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT49), .ZN(new_n974));
  OR2_X1    g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n698), .A2(G326), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n973), .A2(new_n974), .ZN(new_n977));
  INV_X1    g0777(.A(new_n694), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n289), .B1(new_n978), .B2(G116), .ZN(new_n979));
  NAND4_X1  g0779(.A1(new_n975), .A2(new_n976), .A3(new_n977), .A4(new_n979), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n481), .A2(new_n705), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n712), .A2(new_n256), .ZN(new_n982));
  AOI211_X1 g0782(.A(new_n296), .B(new_n982), .C1(G50), .C2(new_n766), .ZN(new_n983));
  INV_X1    g0783(.A(G159), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n983), .B1(new_n984), .B2(new_n769), .ZN(new_n985));
  AOI211_X1 g0785(.A(new_n981), .B(new_n985), .C1(G97), .C2(new_n695), .ZN(new_n986));
  AOI22_X1  g0786(.A1(new_n267), .A2(new_n714), .B1(G68), .B2(new_n777), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT113), .ZN(new_n988));
  OAI211_X1 g0788(.A(new_n986), .B(new_n988), .C1(new_n271), .C2(new_n697), .ZN(new_n989));
  AND2_X1   g0789(.A1(new_n980), .A2(new_n989), .ZN(new_n990));
  OAI221_X1 g0790(.A(new_n968), .B1(new_n636), .B2(new_n745), .C1(new_n742), .C2(new_n990), .ZN(new_n991));
  XOR2_X1   g0791(.A(new_n991), .B(KEYINPUT114), .Z(new_n992));
  OAI211_X1 g0792(.A(new_n957), .B(new_n992), .C1(new_n688), .C2(new_n923), .ZN(G393));
  NAND2_X1  g0793(.A1(new_n920), .A2(new_n921), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT115), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n920), .A2(KEYINPUT115), .A3(new_n921), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n996), .A2(new_n689), .A3(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n994), .A2(new_n955), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n999), .A2(new_n925), .A3(new_n644), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n951), .A2(new_n252), .ZN(new_n1001));
  AOI211_X1 g0801(.A(new_n747), .B(new_n1001), .C1(G97), .C2(new_n227), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n289), .B1(new_n935), .B2(G283), .ZN(new_n1003));
  OAI211_X1 g0803(.A(new_n729), .B(new_n1003), .C1(new_n710), .C2(new_n697), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT117), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(new_n766), .A2(G311), .B1(G317), .B2(new_n702), .ZN(new_n1006));
  XOR2_X1   g0806(.A(KEYINPUT116), .B(KEYINPUT52), .Z(new_n1007));
  AND2_X1   g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n780), .A2(new_n711), .B1(new_n705), .B2(new_n210), .ZN(new_n1010));
  NOR3_X1   g0810(.A1(new_n1008), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  OAI211_X1 g0811(.A(new_n1005), .B(new_n1011), .C1(new_n704), .C2(new_n719), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n712), .A2(new_n214), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n705), .A2(new_n256), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n289), .B1(new_n697), .B2(new_n779), .C1(new_n333), .C2(new_n719), .ZN(new_n1015));
  AOI211_X1 g0815(.A(new_n1014), .B(new_n1015), .C1(G50), .C2(new_n714), .ZN(new_n1016));
  OAI22_X1  g0816(.A1(new_n769), .A2(new_n271), .B1(new_n709), .B2(new_n984), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1017), .B(KEYINPUT51), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1016), .A2(new_n765), .A3(new_n1018), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1012), .B1(new_n1013), .B2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1002), .B1(new_n1020), .B2(new_n735), .ZN(new_n1021));
  OAI211_X1 g0821(.A(new_n690), .B(new_n1021), .C1(new_n885), .C2(new_n745), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n998), .A2(new_n1000), .A3(new_n1022), .ZN(G390));
  NAND3_X1  g0823(.A1(new_n847), .A2(G330), .A3(new_n848), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n867), .A2(new_n1024), .A3(new_n594), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n827), .B1(new_n674), .B2(new_n758), .ZN(new_n1026));
  AND2_X1   g0826(.A1(new_n831), .A2(G330), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n857), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n674), .A2(new_n758), .A3(new_n827), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n682), .A2(new_n628), .A3(new_n853), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1030), .A2(new_n855), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1031), .A2(KEYINPUT118), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT118), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1030), .A2(new_n1033), .A3(new_n855), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n848), .A2(G330), .A3(new_n758), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n827), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1029), .A2(new_n1035), .A3(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1025), .B1(new_n1028), .B2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1032), .A2(new_n827), .A3(new_n1034), .ZN(new_n1041));
  OAI211_X1 g0841(.A(new_n1041), .B(new_n865), .C1(new_n844), .C2(new_n843), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n865), .B1(new_n856), .B2(new_n1037), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1043), .A2(new_n862), .A3(new_n861), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1029), .ZN(new_n1045));
  AND3_X1   g0845(.A1(new_n1042), .A2(new_n1044), .A3(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1027), .B1(new_n1042), .B2(new_n1044), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1040), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  AND2_X1   g0848(.A1(new_n1048), .A2(new_n644), .ZN(new_n1049));
  OR2_X1    g0849(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1049), .B1(new_n1050), .B2(new_n1040), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n709), .A2(new_n210), .B1(new_n697), .B2(new_n704), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n776), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n777), .A2(G97), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n296), .B1(new_n712), .B2(new_n488), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT119), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n769), .A2(new_n939), .ZN(new_n1057));
  AOI211_X1 g0857(.A(new_n1014), .B(new_n1057), .C1(G107), .C2(new_n714), .ZN(new_n1058));
  NAND4_X1  g0858(.A1(new_n1053), .A2(new_n1054), .A3(new_n1056), .A4(new_n1058), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n289), .B1(new_n780), .B2(new_n933), .ZN(new_n1060));
  INV_X1    g0860(.A(G128), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n769), .A2(new_n1061), .B1(new_n705), .B2(new_n984), .ZN(new_n1062));
  AOI211_X1 g0862(.A(new_n1060), .B(new_n1062), .C1(G50), .C2(new_n978), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n698), .A2(G125), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(KEYINPUT54), .B(G143), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n709), .A2(new_n774), .B1(new_n719), .B2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n935), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT53), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1068), .B1(new_n712), .B2(new_n271), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1066), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1063), .A2(new_n1064), .A3(new_n1070), .ZN(new_n1071));
  AND2_X1   g0871(.A1(new_n1059), .A2(new_n1071), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n1072), .A2(new_n742), .B1(new_n267), .B2(new_n788), .ZN(new_n1073));
  AOI211_X1 g0873(.A(new_n691), .B(new_n1073), .C1(new_n863), .C2(new_n744), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1074), .B1(new_n1050), .B2(new_n689), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1051), .A2(new_n1075), .ZN(G378));
  OAI211_X1 g0876(.A(G330), .B(new_n845), .C1(new_n834), .C2(new_n836), .ZN(new_n1077));
  INV_X1    g0877(.A(KEYINPUT55), .ZN(new_n1078));
  AND3_X1   g0878(.A1(new_n593), .A2(new_n1078), .A3(new_n317), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1078), .B1(new_n593), .B2(new_n317), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n1081), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n285), .A2(new_n625), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1083), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1080), .A2(new_n1082), .A3(new_n1084), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1083), .B1(new_n1079), .B2(new_n1081), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(KEYINPUT122), .B(KEYINPUT56), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1088), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1088), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  AND2_X1   g0892(.A1(new_n1077), .A2(new_n1092), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n1077), .A2(new_n1092), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n866), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(new_n1087), .B(new_n1089), .ZN(new_n1096));
  NAND4_X1  g0896(.A1(new_n1096), .A2(new_n837), .A3(G330), .A4(new_n845), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n866), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1077), .A2(new_n1092), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1097), .A2(new_n1098), .A3(new_n1099), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1095), .A2(new_n689), .A3(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n691), .B1(new_n787), .B2(new_n202), .ZN(new_n1102));
  XOR2_X1   g0902(.A(new_n1102), .B(KEYINPUT121), .Z(new_n1103));
  OAI221_X1 g0903(.A(new_n929), .B1(new_n780), .B2(new_n205), .C1(new_n210), .C2(new_n769), .ZN(new_n1104));
  OR4_X1    g0904(.A1(G41), .A2(new_n1104), .A3(new_n289), .A4(new_n982), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n694), .A2(new_n263), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n481), .A2(new_n719), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n709), .A2(new_n206), .B1(new_n697), .B2(new_n939), .ZN(new_n1108));
  NOR4_X1   g0908(.A1(new_n1105), .A2(new_n1106), .A3(new_n1107), .A4(new_n1108), .ZN(new_n1109));
  XOR2_X1   g0909(.A(new_n1109), .B(KEYINPUT58), .Z(new_n1110));
  OAI21_X1  g0910(.A(new_n202), .B1(new_n294), .B2(G41), .ZN(new_n1111));
  OAI22_X1  g0911(.A1(new_n1061), .A2(new_n709), .B1(new_n712), .B2(new_n1065), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1112), .B1(G137), .B2(new_n777), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n928), .A2(G150), .B1(G125), .B2(new_n702), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n1113), .B(new_n1114), .C1(new_n774), .C2(new_n780), .ZN(new_n1115));
  XOR2_X1   g0915(.A(new_n1115), .B(KEYINPUT59), .Z(new_n1116));
  XNOR2_X1  g0916(.A(KEYINPUT120), .B(G124), .ZN(new_n1117));
  AOI21_X1  g0917(.A(G41), .B1(new_n698), .B2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(G33), .B1(new_n978), .B2(G159), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1116), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1120));
  AND3_X1   g0920(.A1(new_n1110), .A2(new_n1111), .A3(new_n1120), .ZN(new_n1121));
  OAI221_X1 g0921(.A(new_n1103), .B1(new_n742), .B2(new_n1121), .C1(new_n1092), .C2(new_n789), .ZN(new_n1122));
  AND3_X1   g0922(.A1(new_n1101), .A2(KEYINPUT123), .A3(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(KEYINPUT123), .B1(new_n1101), .B2(new_n1122), .ZN(new_n1124));
  OR2_X1    g0924(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1025), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1048), .A2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1095), .A2(new_n1100), .A3(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(KEYINPUT57), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n1095), .A2(new_n1100), .A3(new_n1127), .A4(KEYINPUT57), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1130), .A2(new_n644), .A3(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1125), .A2(new_n1132), .ZN(G375));
  INV_X1    g0933(.A(new_n1040), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1028), .A2(new_n1025), .A3(new_n1039), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1134), .A2(new_n908), .A3(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n688), .B1(new_n1028), .B2(new_n1039), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1037), .A2(KEYINPUT124), .A3(new_n743), .ZN(new_n1138));
  INV_X1    g0938(.A(KEYINPUT124), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n743), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1139), .B1(new_n827), .B2(new_n1140), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(G137), .A2(new_n766), .B1(new_n698), .B2(G128), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n769), .A2(new_n774), .ZN(new_n1143));
  INV_X1    g0943(.A(KEYINPUT125), .ZN(new_n1144));
  OAI221_X1 g0944(.A(new_n1142), .B1(new_n271), .B2(new_n719), .C1(new_n1143), .C2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1145), .B1(new_n1144), .B2(new_n1143), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n289), .B1(new_n780), .B2(new_n1065), .ZN(new_n1147));
  AOI211_X1 g0947(.A(new_n1106), .B(new_n1147), .C1(G50), .C2(new_n928), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n1146), .B(new_n1148), .C1(new_n984), .C2(new_n712), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n719), .A2(new_n206), .ZN(new_n1150));
  OAI221_X1 g0950(.A(new_n296), .B1(new_n780), .B2(new_n210), .C1(new_n704), .C2(new_n769), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(G283), .B2(new_n766), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n695), .A2(G77), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n712), .A2(new_n205), .B1(new_n697), .B2(new_n711), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n981), .A2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1152), .A2(new_n1153), .A3(new_n1155), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1149), .B1(new_n1150), .B2(new_n1156), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(new_n1157), .A2(new_n735), .B1(new_n214), .B2(new_n787), .ZN(new_n1158));
  AND3_X1   g0958(.A1(new_n1138), .A2(new_n1141), .A3(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1137), .B1(new_n690), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1136), .A2(new_n1160), .ZN(G381));
  NOR2_X1   g0961(.A1(G375), .A2(G378), .ZN(new_n1162));
  INV_X1    g0962(.A(G381), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(G393), .A2(G396), .ZN(new_n1164));
  NOR3_X1   g0964(.A1(G387), .A2(G384), .A3(G390), .ZN(new_n1165));
  NAND4_X1  g0965(.A1(new_n1162), .A2(new_n1163), .A3(new_n1164), .A4(new_n1165), .ZN(G407));
  NAND2_X1  g0966(.A1(new_n626), .A2(G213), .ZN(new_n1167));
  XOR2_X1   g0967(.A(new_n1167), .B(KEYINPUT126), .Z(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1162), .A2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(G407), .A2(G213), .A3(new_n1170), .ZN(G409));
  INV_X1    g0971(.A(new_n1167), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n1132), .B(G378), .C1(new_n1124), .C2(new_n1123), .ZN(new_n1173));
  INV_X1    g0973(.A(G378), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n1101), .B(new_n1122), .C1(new_n1128), .C2(new_n909), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1172), .B1(new_n1173), .B2(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT60), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n645), .B1(new_n1135), .B2(new_n1178), .ZN(new_n1179));
  OAI211_X1 g0979(.A(new_n1179), .B(new_n1134), .C1(new_n1178), .C2(new_n1135), .ZN(new_n1180));
  AOI21_X1  g0980(.A(G384), .B1(new_n1180), .B2(new_n1160), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1180), .A2(G384), .A3(new_n1160), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1184), .A2(G2897), .A3(new_n1169), .ZN(new_n1185));
  AND2_X1   g0985(.A1(new_n1172), .A2(G2897), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1185), .B1(new_n1184), .B2(new_n1186), .ZN(new_n1187));
  OAI21_X1  g0987(.A(KEYINPUT63), .B1(new_n1177), .B2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1184), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1177), .A2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1188), .A2(new_n1190), .ZN(new_n1191));
  XOR2_X1   g0991(.A(G393), .B(G396), .Z(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(G390), .A2(new_n927), .A3(new_n953), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(G390), .B1(new_n927), .B2(new_n953), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1193), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(G390), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(G387), .A2(new_n1198), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1199), .A2(new_n1192), .A3(new_n1194), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1197), .A2(new_n1200), .ZN(new_n1201));
  AOI211_X1 g1001(.A(new_n1169), .B(new_n1184), .C1(new_n1173), .C2(new_n1176), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1201), .B1(new_n1202), .B2(KEYINPUT63), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT61), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1191), .A2(new_n1203), .A3(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1169), .B1(new_n1173), .B2(new_n1176), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1204), .B1(new_n1206), .B2(new_n1187), .ZN(new_n1207));
  XOR2_X1   g1007(.A(KEYINPUT127), .B(KEYINPUT62), .Z(new_n1208));
  NAND2_X1  g1008(.A1(new_n1190), .A2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1202), .A2(KEYINPUT62), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1207), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1201), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1205), .B1(new_n1211), .B2(new_n1212), .ZN(G405));
  AOI21_X1  g1013(.A(G378), .B1(new_n1125), .B2(new_n1132), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1173), .ZN(new_n1215));
  OR3_X1    g1015(.A1(new_n1214), .A2(new_n1215), .A3(new_n1189), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1189), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1218), .A2(new_n1201), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1216), .A2(new_n1212), .A3(new_n1217), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1219), .A2(new_n1220), .ZN(G402));
endmodule


