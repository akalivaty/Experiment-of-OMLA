//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 1 0 1 0 0 0 0 1 1 1 1 0 0 0 0 0 0 1 1 1 0 1 1 1 0 0 1 0 1 0 0 1 0 0 1 0 0 1 0 1 0 1 1 1 0 1 1 1 1 1 1 0 1 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:58 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1259, new_n1260, new_n1261,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1335,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n210));
  INV_X1    g0010(.A(G77), .ZN(new_n211));
  INV_X1    g0011(.A(G244), .ZN(new_n212));
  INV_X1    g0012(.A(G87), .ZN(new_n213));
  INV_X1    g0013(.A(G250), .ZN(new_n214));
  OAI221_X1 g0014(.A(new_n210), .B1(new_n211), .B2(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n206), .B1(new_n215), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n219), .A2(KEYINPUT1), .ZN(new_n220));
  OR2_X1    g0020(.A1(new_n219), .A2(KEYINPUT1), .ZN(new_n221));
  NAND3_X1  g0021(.A1(new_n209), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G1), .A2(G13), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n223), .A2(new_n204), .ZN(new_n224));
  OAI21_X1  g0024(.A(G50), .B1(G58), .B2(G68), .ZN(new_n225));
  XOR2_X1   g0025(.A(new_n225), .B(KEYINPUT64), .Z(new_n226));
  XOR2_X1   g0026(.A(new_n226), .B(KEYINPUT65), .Z(new_n227));
  AOI21_X1  g0027(.A(new_n222), .B1(new_n224), .B2(new_n227), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT2), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(G226), .ZN(new_n231));
  INV_X1    g0031(.A(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XOR2_X1   g0037(.A(G68), .B(G77), .Z(new_n238));
  XOR2_X1   g0038(.A(G50), .B(G58), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n240), .B(new_n243), .Z(G351));
  INV_X1    g0044(.A(G200), .ZN(new_n245));
  INV_X1    g0045(.A(KEYINPUT66), .ZN(new_n246));
  AND2_X1   g0046(.A1(G33), .A2(G41), .ZN(new_n247));
  OAI21_X1  g0047(.A(G274), .B1(new_n247), .B2(new_n223), .ZN(new_n248));
  OAI21_X1  g0048(.A(new_n203), .B1(G41), .B2(G45), .ZN(new_n249));
  OAI21_X1  g0049(.A(new_n246), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(G274), .ZN(new_n251));
  AND2_X1   g0051(.A1(G1), .A2(G13), .ZN(new_n252));
  NAND2_X1  g0052(.A1(G33), .A2(G41), .ZN(new_n253));
  AOI21_X1  g0053(.A(new_n251), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G41), .ZN(new_n255));
  INV_X1    g0055(.A(G45), .ZN(new_n256));
  AOI21_X1  g0056(.A(G1), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n254), .A2(KEYINPUT66), .A3(new_n257), .ZN(new_n258));
  XNOR2_X1  g0058(.A(KEYINPUT3), .B(G33), .ZN(new_n259));
  INV_X1    g0059(.A(G1698), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(G222), .ZN(new_n261));
  INV_X1    g0061(.A(G223), .ZN(new_n262));
  OAI211_X1 g0062(.A(new_n259), .B(new_n261), .C1(new_n262), .C2(new_n260), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n253), .A2(G1), .A3(G13), .ZN(new_n264));
  INV_X1    g0064(.A(G33), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(KEYINPUT3), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT3), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G33), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n264), .B1(new_n269), .B2(new_n211), .ZN(new_n270));
  AOI22_X1  g0070(.A1(new_n250), .A2(new_n258), .B1(new_n263), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n264), .A2(new_n249), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(KEYINPUT67), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT67), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n272), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n274), .A2(G226), .A3(new_n276), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n245), .B1(new_n271), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n271), .A2(new_n277), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n278), .B1(new_n280), .B2(G190), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT71), .ZN(new_n282));
  AOI21_X1  g0082(.A(KEYINPUT10), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n203), .A2(G20), .ZN(new_n284));
  XNOR2_X1  g0084(.A(new_n284), .B(KEYINPUT68), .ZN(new_n285));
  AND2_X1   g0085(.A1(new_n285), .A2(G50), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n203), .A2(G13), .A3(G20), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(new_n223), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G50), .ZN(new_n292));
  AOI22_X1  g0092(.A1(new_n286), .A2(new_n291), .B1(new_n292), .B2(new_n288), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT9), .ZN(new_n294));
  XNOR2_X1  g0094(.A(KEYINPUT8), .B(G58), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n204), .A2(G33), .ZN(new_n296));
  INV_X1    g0096(.A(G150), .ZN(new_n297));
  NOR2_X1   g0097(.A1(G20), .A2(G33), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  OAI22_X1  g0099(.A1(new_n295), .A2(new_n296), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  NOR2_X1   g0100(.A1(G50), .A2(G58), .ZN(new_n301));
  INV_X1    g0101(.A(G68), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n204), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n290), .B1(new_n300), .B2(new_n303), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n293), .A2(new_n294), .A3(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n294), .B1(new_n293), .B2(new_n304), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n281), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n283), .A2(new_n308), .ZN(new_n309));
  OAI221_X1 g0109(.A(new_n281), .B1(new_n282), .B2(KEYINPUT10), .C1(new_n306), .C2(new_n307), .ZN(new_n310));
  INV_X1    g0110(.A(G179), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n280), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n293), .A2(new_n304), .ZN(new_n313));
  OAI211_X1 g0113(.A(new_n312), .B(new_n313), .C1(G169), .C2(new_n280), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n309), .A2(new_n310), .A3(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n274), .A2(G244), .A3(new_n276), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n250), .A2(new_n258), .ZN(new_n317));
  NAND2_X1  g0117(.A1(G238), .A2(G1698), .ZN(new_n318));
  OAI211_X1 g0118(.A(new_n259), .B(new_n318), .C1(new_n232), .C2(G1698), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n247), .A2(new_n223), .ZN(new_n320));
  OAI211_X1 g0120(.A(new_n319), .B(new_n320), .C1(G107), .C2(new_n259), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n316), .A2(new_n317), .A3(new_n321), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n322), .A2(G179), .ZN(new_n323));
  INV_X1    g0123(.A(G169), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n323), .B1(new_n324), .B2(new_n322), .ZN(new_n325));
  XNOR2_X1  g0125(.A(KEYINPUT15), .B(G87), .ZN(new_n326));
  OAI22_X1  g0126(.A1(new_n326), .A2(new_n296), .B1(new_n204), .B2(new_n211), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n295), .A2(new_n299), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n290), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  OR2_X1    g0129(.A1(new_n329), .A2(KEYINPUT69), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(KEYINPUT69), .ZN(new_n331));
  AOI22_X1  g0131(.A1(new_n330), .A2(new_n331), .B1(new_n211), .B2(new_n288), .ZN(new_n332));
  AND2_X1   g0132(.A1(new_n289), .A2(new_n223), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n333), .A2(KEYINPUT70), .A3(new_n287), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT70), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n335), .B1(new_n288), .B2(new_n290), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n285), .A2(new_n334), .A3(new_n336), .ZN(new_n337));
  OR2_X1    g0137(.A1(new_n337), .A2(new_n211), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n332), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n325), .A2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(G190), .ZN(new_n341));
  OR2_X1    g0141(.A1(new_n322), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n322), .A2(G200), .ZN(new_n343));
  NAND4_X1  g0143(.A1(new_n342), .A2(new_n332), .A3(new_n338), .A4(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n340), .A2(new_n344), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n315), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(KEYINPUT72), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT17), .ZN(new_n348));
  INV_X1    g0148(.A(new_n295), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n285), .A2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(new_n291), .ZN(new_n351));
  OAI22_X1  g0151(.A1(new_n350), .A2(new_n351), .B1(new_n349), .B2(new_n287), .ZN(new_n352));
  XNOR2_X1  g0152(.A(G58), .B(G68), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(G20), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n298), .A2(G159), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT7), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n357), .B1(new_n259), .B2(G20), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n269), .A2(KEYINPUT7), .A3(new_n204), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n356), .B1(new_n360), .B2(G68), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n333), .B1(new_n361), .B2(KEYINPUT16), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT16), .ZN(new_n363));
  OAI21_X1  g0163(.A(KEYINPUT73), .B1(new_n265), .B2(KEYINPUT3), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT73), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n365), .A2(new_n267), .A3(G33), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n364), .A2(new_n366), .A3(new_n266), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n357), .A2(G20), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n302), .B1(new_n369), .B2(new_n358), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n363), .B1(new_n370), .B2(new_n356), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n352), .B1(new_n362), .B2(new_n371), .ZN(new_n372));
  NOR3_X1   g0172(.A1(new_n248), .A2(new_n246), .A3(new_n249), .ZN(new_n373));
  AOI21_X1  g0173(.A(KEYINPUT66), .B1(new_n254), .B2(new_n257), .ZN(new_n374));
  OAI22_X1  g0174(.A1(new_n373), .A2(new_n374), .B1(new_n232), .B2(new_n272), .ZN(new_n375));
  NOR2_X1   g0175(.A1(G223), .A2(G1698), .ZN(new_n376));
  INV_X1    g0176(.A(G226), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n376), .B1(new_n377), .B2(G1698), .ZN(new_n378));
  AOI22_X1  g0178(.A1(new_n378), .A2(new_n259), .B1(G33), .B2(G87), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n379), .A2(new_n264), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n245), .B1(new_n375), .B2(new_n380), .ZN(new_n381));
  OAI21_X1  g0181(.A(KEYINPUT74), .B1(new_n379), .B2(new_n264), .ZN(new_n382));
  AND3_X1   g0182(.A1(new_n264), .A2(G232), .A3(new_n249), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n383), .B1(new_n250), .B2(new_n258), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n262), .A2(new_n260), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n377), .A2(G1698), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  OAI22_X1  g0187(.A1(new_n269), .A2(new_n387), .B1(new_n265), .B2(new_n213), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT74), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n388), .A2(new_n389), .A3(new_n320), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n382), .A2(new_n384), .A3(new_n390), .A4(new_n341), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n381), .A2(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n348), .B1(new_n372), .B2(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(KEYINPUT7), .B1(new_n269), .B2(new_n204), .ZN(new_n394));
  AOI211_X1 g0194(.A(new_n357), .B(G20), .C1(new_n266), .C2(new_n268), .ZN(new_n395));
  OAI21_X1  g0195(.A(G68), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(new_n356), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n396), .A2(KEYINPUT16), .A3(new_n397), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n371), .A2(new_n290), .A3(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(new_n352), .ZN(new_n400));
  AND4_X1   g0200(.A1(new_n348), .A2(new_n392), .A3(new_n399), .A4(new_n400), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n393), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n399), .A2(new_n400), .ZN(new_n403));
  AND2_X1   g0203(.A1(new_n382), .A2(new_n390), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n375), .A2(G179), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n384), .B1(new_n264), .B2(new_n379), .ZN(new_n406));
  AOI22_X1  g0206(.A1(new_n404), .A2(new_n405), .B1(new_n406), .B2(new_n324), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n403), .A2(KEYINPUT18), .A3(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(KEYINPUT18), .B1(new_n403), .B2(new_n407), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n408), .B1(new_n409), .B2(KEYINPUT75), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT18), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n382), .A2(new_n384), .A3(new_n390), .A4(new_n311), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n375), .A2(new_n380), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n412), .B1(new_n413), .B2(G169), .ZN(new_n414));
  NOR3_X1   g0214(.A1(new_n372), .A2(new_n411), .A3(new_n414), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n411), .B1(new_n372), .B2(new_n414), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT75), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n415), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n402), .B1(new_n410), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n347), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n302), .A2(G20), .ZN(new_n421));
  OAI221_X1 g0221(.A(new_n421), .B1(new_n296), .B2(new_n211), .C1(new_n299), .C2(new_n292), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n422), .A2(KEYINPUT11), .A3(new_n290), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT12), .ZN(new_n424));
  INV_X1    g0224(.A(G13), .ZN(new_n425));
  NOR3_X1   g0225(.A1(new_n424), .A2(new_n425), .A3(G1), .ZN(new_n426));
  INV_X1    g0226(.A(new_n421), .ZN(new_n427));
  AOI22_X1  g0227(.A1(new_n426), .A2(new_n427), .B1(new_n424), .B2(new_n287), .ZN(new_n428));
  AND2_X1   g0228(.A1(new_n423), .A2(new_n428), .ZN(new_n429));
  AND2_X1   g0229(.A1(new_n422), .A2(new_n290), .ZN(new_n430));
  AND2_X1   g0230(.A1(new_n337), .A2(KEYINPUT12), .ZN(new_n431));
  OAI221_X1 g0231(.A(new_n429), .B1(KEYINPUT11), .B2(new_n430), .C1(new_n431), .C2(new_n302), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT13), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n232), .A2(G1698), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n434), .B1(G226), .B2(G1698), .ZN(new_n435));
  INV_X1    g0235(.A(G97), .ZN(new_n436));
  OAI22_X1  g0236(.A1(new_n435), .A2(new_n269), .B1(new_n265), .B2(new_n436), .ZN(new_n437));
  AOI22_X1  g0237(.A1(new_n437), .A2(new_n320), .B1(new_n250), .B2(new_n258), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n274), .A2(G238), .A3(new_n276), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n433), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n438), .A2(new_n433), .A3(new_n439), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n324), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT14), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n442), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n444), .B(G169), .C1(new_n446), .C2(new_n440), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n441), .A2(G179), .A3(new_n442), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n432), .B1(new_n445), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n441), .A2(new_n442), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n432), .B1(new_n451), .B2(G200), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n452), .B1(new_n341), .B2(new_n451), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n450), .B(new_n453), .C1(new_n346), .C2(KEYINPUT72), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n420), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n288), .A2(new_n436), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n203), .A2(G33), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n291), .A2(new_n457), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n456), .B1(new_n458), .B2(new_n436), .ZN(new_n459));
  XOR2_X1   g0259(.A(G97), .B(G107), .Z(new_n460));
  XNOR2_X1  g0260(.A(KEYINPUT76), .B(KEYINPUT6), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n436), .A2(G107), .ZN(new_n463));
  AND2_X1   g0263(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  OAI21_X1  g0264(.A(G20), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n298), .A2(G77), .ZN(new_n466));
  INV_X1    g0266(.A(G107), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n269), .A2(new_n204), .ZN(new_n468));
  AOI22_X1  g0268(.A1(new_n468), .A2(new_n357), .B1(new_n367), .B2(new_n368), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n465), .B(new_n466), .C1(new_n467), .C2(new_n469), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n459), .B1(new_n470), .B2(new_n290), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n203), .A2(G45), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n255), .A2(KEYINPUT5), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT5), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(G41), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n473), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n477), .A2(G257), .A3(new_n264), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n254), .A2(new_n474), .A3(new_n473), .A4(new_n476), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n266), .A2(new_n268), .A3(G244), .A4(new_n260), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(KEYINPUT77), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(KEYINPUT4), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n266), .A2(new_n268), .A3(G250), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT77), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n485), .A2(KEYINPUT4), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(G1698), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n266), .A2(new_n268), .A3(G244), .ZN(new_n490));
  AOI22_X1  g0290(.A1(new_n490), .A2(new_n486), .B1(G33), .B2(G283), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n483), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n480), .B1(new_n492), .B2(new_n320), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(G190), .ZN(new_n494));
  AND2_X1   g0294(.A1(new_n471), .A2(new_n494), .ZN(new_n495));
  OAI21_X1  g0295(.A(KEYINPUT78), .B1(new_n493), .B2(new_n245), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT78), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n490), .A2(new_n486), .ZN(new_n498));
  NAND2_X1  g0298(.A1(G33), .A2(G283), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n260), .B1(new_n484), .B2(new_n487), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n264), .B1(new_n502), .B2(new_n483), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n497), .B(G200), .C1(new_n503), .C2(new_n480), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n496), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n495), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n492), .A2(new_n320), .ZN(new_n507));
  INV_X1    g0307(.A(new_n480), .ZN(new_n508));
  AOI21_X1  g0308(.A(G169), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  AOI211_X1 g0309(.A(G179), .B(new_n480), .C1(new_n492), .C2(new_n320), .ZN(new_n510));
  OR3_X1    g0310(.A1(new_n471), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(G116), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n265), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n259), .A2(G244), .A3(G1698), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n513), .B1(new_n514), .B2(KEYINPUT80), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n260), .A2(G238), .ZN(new_n516));
  OAI21_X1  g0316(.A(KEYINPUT79), .B1(new_n269), .B2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT79), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n259), .A2(new_n518), .A3(G238), .A4(new_n260), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  OR3_X1    g0320(.A1(new_n490), .A2(KEYINPUT80), .A3(new_n260), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n515), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(new_n320), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n473), .A2(new_n251), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n472), .A2(new_n214), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n524), .A2(new_n264), .A3(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n523), .A2(new_n311), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(KEYINPUT81), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n523), .A2(new_n526), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(new_n324), .ZN(new_n530));
  INV_X1    g0330(.A(new_n458), .ZN(new_n531));
  INV_X1    g0331(.A(new_n326), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT82), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n259), .A2(new_n204), .A3(G68), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n204), .B1(new_n265), .B2(new_n436), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n213), .A2(new_n436), .A3(new_n467), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n536), .A2(KEYINPUT19), .A3(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT19), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n539), .B1(new_n296), .B2(new_n436), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n535), .A2(new_n538), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(new_n290), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n532), .A2(new_n287), .ZN(new_n543));
  INV_X1    g0343(.A(new_n543), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n534), .B1(new_n542), .B2(new_n544), .ZN(new_n545));
  AOI211_X1 g0345(.A(KEYINPUT82), .B(new_n543), .C1(new_n541), .C2(new_n290), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n533), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(new_n526), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n548), .B1(new_n522), .B2(new_n320), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT81), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n549), .A2(new_n550), .A3(new_n311), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n528), .A2(new_n530), .A3(new_n547), .A4(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n542), .A2(new_n544), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(KEYINPUT82), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n542), .A2(new_n534), .A3(new_n544), .ZN(new_n555));
  AOI22_X1  g0355(.A1(new_n554), .A2(new_n555), .B1(G87), .B2(new_n531), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n529), .A2(G200), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n549), .A2(G190), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n506), .A2(new_n511), .A3(new_n552), .A4(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT25), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n561), .B1(new_n287), .B2(G107), .ZN(new_n562));
  NOR3_X1   g0362(.A1(new_n287), .A2(new_n561), .A3(G107), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  AOI22_X1  g0364(.A1(new_n531), .A2(G107), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT83), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT24), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n266), .A2(new_n268), .A3(new_n204), .A4(G87), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(KEYINPUT22), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT22), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n259), .A2(new_n571), .A3(new_n204), .A4(G87), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n296), .A2(new_n512), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT23), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n575), .B1(new_n204), .B2(G107), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n467), .A2(KEYINPUT23), .A3(G20), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n574), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n573), .A2(new_n578), .ZN(new_n579));
  NOR2_X1   g0379(.A1(KEYINPUT83), .A2(KEYINPUT24), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(new_n580), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n573), .A2(new_n582), .A3(new_n578), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n568), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n565), .B1(new_n584), .B2(new_n333), .ZN(new_n585));
  AND2_X1   g0385(.A1(G257), .A2(G1698), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n266), .A2(new_n268), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(KEYINPUT84), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n259), .A2(G250), .A3(new_n260), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT84), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n259), .A2(new_n590), .A3(new_n586), .ZN(new_n591));
  NAND2_X1  g0391(.A1(G33), .A2(G294), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n588), .A2(new_n589), .A3(new_n591), .A4(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(new_n320), .ZN(new_n594));
  INV_X1    g0394(.A(new_n474), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n203), .B(G45), .C1(new_n255), .C2(KEYINPUT5), .ZN(new_n596));
  OAI211_X1 g0396(.A(G264), .B(new_n264), .C1(new_n595), .C2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT85), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n477), .A2(KEYINPUT85), .A3(G264), .A4(new_n264), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n594), .A2(new_n479), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(G169), .ZN(new_n603));
  AOI22_X1  g0403(.A1(new_n593), .A2(new_n320), .B1(new_n599), .B2(new_n600), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n604), .A2(G179), .A3(new_n479), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n585), .A2(new_n606), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n512), .B1(new_n203), .B2(G33), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n334), .A2(new_n336), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n288), .A2(new_n512), .ZN(new_n610));
  AOI22_X1  g0410(.A1(new_n289), .A2(new_n223), .B1(G20), .B2(new_n512), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n499), .B(new_n204), .C1(G33), .C2(new_n436), .ZN(new_n612));
  AOI21_X1  g0412(.A(KEYINPUT20), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  AND3_X1   g0413(.A1(new_n611), .A2(KEYINPUT20), .A3(new_n612), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n609), .B(new_n610), .C1(new_n613), .C2(new_n614), .ZN(new_n615));
  OAI211_X1 g0415(.A(G270), .B(new_n264), .C1(new_n595), .C2(new_n596), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n260), .A2(G257), .ZN(new_n617));
  NAND2_X1  g0417(.A1(G264), .A2(G1698), .ZN(new_n618));
  AND3_X1   g0418(.A1(new_n259), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n320), .B1(new_n259), .B2(G303), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n479), .B(new_n616), .C1(new_n619), .C2(new_n620), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n615), .A2(KEYINPUT21), .A3(G169), .A4(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT21), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n610), .B1(new_n614), .B2(new_n613), .ZN(new_n624));
  AND3_X1   g0424(.A1(new_n334), .A2(new_n336), .A3(new_n608), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n621), .A2(G169), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n623), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n621), .A2(new_n311), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(new_n615), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n621), .A2(G200), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n259), .A2(new_n617), .A3(new_n618), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n632), .B(new_n320), .C1(G303), .C2(new_n259), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n633), .A2(G190), .A3(new_n479), .A4(new_n616), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n626), .A2(new_n631), .A3(new_n634), .ZN(new_n635));
  AND4_X1   g0435(.A1(new_n622), .A2(new_n628), .A3(new_n630), .A4(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n565), .ZN(new_n637));
  AND3_X1   g0437(.A1(new_n573), .A2(new_n582), .A3(new_n578), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n582), .B1(new_n573), .B2(new_n578), .ZN(new_n639));
  OAI22_X1  g0439(.A1(new_n638), .A2(new_n639), .B1(new_n566), .B2(new_n567), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n637), .B1(new_n640), .B2(new_n290), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n602), .A2(new_n245), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n604), .A2(new_n341), .A3(new_n479), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n607), .A2(new_n636), .A3(new_n645), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n560), .A2(new_n646), .ZN(new_n647));
  AND2_X1   g0447(.A1(new_n455), .A2(new_n647), .ZN(G372));
  INV_X1    g0448(.A(new_n314), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n453), .A2(new_n339), .A3(new_n325), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n402), .B1(new_n650), .B2(new_n450), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n415), .A2(new_n409), .ZN(new_n652));
  OR2_X1    g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  AND2_X1   g0453(.A1(new_n309), .A2(new_n310), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n649), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n455), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT26), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n559), .A2(new_n657), .ZN(new_n658));
  AOI22_X1  g0458(.A1(new_n495), .A2(new_n505), .B1(new_n641), .B2(new_n644), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n628), .A2(new_n630), .ZN(new_n660));
  AND2_X1   g0460(.A1(new_n603), .A2(new_n605), .ZN(new_n661));
  OAI211_X1 g0461(.A(new_n660), .B(new_n622), .C1(new_n661), .C2(new_n641), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n658), .B1(new_n663), .B2(new_n511), .ZN(new_n664));
  NOR3_X1   g0464(.A1(new_n471), .A2(new_n509), .A3(new_n510), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n552), .A2(new_n665), .A3(new_n559), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(KEYINPUT26), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n554), .A2(new_n555), .ZN(new_n668));
  AOI22_X1  g0468(.A1(new_n668), .A2(new_n533), .B1(new_n529), .B2(new_n324), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(new_n527), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n664), .A2(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n655), .B1(new_n656), .B2(new_n672), .ZN(G369));
  NAND3_X1  g0473(.A1(new_n203), .A2(new_n204), .A3(G13), .ZN(new_n674));
  OR2_X1    g0474(.A1(new_n674), .A2(KEYINPUT27), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(KEYINPUT27), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n675), .A2(G213), .A3(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(G343), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n585), .A2(new_n606), .A3(new_n679), .ZN(new_n680));
  XNOR2_X1  g0480(.A(new_n680), .B(KEYINPUT87), .ZN(new_n681));
  INV_X1    g0481(.A(new_n679), .ZN(new_n682));
  OAI211_X1 g0482(.A(new_n607), .B(new_n645), .C1(new_n641), .C2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n660), .A2(new_n622), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n626), .A2(new_n682), .ZN(new_n687));
  MUX2_X1   g0487(.A(new_n636), .B(new_n686), .S(new_n687), .Z(new_n688));
  XOR2_X1   g0488(.A(KEYINPUT86), .B(G330), .Z(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n685), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n686), .A2(new_n682), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n694), .B1(new_n681), .B2(new_n683), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n607), .A2(new_n679), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n693), .A2(new_n697), .ZN(G399));
  NAND2_X1  g0498(.A1(new_n207), .A2(new_n255), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n537), .A2(G116), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n699), .A2(G1), .A3(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n226), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n701), .B1(new_n702), .B2(new_n699), .ZN(new_n703));
  XNOR2_X1  g0503(.A(new_n703), .B(KEYINPUT28), .ZN(new_n704));
  AND3_X1   g0504(.A1(new_n607), .A2(new_n636), .A3(new_n645), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n665), .B1(new_n505), .B2(new_n495), .ZN(new_n706));
  AND3_X1   g0506(.A1(new_n549), .A2(new_n550), .A3(new_n311), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n550), .B1(new_n549), .B2(new_n311), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n549), .A2(new_n245), .ZN(new_n710));
  AOI211_X1 g0510(.A(new_n341), .B(new_n548), .C1(new_n522), .C2(new_n320), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  AOI22_X1  g0512(.A1(new_n709), .A2(new_n669), .B1(new_n556), .B2(new_n712), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n705), .A2(new_n706), .A3(new_n713), .A4(new_n682), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(KEYINPUT88), .ZN(new_n715));
  INV_X1    g0515(.A(new_n560), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT88), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n716), .A2(new_n717), .A3(new_n705), .A4(new_n682), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n715), .A2(new_n718), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n549), .A2(new_n493), .A3(new_n604), .A4(new_n629), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT30), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  AND2_X1   g0522(.A1(new_n629), .A2(new_n604), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n723), .A2(KEYINPUT30), .A3(new_n493), .A4(new_n549), .ZN(new_n724));
  INV_X1    g0524(.A(new_n493), .ZN(new_n725));
  AND2_X1   g0525(.A1(new_n621), .A2(new_n311), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n725), .A2(new_n529), .A3(new_n602), .A4(new_n726), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n722), .A2(new_n724), .A3(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(new_n679), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT31), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n728), .A2(KEYINPUT31), .A3(new_n679), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n689), .B1(new_n719), .B2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n670), .A2(new_n559), .ZN(new_n737));
  NOR3_X1   g0537(.A1(new_n663), .A2(new_n665), .A3(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n559), .ZN(new_n739));
  OAI21_X1  g0539(.A(KEYINPUT26), .B1(new_n739), .B2(new_n511), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n552), .A2(new_n559), .A3(new_n665), .A4(new_n657), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n740), .A2(new_n670), .A3(new_n741), .ZN(new_n742));
  OAI211_X1 g0542(.A(KEYINPUT29), .B(new_n682), .C1(new_n738), .C2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n672), .A2(new_n679), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n743), .B1(new_n744), .B2(KEYINPUT29), .ZN(new_n745));
  AND2_X1   g0545(.A1(new_n736), .A2(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n704), .B1(new_n746), .B2(G1), .ZN(G364));
  INV_X1    g0547(.A(new_n691), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n204), .A2(G13), .A3(G45), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n699), .A2(G1), .A3(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT89), .ZN(new_n751));
  OR2_X1    g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n750), .A2(new_n751), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n748), .A2(new_n755), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n756), .B1(new_n690), .B2(new_n688), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n207), .A2(new_n259), .ZN(new_n758));
  INV_X1    g0558(.A(G355), .ZN(new_n759));
  OAI22_X1  g0559(.A1(new_n758), .A2(new_n759), .B1(G116), .B2(new_n207), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n227), .A2(new_n256), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n207), .A2(new_n269), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n762), .B1(new_n240), .B2(G45), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n760), .B1(new_n761), .B2(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(G13), .A2(G33), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(G20), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n223), .B1(G20), .B2(new_n324), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n755), .B1(new_n764), .B2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n204), .A2(new_n311), .ZN(new_n772));
  NOR2_X1   g0572(.A1(G190), .A2(G200), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n772), .ZN(new_n775));
  NOR3_X1   g0575(.A1(new_n775), .A2(new_n341), .A3(G200), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(G58), .ZN(new_n778));
  OAI221_X1 g0578(.A(new_n259), .B1(new_n211), .B2(new_n774), .C1(new_n777), .C2(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n204), .A2(G179), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n780), .A2(new_n341), .A3(G200), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(new_n467), .ZN(new_n782));
  NOR3_X1   g0582(.A1(new_n341), .A2(G179), .A3(G200), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(new_n204), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n784), .A2(new_n436), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n780), .A2(G190), .A3(G200), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(new_n213), .ZN(new_n787));
  NOR4_X1   g0587(.A1(new_n779), .A2(new_n782), .A3(new_n785), .A4(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n772), .A2(G200), .ZN(new_n789));
  XNOR2_X1  g0589(.A(new_n789), .B(KEYINPUT90), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(new_n341), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n790), .A2(G190), .ZN(new_n792));
  AOI22_X1  g0592(.A1(G50), .A2(new_n791), .B1(new_n792), .B2(G68), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n780), .A2(new_n773), .ZN(new_n794));
  INV_X1    g0594(.A(G159), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  XNOR2_X1  g0596(.A(new_n796), .B(KEYINPUT91), .ZN(new_n797));
  XNOR2_X1  g0597(.A(new_n797), .B(KEYINPUT32), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n788), .A2(new_n793), .A3(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n774), .ZN(new_n800));
  AOI22_X1  g0600(.A1(new_n776), .A2(G322), .B1(G311), .B2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n794), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(G329), .ZN(new_n803));
  INV_X1    g0603(.A(G283), .ZN(new_n804));
  OAI211_X1 g0604(.A(new_n801), .B(new_n803), .C1(new_n804), .C2(new_n781), .ZN(new_n805));
  INV_X1    g0605(.A(new_n786), .ZN(new_n806));
  AOI211_X1 g0606(.A(new_n259), .B(new_n805), .C1(G303), .C2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n792), .ZN(new_n808));
  XOR2_X1   g0608(.A(KEYINPUT33), .B(G317), .Z(new_n809));
  OAI21_X1  g0609(.A(new_n807), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n784), .ZN(new_n811));
  AOI22_X1  g0611(.A1(new_n791), .A2(G326), .B1(G294), .B2(new_n811), .ZN(new_n812));
  XOR2_X1   g0612(.A(new_n812), .B(KEYINPUT92), .Z(new_n813));
  OAI21_X1  g0613(.A(new_n799), .B1(new_n810), .B2(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n771), .B1(new_n814), .B2(new_n768), .ZN(new_n815));
  INV_X1    g0615(.A(new_n767), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n815), .B1(new_n688), .B2(new_n816), .ZN(new_n817));
  AND2_X1   g0617(.A1(new_n757), .A2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(G396));
  INV_X1    g0619(.A(new_n345), .ZN(new_n820));
  OAI211_X1 g0620(.A(new_n820), .B(new_n682), .C1(new_n664), .C2(new_n671), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n340), .A2(new_n679), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n339), .A2(new_n679), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(new_n344), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n822), .B1(new_n340), .B2(new_n824), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n821), .B1(new_n744), .B2(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n755), .B1(new_n736), .B2(new_n826), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n827), .B1(new_n736), .B2(new_n826), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n768), .A2(new_n765), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n754), .B1(new_n211), .B2(new_n829), .ZN(new_n830));
  XNOR2_X1  g0630(.A(new_n830), .B(KEYINPUT93), .ZN(new_n831));
  AOI22_X1  g0631(.A1(new_n776), .A2(G143), .B1(G159), .B2(new_n800), .ZN(new_n832));
  INV_X1    g0632(.A(new_n791), .ZN(new_n833));
  INV_X1    g0633(.A(G137), .ZN(new_n834));
  OAI221_X1 g0634(.A(new_n832), .B1(new_n833), .B2(new_n834), .C1(new_n297), .C2(new_n808), .ZN(new_n835));
  XOR2_X1   g0635(.A(new_n835), .B(KEYINPUT34), .Z(new_n836));
  AOI22_X1  g0636(.A1(new_n811), .A2(G58), .B1(new_n806), .B2(G50), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n269), .B1(new_n802), .B2(G132), .ZN(new_n838));
  OAI211_X1 g0638(.A(new_n837), .B(new_n838), .C1(new_n302), .C2(new_n781), .ZN(new_n839));
  INV_X1    g0639(.A(G311), .ZN(new_n840));
  OAI22_X1  g0640(.A1(new_n774), .A2(new_n512), .B1(new_n794), .B2(new_n840), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n841), .B1(G294), .B2(new_n776), .ZN(new_n842));
  INV_X1    g0642(.A(new_n781), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n785), .B1(G87), .B2(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n259), .B1(new_n806), .B2(G107), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n842), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n791), .A2(G303), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n847), .B1(new_n808), .B2(new_n804), .ZN(new_n848));
  OAI22_X1  g0648(.A1(new_n836), .A2(new_n839), .B1(new_n846), .B2(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n831), .B1(new_n849), .B2(new_n768), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n850), .B1(new_n825), .B2(new_n766), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n828), .A2(new_n851), .ZN(G384));
  OR2_X1    g0652(.A1(new_n462), .A2(new_n464), .ZN(new_n853));
  OR2_X1    g0653(.A1(new_n853), .A2(KEYINPUT35), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n853), .A2(KEYINPUT35), .ZN(new_n855));
  NAND4_X1  g0655(.A1(new_n854), .A2(G116), .A3(new_n224), .A4(new_n855), .ZN(new_n856));
  XOR2_X1   g0656(.A(new_n856), .B(KEYINPUT36), .Z(new_n857));
  OAI211_X1 g0657(.A(new_n226), .B(G77), .C1(new_n778), .C2(new_n302), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n292), .A2(G68), .ZN(new_n859));
  AOI211_X1 g0659(.A(new_n203), .B(G13), .C1(new_n858), .C2(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT38), .ZN(new_n862));
  OR2_X1    g0662(.A1(new_n361), .A2(KEYINPUT16), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n352), .B1(new_n863), .B2(new_n362), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n677), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n410), .A2(new_n418), .ZN(new_n868));
  INV_X1    g0668(.A(new_n393), .ZN(new_n869));
  INV_X1    g0669(.A(new_n401), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n867), .B1(new_n868), .B2(new_n871), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n392), .A2(new_n399), .A3(new_n400), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n873), .B1(new_n864), .B2(new_n677), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n864), .A2(new_n414), .ZN(new_n875));
  OAI21_X1  g0675(.A(KEYINPUT37), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n403), .A2(new_n407), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n403), .A2(new_n866), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT37), .ZN(new_n879));
  NAND4_X1  g0679(.A1(new_n877), .A2(new_n878), .A3(new_n879), .A4(new_n873), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n876), .A2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n862), .B1(new_n872), .B2(new_n882), .ZN(new_n883));
  OAI211_X1 g0683(.A(KEYINPUT38), .B(new_n881), .C1(new_n419), .C2(new_n867), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n717), .B1(new_n647), .B2(new_n682), .ZN(new_n886));
  NOR4_X1   g0686(.A1(new_n560), .A2(new_n646), .A3(KEYINPUT88), .A4(new_n679), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n734), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  OR2_X1    g0688(.A1(new_n445), .A2(new_n449), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n889), .A2(new_n432), .A3(new_n679), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n432), .A2(new_n679), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n450), .A2(new_n453), .A3(new_n891), .ZN(new_n892));
  AND2_X1   g0692(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(new_n825), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n885), .A2(new_n888), .A3(new_n895), .ZN(new_n896));
  XNOR2_X1  g0696(.A(KEYINPUT96), .B(KEYINPUT40), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(KEYINPUT97), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT97), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n896), .A2(new_n900), .A3(new_n897), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n733), .B1(new_n715), .B2(new_n718), .ZN(new_n903));
  NOR3_X1   g0703(.A1(new_n903), .A2(new_n894), .A3(new_n893), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT40), .ZN(new_n905));
  AOI22_X1  g0705(.A1(new_n869), .A2(new_n870), .B1(new_n416), .B2(new_n408), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n877), .A2(new_n878), .A3(new_n873), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(KEYINPUT37), .ZN(new_n908));
  OAI22_X1  g0708(.A1(new_n906), .A2(new_n878), .B1(new_n908), .B2(KEYINPUT95), .ZN(new_n909));
  AND3_X1   g0709(.A1(new_n908), .A2(KEYINPUT95), .A3(new_n880), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n862), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n905), .B1(new_n911), .B2(new_n884), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n904), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n902), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n455), .A2(new_n888), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n690), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n916), .B1(new_n914), .B2(new_n915), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n822), .B(KEYINPUT94), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n893), .B1(new_n821), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(new_n885), .ZN(new_n920));
  INV_X1    g0720(.A(new_n652), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n920), .B1(new_n921), .B2(new_n866), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n889), .A2(new_n432), .A3(new_n682), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n415), .B1(new_n417), .B2(new_n416), .ZN(new_n924));
  NOR3_X1   g0724(.A1(new_n877), .A2(KEYINPUT75), .A3(new_n411), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n871), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n867), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(KEYINPUT38), .B1(new_n928), .B2(new_n881), .ZN(new_n929));
  INV_X1    g0729(.A(new_n884), .ZN(new_n930));
  OAI21_X1  g0730(.A(KEYINPUT39), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT39), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n911), .A2(new_n932), .A3(new_n884), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n923), .B1(new_n931), .B2(new_n933), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n922), .A2(new_n934), .ZN(new_n935));
  OAI211_X1 g0735(.A(new_n455), .B(new_n743), .C1(new_n744), .C2(KEYINPUT29), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(new_n655), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n935), .B(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n917), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(G1), .B1(new_n425), .B2(G20), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n939), .A2(KEYINPUT98), .A3(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n941), .B1(new_n938), .B2(new_n917), .ZN(new_n942));
  AOI21_X1  g0742(.A(KEYINPUT98), .B1(new_n939), .B2(new_n940), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n861), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  XOR2_X1   g0744(.A(new_n944), .B(KEYINPUT99), .Z(G367));
  OAI21_X1  g0745(.A(new_n706), .B1(new_n471), .B2(new_n682), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n665), .A2(new_n679), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n692), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n949), .A2(KEYINPUT102), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n556), .A2(new_n682), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n952), .A2(new_n669), .A3(new_n527), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n953), .B1(new_n737), .B2(new_n952), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n954), .A2(KEYINPUT43), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n955), .A2(KEYINPUT101), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n949), .A2(KEYINPUT102), .ZN(new_n957));
  OR3_X1    g0757(.A1(new_n951), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n956), .B1(new_n951), .B2(new_n957), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n695), .A2(new_n948), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(KEYINPUT42), .ZN(new_n962));
  OR2_X1    g0762(.A1(new_n946), .A2(new_n607), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n679), .B1(new_n963), .B2(new_n511), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  AND2_X1   g0765(.A1(new_n955), .A2(KEYINPUT101), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n954), .A2(KEYINPUT43), .ZN(new_n967));
  XOR2_X1   g0767(.A(new_n967), .B(KEYINPUT100), .Z(new_n968));
  NOR3_X1   g0768(.A1(new_n965), .A2(new_n966), .A3(new_n968), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n960), .B(new_n969), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n699), .B(KEYINPUT41), .ZN(new_n971));
  INV_X1    g0771(.A(new_n697), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT45), .ZN(new_n973));
  INV_X1    g0773(.A(new_n948), .ZN(new_n974));
  NOR3_X1   g0774(.A1(new_n972), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  AOI21_X1  g0775(.A(KEYINPUT45), .B1(new_n697), .B2(new_n948), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  OR3_X1    g0777(.A1(new_n697), .A2(KEYINPUT44), .A3(new_n948), .ZN(new_n978));
  OAI21_X1  g0778(.A(KEYINPUT44), .B1(new_n697), .B2(new_n948), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  OR3_X1    g0780(.A1(new_n977), .A2(new_n980), .A3(new_n692), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n692), .B1(new_n977), .B2(new_n980), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n685), .A2(new_n694), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n691), .B1(new_n984), .B2(new_n695), .ZN(new_n985));
  INV_X1    g0785(.A(new_n695), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n983), .A2(new_n748), .A3(new_n986), .ZN(new_n987));
  AND2_X1   g0787(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n988), .A2(new_n746), .ZN(new_n989));
  INV_X1    g0789(.A(new_n989), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n981), .A2(new_n982), .A3(new_n990), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n971), .B1(new_n991), .B2(new_n746), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n749), .A2(G1), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n970), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(new_n236), .ZN(new_n995));
  OAI221_X1 g0795(.A(new_n769), .B1(new_n207), .B2(new_n326), .C1(new_n995), .C2(new_n762), .ZN(new_n996));
  AND2_X1   g0796(.A1(new_n755), .A2(new_n996), .ZN(new_n997));
  AOI22_X1  g0797(.A1(G143), .A2(new_n791), .B1(new_n792), .B2(G159), .ZN(new_n998));
  OAI22_X1  g0798(.A1(new_n774), .A2(new_n292), .B1(new_n794), .B2(new_n834), .ZN(new_n999));
  AOI211_X1 g0799(.A(new_n269), .B(new_n999), .C1(G150), .C2(new_n776), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n786), .A2(new_n778), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n781), .A2(new_n211), .ZN(new_n1002));
  AOI211_X1 g0802(.A(new_n1001), .B(new_n1002), .C1(G68), .C2(new_n811), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n998), .A2(new_n1000), .A3(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n806), .A2(G116), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1005), .B(KEYINPUT46), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n259), .B1(new_n776), .B2(G303), .ZN(new_n1007));
  XOR2_X1   g0807(.A(KEYINPUT103), .B(G317), .Z(new_n1008));
  INV_X1    g0808(.A(new_n1008), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(new_n802), .A2(new_n1009), .B1(new_n800), .B2(G283), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(new_n811), .A2(G107), .B1(new_n843), .B2(G97), .ZN(new_n1011));
  NAND4_X1  g0811(.A1(new_n1006), .A2(new_n1007), .A3(new_n1010), .A4(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(G294), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n1013), .A2(new_n808), .B1(new_n833), .B2(new_n840), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1004), .B1(new_n1012), .B2(new_n1014), .ZN(new_n1015));
  XOR2_X1   g0815(.A(new_n1015), .B(KEYINPUT47), .Z(new_n1016));
  INV_X1    g0816(.A(new_n768), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n997), .B1(new_n954), .B2(new_n816), .C1(new_n1016), .C2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n994), .A2(new_n1018), .ZN(G387));
  OAI22_X1  g0819(.A1(new_n758), .A2(new_n700), .B1(G107), .B2(new_n207), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n233), .A2(G45), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n700), .ZN(new_n1022));
  AOI211_X1 g0822(.A(G45), .B(new_n1022), .C1(G68), .C2(G77), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n295), .A2(G50), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1024), .B(KEYINPUT50), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n762), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1020), .B1(new_n1021), .B2(new_n1026), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n755), .B1(new_n770), .B2(new_n1027), .C1(new_n684), .C2(new_n816), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n792), .A2(new_n349), .B1(G68), .B2(new_n800), .ZN(new_n1029));
  XOR2_X1   g0829(.A(new_n1029), .B(KEYINPUT105), .Z(new_n1030));
  AOI21_X1  g0830(.A(new_n269), .B1(new_n802), .B2(G150), .ZN(new_n1031));
  OAI221_X1 g0831(.A(new_n1031), .B1(new_n211), .B2(new_n786), .C1(new_n436), .C2(new_n781), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1032), .B(KEYINPUT104), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n784), .A2(new_n326), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n777), .A2(new_n292), .ZN(new_n1035));
  AOI211_X1 g0835(.A(new_n1034), .B(new_n1035), .C1(new_n791), .C2(G159), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1030), .A2(new_n1033), .A3(new_n1036), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n784), .A2(new_n804), .B1(new_n786), .B2(new_n1013), .ZN(new_n1038));
  OR2_X1    g0838(.A1(new_n1038), .A2(KEYINPUT106), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1038), .A2(KEYINPUT106), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n776), .A2(new_n1009), .B1(new_n800), .B2(G303), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1041), .B1(new_n808), .B2(new_n840), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(KEYINPUT107), .B(G322), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n1043), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1042), .B1(new_n791), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT48), .ZN(new_n1047));
  OAI211_X1 g0847(.A(new_n1039), .B(new_n1040), .C1(new_n1046), .C2(new_n1047), .ZN(new_n1048));
  XOR2_X1   g0848(.A(new_n1048), .B(KEYINPUT108), .Z(new_n1049));
  NAND2_X1  g0849(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1049), .A2(KEYINPUT49), .A3(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n259), .B1(new_n802), .B2(G326), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1052), .B1(new_n512), .B2(new_n781), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(KEYINPUT109), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1051), .A2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g0855(.A(KEYINPUT49), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1037), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1028), .B1(new_n1057), .B2(new_n768), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(new_n993), .B2(new_n988), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n699), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n989), .A2(new_n1060), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n988), .A2(new_n746), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1059), .B1(new_n1061), .B2(new_n1062), .ZN(G393));
  NAND3_X1  g0863(.A1(new_n981), .A2(new_n982), .A3(new_n993), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n769), .B1(new_n436), .B2(new_n207), .C1(new_n243), .C2(new_n762), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n791), .A2(G150), .B1(G159), .B2(new_n776), .ZN(new_n1066));
  XOR2_X1   g0866(.A(new_n1066), .B(KEYINPUT51), .Z(new_n1067));
  NOR2_X1   g0867(.A1(new_n808), .A2(new_n292), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n806), .A2(G68), .B1(new_n802), .B2(G143), .ZN(new_n1069));
  XOR2_X1   g0869(.A(new_n1069), .B(KEYINPUT110), .Z(new_n1070));
  NOR2_X1   g0870(.A1(new_n784), .A2(new_n211), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n259), .B1(new_n774), .B2(new_n295), .C1(new_n213), .C2(new_n781), .ZN(new_n1072));
  NOR4_X1   g0872(.A1(new_n1068), .A2(new_n1070), .A3(new_n1071), .A4(new_n1072), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n791), .A2(G317), .B1(G311), .B2(new_n776), .ZN(new_n1074));
  XOR2_X1   g0874(.A(new_n1074), .B(KEYINPUT52), .Z(new_n1075));
  OAI221_X1 g0875(.A(new_n269), .B1(new_n794), .B2(new_n1043), .C1(new_n1013), .C2(new_n774), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n782), .B1(G116), .B2(new_n811), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1077), .B1(new_n804), .B2(new_n786), .ZN(new_n1078));
  AOI211_X1 g0878(.A(new_n1076), .B(new_n1078), .C1(G303), .C2(new_n792), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n1067), .A2(new_n1073), .B1(new_n1075), .B2(new_n1079), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n755), .B(new_n1065), .C1(new_n1080), .C2(new_n1017), .ZN(new_n1081));
  XOR2_X1   g0881(.A(new_n1081), .B(KEYINPUT111), .Z(new_n1082));
  OAI21_X1  g0882(.A(new_n1082), .B1(new_n816), .B2(new_n948), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1064), .A2(new_n1083), .ZN(new_n1084));
  AND2_X1   g0884(.A1(new_n991), .A2(new_n1060), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n981), .A2(new_n982), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1086), .A2(new_n989), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1084), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1088), .ZN(G390));
  INV_X1    g0889(.A(new_n923), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n931), .B(new_n933), .C1(new_n1090), .C2(new_n919), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1090), .B1(new_n911), .B2(new_n884), .ZN(new_n1092));
  OAI211_X1 g0892(.A(new_n682), .B(new_n825), .C1(new_n738), .C2(new_n742), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1093), .A2(new_n918), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1094), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1092), .B1(new_n1095), .B2(new_n893), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n893), .ZN(new_n1097));
  NAND4_X1  g0897(.A1(new_n888), .A2(new_n690), .A3(new_n825), .A4(new_n1097), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1091), .A2(new_n1096), .A3(new_n1098), .ZN(new_n1099));
  AND2_X1   g0899(.A1(new_n1091), .A2(new_n1096), .ZN(new_n1100));
  INV_X1    g0900(.A(G330), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(new_n719), .B2(new_n734), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1102), .A2(new_n895), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n993), .B(new_n1099), .C1(new_n1100), .C2(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(KEYINPUT116), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n791), .A2(G128), .B1(G132), .B2(new_n776), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(new_n1106), .B(KEYINPUT113), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n786), .A2(new_n297), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(new_n1108), .B(KEYINPUT53), .ZN(new_n1109));
  INV_X1    g0909(.A(G125), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(KEYINPUT54), .B(G143), .ZN(new_n1111));
  OAI221_X1 g0911(.A(new_n259), .B1(new_n794), .B2(new_n1110), .C1(new_n774), .C2(new_n1111), .ZN(new_n1112));
  OAI22_X1  g0912(.A1(new_n784), .A2(new_n795), .B1(new_n781), .B2(new_n292), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n1109), .B(new_n1114), .C1(new_n808), .C2(new_n834), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n269), .B1(new_n774), .B2(new_n436), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1116), .B1(G294), .B2(new_n802), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n787), .B1(G68), .B2(new_n843), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n1117), .B(new_n1118), .C1(new_n808), .C2(new_n467), .ZN(new_n1119));
  OAI22_X1  g0919(.A1(new_n777), .A2(new_n512), .B1(new_n211), .B2(new_n784), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(G283), .A2(new_n791), .B1(new_n1120), .B2(KEYINPUT114), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1121), .B1(KEYINPUT114), .B2(new_n1120), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n1107), .A2(new_n1115), .B1(new_n1119), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1123), .A2(new_n768), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n829), .ZN(new_n1125));
  OAI211_X1 g0925(.A(new_n1124), .B(new_n755), .C1(new_n349), .C2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n931), .A2(new_n933), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1127), .B1(new_n1128), .B2(new_n766), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1129), .A2(KEYINPUT115), .ZN(new_n1130));
  INV_X1    g0930(.A(KEYINPUT115), .ZN(new_n1131));
  OAI211_X1 g0931(.A(new_n1131), .B(new_n1127), .C1(new_n1128), .C2(new_n766), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1133));
  AND3_X1   g0933(.A1(new_n1104), .A2(new_n1105), .A3(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1105), .B1(new_n1104), .B2(new_n1133), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  AND3_X1   g0936(.A1(new_n1091), .A2(new_n1096), .A3(new_n1098), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1103), .B1(new_n1091), .B2(new_n1096), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1102), .A2(new_n455), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n936), .A2(new_n655), .A3(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n821), .A2(new_n918), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1097), .B1(new_n735), .B2(new_n825), .ZN(new_n1143));
  AND3_X1   g0943(.A1(new_n888), .A2(new_n895), .A3(G330), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1142), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  NOR3_X1   g0945(.A1(new_n903), .A2(new_n1101), .A3(new_n894), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n1098), .B(new_n1095), .C1(new_n1146), .C2(new_n1097), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1141), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1139), .A2(new_n1148), .ZN(new_n1149));
  NOR3_X1   g0949(.A1(new_n903), .A2(new_n689), .A3(new_n894), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1103), .B1(new_n1150), .B2(new_n1097), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1094), .B1(new_n1150), .B2(new_n1097), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1102), .A2(new_n825), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(new_n893), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n1142), .A2(new_n1151), .B1(new_n1152), .B2(new_n1154), .ZN(new_n1155));
  OAI22_X1  g0955(.A1(new_n1155), .A2(new_n1141), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1149), .A2(new_n1060), .A3(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(KEYINPUT112), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n1149), .A2(new_n1156), .A3(KEYINPUT112), .A4(new_n1060), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1136), .A2(new_n1159), .A3(new_n1160), .ZN(G378));
  INV_X1    g0961(.A(new_n935), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(new_n315), .B(KEYINPUT118), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(new_n1164), .B(KEYINPUT119), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n1163), .A2(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1163), .A2(new_n1165), .ZN(new_n1168));
  NAND4_X1  g0968(.A1(new_n1167), .A2(new_n313), .A3(new_n866), .A4(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n313), .A2(new_n866), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1168), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1170), .B1(new_n1171), .B2(new_n1166), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1169), .A2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1101), .B1(new_n904), .B2(new_n912), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1173), .B1(new_n902), .B2(new_n1174), .ZN(new_n1175));
  AND3_X1   g0975(.A1(new_n896), .A2(new_n900), .A3(new_n897), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n900), .B1(new_n896), .B2(new_n897), .ZN(new_n1177));
  OAI211_X1 g0977(.A(new_n1174), .B(new_n1173), .C1(new_n1176), .C2(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1162), .B1(new_n1175), .B2(new_n1179), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1174), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1173), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1183), .A2(new_n935), .A3(new_n1178), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1180), .A2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1182), .A2(new_n765), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n755), .B1(G50), .B2(new_n1125), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(G33), .A2(G41), .ZN(new_n1188));
  AOI211_X1 g0988(.A(G50), .B(new_n1188), .C1(new_n269), .C2(new_n255), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n781), .A2(new_n778), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  OAI221_X1 g0991(.A(new_n1191), .B1(new_n302), .B2(new_n784), .C1(new_n211), .C2(new_n786), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n777), .A2(new_n467), .B1(new_n794), .B2(new_n804), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n255), .B(new_n269), .C1(new_n774), .C2(new_n326), .ZN(new_n1194));
  NOR3_X1   g0994(.A1(new_n1192), .A2(new_n1193), .A3(new_n1194), .ZN(new_n1195));
  OAI221_X1 g0995(.A(new_n1195), .B1(new_n436), .B2(new_n808), .C1(new_n512), .C2(new_n833), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT58), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1189), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n784), .A2(new_n297), .ZN(new_n1199));
  INV_X1    g0999(.A(G128), .ZN(new_n1200));
  OAI22_X1  g1000(.A1(new_n777), .A2(new_n1200), .B1(new_n774), .B2(new_n834), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1111), .ZN(new_n1202));
  AOI211_X1 g1002(.A(new_n1199), .B(new_n1201), .C1(new_n806), .C2(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(G132), .ZN(new_n1204));
  OAI221_X1 g1004(.A(new_n1203), .B1(new_n1110), .B2(new_n833), .C1(new_n1204), .C2(new_n808), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1205), .A2(KEYINPUT59), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1188), .ZN(new_n1207));
  XNOR2_X1  g1007(.A(KEYINPUT117), .B(G124), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1207), .B1(new_n802), .B2(new_n1208), .ZN(new_n1209));
  OAI211_X1 g1009(.A(new_n1206), .B(new_n1209), .C1(new_n795), .C2(new_n781), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n1205), .A2(KEYINPUT59), .ZN(new_n1211));
  OAI221_X1 g1011(.A(new_n1198), .B1(new_n1197), .B2(new_n1196), .C1(new_n1210), .C2(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1187), .B1(new_n1212), .B2(new_n768), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n1185), .A2(new_n993), .B1(new_n1186), .B2(new_n1213), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n888), .A2(new_n690), .A3(new_n825), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n1215), .A2(new_n893), .B1(new_n1102), .B2(new_n895), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1142), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1147), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1141), .B1(new_n1139), .B2(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1219), .B1(new_n1180), .B2(new_n1184), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1060), .B1(new_n1220), .B2(KEYINPUT57), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1141), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1149), .A2(new_n1222), .ZN(new_n1223));
  AND3_X1   g1023(.A1(new_n1183), .A2(new_n935), .A3(new_n1178), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n935), .B1(new_n1183), .B2(new_n1178), .ZN(new_n1225));
  OAI211_X1 g1025(.A(new_n1223), .B(KEYINPUT57), .C1(new_n1224), .C2(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1226), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1214), .B1(new_n1221), .B2(new_n1227), .ZN(G375));
  NOR2_X1   g1028(.A1(new_n1148), .A2(new_n971), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1145), .A2(new_n1141), .A3(new_n1147), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  OAI221_X1 g1031(.A(new_n259), .B1(new_n794), .B2(new_n1200), .C1(new_n297), .C2(new_n774), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1191), .B1(new_n292), .B2(new_n784), .ZN(new_n1233));
  AOI211_X1 g1033(.A(new_n1232), .B(new_n1233), .C1(G159), .C2(new_n806), .ZN(new_n1234));
  OR2_X1    g1034(.A1(new_n1234), .A2(KEYINPUT120), .ZN(new_n1235));
  OAI22_X1  g1035(.A1(new_n833), .A2(new_n1204), .B1(new_n834), .B2(new_n777), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1236), .B1(new_n792), .B2(new_n1202), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1234), .A2(KEYINPUT120), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1235), .A2(new_n1237), .A3(new_n1238), .ZN(new_n1239));
  AOI22_X1  g1039(.A1(G116), .A2(new_n792), .B1(new_n791), .B2(G294), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n259), .B1(new_n802), .B2(G303), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(new_n776), .A2(G283), .B1(G107), .B2(new_n800), .ZN(new_n1242));
  AOI211_X1 g1042(.A(new_n1002), .B(new_n1034), .C1(G97), .C2(new_n806), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1240), .A2(new_n1241), .A3(new_n1242), .A4(new_n1243), .ZN(new_n1244));
  AND2_X1   g1044(.A1(new_n1239), .A2(new_n1244), .ZN(new_n1245));
  OR2_X1    g1045(.A1(new_n1245), .A2(KEYINPUT121), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1245), .A2(KEYINPUT121), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1246), .A2(new_n768), .A3(new_n1247), .ZN(new_n1248));
  OAI211_X1 g1048(.A(new_n1248), .B(new_n755), .C1(G68), .C2(new_n1125), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1249), .B1(new_n893), .B2(new_n765), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1250), .B1(new_n1218), .B2(new_n993), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1231), .A2(new_n1251), .ZN(G381));
  INV_X1    g1052(.A(G375), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1088), .A2(new_n994), .A3(new_n1018), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  AND3_X1   g1055(.A1(new_n1157), .A2(new_n1133), .A3(new_n1104), .ZN(new_n1256));
  NOR4_X1   g1056(.A1(G381), .A2(G393), .A3(G396), .A4(G384), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1253), .A2(new_n1255), .A3(new_n1256), .A4(new_n1257), .ZN(G407));
  NAND2_X1  g1058(.A1(new_n678), .A2(G213), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1253), .A2(new_n1256), .A3(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(G407), .A2(new_n1261), .A3(G213), .ZN(G409));
  OAI211_X1 g1062(.A(G378), .B(new_n1214), .C1(new_n1221), .C2(new_n1227), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n993), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1186), .A2(new_n1213), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1223), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1266));
  OAI211_X1 g1066(.A(new_n1264), .B(new_n1265), .C1(new_n1266), .C2(new_n971), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1267), .A2(new_n1256), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1260), .B1(new_n1263), .B2(new_n1268), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1155), .A2(KEYINPUT122), .A3(KEYINPUT60), .A4(new_n1141), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1145), .A2(KEYINPUT60), .A3(new_n1141), .A4(new_n1147), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT122), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT60), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1230), .A2(new_n1274), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n699), .B1(new_n1218), .B2(new_n1222), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1270), .A2(new_n1273), .A3(new_n1275), .A4(new_n1276), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1277), .A2(G384), .A3(new_n1251), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(G384), .B1(new_n1277), .B2(new_n1251), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(KEYINPUT62), .B1(new_n1269), .B2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1277), .A2(new_n1251), .ZN(new_n1284));
  INV_X1    g1084(.A(G384), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1286), .A2(new_n1278), .ZN(new_n1287));
  AOI211_X1 g1087(.A(new_n1260), .B(new_n1287), .C1(new_n1263), .C2(new_n1268), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1288), .A2(KEYINPUT62), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1283), .A2(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1263), .A2(new_n1268), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1291), .A2(new_n1259), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1260), .A2(G2897), .ZN(new_n1293));
  XOR2_X1   g1093(.A(new_n1293), .B(KEYINPUT124), .Z(new_n1294));
  NAND2_X1  g1094(.A1(new_n1260), .A2(KEYINPUT123), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1294), .B1(new_n1281), .B2(new_n1295), .ZN(new_n1296));
  NAND4_X1  g1096(.A1(new_n1286), .A2(new_n1278), .A3(new_n1295), .A4(new_n1294), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1297), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(new_n1296), .A2(new_n1298), .ZN(new_n1299));
  AOI21_X1  g1099(.A(KEYINPUT61), .B1(new_n1292), .B2(new_n1299), .ZN(new_n1300));
  AOI21_X1  g1100(.A(KEYINPUT127), .B1(new_n1290), .B2(new_n1300), .ZN(new_n1301));
  AND3_X1   g1101(.A1(new_n1269), .A2(KEYINPUT62), .A3(new_n1281), .ZN(new_n1302));
  OAI211_X1 g1102(.A(new_n1300), .B(KEYINPUT127), .C1(new_n1302), .C2(new_n1282), .ZN(new_n1303));
  XNOR2_X1  g1103(.A(G393), .B(new_n818), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1088), .B1(new_n994), .B2(new_n1018), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1304), .B1(new_n1255), .B2(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(G387), .A2(G390), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1304), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1307), .A2(new_n1254), .A3(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1306), .A2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1303), .A2(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT125), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1312), .B1(new_n1296), .B2(new_n1298), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1286), .A2(new_n1278), .A3(new_n1295), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1294), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1314), .A2(new_n1315), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1316), .A2(KEYINPUT125), .A3(new_n1297), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1292), .A2(new_n1313), .A3(new_n1317), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1269), .A2(KEYINPUT63), .A3(new_n1281), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1318), .A2(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT61), .ZN(new_n1321));
  AND3_X1   g1121(.A1(new_n1306), .A2(new_n1321), .A3(new_n1309), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1322), .B1(new_n1288), .B2(KEYINPUT63), .ZN(new_n1323));
  NOR3_X1   g1123(.A1(new_n1320), .A2(new_n1323), .A3(KEYINPUT126), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT126), .ZN(new_n1325));
  AOI21_X1  g1125(.A(KEYINPUT125), .B1(new_n1316), .B2(new_n1297), .ZN(new_n1326));
  NOR2_X1   g1126(.A1(new_n1269), .A2(new_n1326), .ZN(new_n1327));
  AOI22_X1  g1127(.A1(new_n1327), .A2(new_n1317), .B1(new_n1288), .B2(KEYINPUT63), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1306), .A2(new_n1309), .A3(new_n1321), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1269), .A2(new_n1281), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT63), .ZN(new_n1331));
  AOI21_X1  g1131(.A(new_n1329), .B1(new_n1330), .B2(new_n1331), .ZN(new_n1332));
  AOI21_X1  g1132(.A(new_n1325), .B1(new_n1328), .B2(new_n1332), .ZN(new_n1333));
  OAI22_X1  g1133(.A1(new_n1301), .A2(new_n1311), .B1(new_n1324), .B2(new_n1333), .ZN(G405));
  INV_X1    g1134(.A(new_n1263), .ZN(new_n1335));
  AOI21_X1  g1135(.A(new_n1335), .B1(G375), .B2(new_n1256), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1336), .A2(new_n1287), .ZN(new_n1337));
  INV_X1    g1137(.A(new_n1337), .ZN(new_n1338));
  NOR2_X1   g1138(.A1(new_n1336), .A2(new_n1287), .ZN(new_n1339));
  OR3_X1    g1139(.A1(new_n1338), .A2(new_n1310), .A3(new_n1339), .ZN(new_n1340));
  OAI21_X1  g1140(.A(new_n1310), .B1(new_n1338), .B2(new_n1339), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1340), .A2(new_n1341), .ZN(G402));
endmodule


