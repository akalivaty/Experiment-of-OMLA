//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 0 0 1 1 1 1 0 0 0 1 1 0 0 0 0 0 0 0 0 1 1 1 0 0 0 0 0 0 0 1 0 0 1 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 1 0 1 1 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:00 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n447, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n558, new_n559, new_n560, new_n561, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n572, new_n574,
    new_n575, new_n577, new_n578, new_n579, new_n580, new_n581, new_n582,
    new_n583, new_n584, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n624, new_n625, new_n628, new_n630, new_n631, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n860, new_n861, new_n862, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1210, new_n1211, new_n1212;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT65), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XOR2_X1   g011(.A(new_n436), .B(KEYINPUT66), .Z(new_n437));
  INV_X1    g012(.A(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  NAND2_X1  g021(.A1(G94), .A2(G452), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n447), .B(KEYINPUT67), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g027(.A1(new_n437), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT68), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  INV_X1    g033(.A(G2106), .ZN(new_n459));
  INV_X1    g034(.A(G567), .ZN(new_n460));
  OAI22_X1  g035(.A1(new_n454), .A2(new_n459), .B1(new_n460), .B2(new_n455), .ZN(new_n461));
  XNOR2_X1  g036(.A(new_n461), .B(KEYINPUT69), .ZN(G319));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  OAI21_X1  g038(.A(KEYINPUT72), .B1(new_n463), .B2(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n463), .A2(KEYINPUT72), .A3(G2104), .ZN(new_n468));
  NAND4_X1  g043(.A1(new_n466), .A2(G137), .A3(new_n467), .A4(new_n468), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n467), .A2(G101), .A3(G2104), .ZN(new_n470));
  XNOR2_X1  g045(.A(new_n470), .B(KEYINPUT73), .ZN(new_n471));
  AND2_X1   g046(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(KEYINPUT3), .ZN(new_n474));
  AND3_X1   g049(.A1(new_n465), .A2(new_n474), .A3(G125), .ZN(new_n475));
  INV_X1    g050(.A(G113), .ZN(new_n476));
  OAI21_X1  g051(.A(KEYINPUT70), .B1(new_n476), .B2(new_n473), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT70), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n478), .A2(G113), .A3(G2104), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  OAI21_X1  g055(.A(G2105), .B1(new_n475), .B2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT71), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  OAI211_X1 g058(.A(KEYINPUT71), .B(G2105), .C1(new_n475), .C2(new_n480), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n472), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G160));
  AND2_X1   g061(.A1(new_n466), .A2(new_n468), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(new_n467), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT74), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n487), .A2(KEYINPUT74), .A3(new_n467), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n487), .A2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  AOI22_X1  g069(.A1(new_n492), .A2(G136), .B1(G124), .B2(new_n494), .ZN(new_n495));
  OAI21_X1  g070(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n467), .A2(G112), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT75), .ZN(new_n499));
  AND2_X1   g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n498), .A2(new_n499), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n500), .A2(new_n501), .ZN(G162));
  NAND4_X1  g077(.A1(new_n466), .A2(G126), .A3(G2105), .A4(new_n468), .ZN(new_n503));
  OR2_X1    g078(.A1(G102), .A2(G2105), .ZN(new_n504));
  OAI211_X1 g079(.A(new_n504), .B(G2104), .C1(G114), .C2(new_n467), .ZN(new_n505));
  AND3_X1   g080(.A1(new_n503), .A2(KEYINPUT76), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g081(.A(KEYINPUT76), .B1(new_n503), .B2(new_n505), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AND2_X1   g083(.A1(new_n467), .A2(G138), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT72), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n510), .B1(KEYINPUT3), .B2(new_n473), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n473), .A2(KEYINPUT3), .ZN(new_n512));
  OAI211_X1 g087(.A(new_n468), .B(new_n509), .C1(new_n511), .C2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(KEYINPUT77), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT77), .ZN(new_n515));
  NAND4_X1  g090(.A1(new_n466), .A2(new_n515), .A3(new_n468), .A4(new_n509), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n514), .A2(KEYINPUT4), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n465), .A2(new_n474), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n518), .A2(KEYINPUT4), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(new_n509), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n517), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n508), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(new_n522), .ZN(G164));
  XNOR2_X1  g098(.A(KEYINPUT5), .B(G543), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n524), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n525));
  INV_X1    g100(.A(G651), .ZN(new_n526));
  OR2_X1    g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT6), .ZN(new_n528));
  OAI21_X1  g103(.A(KEYINPUT78), .B1(new_n528), .B2(G651), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT78), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n530), .A2(new_n526), .A3(KEYINPUT6), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n528), .A2(G651), .ZN(new_n533));
  NAND4_X1  g108(.A1(new_n532), .A2(G88), .A3(new_n524), .A4(new_n533), .ZN(new_n534));
  NAND4_X1  g109(.A1(new_n532), .A2(G50), .A3(G543), .A4(new_n533), .ZN(new_n535));
  AND3_X1   g110(.A1(new_n534), .A2(new_n535), .A3(KEYINPUT79), .ZN(new_n536));
  AOI21_X1  g111(.A(KEYINPUT79), .B1(new_n534), .B2(new_n535), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n527), .B1(new_n536), .B2(new_n537), .ZN(G303));
  INV_X1    g113(.A(G303), .ZN(G166));
  AND2_X1   g114(.A1(new_n532), .A2(new_n533), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G543), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT80), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n532), .A2(new_n533), .ZN(new_n544));
  INV_X1    g119(.A(G543), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(KEYINPUT80), .ZN(new_n547));
  AND2_X1   g122(.A1(new_n543), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G51), .ZN(new_n549));
  AND3_X1   g124(.A1(new_n524), .A2(G63), .A3(G651), .ZN(new_n550));
  NAND3_X1  g125(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n551));
  XOR2_X1   g126(.A(new_n551), .B(KEYINPUT7), .Z(new_n552));
  INV_X1    g127(.A(new_n524), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n544), .A2(new_n553), .ZN(new_n554));
  AOI211_X1 g129(.A(new_n550), .B(new_n552), .C1(new_n554), .C2(G89), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n549), .A2(new_n555), .ZN(G286));
  INV_X1    g131(.A(G286), .ZN(G168));
  NAND3_X1  g132(.A1(new_n543), .A2(G52), .A3(new_n547), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n524), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n559));
  OR2_X1    g134(.A1(new_n559), .A2(new_n526), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n554), .A2(G90), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n558), .A2(new_n560), .A3(new_n561), .ZN(G301));
  INV_X1    g137(.A(G301), .ZN(G171));
  AOI22_X1  g138(.A1(new_n524), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n564));
  OR2_X1    g139(.A1(new_n564), .A2(new_n526), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n554), .A2(G81), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n543), .A2(new_n547), .ZN(new_n567));
  INV_X1    g142(.A(G43), .ZN(new_n568));
  OAI211_X1 g143(.A(new_n565), .B(new_n566), .C1(new_n567), .C2(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(G860), .ZN(G153));
  AND3_X1   g146(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(G36), .ZN(G176));
  NAND2_X1  g148(.A1(G1), .A2(G3), .ZN(new_n574));
  XNOR2_X1  g149(.A(new_n574), .B(KEYINPUT8), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n572), .A2(new_n575), .ZN(G188));
  INV_X1    g151(.A(G53), .ZN(new_n577));
  OAI21_X1  g152(.A(KEYINPUT9), .B1(new_n541), .B2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT9), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n546), .A2(new_n579), .A3(G53), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n578), .A2(new_n580), .B1(G91), .B2(new_n554), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n524), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n582), .A2(new_n526), .ZN(new_n583));
  XNOR2_X1  g158(.A(new_n583), .B(KEYINPUT81), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n581), .A2(new_n584), .ZN(G299));
  NAND2_X1  g160(.A1(new_n546), .A2(G49), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n554), .A2(G87), .ZN(new_n587));
  OAI21_X1  g162(.A(G651), .B1(new_n524), .B2(G74), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(G288));
  NAND3_X1  g164(.A1(new_n540), .A2(G86), .A3(new_n524), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n540), .A2(G48), .A3(G543), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n524), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT82), .ZN(new_n593));
  NOR3_X1   g168(.A1(new_n592), .A2(new_n593), .A3(new_n526), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n545), .A2(KEYINPUT5), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT5), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n596), .A2(G543), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n595), .A2(new_n597), .A3(G61), .ZN(new_n598));
  NAND2_X1  g173(.A1(G73), .A2(G543), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AOI21_X1  g175(.A(KEYINPUT82), .B1(new_n600), .B2(G651), .ZN(new_n601));
  OAI211_X1 g176(.A(new_n590), .B(new_n591), .C1(new_n594), .C2(new_n601), .ZN(G305));
  NAND2_X1  g177(.A1(new_n548), .A2(G47), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n554), .A2(G85), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n524), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n605));
  NOR2_X1   g180(.A1(new_n605), .A2(new_n526), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(KEYINPUT83), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n603), .A2(new_n604), .A3(new_n607), .ZN(G290));
  NAND2_X1  g183(.A1(G301), .A2(G868), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n554), .A2(G92), .ZN(new_n610));
  INV_X1    g185(.A(KEYINPUT84), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n610), .B(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(KEYINPUT10), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n610), .B(KEYINPUT84), .ZN(new_n614));
  INV_X1    g189(.A(KEYINPUT10), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g191(.A1(G79), .A2(G543), .ZN(new_n617));
  INV_X1    g192(.A(G66), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n553), .B2(new_n618), .ZN(new_n619));
  AOI22_X1  g194(.A1(new_n548), .A2(G54), .B1(G651), .B2(new_n619), .ZN(new_n620));
  AND3_X1   g195(.A1(new_n613), .A2(new_n616), .A3(new_n620), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n609), .B1(new_n621), .B2(G868), .ZN(G284));
  OAI21_X1  g197(.A(new_n609), .B1(new_n621), .B2(G868), .ZN(G321));
  INV_X1    g198(.A(G868), .ZN(new_n624));
  NAND2_X1  g199(.A1(G299), .A2(new_n624), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n625), .B1(G168), .B2(new_n624), .ZN(G297));
  XOR2_X1   g201(.A(G297), .B(KEYINPUT85), .Z(G280));
  INV_X1    g202(.A(G559), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n621), .B1(new_n628), .B2(G860), .ZN(G148));
  NAND2_X1  g204(.A1(new_n621), .A2(new_n628), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n630), .A2(G868), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n631), .B1(G868), .B2(new_n570), .ZN(G323));
  XNOR2_X1  g207(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AOI22_X1  g208(.A1(new_n492), .A2(G135), .B1(G123), .B2(new_n494), .ZN(new_n634));
  OAI21_X1  g209(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n635));
  INV_X1    g210(.A(G111), .ZN(new_n636));
  AOI21_X1  g211(.A(new_n635), .B1(new_n636), .B2(G2105), .ZN(new_n637));
  INV_X1    g212(.A(new_n637), .ZN(new_n638));
  AND2_X1   g213(.A1(new_n634), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2096), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n467), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n641));
  XOR2_X1   g216(.A(new_n641), .B(KEYINPUT12), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT13), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(G2100), .Z(new_n644));
  NAND2_X1  g219(.A1(new_n640), .A2(new_n644), .ZN(G156));
  XNOR2_X1  g220(.A(G2427), .B(G2438), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(G2430), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT15), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(G2435), .Z(new_n649));
  NAND2_X1  g224(.A1(new_n649), .A2(KEYINPUT14), .ZN(new_n650));
  XOR2_X1   g225(.A(G2443), .B(G2446), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G1341), .B(G1348), .ZN(new_n653));
  XNOR2_X1  g228(.A(KEYINPUT86), .B(KEYINPUT16), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n652), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2451), .B(G2454), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  INV_X1    g233(.A(G14), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n658), .A2(new_n659), .ZN(G401));
  XOR2_X1   g235(.A(G2072), .B(G2078), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT17), .ZN(new_n662));
  XOR2_X1   g237(.A(G2084), .B(G2090), .Z(new_n663));
  XOR2_X1   g238(.A(G2067), .B(G2678), .Z(new_n664));
  NAND3_X1  g239(.A1(new_n662), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n665), .B(KEYINPUT87), .Z(new_n666));
  INV_X1    g241(.A(new_n663), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n661), .A2(new_n664), .ZN(new_n668));
  OAI211_X1 g243(.A(new_n667), .B(new_n668), .C1(new_n662), .C2(new_n664), .ZN(new_n669));
  NOR3_X1   g244(.A1(new_n667), .A2(new_n661), .A3(new_n664), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT18), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n666), .A2(new_n669), .A3(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G2096), .B(G2100), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(G227));
  XOR2_X1   g250(.A(G1956), .B(G2474), .Z(new_n676));
  XOR2_X1   g251(.A(G1961), .B(G1966), .Z(new_n677));
  NOR2_X1   g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1971), .B(G1976), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT19), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n676), .A2(new_n677), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  INV_X1    g259(.A(KEYINPUT20), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n682), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n679), .A2(new_n681), .A3(new_n683), .ZN(new_n687));
  OAI211_X1 g262(.A(new_n686), .B(new_n687), .C1(new_n685), .C2(new_n684), .ZN(new_n688));
  XOR2_X1   g263(.A(G1981), .B(G1986), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(KEYINPUT88), .B(KEYINPUT89), .Z(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XOR2_X1   g268(.A(G1991), .B(G1996), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n690), .B(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(G229));
  OR2_X1    g272(.A1(G5), .A2(G16), .ZN(new_n698));
  INV_X1    g273(.A(G16), .ZN(new_n699));
  OAI211_X1 g274(.A(G1961), .B(new_n698), .C1(G301), .C2(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT101), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n698), .B1(G301), .B2(new_n699), .ZN(new_n702));
  INV_X1    g277(.A(G1961), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  AOI21_X1  g279(.A(KEYINPUT23), .B1(new_n699), .B2(G20), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n705), .B1(G299), .B2(G16), .ZN(new_n706));
  AND3_X1   g281(.A1(new_n699), .A2(KEYINPUT23), .A3(G20), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  AND3_X1   g283(.A1(new_n706), .A2(G1956), .A3(new_n708), .ZN(new_n709));
  AOI21_X1  g284(.A(G1956), .B1(new_n706), .B2(new_n708), .ZN(new_n710));
  OAI211_X1 g285(.A(new_n701), .B(new_n704), .C1(new_n709), .C2(new_n710), .ZN(new_n711));
  NAND4_X1  g286(.A1(new_n613), .A2(new_n616), .A3(new_n620), .A4(G16), .ZN(new_n712));
  OR2_X1    g287(.A1(G4), .A2(G16), .ZN(new_n713));
  XNOR2_X1  g288(.A(KEYINPUT93), .B(G1348), .ZN(new_n714));
  AND3_X1   g289(.A1(new_n712), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n714), .B1(new_n712), .B2(new_n713), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(G168), .A2(G16), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(G16), .B2(G21), .ZN(new_n719));
  INV_X1    g294(.A(G1966), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(G29), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n722), .A2(G27), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(G164), .B2(new_n722), .ZN(new_n724));
  XOR2_X1   g299(.A(KEYINPUT102), .B(G2078), .Z(new_n725));
  AND2_X1   g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NOR4_X1   g301(.A1(new_n711), .A2(new_n717), .A3(new_n721), .A4(new_n726), .ZN(new_n727));
  XNOR2_X1  g302(.A(KEYINPUT31), .B(G11), .ZN(new_n728));
  INV_X1    g303(.A(KEYINPUT97), .ZN(new_n729));
  NOR2_X1   g304(.A1(KEYINPUT24), .A2(G34), .ZN(new_n730));
  INV_X1    g305(.A(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(KEYINPUT24), .A2(G34), .ZN(new_n732));
  AOI21_X1  g307(.A(G29), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  AOI22_X1  g308(.A1(G160), .A2(G29), .B1(new_n729), .B2(new_n733), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(new_n729), .B2(new_n733), .ZN(new_n735));
  INV_X1    g310(.A(G2084), .ZN(new_n736));
  AND2_X1   g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(KEYINPUT30), .ZN(new_n738));
  OR2_X1    g313(.A1(new_n738), .A2(G28), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n738), .A2(G28), .ZN(new_n740));
  AND3_X1   g315(.A1(new_n739), .A2(new_n740), .A3(new_n722), .ZN(new_n741));
  AOI211_X1 g316(.A(new_n737), .B(new_n741), .C1(new_n719), .C2(new_n720), .ZN(new_n742));
  OR2_X1    g317(.A1(new_n724), .A2(new_n725), .ZN(new_n743));
  NAND4_X1  g318(.A1(new_n727), .A2(new_n728), .A3(new_n742), .A4(new_n743), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n735), .A2(new_n736), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n492), .A2(G141), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n746), .A2(KEYINPUT98), .ZN(new_n747));
  INV_X1    g322(.A(KEYINPUT98), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n492), .A2(new_n748), .A3(G141), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(G105), .ZN(new_n751));
  NOR3_X1   g326(.A1(new_n751), .A2(new_n473), .A3(G2105), .ZN(new_n752));
  NAND3_X1  g327(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT26), .ZN(new_n754));
  AOI211_X1 g329(.A(new_n752), .B(new_n754), .C1(new_n494), .C2(G129), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n722), .B1(new_n750), .B2(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n722), .A2(G32), .ZN(new_n757));
  INV_X1    g332(.A(new_n757), .ZN(new_n758));
  NOR3_X1   g333(.A1(new_n756), .A2(KEYINPUT99), .A3(new_n758), .ZN(new_n759));
  INV_X1    g334(.A(new_n759), .ZN(new_n760));
  OAI21_X1  g335(.A(KEYINPUT99), .B1(new_n756), .B2(new_n758), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  XOR2_X1   g337(.A(KEYINPUT27), .B(G1996), .Z(new_n763));
  INV_X1    g338(.A(new_n763), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n745), .B1(new_n762), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n492), .A2(G139), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n467), .A2(G103), .A3(G2104), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT25), .ZN(new_n768));
  INV_X1    g343(.A(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(G115), .A2(G2104), .ZN(new_n770));
  INV_X1    g345(.A(G127), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n770), .B1(new_n518), .B2(new_n771), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT95), .ZN(new_n773));
  OAI211_X1 g348(.A(new_n766), .B(new_n769), .C1(new_n467), .C2(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n774), .A2(G29), .ZN(new_n775));
  NAND2_X1  g350(.A1(KEYINPUT96), .A2(G2072), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n722), .A2(G33), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n775), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  NOR2_X1   g353(.A1(KEYINPUT96), .A2(G2072), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  AOI21_X1  g355(.A(KEYINPUT100), .B1(new_n765), .B2(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(new_n761), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n764), .B1(new_n782), .B2(new_n759), .ZN(new_n783));
  INV_X1    g358(.A(new_n745), .ZN(new_n784));
  AND4_X1   g359(.A1(KEYINPUT100), .A2(new_n783), .A3(new_n784), .A4(new_n780), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n762), .A2(new_n764), .ZN(new_n786));
  NOR4_X1   g361(.A1(new_n744), .A2(new_n781), .A3(new_n785), .A4(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n699), .A2(G19), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(new_n570), .B2(new_n699), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(G1341), .Z(new_n790));
  INV_X1    g365(.A(KEYINPUT91), .ZN(new_n791));
  AND2_X1   g366(.A1(new_n699), .A2(G23), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(G288), .B2(G16), .ZN(new_n793));
  INV_X1    g368(.A(KEYINPUT33), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(new_n795), .ZN(new_n796));
  AOI211_X1 g371(.A(KEYINPUT33), .B(new_n792), .C1(G288), .C2(G16), .ZN(new_n797));
  INV_X1    g372(.A(new_n797), .ZN(new_n798));
  NAND3_X1  g373(.A1(new_n796), .A2(G1976), .A3(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(G1976), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(new_n795), .B2(new_n797), .ZN(new_n801));
  AND2_X1   g376(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(KEYINPUT34), .ZN(new_n803));
  MUX2_X1   g378(.A(G6), .B(G305), .S(G16), .Z(new_n804));
  XOR2_X1   g379(.A(KEYINPUT32), .B(G1981), .Z(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n699), .A2(G22), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(G166), .B2(new_n699), .ZN(new_n808));
  INV_X1    g383(.A(G1971), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  NAND4_X1  g385(.A1(new_n802), .A2(new_n803), .A3(new_n806), .A4(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n722), .A2(G25), .ZN(new_n812));
  AOI22_X1  g387(.A1(new_n492), .A2(G131), .B1(G119), .B2(new_n494), .ZN(new_n813));
  OR2_X1    g388(.A1(G95), .A2(G2105), .ZN(new_n814));
  OAI211_X1 g389(.A(new_n814), .B(G2104), .C1(G107), .C2(new_n467), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT90), .ZN(new_n816));
  AND2_X1   g391(.A1(new_n813), .A2(new_n816), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n812), .B1(new_n817), .B2(new_n722), .ZN(new_n818));
  XNOR2_X1  g393(.A(KEYINPUT35), .B(G1991), .ZN(new_n819));
  XOR2_X1   g394(.A(new_n818), .B(new_n819), .Z(new_n820));
  NAND4_X1  g395(.A1(new_n810), .A2(new_n806), .A3(new_n799), .A4(new_n801), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n821), .A2(KEYINPUT34), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n699), .A2(G24), .ZN(new_n823));
  INV_X1    g398(.A(G290), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n823), .B1(new_n824), .B2(new_n699), .ZN(new_n825));
  INV_X1    g400(.A(G1986), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(new_n827));
  NAND4_X1  g402(.A1(new_n811), .A2(new_n820), .A3(new_n822), .A4(new_n827), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n791), .B1(new_n828), .B2(KEYINPUT92), .ZN(new_n829));
  OAI21_X1  g404(.A(KEYINPUT36), .B1(new_n828), .B2(new_n791), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  OAI211_X1 g406(.A(new_n791), .B(KEYINPUT36), .C1(new_n828), .C2(KEYINPUT92), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NOR2_X1   g408(.A1(G29), .A2(G35), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n834), .B1(G162), .B2(G29), .ZN(new_n835));
  XOR2_X1   g410(.A(KEYINPUT104), .B(G2090), .Z(new_n836));
  INV_X1    g411(.A(new_n836), .ZN(new_n837));
  OR2_X1    g412(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n835), .A2(new_n837), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(KEYINPUT103), .B(KEYINPUT29), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(new_n842));
  NAND4_X1  g417(.A1(new_n787), .A2(new_n790), .A3(new_n833), .A4(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT28), .ZN(new_n844));
  AND2_X1   g419(.A1(new_n492), .A2(G140), .ZN(new_n845));
  NOR2_X1   g420(.A1(G104), .A2(G2105), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT94), .ZN(new_n847));
  OAI211_X1 g422(.A(new_n847), .B(G2104), .C1(G116), .C2(new_n467), .ZN(new_n848));
  INV_X1    g423(.A(G128), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n848), .B1(new_n493), .B2(new_n849), .ZN(new_n850));
  OAI21_X1  g425(.A(G29), .B1(new_n845), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n722), .A2(G26), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n844), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n853), .B1(new_n844), .B2(new_n852), .ZN(new_n854));
  INV_X1    g429(.A(G2067), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n854), .B(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(new_n639), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n857), .A2(new_n722), .ZN(new_n858));
  NOR3_X1   g433(.A1(new_n843), .A2(new_n856), .A3(new_n858), .ZN(G311));
  AND3_X1   g434(.A1(new_n787), .A2(new_n833), .A3(new_n842), .ZN(new_n860));
  INV_X1    g435(.A(new_n856), .ZN(new_n861));
  INV_X1    g436(.A(new_n858), .ZN(new_n862));
  NAND4_X1  g437(.A1(new_n860), .A2(new_n861), .A3(new_n862), .A4(new_n790), .ZN(G150));
  NAND2_X1  g438(.A1(new_n554), .A2(G93), .ZN(new_n864));
  AOI22_X1  g439(.A1(new_n524), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n865));
  INV_X1    g440(.A(G55), .ZN(new_n866));
  OAI221_X1 g441(.A(new_n864), .B1(new_n526), .B2(new_n865), .C1(new_n567), .C2(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n867), .A2(G860), .ZN(new_n868));
  XOR2_X1   g443(.A(new_n868), .B(KEYINPUT37), .Z(new_n869));
  NAND3_X1  g444(.A1(new_n613), .A2(new_n616), .A3(new_n620), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n870), .A2(new_n628), .ZN(new_n871));
  XOR2_X1   g446(.A(KEYINPUT105), .B(KEYINPUT38), .Z(new_n872));
  XNOR2_X1  g447(.A(new_n871), .B(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n867), .B(new_n569), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(KEYINPUT39), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n873), .B(new_n875), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n869), .B1(new_n876), .B2(G860), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(KEYINPUT106), .ZN(G145));
  INV_X1    g453(.A(G37), .ZN(new_n879));
  NOR3_X1   g454(.A1(new_n500), .A2(new_n501), .A3(new_n639), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n639), .B1(new_n500), .B2(new_n501), .ZN(new_n882));
  AND3_X1   g457(.A1(new_n881), .A2(G160), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g458(.A(G160), .B1(new_n881), .B2(new_n882), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n642), .ZN(new_n886));
  AOI22_X1  g461(.A1(new_n492), .A2(G142), .B1(G130), .B2(new_n494), .ZN(new_n887));
  OAI21_X1  g462(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n888));
  INV_X1    g463(.A(G118), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n888), .B1(new_n889), .B2(G2105), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n887), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n817), .A2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT107), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n813), .A2(new_n816), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n895), .A2(new_n887), .A3(new_n891), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n893), .A2(new_n894), .A3(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n894), .B1(new_n893), .B2(new_n896), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n886), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n899), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n901), .A2(new_n642), .A3(new_n897), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n845), .A2(new_n850), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n904), .B(new_n774), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n750), .A2(new_n755), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n503), .A2(new_n505), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n907), .B1(new_n517), .B2(new_n520), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n907), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n521), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n911), .B1(new_n750), .B2(new_n755), .ZN(new_n912));
  OR3_X1    g487(.A1(new_n905), .A2(new_n909), .A3(new_n912), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n905), .B1(new_n909), .B2(new_n912), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n903), .A2(new_n915), .ZN(new_n916));
  NAND4_X1  g491(.A1(new_n900), .A2(new_n913), .A3(new_n902), .A4(new_n914), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n885), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT108), .ZN(new_n919));
  OAI211_X1 g494(.A(new_n913), .B(new_n914), .C1(new_n903), .C2(new_n919), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n915), .A2(KEYINPUT108), .A3(new_n902), .A4(new_n900), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  OAI211_X1 g497(.A(new_n879), .B(new_n918), .C1(new_n922), .C2(new_n885), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n923), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g499(.A1(new_n867), .A2(new_n624), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n630), .B(new_n874), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n621), .A2(G299), .ZN(new_n927));
  INV_X1    g502(.A(G299), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n870), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n926), .A2(new_n930), .ZN(new_n931));
  OR2_X1    g506(.A1(new_n931), .A2(KEYINPUT109), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(KEYINPUT109), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n927), .A2(KEYINPUT41), .A3(new_n929), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(KEYINPUT41), .B1(new_n927), .B2(new_n929), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  OAI211_X1 g512(.A(new_n932), .B(new_n933), .C1(new_n937), .C2(new_n926), .ZN(new_n938));
  XNOR2_X1  g513(.A(G303), .B(G288), .ZN(new_n939));
  XNOR2_X1  g514(.A(new_n939), .B(G290), .ZN(new_n940));
  XNOR2_X1  g515(.A(G305), .B(KEYINPUT110), .ZN(new_n941));
  INV_X1    g516(.A(new_n941), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n940), .B(new_n942), .ZN(new_n943));
  XNOR2_X1  g518(.A(new_n943), .B(KEYINPUT42), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n938), .B(new_n944), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n925), .B1(new_n945), .B2(new_n624), .ZN(G295));
  OAI21_X1  g521(.A(new_n925), .B1(new_n945), .B2(new_n624), .ZN(G331));
  INV_X1    g522(.A(KEYINPUT43), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n940), .B(new_n941), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT41), .ZN(new_n950));
  INV_X1    g525(.A(new_n929), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n870), .A2(new_n928), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n950), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  XNOR2_X1  g528(.A(G286), .B(G171), .ZN(new_n954));
  XNOR2_X1  g529(.A(new_n570), .B(new_n867), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  XNOR2_X1  g531(.A(G286), .B(G301), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(new_n874), .ZN(new_n958));
  AOI22_X1  g533(.A1(new_n953), .A2(new_n934), .B1(new_n956), .B2(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n956), .A2(new_n930), .A3(new_n958), .ZN(new_n960));
  INV_X1    g535(.A(new_n960), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n949), .B1(new_n959), .B2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT113), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  OAI211_X1 g539(.A(KEYINPUT113), .B(new_n949), .C1(new_n959), .C2(new_n961), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n956), .A2(new_n958), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n967), .B1(new_n935), .B2(new_n936), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n960), .A2(KEYINPUT112), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT112), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n930), .A2(new_n956), .A3(new_n958), .A4(new_n970), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n968), .A2(new_n969), .A3(new_n943), .A4(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(new_n879), .ZN(new_n973));
  INV_X1    g548(.A(new_n973), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n948), .B1(new_n966), .B2(new_n974), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n968), .A2(new_n969), .A3(new_n971), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(new_n949), .ZN(new_n977));
  INV_X1    g552(.A(new_n977), .ZN(new_n978));
  XNOR2_X1  g553(.A(KEYINPUT111), .B(KEYINPUT43), .ZN(new_n979));
  NOR3_X1   g554(.A1(new_n978), .A2(new_n973), .A3(new_n979), .ZN(new_n980));
  OAI21_X1  g555(.A(KEYINPUT44), .B1(new_n975), .B2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT44), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n979), .B1(new_n966), .B2(new_n974), .ZN(new_n983));
  INV_X1    g558(.A(new_n979), .ZN(new_n984));
  NOR3_X1   g559(.A1(new_n978), .A2(new_n973), .A3(new_n984), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n982), .B1(new_n983), .B2(new_n985), .ZN(new_n986));
  AND2_X1   g561(.A1(new_n981), .A2(new_n986), .ZN(G397));
  NAND4_X1  g562(.A1(new_n472), .A2(new_n483), .A3(G40), .A4(new_n484), .ZN(new_n988));
  INV_X1    g563(.A(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(G1384), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n989), .A2(new_n911), .A3(new_n990), .ZN(new_n991));
  XOR2_X1   g566(.A(KEYINPUT58), .B(G1341), .Z(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  AND2_X1   g568(.A1(new_n517), .A2(new_n520), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT76), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n907), .A2(new_n995), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n503), .A2(KEYINPUT76), .A3(new_n505), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n990), .B1(new_n994), .B2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT45), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g576(.A(G1384), .B1(new_n521), .B2(new_n910), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n988), .B1(new_n1002), .B2(KEYINPUT45), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n993), .B1(new_n1004), .B2(G1996), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(KEYINPUT121), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT121), .ZN(new_n1007));
  OAI211_X1 g582(.A(new_n1007), .B(new_n993), .C1(new_n1004), .C2(G1996), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1006), .A2(new_n570), .A3(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(KEYINPUT59), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT59), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n1006), .A2(new_n1011), .A3(new_n570), .A4(new_n1008), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n991), .A2(G2067), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT50), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n911), .A2(new_n1015), .A3(new_n990), .ZN(new_n1016));
  AOI21_X1  g591(.A(G1384), .B1(new_n508), .B2(new_n521), .ZN(new_n1017));
  OAI211_X1 g592(.A(new_n1016), .B(new_n989), .C1(new_n1015), .C2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(G1348), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1014), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(KEYINPUT60), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT123), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT60), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n988), .B1(new_n999), .B2(KEYINPUT50), .ZN(new_n1024));
  AOI21_X1  g599(.A(G1348), .B1(new_n1024), .B2(new_n1016), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1023), .B1(new_n1025), .B2(new_n1014), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1022), .B1(new_n1026), .B2(new_n621), .ZN(new_n1027));
  OAI211_X1 g602(.A(new_n1022), .B(new_n621), .C1(new_n1020), .C2(KEYINPUT60), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1028), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1021), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1030));
  NOR2_X1   g605(.A1(KEYINPUT122), .A2(KEYINPUT61), .ZN(new_n1031));
  NAND2_X1  g606(.A1(KEYINPUT122), .A2(KEYINPUT61), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1032), .ZN(new_n1033));
  XOR2_X1   g608(.A(KEYINPUT119), .B(G1956), .Z(new_n1034));
  OAI21_X1  g609(.A(new_n989), .B1(new_n1002), .B2(new_n1015), .ZN(new_n1035));
  AOI211_X1 g610(.A(KEYINPUT50), .B(G1384), .C1(new_n508), .C2(new_n521), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1034), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT57), .ZN(new_n1038));
  NAND2_X1  g613(.A1(G299), .A2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n581), .A2(KEYINPUT57), .A3(new_n584), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  XNOR2_X1  g616(.A(KEYINPUT56), .B(G2072), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1001), .A2(new_n1003), .A3(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1037), .A2(new_n1041), .A3(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1041), .B1(new_n1043), .B2(new_n1037), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1033), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1037), .A2(new_n1043), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1041), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1050), .A2(new_n1044), .A3(new_n1032), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1031), .B1(new_n1047), .B2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n621), .B1(new_n1020), .B2(KEYINPUT60), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(KEYINPUT123), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1054), .A2(KEYINPUT60), .A3(new_n1020), .A4(new_n1028), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1013), .A2(new_n1030), .A3(new_n1052), .A4(new_n1055), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1020), .A2(new_n870), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1046), .B1(new_n1057), .B2(KEYINPUT120), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1058), .B1(KEYINPUT120), .B2(new_n1057), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(new_n1044), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1056), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(G303), .A2(G8), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT115), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1063), .A2(KEYINPUT55), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1064), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1062), .A2(new_n1065), .ZN(new_n1066));
  XNOR2_X1  g641(.A(KEYINPUT115), .B(KEYINPUT55), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1066), .B1(new_n1062), .B2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1015), .B1(new_n522), .B2(new_n990), .ZN(new_n1069));
  NOR3_X1   g644(.A1(new_n908), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1070));
  NOR4_X1   g645(.A1(new_n1069), .A2(new_n1070), .A3(G2090), .A4(new_n988), .ZN(new_n1071));
  AOI21_X1  g646(.A(G1971), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1072));
  OAI211_X1 g647(.A(G8), .B(new_n1068), .C1(new_n1071), .C2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(G288), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(G1976), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n991), .A2(G8), .A3(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(KEYINPUT52), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT49), .ZN(new_n1078));
  NOR2_X1   g653(.A1(G305), .A2(G1981), .ZN(new_n1079));
  INV_X1    g654(.A(G1981), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n593), .B1(new_n592), .B2(new_n526), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n600), .A2(KEYINPUT82), .A3(G651), .ZN(new_n1082));
  AOI22_X1  g657(.A1(new_n1081), .A2(new_n1082), .B1(new_n546), .B2(G48), .ZN(new_n1083));
  XOR2_X1   g658(.A(KEYINPUT116), .B(G86), .Z(new_n1084));
  NAND2_X1  g659(.A1(new_n554), .A2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1080), .B1(new_n1083), .B2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1078), .B1(new_n1079), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(G8), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1088), .B1(new_n1002), .B2(new_n989), .ZN(new_n1089));
  OAI211_X1 g664(.A(new_n1085), .B(new_n591), .C1(new_n601), .C2(new_n594), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(G1981), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1083), .A2(new_n1080), .A3(new_n590), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1091), .A2(KEYINPUT49), .A3(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1087), .A2(new_n1089), .A3(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(KEYINPUT52), .B1(G288), .B2(new_n800), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1089), .A2(new_n1075), .A3(new_n1095), .ZN(new_n1096));
  AND3_X1   g671(.A1(new_n1077), .A2(new_n1094), .A3(new_n1096), .ZN(new_n1097));
  OR3_X1    g672(.A1(new_n1035), .A2(new_n1036), .A3(G2090), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n911), .A2(KEYINPUT45), .A3(new_n990), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(new_n989), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1017), .A2(KEYINPUT45), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n809), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1088), .B1(new_n1098), .B2(new_n1102), .ZN(new_n1103));
  OAI211_X1 g678(.A(new_n1073), .B(new_n1097), .C1(new_n1103), .C2(new_n1068), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT117), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1105), .B1(new_n1018), .B2(G2084), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n999), .A2(new_n1000), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n989), .B1(new_n1002), .B2(KEYINPUT45), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n720), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1024), .A2(KEYINPUT117), .A3(new_n736), .A4(new_n1016), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1106), .A2(new_n1109), .A3(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1111), .A2(G8), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT51), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1113), .A2(KEYINPUT124), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(G286), .A2(G8), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1112), .A2(new_n1115), .A3(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1113), .A2(KEYINPUT124), .ZN(new_n1118));
  OAI211_X1 g693(.A(G8), .B(new_n1114), .C1(new_n1111), .C2(G286), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1117), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1111), .A2(G8), .A3(G286), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1104), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1002), .ZN(new_n1123));
  OR2_X1    g698(.A1(new_n1123), .A2(KEYINPUT114), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(KEYINPUT114), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1124), .A2(new_n1000), .A3(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(G2078), .ZN(new_n1127));
  AND4_X1   g702(.A1(KEYINPUT53), .A2(new_n1099), .A3(new_n1127), .A4(new_n481), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1126), .A2(G40), .A3(new_n472), .A4(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1001), .A2(new_n1003), .A3(new_n1127), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT53), .ZN(new_n1131));
  AOI22_X1  g706(.A1(new_n1130), .A2(new_n1131), .B1(new_n1018), .B2(new_n703), .ZN(new_n1132));
  XNOR2_X1  g707(.A(KEYINPUT125), .B(KEYINPUT54), .ZN(new_n1133));
  NAND2_X1  g708(.A1(G301), .A2(new_n1133), .ZN(new_n1134));
  AND3_X1   g709(.A1(new_n1129), .A2(new_n1132), .A3(new_n1134), .ZN(new_n1135));
  OR2_X1    g710(.A1(G301), .A2(KEYINPUT54), .ZN(new_n1136));
  OR2_X1    g711(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1127), .A2(KEYINPUT53), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1132), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  NOR2_X1   g714(.A1(G171), .A2(KEYINPUT54), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1140), .B1(G171), .B2(new_n1133), .ZN(new_n1141));
  AOI22_X1  g716(.A1(new_n1135), .A2(new_n1136), .B1(new_n1139), .B2(new_n1141), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1061), .A2(new_n1122), .A3(new_n1142), .ZN(new_n1143));
  AND2_X1   g718(.A1(new_n1094), .A2(new_n800), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1079), .B1(new_n1144), .B2(new_n1074), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1089), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1097), .ZN(new_n1147));
  OAI22_X1  g722(.A1(new_n1145), .A2(new_n1146), .B1(new_n1147), .B2(new_n1073), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT118), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1111), .A2(G8), .A3(G168), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1073), .A2(new_n1097), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n999), .A2(KEYINPUT50), .ZN(new_n1153));
  INV_X1    g728(.A(G2090), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1153), .A2(new_n1154), .A3(new_n989), .A4(new_n1016), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1088), .B1(new_n1102), .B2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g731(.A(KEYINPUT63), .B1(new_n1156), .B2(new_n1068), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1157), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1149), .B1(new_n1152), .B2(new_n1158), .ZN(new_n1159));
  NOR4_X1   g734(.A1(new_n1150), .A2(new_n1157), .A3(new_n1151), .A4(KEYINPUT118), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT63), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1162), .B1(new_n1104), .B2(new_n1150), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1148), .B1(new_n1161), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1165), .A2(KEYINPUT62), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1139), .A2(G171), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n1104), .A2(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT62), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1120), .A2(new_n1169), .A3(new_n1121), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1166), .A2(new_n1168), .A3(new_n1170), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1143), .A2(new_n1164), .A3(new_n1171), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1126), .A2(new_n988), .ZN(new_n1173));
  XNOR2_X1  g748(.A(new_n906), .B(G1996), .ZN(new_n1174));
  XNOR2_X1  g749(.A(new_n904), .B(G2067), .ZN(new_n1175));
  INV_X1    g750(.A(new_n1175), .ZN(new_n1176));
  NOR2_X1   g751(.A1(new_n1174), .A2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n895), .A2(new_n819), .ZN(new_n1178));
  NOR2_X1   g753(.A1(new_n895), .A2(new_n819), .ZN(new_n1179));
  INV_X1    g754(.A(new_n1179), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1177), .A2(new_n1178), .A3(new_n1180), .ZN(new_n1181));
  NOR2_X1   g756(.A1(new_n824), .A2(new_n826), .ZN(new_n1182));
  OR2_X1    g757(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  NOR2_X1   g758(.A1(G290), .A2(G1986), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n1173), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1172), .A2(new_n1185), .ZN(new_n1186));
  INV_X1    g761(.A(new_n1173), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1177), .A2(new_n1179), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n904), .A2(new_n855), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n1187), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1181), .A2(new_n1173), .ZN(new_n1191));
  XNOR2_X1  g766(.A(new_n1191), .B(KEYINPUT127), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1173), .A2(new_n1184), .ZN(new_n1193));
  XNOR2_X1  g768(.A(new_n1193), .B(KEYINPUT48), .ZN(new_n1194));
  AOI21_X1  g769(.A(new_n1190), .B1(new_n1192), .B2(new_n1194), .ZN(new_n1195));
  INV_X1    g770(.A(KEYINPUT46), .ZN(new_n1196));
  OR3_X1    g771(.A1(new_n1187), .A2(new_n1196), .A3(G1996), .ZN(new_n1197));
  OAI21_X1  g772(.A(new_n1173), .B1(new_n1176), .B2(new_n906), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n1196), .B1(new_n1187), .B2(G1996), .ZN(new_n1199));
  NAND3_X1  g774(.A1(new_n1197), .A2(new_n1198), .A3(new_n1199), .ZN(new_n1200));
  XOR2_X1   g775(.A(KEYINPUT126), .B(KEYINPUT47), .Z(new_n1201));
  XNOR2_X1  g776(.A(new_n1200), .B(new_n1201), .ZN(new_n1202));
  NAND3_X1  g777(.A1(new_n1186), .A2(new_n1195), .A3(new_n1202), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g778(.A1(new_n974), .A2(new_n977), .A3(new_n979), .ZN(new_n1205));
  AOI21_X1  g779(.A(new_n973), .B1(new_n964), .B2(new_n965), .ZN(new_n1206));
  OAI211_X1 g780(.A(new_n1205), .B(G319), .C1(new_n1206), .C2(new_n979), .ZN(new_n1207));
  NAND3_X1  g781(.A1(new_n923), .A2(new_n674), .A3(new_n696), .ZN(new_n1208));
  NOR3_X1   g782(.A1(new_n1207), .A2(new_n1208), .A3(G401), .ZN(G308));
  INV_X1    g783(.A(new_n1208), .ZN(new_n1210));
  INV_X1    g784(.A(G401), .ZN(new_n1211));
  NOR2_X1   g785(.A1(new_n983), .A2(new_n985), .ZN(new_n1212));
  NAND4_X1  g786(.A1(new_n1210), .A2(G319), .A3(new_n1211), .A4(new_n1212), .ZN(G225));
endmodule


