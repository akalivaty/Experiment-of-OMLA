

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038, n1039, n1040;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U553 ( .A1(n727), .A2(n726), .ZN(n743) );
  BUF_X1 U554 ( .A(n731), .Z(n732) );
  INV_X4 U555 ( .A(n729), .ZN(n708) );
  NOR2_X1 U556 ( .A1(n717), .A2(n747), .ZN(n719) );
  NOR2_X1 U557 ( .A1(G1966), .A2(n731), .ZN(n744) );
  XOR2_X1 U558 ( .A(n815), .B(KEYINPUT89), .Z(n520) );
  INV_X1 U559 ( .A(KEYINPUT30), .ZN(n718) );
  XNOR2_X1 U560 ( .A(n719), .B(n718), .ZN(n720) );
  NOR2_X1 U561 ( .A1(n714), .A2(n713), .ZN(n727) );
  INV_X1 U562 ( .A(KEYINPUT99), .ZN(n738) );
  INV_X1 U563 ( .A(KEYINPUT97), .ZN(n745) );
  XNOR2_X1 U564 ( .A(KEYINPUT32), .B(KEYINPUT100), .ZN(n741) );
  XNOR2_X1 U565 ( .A(n742), .B(n741), .ZN(n770) );
  OR2_X1 U566 ( .A1(n676), .A2(n675), .ZN(n781) );
  NOR2_X1 U567 ( .A1(n672), .A2(G1384), .ZN(n782) );
  NAND2_X1 U568 ( .A1(n520), .A2(n816), .ZN(n817) );
  NOR2_X1 U569 ( .A1(G651), .A2(n631), .ZN(n638) );
  XOR2_X1 U570 ( .A(KEYINPUT17), .B(n521), .Z(n991) );
  XNOR2_X1 U571 ( .A(KEYINPUT1), .B(n535), .ZN(n642) );
  AND2_X1 U572 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U573 ( .A(G57), .ZN(G237) );
  INV_X1 U574 ( .A(G132), .ZN(G219) );
  INV_X1 U575 ( .A(G82), .ZN(G220) );
  NOR2_X1 U576 ( .A1(G2105), .A2(G2104), .ZN(n521) );
  NAND2_X1 U577 ( .A1(G138), .A2(n991), .ZN(n523) );
  INV_X1 U578 ( .A(G2104), .ZN(n525) );
  NOR2_X2 U579 ( .A1(G2105), .A2(n525), .ZN(n992) );
  NAND2_X1 U580 ( .A1(G102), .A2(n992), .ZN(n522) );
  NAND2_X1 U581 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U582 ( .A(KEYINPUT80), .B(n524), .ZN(n529) );
  AND2_X1 U583 ( .A1(n525), .A2(G2105), .ZN(n987) );
  NAND2_X1 U584 ( .A1(G126), .A2(n987), .ZN(n527) );
  AND2_X1 U585 ( .A1(G2104), .A2(G2105), .ZN(n988) );
  NAND2_X1 U586 ( .A1(G114), .A2(n988), .ZN(n526) );
  NAND2_X1 U587 ( .A1(n527), .A2(n526), .ZN(n528) );
  NOR2_X1 U588 ( .A1(n529), .A2(n528), .ZN(n672) );
  BUF_X1 U589 ( .A(n672), .Z(G164) );
  XOR2_X1 U590 ( .A(G543), .B(KEYINPUT0), .Z(n631) );
  XNOR2_X1 U591 ( .A(G651), .B(KEYINPUT65), .ZN(n533) );
  NOR2_X1 U592 ( .A1(n631), .A2(n533), .ZN(n646) );
  NAND2_X1 U593 ( .A1(n646), .A2(G75), .ZN(n532) );
  NOR2_X1 U594 ( .A1(G651), .A2(G543), .ZN(n530) );
  XNOR2_X1 U595 ( .A(n530), .B(KEYINPUT64), .ZN(n639) );
  NAND2_X1 U596 ( .A1(G88), .A2(n639), .ZN(n531) );
  NAND2_X1 U597 ( .A1(n532), .A2(n531), .ZN(n539) );
  NAND2_X1 U598 ( .A1(G50), .A2(n638), .ZN(n537) );
  NOR2_X1 U599 ( .A1(G543), .A2(n533), .ZN(n534) );
  XOR2_X1 U600 ( .A(KEYINPUT66), .B(n534), .Z(n535) );
  NAND2_X1 U601 ( .A1(G62), .A2(n642), .ZN(n536) );
  NAND2_X1 U602 ( .A1(n537), .A2(n536), .ZN(n538) );
  NOR2_X1 U603 ( .A1(n539), .A2(n538), .ZN(G166) );
  NAND2_X1 U604 ( .A1(n991), .A2(G137), .ZN(n542) );
  NAND2_X1 U605 ( .A1(G101), .A2(n992), .ZN(n540) );
  XOR2_X1 U606 ( .A(KEYINPUT23), .B(n540), .Z(n541) );
  NAND2_X1 U607 ( .A1(n542), .A2(n541), .ZN(n676) );
  NAND2_X1 U608 ( .A1(G125), .A2(n987), .ZN(n544) );
  NAND2_X1 U609 ( .A1(G113), .A2(n988), .ZN(n543) );
  NAND2_X1 U610 ( .A1(n544), .A2(n543), .ZN(n673) );
  NOR2_X1 U611 ( .A1(n676), .A2(n673), .ZN(G160) );
  NAND2_X1 U612 ( .A1(G7), .A2(G661), .ZN(n545) );
  XNOR2_X1 U613 ( .A(n545), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U614 ( .A(G223), .ZN(n833) );
  NAND2_X1 U615 ( .A1(n833), .A2(G567), .ZN(n546) );
  XOR2_X1 U616 ( .A(KEYINPUT11), .B(n546), .Z(G234) );
  NAND2_X1 U617 ( .A1(G56), .A2(n642), .ZN(n547) );
  XNOR2_X1 U618 ( .A(n547), .B(KEYINPUT14), .ZN(n549) );
  NAND2_X1 U619 ( .A1(G43), .A2(n638), .ZN(n548) );
  NAND2_X1 U620 ( .A1(n549), .A2(n548), .ZN(n556) );
  NAND2_X1 U621 ( .A1(G81), .A2(n639), .ZN(n550) );
  XNOR2_X1 U622 ( .A(n550), .B(KEYINPUT12), .ZN(n552) );
  NAND2_X1 U623 ( .A1(G68), .A2(n646), .ZN(n551) );
  NAND2_X1 U624 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U625 ( .A(KEYINPUT69), .B(n553), .ZN(n554) );
  XNOR2_X1 U626 ( .A(KEYINPUT13), .B(n554), .ZN(n555) );
  NOR2_X1 U627 ( .A1(n556), .A2(n555), .ZN(n1019) );
  NAND2_X1 U628 ( .A1(G860), .A2(n1019), .ZN(n557) );
  XNOR2_X1 U629 ( .A(n557), .B(KEYINPUT70), .ZN(G153) );
  NAND2_X1 U630 ( .A1(G52), .A2(n638), .ZN(n559) );
  NAND2_X1 U631 ( .A1(G64), .A2(n642), .ZN(n558) );
  NAND2_X1 U632 ( .A1(n559), .A2(n558), .ZN(n564) );
  NAND2_X1 U633 ( .A1(n646), .A2(G77), .ZN(n561) );
  NAND2_X1 U634 ( .A1(G90), .A2(n639), .ZN(n560) );
  NAND2_X1 U635 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U636 ( .A(KEYINPUT9), .B(n562), .Z(n563) );
  NOR2_X1 U637 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U638 ( .A(KEYINPUT68), .B(n565), .ZN(G171) );
  XNOR2_X1 U639 ( .A(KEYINPUT71), .B(G171), .ZN(G301) );
  NAND2_X1 U640 ( .A1(G868), .A2(G301), .ZN(n575) );
  NAND2_X1 U641 ( .A1(G66), .A2(n642), .ZN(n572) );
  NAND2_X1 U642 ( .A1(n646), .A2(G79), .ZN(n567) );
  NAND2_X1 U643 ( .A1(G92), .A2(n639), .ZN(n566) );
  NAND2_X1 U644 ( .A1(n567), .A2(n566), .ZN(n570) );
  NAND2_X1 U645 ( .A1(n638), .A2(G54), .ZN(n568) );
  XOR2_X1 U646 ( .A(KEYINPUT72), .B(n568), .Z(n569) );
  NOR2_X1 U647 ( .A1(n570), .A2(n569), .ZN(n571) );
  NAND2_X1 U648 ( .A1(n572), .A2(n571), .ZN(n573) );
  XOR2_X2 U649 ( .A(KEYINPUT15), .B(n573), .Z(n1016) );
  INV_X1 U650 ( .A(G868), .ZN(n656) );
  NAND2_X1 U651 ( .A1(n1016), .A2(n656), .ZN(n574) );
  NAND2_X1 U652 ( .A1(n575), .A2(n574), .ZN(G284) );
  NAND2_X1 U653 ( .A1(n646), .A2(G78), .ZN(n577) );
  NAND2_X1 U654 ( .A1(G91), .A2(n639), .ZN(n576) );
  NAND2_X1 U655 ( .A1(n577), .A2(n576), .ZN(n581) );
  NAND2_X1 U656 ( .A1(G53), .A2(n638), .ZN(n579) );
  NAND2_X1 U657 ( .A1(G65), .A2(n642), .ZN(n578) );
  NAND2_X1 U658 ( .A1(n579), .A2(n578), .ZN(n580) );
  NOR2_X1 U659 ( .A1(n581), .A2(n580), .ZN(n914) );
  INV_X1 U660 ( .A(n914), .ZN(G299) );
  NAND2_X1 U661 ( .A1(n639), .A2(G89), .ZN(n582) );
  XOR2_X1 U662 ( .A(KEYINPUT73), .B(n582), .Z(n583) );
  XNOR2_X1 U663 ( .A(n583), .B(KEYINPUT4), .ZN(n585) );
  NAND2_X1 U664 ( .A1(G76), .A2(n646), .ZN(n584) );
  NAND2_X1 U665 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U666 ( .A(n586), .B(KEYINPUT5), .ZN(n591) );
  NAND2_X1 U667 ( .A1(G51), .A2(n638), .ZN(n588) );
  NAND2_X1 U668 ( .A1(G63), .A2(n642), .ZN(n587) );
  NAND2_X1 U669 ( .A1(n588), .A2(n587), .ZN(n589) );
  XOR2_X1 U670 ( .A(KEYINPUT6), .B(n589), .Z(n590) );
  NAND2_X1 U671 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U672 ( .A(n592), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U673 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NOR2_X1 U674 ( .A1(G868), .A2(G299), .ZN(n594) );
  NOR2_X1 U675 ( .A1(G286), .A2(n656), .ZN(n593) );
  NOR2_X1 U676 ( .A1(n594), .A2(n593), .ZN(G297) );
  INV_X1 U677 ( .A(G860), .ZN(n595) );
  NAND2_X1 U678 ( .A1(n595), .A2(G559), .ZN(n596) );
  INV_X1 U679 ( .A(n1016), .ZN(n612) );
  NAND2_X1 U680 ( .A1(n596), .A2(n612), .ZN(n597) );
  XNOR2_X1 U681 ( .A(n597), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U682 ( .A1(n1019), .A2(n656), .ZN(n598) );
  XOR2_X1 U683 ( .A(KEYINPUT74), .B(n598), .Z(n601) );
  NAND2_X1 U684 ( .A1(G868), .A2(n612), .ZN(n599) );
  NOR2_X1 U685 ( .A1(G559), .A2(n599), .ZN(n600) );
  NOR2_X1 U686 ( .A1(n601), .A2(n600), .ZN(G282) );
  NAND2_X1 U687 ( .A1(G123), .A2(n987), .ZN(n602) );
  XOR2_X1 U688 ( .A(KEYINPUT18), .B(n602), .Z(n603) );
  XNOR2_X1 U689 ( .A(n603), .B(KEYINPUT75), .ZN(n605) );
  NAND2_X1 U690 ( .A1(G99), .A2(n992), .ZN(n604) );
  NAND2_X1 U691 ( .A1(n605), .A2(n604), .ZN(n609) );
  NAND2_X1 U692 ( .A1(G111), .A2(n988), .ZN(n607) );
  NAND2_X1 U693 ( .A1(G135), .A2(n991), .ZN(n606) );
  NAND2_X1 U694 ( .A1(n607), .A2(n606), .ZN(n608) );
  NOR2_X1 U695 ( .A1(n609), .A2(n608), .ZN(n1001) );
  XNOR2_X1 U696 ( .A(n1001), .B(G2096), .ZN(n611) );
  INV_X1 U697 ( .A(G2100), .ZN(n610) );
  NAND2_X1 U698 ( .A1(n611), .A2(n610), .ZN(G156) );
  NAND2_X1 U699 ( .A1(G559), .A2(n612), .ZN(n613) );
  XOR2_X1 U700 ( .A(n1019), .B(n613), .Z(n654) );
  NOR2_X1 U701 ( .A1(G860), .A2(n654), .ZN(n621) );
  NAND2_X1 U702 ( .A1(n646), .A2(G80), .ZN(n615) );
  NAND2_X1 U703 ( .A1(G93), .A2(n639), .ZN(n614) );
  NAND2_X1 U704 ( .A1(n615), .A2(n614), .ZN(n619) );
  NAND2_X1 U705 ( .A1(G55), .A2(n638), .ZN(n617) );
  NAND2_X1 U706 ( .A1(G67), .A2(n642), .ZN(n616) );
  NAND2_X1 U707 ( .A1(n617), .A2(n616), .ZN(n618) );
  OR2_X1 U708 ( .A1(n619), .A2(n618), .ZN(n657) );
  XOR2_X1 U709 ( .A(n657), .B(KEYINPUT76), .Z(n620) );
  XNOR2_X1 U710 ( .A(n621), .B(n620), .ZN(G145) );
  NAND2_X1 U711 ( .A1(G48), .A2(n638), .ZN(n622) );
  XNOR2_X1 U712 ( .A(n622), .B(KEYINPUT78), .ZN(n629) );
  NAND2_X1 U713 ( .A1(G86), .A2(n639), .ZN(n624) );
  NAND2_X1 U714 ( .A1(G61), .A2(n642), .ZN(n623) );
  NAND2_X1 U715 ( .A1(n624), .A2(n623), .ZN(n627) );
  NAND2_X1 U716 ( .A1(n646), .A2(G73), .ZN(n625) );
  XOR2_X1 U717 ( .A(KEYINPUT2), .B(n625), .Z(n626) );
  NOR2_X1 U718 ( .A1(n627), .A2(n626), .ZN(n628) );
  NAND2_X1 U719 ( .A1(n629), .A2(n628), .ZN(n630) );
  XOR2_X1 U720 ( .A(KEYINPUT79), .B(n630), .Z(G305) );
  NAND2_X1 U721 ( .A1(G49), .A2(n638), .ZN(n633) );
  NAND2_X1 U722 ( .A1(G87), .A2(n631), .ZN(n632) );
  NAND2_X1 U723 ( .A1(n633), .A2(n632), .ZN(n634) );
  NOR2_X1 U724 ( .A1(n642), .A2(n634), .ZN(n637) );
  NAND2_X1 U725 ( .A1(G74), .A2(G651), .ZN(n635) );
  XOR2_X1 U726 ( .A(KEYINPUT77), .B(n635), .Z(n636) );
  NAND2_X1 U727 ( .A1(n637), .A2(n636), .ZN(G288) );
  NAND2_X1 U728 ( .A1(n638), .A2(G47), .ZN(n641) );
  NAND2_X1 U729 ( .A1(G85), .A2(n639), .ZN(n640) );
  NAND2_X1 U730 ( .A1(n641), .A2(n640), .ZN(n645) );
  NAND2_X1 U731 ( .A1(G60), .A2(n642), .ZN(n643) );
  XNOR2_X1 U732 ( .A(KEYINPUT67), .B(n643), .ZN(n644) );
  NOR2_X1 U733 ( .A1(n645), .A2(n644), .ZN(n648) );
  NAND2_X1 U734 ( .A1(n646), .A2(G72), .ZN(n647) );
  NAND2_X1 U735 ( .A1(n648), .A2(n647), .ZN(G290) );
  XNOR2_X1 U736 ( .A(KEYINPUT19), .B(n657), .ZN(n649) );
  XNOR2_X1 U737 ( .A(G288), .B(n649), .ZN(n650) );
  XNOR2_X1 U738 ( .A(G305), .B(n650), .ZN(n652) );
  XNOR2_X1 U739 ( .A(G166), .B(n914), .ZN(n651) );
  XNOR2_X1 U740 ( .A(n652), .B(n651), .ZN(n653) );
  XOR2_X1 U741 ( .A(n653), .B(G290), .Z(n1017) );
  XNOR2_X1 U742 ( .A(n654), .B(n1017), .ZN(n655) );
  NAND2_X1 U743 ( .A1(n655), .A2(G868), .ZN(n659) );
  NAND2_X1 U744 ( .A1(n657), .A2(n656), .ZN(n658) );
  NAND2_X1 U745 ( .A1(n659), .A2(n658), .ZN(G295) );
  NAND2_X1 U746 ( .A1(G2078), .A2(G2084), .ZN(n660) );
  XOR2_X1 U747 ( .A(KEYINPUT20), .B(n660), .Z(n661) );
  NAND2_X1 U748 ( .A1(G2090), .A2(n661), .ZN(n662) );
  XNOR2_X1 U749 ( .A(KEYINPUT21), .B(n662), .ZN(n663) );
  NAND2_X1 U750 ( .A1(n663), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U751 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U752 ( .A1(G220), .A2(G219), .ZN(n664) );
  XOR2_X1 U753 ( .A(KEYINPUT22), .B(n664), .Z(n665) );
  NOR2_X1 U754 ( .A1(G218), .A2(n665), .ZN(n666) );
  NAND2_X1 U755 ( .A1(G96), .A2(n666), .ZN(n965) );
  NAND2_X1 U756 ( .A1(n965), .A2(G2106), .ZN(n670) );
  NAND2_X1 U757 ( .A1(G69), .A2(G120), .ZN(n667) );
  NOR2_X1 U758 ( .A1(G237), .A2(n667), .ZN(n668) );
  NAND2_X1 U759 ( .A1(G108), .A2(n668), .ZN(n964) );
  NAND2_X1 U760 ( .A1(n964), .A2(G567), .ZN(n669) );
  NAND2_X1 U761 ( .A1(n670), .A2(n669), .ZN(n967) );
  NAND2_X1 U762 ( .A1(G483), .A2(G661), .ZN(n671) );
  NOR2_X1 U763 ( .A1(n967), .A2(n671), .ZN(n838) );
  NAND2_X1 U764 ( .A1(n838), .A2(G36), .ZN(G176) );
  INV_X1 U765 ( .A(G166), .ZN(G303) );
  INV_X1 U766 ( .A(G40), .ZN(n674) );
  OR2_X1 U767 ( .A1(n674), .A2(n673), .ZN(n675) );
  XOR2_X1 U768 ( .A(KEYINPUT90), .B(n781), .Z(n677) );
  NAND2_X1 U769 ( .A1(n782), .A2(n677), .ZN(n729) );
  NAND2_X1 U770 ( .A1(n708), .A2(G2072), .ZN(n678) );
  XNOR2_X1 U771 ( .A(n678), .B(KEYINPUT27), .ZN(n680) );
  XOR2_X1 U772 ( .A(G1956), .B(KEYINPUT94), .Z(n931) );
  NOR2_X1 U773 ( .A1(n708), .A2(n931), .ZN(n679) );
  NOR2_X1 U774 ( .A1(n680), .A2(n679), .ZN(n702) );
  NOR2_X1 U775 ( .A1(n702), .A2(n914), .ZN(n682) );
  INV_X1 U776 ( .A(KEYINPUT28), .ZN(n681) );
  XNOR2_X1 U777 ( .A(n682), .B(n681), .ZN(n706) );
  INV_X1 U778 ( .A(G1341), .ZN(n684) );
  NAND2_X1 U779 ( .A1(G1348), .A2(n1016), .ZN(n683) );
  NAND2_X1 U780 ( .A1(n684), .A2(n683), .ZN(n685) );
  NAND2_X1 U781 ( .A1(n729), .A2(n685), .ZN(n688) );
  NAND2_X1 U782 ( .A1(n708), .A2(G1996), .ZN(n686) );
  XNOR2_X1 U783 ( .A(KEYINPUT26), .B(KEYINPUT95), .ZN(n689) );
  NAND2_X1 U784 ( .A1(n686), .A2(n689), .ZN(n687) );
  NAND2_X1 U785 ( .A1(n688), .A2(n687), .ZN(n696) );
  NAND2_X1 U786 ( .A1(G2067), .A2(n1016), .ZN(n692) );
  INV_X1 U787 ( .A(n689), .ZN(n690) );
  NAND2_X1 U788 ( .A1(G1996), .A2(n690), .ZN(n691) );
  NAND2_X1 U789 ( .A1(n692), .A2(n691), .ZN(n693) );
  NAND2_X1 U790 ( .A1(n693), .A2(n708), .ZN(n694) );
  NAND2_X1 U791 ( .A1(n694), .A2(n1019), .ZN(n695) );
  NOR2_X1 U792 ( .A1(n696), .A2(n695), .ZN(n701) );
  NAND2_X1 U793 ( .A1(G1348), .A2(n729), .ZN(n698) );
  NAND2_X1 U794 ( .A1(G2067), .A2(n708), .ZN(n697) );
  NAND2_X1 U795 ( .A1(n698), .A2(n697), .ZN(n699) );
  NOR2_X1 U796 ( .A1(n699), .A2(n1016), .ZN(n700) );
  NOR2_X1 U797 ( .A1(n701), .A2(n700), .ZN(n704) );
  NAND2_X1 U798 ( .A1(n702), .A2(n914), .ZN(n703) );
  NAND2_X1 U799 ( .A1(n704), .A2(n703), .ZN(n705) );
  NAND2_X1 U800 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U801 ( .A(n707), .B(KEYINPUT29), .ZN(n714) );
  INV_X1 U802 ( .A(G171), .ZN(n1021) );
  NOR2_X1 U803 ( .A1(n708), .A2(G1961), .ZN(n709) );
  XNOR2_X1 U804 ( .A(n709), .B(KEYINPUT92), .ZN(n712) );
  XNOR2_X1 U805 ( .A(G2078), .B(KEYINPUT25), .ZN(n710) );
  XNOR2_X1 U806 ( .A(n710), .B(KEYINPUT93), .ZN(n886) );
  NOR2_X1 U807 ( .A1(n729), .A2(n886), .ZN(n711) );
  NOR2_X1 U808 ( .A1(n712), .A2(n711), .ZN(n721) );
  NOR2_X1 U809 ( .A1(n1021), .A2(n721), .ZN(n713) );
  INV_X1 U810 ( .A(G8), .ZN(n715) );
  NAND2_X1 U811 ( .A1(G8), .A2(n729), .ZN(n731) );
  OR2_X1 U812 ( .A1(n715), .A2(n744), .ZN(n717) );
  NOR2_X1 U813 ( .A1(G2084), .A2(n729), .ZN(n716) );
  XOR2_X1 U814 ( .A(KEYINPUT91), .B(n716), .Z(n747) );
  NOR2_X1 U815 ( .A1(G168), .A2(n720), .ZN(n724) );
  AND2_X1 U816 ( .A1(n1021), .A2(n721), .ZN(n722) );
  XNOR2_X1 U817 ( .A(n722), .B(KEYINPUT96), .ZN(n723) );
  NOR2_X1 U818 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U819 ( .A(n725), .B(KEYINPUT31), .ZN(n726) );
  INV_X1 U820 ( .A(n743), .ZN(n728) );
  NAND2_X1 U821 ( .A1(G286), .A2(n728), .ZN(n737) );
  NOR2_X1 U822 ( .A1(G2090), .A2(n729), .ZN(n730) );
  XNOR2_X1 U823 ( .A(n730), .B(KEYINPUT98), .ZN(n734) );
  NOR2_X1 U824 ( .A1(n732), .A2(G1971), .ZN(n733) );
  NOR2_X1 U825 ( .A1(n734), .A2(n733), .ZN(n735) );
  NAND2_X1 U826 ( .A1(n735), .A2(G303), .ZN(n736) );
  NAND2_X1 U827 ( .A1(n737), .A2(n736), .ZN(n739) );
  XNOR2_X1 U828 ( .A(n739), .B(n738), .ZN(n740) );
  NAND2_X1 U829 ( .A1(n740), .A2(G8), .ZN(n742) );
  NOR2_X1 U830 ( .A1(n744), .A2(n743), .ZN(n746) );
  XNOR2_X1 U831 ( .A(n746), .B(n745), .ZN(n749) );
  NAND2_X1 U832 ( .A1(n747), .A2(G8), .ZN(n748) );
  NAND2_X1 U833 ( .A1(n749), .A2(n748), .ZN(n771) );
  AND2_X1 U834 ( .A1(G1976), .A2(G288), .ZN(n917) );
  NOR2_X1 U835 ( .A1(n917), .A2(n732), .ZN(n752) );
  AND2_X1 U836 ( .A1(n771), .A2(n752), .ZN(n750) );
  AND2_X1 U837 ( .A1(n750), .A2(n760), .ZN(n751) );
  NAND2_X1 U838 ( .A1(n770), .A2(n751), .ZN(n757) );
  INV_X1 U839 ( .A(n752), .ZN(n754) );
  NOR2_X1 U840 ( .A1(G1976), .A2(G288), .ZN(n761) );
  NOR2_X1 U841 ( .A1(G1971), .A2(G303), .ZN(n753) );
  NOR2_X1 U842 ( .A1(n761), .A2(n753), .ZN(n923) );
  OR2_X1 U843 ( .A1(n754), .A2(n923), .ZN(n755) );
  OR2_X1 U844 ( .A1(KEYINPUT101), .A2(n755), .ZN(n756) );
  NAND2_X1 U845 ( .A1(n757), .A2(n756), .ZN(n758) );
  NOR2_X1 U846 ( .A1(KEYINPUT33), .A2(n758), .ZN(n766) );
  INV_X1 U847 ( .A(KEYINPUT101), .ZN(n760) );
  NAND2_X1 U848 ( .A1(n761), .A2(KEYINPUT33), .ZN(n759) );
  NAND2_X1 U849 ( .A1(n760), .A2(n759), .ZN(n763) );
  NAND2_X1 U850 ( .A1(n761), .A2(KEYINPUT101), .ZN(n762) );
  NAND2_X1 U851 ( .A1(n763), .A2(n762), .ZN(n764) );
  NOR2_X1 U852 ( .A1(n732), .A2(n764), .ZN(n765) );
  NOR2_X1 U853 ( .A1(n766), .A2(n765), .ZN(n767) );
  XOR2_X1 U854 ( .A(G1981), .B(G305), .Z(n908) );
  NAND2_X1 U855 ( .A1(n767), .A2(n908), .ZN(n776) );
  NOR2_X1 U856 ( .A1(G2090), .A2(G303), .ZN(n768) );
  XNOR2_X1 U857 ( .A(n768), .B(KEYINPUT102), .ZN(n769) );
  NAND2_X1 U858 ( .A1(n769), .A2(G8), .ZN(n773) );
  NAND2_X1 U859 ( .A1(n771), .A2(n770), .ZN(n772) );
  NAND2_X1 U860 ( .A1(n773), .A2(n772), .ZN(n774) );
  NAND2_X1 U861 ( .A1(n774), .A2(n732), .ZN(n775) );
  NAND2_X1 U862 ( .A1(n776), .A2(n775), .ZN(n780) );
  NOR2_X1 U863 ( .A1(G1981), .A2(G305), .ZN(n777) );
  XOR2_X1 U864 ( .A(n777), .B(KEYINPUT24), .Z(n778) );
  NOR2_X1 U865 ( .A1(n732), .A2(n778), .ZN(n779) );
  NOR2_X1 U866 ( .A1(n780), .A2(n779), .ZN(n818) );
  NOR2_X1 U867 ( .A1(n782), .A2(n781), .ZN(n828) );
  NAND2_X1 U868 ( .A1(G105), .A2(n992), .ZN(n783) );
  XNOR2_X1 U869 ( .A(n783), .B(KEYINPUT38), .ZN(n791) );
  NAND2_X1 U870 ( .A1(G117), .A2(n988), .ZN(n784) );
  XNOR2_X1 U871 ( .A(n784), .B(KEYINPUT86), .ZN(n786) );
  NAND2_X1 U872 ( .A1(n987), .A2(G129), .ZN(n785) );
  NAND2_X1 U873 ( .A1(n786), .A2(n785), .ZN(n789) );
  NAND2_X1 U874 ( .A1(G141), .A2(n991), .ZN(n787) );
  XNOR2_X1 U875 ( .A(KEYINPUT87), .B(n787), .ZN(n788) );
  NOR2_X1 U876 ( .A1(n789), .A2(n788), .ZN(n790) );
  NAND2_X1 U877 ( .A1(n791), .A2(n790), .ZN(n1008) );
  NAND2_X1 U878 ( .A1(G1996), .A2(n1008), .ZN(n792) );
  XNOR2_X1 U879 ( .A(n792), .B(KEYINPUT88), .ZN(n802) );
  XOR2_X1 U880 ( .A(G1991), .B(KEYINPUT85), .Z(n892) );
  NAND2_X1 U881 ( .A1(G95), .A2(n992), .ZN(n799) );
  NAND2_X1 U882 ( .A1(G119), .A2(n987), .ZN(n794) );
  NAND2_X1 U883 ( .A1(G131), .A2(n991), .ZN(n793) );
  NAND2_X1 U884 ( .A1(n794), .A2(n793), .ZN(n797) );
  NAND2_X1 U885 ( .A1(G107), .A2(n988), .ZN(n795) );
  XNOR2_X1 U886 ( .A(KEYINPUT83), .B(n795), .ZN(n796) );
  NOR2_X1 U887 ( .A1(n797), .A2(n796), .ZN(n798) );
  NAND2_X1 U888 ( .A1(n799), .A2(n798), .ZN(n800) );
  XNOR2_X1 U889 ( .A(n800), .B(KEYINPUT84), .ZN(n1003) );
  NAND2_X1 U890 ( .A1(n892), .A2(n1003), .ZN(n801) );
  NAND2_X1 U891 ( .A1(n802), .A2(n801), .ZN(n822) );
  INV_X1 U892 ( .A(n822), .ZN(n854) );
  NAND2_X1 U893 ( .A1(G128), .A2(n987), .ZN(n804) );
  NAND2_X1 U894 ( .A1(G116), .A2(n988), .ZN(n803) );
  NAND2_X1 U895 ( .A1(n804), .A2(n803), .ZN(n805) );
  XNOR2_X1 U896 ( .A(KEYINPUT35), .B(n805), .ZN(n811) );
  NAND2_X1 U897 ( .A1(G140), .A2(n991), .ZN(n807) );
  NAND2_X1 U898 ( .A1(G104), .A2(n992), .ZN(n806) );
  NAND2_X1 U899 ( .A1(n807), .A2(n806), .ZN(n809) );
  XOR2_X1 U900 ( .A(KEYINPUT34), .B(KEYINPUT82), .Z(n808) );
  XNOR2_X1 U901 ( .A(n809), .B(n808), .ZN(n810) );
  NAND2_X1 U902 ( .A1(n811), .A2(n810), .ZN(n812) );
  XOR2_X1 U903 ( .A(KEYINPUT36), .B(n812), .Z(n1004) );
  XNOR2_X1 U904 ( .A(G2067), .B(KEYINPUT37), .ZN(n813) );
  XOR2_X1 U905 ( .A(n813), .B(KEYINPUT81), .Z(n826) );
  OR2_X1 U906 ( .A1(n1004), .A2(n826), .ZN(n849) );
  NAND2_X1 U907 ( .A1(n854), .A2(n849), .ZN(n814) );
  NAND2_X1 U908 ( .A1(n828), .A2(n814), .ZN(n815) );
  XNOR2_X1 U909 ( .A(G1986), .B(G290), .ZN(n921) );
  NAND2_X1 U910 ( .A1(n921), .A2(n828), .ZN(n816) );
  OR2_X1 U911 ( .A1(n818), .A2(n817), .ZN(n831) );
  NOR2_X1 U912 ( .A1(G1996), .A2(n1008), .ZN(n873) );
  NOR2_X1 U913 ( .A1(G1986), .A2(G290), .ZN(n819) );
  NOR2_X1 U914 ( .A1(n1003), .A2(n892), .ZN(n852) );
  NOR2_X1 U915 ( .A1(n819), .A2(n852), .ZN(n820) );
  XOR2_X1 U916 ( .A(KEYINPUT103), .B(n820), .Z(n821) );
  NOR2_X1 U917 ( .A1(n822), .A2(n821), .ZN(n823) );
  NOR2_X1 U918 ( .A1(n873), .A2(n823), .ZN(n824) );
  XNOR2_X1 U919 ( .A(n824), .B(KEYINPUT39), .ZN(n825) );
  NAND2_X1 U920 ( .A1(n825), .A2(n849), .ZN(n827) );
  NAND2_X1 U921 ( .A1(n1004), .A2(n826), .ZN(n853) );
  NAND2_X1 U922 ( .A1(n827), .A2(n853), .ZN(n829) );
  NAND2_X1 U923 ( .A1(n829), .A2(n828), .ZN(n830) );
  NAND2_X1 U924 ( .A1(n831), .A2(n830), .ZN(n832) );
  XNOR2_X1 U925 ( .A(n832), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U926 ( .A1(G2106), .A2(n833), .ZN(G217) );
  NAND2_X1 U927 ( .A1(G15), .A2(G2), .ZN(n835) );
  INV_X1 U928 ( .A(G661), .ZN(n834) );
  NOR2_X1 U929 ( .A1(n835), .A2(n834), .ZN(n836) );
  XNOR2_X1 U930 ( .A(n836), .B(KEYINPUT105), .ZN(G259) );
  NAND2_X1 U931 ( .A1(G3), .A2(G1), .ZN(n837) );
  NAND2_X1 U932 ( .A1(n838), .A2(n837), .ZN(G188) );
  NAND2_X1 U934 ( .A1(G124), .A2(n987), .ZN(n839) );
  XOR2_X1 U935 ( .A(KEYINPUT44), .B(n839), .Z(n840) );
  XNOR2_X1 U936 ( .A(n840), .B(KEYINPUT109), .ZN(n842) );
  NAND2_X1 U937 ( .A1(G136), .A2(n991), .ZN(n841) );
  NAND2_X1 U938 ( .A1(n842), .A2(n841), .ZN(n843) );
  XNOR2_X1 U939 ( .A(KEYINPUT110), .B(n843), .ZN(n847) );
  NAND2_X1 U940 ( .A1(G112), .A2(n988), .ZN(n845) );
  NAND2_X1 U941 ( .A1(G100), .A2(n992), .ZN(n844) );
  NAND2_X1 U942 ( .A1(n845), .A2(n844), .ZN(n846) );
  NOR2_X1 U943 ( .A1(n847), .A2(n846), .ZN(G162) );
  XOR2_X1 U944 ( .A(G2084), .B(G160), .Z(n848) );
  NOR2_X1 U945 ( .A1(n1001), .A2(n848), .ZN(n850) );
  NAND2_X1 U946 ( .A1(n850), .A2(n849), .ZN(n851) );
  NOR2_X1 U947 ( .A1(n852), .A2(n851), .ZN(n870) );
  NAND2_X1 U948 ( .A1(n854), .A2(n853), .ZN(n868) );
  NAND2_X1 U949 ( .A1(G127), .A2(n987), .ZN(n856) );
  NAND2_X1 U950 ( .A1(G115), .A2(n988), .ZN(n855) );
  NAND2_X1 U951 ( .A1(n856), .A2(n855), .ZN(n857) );
  XNOR2_X1 U952 ( .A(n857), .B(KEYINPUT47), .ZN(n862) );
  NAND2_X1 U953 ( .A1(G139), .A2(n991), .ZN(n859) );
  NAND2_X1 U954 ( .A1(G103), .A2(n992), .ZN(n858) );
  NAND2_X1 U955 ( .A1(n859), .A2(n858), .ZN(n860) );
  XOR2_X1 U956 ( .A(KEYINPUT112), .B(n860), .Z(n861) );
  NAND2_X1 U957 ( .A1(n862), .A2(n861), .ZN(n863) );
  XNOR2_X1 U958 ( .A(n863), .B(KEYINPUT113), .ZN(n1013) );
  XOR2_X1 U959 ( .A(G2072), .B(n1013), .Z(n865) );
  XOR2_X1 U960 ( .A(G164), .B(G2078), .Z(n864) );
  NOR2_X1 U961 ( .A1(n865), .A2(n864), .ZN(n866) );
  XOR2_X1 U962 ( .A(KEYINPUT50), .B(n866), .Z(n867) );
  NOR2_X1 U963 ( .A1(n868), .A2(n867), .ZN(n869) );
  NAND2_X1 U964 ( .A1(n870), .A2(n869), .ZN(n876) );
  XOR2_X1 U965 ( .A(G2090), .B(G162), .Z(n871) );
  XNOR2_X1 U966 ( .A(KEYINPUT116), .B(n871), .ZN(n872) );
  NOR2_X1 U967 ( .A1(n873), .A2(n872), .ZN(n874) );
  XNOR2_X1 U968 ( .A(KEYINPUT51), .B(n874), .ZN(n875) );
  NOR2_X1 U969 ( .A1(n876), .A2(n875), .ZN(n877) );
  XOR2_X1 U970 ( .A(KEYINPUT52), .B(n877), .Z(n878) );
  NOR2_X1 U971 ( .A1(KEYINPUT55), .A2(n878), .ZN(n879) );
  XNOR2_X1 U972 ( .A(KEYINPUT117), .B(n879), .ZN(n880) );
  NAND2_X1 U973 ( .A1(n880), .A2(G29), .ZN(n962) );
  XNOR2_X1 U974 ( .A(KEYINPUT54), .B(G34), .ZN(n881) );
  XNOR2_X1 U975 ( .A(n881), .B(KEYINPUT120), .ZN(n882) );
  XNOR2_X1 U976 ( .A(G2084), .B(n882), .ZN(n900) );
  XNOR2_X1 U977 ( .A(G2090), .B(G35), .ZN(n897) );
  XNOR2_X1 U978 ( .A(G2067), .B(G26), .ZN(n884) );
  XNOR2_X1 U979 ( .A(G33), .B(G2072), .ZN(n883) );
  NOR2_X1 U980 ( .A1(n884), .A2(n883), .ZN(n891) );
  XOR2_X1 U981 ( .A(G1996), .B(G32), .Z(n885) );
  NAND2_X1 U982 ( .A1(n885), .A2(G28), .ZN(n889) );
  XNOR2_X1 U983 ( .A(G27), .B(n886), .ZN(n887) );
  XNOR2_X1 U984 ( .A(KEYINPUT118), .B(n887), .ZN(n888) );
  NOR2_X1 U985 ( .A1(n889), .A2(n888), .ZN(n890) );
  NAND2_X1 U986 ( .A1(n891), .A2(n890), .ZN(n894) );
  XNOR2_X1 U987 ( .A(G25), .B(n892), .ZN(n893) );
  NOR2_X1 U988 ( .A1(n894), .A2(n893), .ZN(n895) );
  XNOR2_X1 U989 ( .A(KEYINPUT53), .B(n895), .ZN(n896) );
  NOR2_X1 U990 ( .A1(n897), .A2(n896), .ZN(n898) );
  XNOR2_X1 U991 ( .A(KEYINPUT119), .B(n898), .ZN(n899) );
  NOR2_X1 U992 ( .A1(n900), .A2(n899), .ZN(n901) );
  XNOR2_X1 U993 ( .A(KEYINPUT55), .B(n901), .ZN(n903) );
  INV_X1 U994 ( .A(G29), .ZN(n902) );
  NAND2_X1 U995 ( .A1(n903), .A2(n902), .ZN(n904) );
  NAND2_X1 U996 ( .A1(n904), .A2(G11), .ZN(n960) );
  INV_X1 U997 ( .A(G16), .ZN(n956) );
  XNOR2_X1 U998 ( .A(KEYINPUT56), .B(KEYINPUT121), .ZN(n905) );
  XNOR2_X1 U999 ( .A(n956), .B(n905), .ZN(n930) );
  XOR2_X1 U1000 ( .A(n1019), .B(G1341), .Z(n907) );
  XNOR2_X1 U1001 ( .A(n1021), .B(G1961), .ZN(n906) );
  NOR2_X1 U1002 ( .A1(n907), .A2(n906), .ZN(n928) );
  XOR2_X1 U1003 ( .A(n1016), .B(G1348), .Z(n913) );
  XNOR2_X1 U1004 ( .A(G168), .B(G1966), .ZN(n909) );
  NAND2_X1 U1005 ( .A1(n909), .A2(n908), .ZN(n910) );
  XNOR2_X1 U1006 ( .A(n910), .B(KEYINPUT57), .ZN(n911) );
  XNOR2_X1 U1007 ( .A(KEYINPUT122), .B(n911), .ZN(n912) );
  NAND2_X1 U1008 ( .A1(n913), .A2(n912), .ZN(n926) );
  XNOR2_X1 U1009 ( .A(n914), .B(G1956), .ZN(n919) );
  INV_X1 U1010 ( .A(G1971), .ZN(n915) );
  NOR2_X1 U1011 ( .A1(G166), .A2(n915), .ZN(n916) );
  NOR2_X1 U1012 ( .A1(n917), .A2(n916), .ZN(n918) );
  NAND2_X1 U1013 ( .A1(n919), .A2(n918), .ZN(n920) );
  NOR2_X1 U1014 ( .A1(n921), .A2(n920), .ZN(n922) );
  NAND2_X1 U1015 ( .A1(n923), .A2(n922), .ZN(n924) );
  XOR2_X1 U1016 ( .A(KEYINPUT123), .B(n924), .Z(n925) );
  NOR2_X1 U1017 ( .A1(n926), .A2(n925), .ZN(n927) );
  NAND2_X1 U1018 ( .A1(n928), .A2(n927), .ZN(n929) );
  NAND2_X1 U1019 ( .A1(n930), .A2(n929), .ZN(n958) );
  XOR2_X1 U1020 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n954) );
  XOR2_X1 U1021 ( .A(G1981), .B(G6), .Z(n933) );
  XNOR2_X1 U1022 ( .A(n931), .B(G20), .ZN(n932) );
  NAND2_X1 U1023 ( .A1(n933), .A2(n932), .ZN(n935) );
  XNOR2_X1 U1024 ( .A(G19), .B(G1341), .ZN(n934) );
  NOR2_X1 U1025 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1026 ( .A(KEYINPUT124), .B(n936), .ZN(n940) );
  XOR2_X1 U1027 ( .A(G4), .B(KEYINPUT125), .Z(n938) );
  XNOR2_X1 U1028 ( .A(G1348), .B(KEYINPUT59), .ZN(n937) );
  XNOR2_X1 U1029 ( .A(n938), .B(n937), .ZN(n939) );
  NAND2_X1 U1030 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1031 ( .A(n941), .B(KEYINPUT60), .ZN(n948) );
  XNOR2_X1 U1032 ( .A(G1971), .B(G22), .ZN(n943) );
  XNOR2_X1 U1033 ( .A(G23), .B(G1976), .ZN(n942) );
  NOR2_X1 U1034 ( .A1(n943), .A2(n942), .ZN(n945) );
  XOR2_X1 U1035 ( .A(G1986), .B(G24), .Z(n944) );
  NAND2_X1 U1036 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1037 ( .A(KEYINPUT58), .B(n946), .ZN(n947) );
  NOR2_X1 U1038 ( .A1(n948), .A2(n947), .ZN(n952) );
  XNOR2_X1 U1039 ( .A(G1961), .B(G5), .ZN(n950) );
  XNOR2_X1 U1040 ( .A(G1966), .B(G21), .ZN(n949) );
  NOR2_X1 U1041 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1042 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1043 ( .A(n954), .B(n953), .ZN(n955) );
  NAND2_X1 U1044 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1045 ( .A1(n958), .A2(n957), .ZN(n959) );
  NOR2_X1 U1046 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1047 ( .A1(n962), .A2(n961), .ZN(n963) );
  XOR2_X1 U1048 ( .A(KEYINPUT62), .B(n963), .Z(G311) );
  XNOR2_X1 U1049 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1050 ( .A(G120), .ZN(G236) );
  INV_X1 U1051 ( .A(G96), .ZN(G221) );
  INV_X1 U1052 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1053 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1054 ( .A(n966), .B(KEYINPUT106), .ZN(G325) );
  INV_X1 U1055 ( .A(G325), .ZN(G261) );
  INV_X1 U1056 ( .A(n967), .ZN(G319) );
  XOR2_X1 U1057 ( .A(KEYINPUT108), .B(KEYINPUT107), .Z(n969) );
  XNOR2_X1 U1058 ( .A(G2090), .B(G2072), .ZN(n968) );
  XNOR2_X1 U1059 ( .A(n969), .B(n968), .ZN(n973) );
  XOR2_X1 U1060 ( .A(KEYINPUT43), .B(G2678), .Z(n971) );
  XNOR2_X1 U1061 ( .A(G2067), .B(KEYINPUT42), .ZN(n970) );
  XNOR2_X1 U1062 ( .A(n971), .B(n970), .ZN(n972) );
  XOR2_X1 U1063 ( .A(n973), .B(n972), .Z(n975) );
  XNOR2_X1 U1064 ( .A(G2096), .B(G2100), .ZN(n974) );
  XNOR2_X1 U1065 ( .A(n975), .B(n974), .ZN(n977) );
  XOR2_X1 U1066 ( .A(G2078), .B(G2084), .Z(n976) );
  XNOR2_X1 U1067 ( .A(n977), .B(n976), .ZN(G227) );
  XOR2_X1 U1068 ( .A(KEYINPUT41), .B(G1966), .Z(n979) );
  XNOR2_X1 U1069 ( .A(G1996), .B(G1956), .ZN(n978) );
  XNOR2_X1 U1070 ( .A(n979), .B(n978), .ZN(n980) );
  XOR2_X1 U1071 ( .A(n980), .B(G2474), .Z(n982) );
  XNOR2_X1 U1072 ( .A(G1986), .B(G1981), .ZN(n981) );
  XNOR2_X1 U1073 ( .A(n982), .B(n981), .ZN(n986) );
  XOR2_X1 U1074 ( .A(G1976), .B(G1961), .Z(n984) );
  XNOR2_X1 U1075 ( .A(G1991), .B(G1971), .ZN(n983) );
  XNOR2_X1 U1076 ( .A(n984), .B(n983), .ZN(n985) );
  XNOR2_X1 U1077 ( .A(n986), .B(n985), .ZN(G229) );
  NAND2_X1 U1078 ( .A1(G130), .A2(n987), .ZN(n990) );
  NAND2_X1 U1079 ( .A1(G118), .A2(n988), .ZN(n989) );
  NAND2_X1 U1080 ( .A1(n990), .A2(n989), .ZN(n997) );
  NAND2_X1 U1081 ( .A1(G142), .A2(n991), .ZN(n994) );
  NAND2_X1 U1082 ( .A1(G106), .A2(n992), .ZN(n993) );
  NAND2_X1 U1083 ( .A1(n994), .A2(n993), .ZN(n995) );
  XOR2_X1 U1084 ( .A(KEYINPUT45), .B(n995), .Z(n996) );
  NOR2_X1 U1085 ( .A1(n997), .A2(n996), .ZN(n998) );
  XNOR2_X1 U1086 ( .A(G162), .B(n998), .ZN(n1012) );
  XOR2_X1 U1087 ( .A(KEYINPUT46), .B(KEYINPUT111), .Z(n1000) );
  XNOR2_X1 U1088 ( .A(KEYINPUT114), .B(KEYINPUT48), .ZN(n999) );
  XNOR2_X1 U1089 ( .A(n1000), .B(n999), .ZN(n1002) );
  XOR2_X1 U1090 ( .A(n1002), .B(n1001), .Z(n1006) );
  XOR2_X1 U1091 ( .A(n1004), .B(n1003), .Z(n1005) );
  XNOR2_X1 U1092 ( .A(n1006), .B(n1005), .ZN(n1007) );
  XNOR2_X1 U1093 ( .A(G160), .B(n1007), .ZN(n1010) );
  XNOR2_X1 U1094 ( .A(n1008), .B(G164), .ZN(n1009) );
  XNOR2_X1 U1095 ( .A(n1010), .B(n1009), .ZN(n1011) );
  XNOR2_X1 U1096 ( .A(n1012), .B(n1011), .ZN(n1014) );
  XNOR2_X1 U1097 ( .A(n1014), .B(n1013), .ZN(n1015) );
  NOR2_X1 U1098 ( .A1(G37), .A2(n1015), .ZN(G395) );
  XNOR2_X1 U1099 ( .A(KEYINPUT115), .B(n1016), .ZN(n1018) );
  XNOR2_X1 U1100 ( .A(n1018), .B(n1017), .ZN(n1020) );
  XOR2_X1 U1101 ( .A(n1020), .B(n1019), .Z(n1023) );
  XNOR2_X1 U1102 ( .A(G286), .B(n1021), .ZN(n1022) );
  XNOR2_X1 U1103 ( .A(n1023), .B(n1022), .ZN(n1024) );
  NOR2_X1 U1104 ( .A1(G37), .A2(n1024), .ZN(G397) );
  XOR2_X1 U1105 ( .A(G2438), .B(G2435), .Z(n1026) );
  XNOR2_X1 U1106 ( .A(G1341), .B(G2430), .ZN(n1025) );
  XNOR2_X1 U1107 ( .A(n1026), .B(n1025), .ZN(n1027) );
  XOR2_X1 U1108 ( .A(n1027), .B(G2454), .Z(n1029) );
  XNOR2_X1 U1109 ( .A(KEYINPUT104), .B(G2446), .ZN(n1028) );
  XNOR2_X1 U1110 ( .A(n1029), .B(n1028), .ZN(n1033) );
  XOR2_X1 U1111 ( .A(G2443), .B(G2451), .Z(n1031) );
  XNOR2_X1 U1112 ( .A(G1348), .B(G2427), .ZN(n1030) );
  XNOR2_X1 U1113 ( .A(n1031), .B(n1030), .ZN(n1032) );
  XOR2_X1 U1114 ( .A(n1033), .B(n1032), .Z(n1034) );
  NAND2_X1 U1115 ( .A1(G14), .A2(n1034), .ZN(n1040) );
  NAND2_X1 U1116 ( .A1(G319), .A2(n1040), .ZN(n1037) );
  NOR2_X1 U1117 ( .A1(G227), .A2(G229), .ZN(n1035) );
  XNOR2_X1 U1118 ( .A(KEYINPUT49), .B(n1035), .ZN(n1036) );
  NOR2_X1 U1119 ( .A1(n1037), .A2(n1036), .ZN(n1039) );
  NOR2_X1 U1120 ( .A1(G395), .A2(G397), .ZN(n1038) );
  NAND2_X1 U1121 ( .A1(n1039), .A2(n1038), .ZN(G225) );
  INV_X1 U1122 ( .A(G225), .ZN(G308) );
  INV_X1 U1123 ( .A(G108), .ZN(G238) );
  INV_X1 U1124 ( .A(n1040), .ZN(G401) );
endmodule

