//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 1 0 0 1 0 0 0 0 1 1 1 1 0 0 0 0 0 0 1 1 0 1 0 0 0 0 0 1 0 0 0 0 0 0 0 1 0 0 0 0 1 1 0 1 0 1 1 1 0 1 1 1 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:15 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n564, new_n565, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n575, new_n576,
    new_n577, new_n578, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n622, new_n624, new_n625, new_n626,
    new_n627, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n858, new_n859, new_n860, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT65), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n446));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  INV_X1    g023(.A(new_n447), .ZN(new_n449));
  NAND2_X1  g024(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n449), .A2(G2106), .ZN(G217));
  OR4_X1    g026(.A1(G221), .A2(G218), .A3(G220), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(new_n453), .ZN(new_n457));
  INV_X1    g032(.A(new_n454), .ZN(new_n458));
  AOI22_X1  g033(.A1(new_n457), .A2(G2106), .B1(G567), .B2(new_n458), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT67), .ZN(G319));
  NOR2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(G2105), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G137), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  AND2_X1   g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G101), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  XNOR2_X1  g044(.A(KEYINPUT3), .B(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G125), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n466), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n469), .A2(new_n473), .ZN(G160));
  NAND2_X1  g049(.A1(new_n470), .A2(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(KEYINPUT69), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT69), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n470), .A2(new_n477), .A3(G2105), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n476), .A2(G124), .A3(new_n478), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n466), .A2(G112), .ZN(new_n480));
  OAI21_X1  g055(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n464), .B(KEYINPUT68), .ZN(new_n482));
  INV_X1    g057(.A(G136), .ZN(new_n483));
  OAI221_X1 g058(.A(new_n479), .B1(new_n480), .B2(new_n481), .C1(new_n482), .C2(new_n483), .ZN(new_n484));
  XOR2_X1   g059(.A(new_n484), .B(KEYINPUT70), .Z(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  OR2_X1    g061(.A1(G102), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G114), .C2(new_n466), .ZN(new_n488));
  AND2_X1   g063(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n489));
  OAI211_X1 g064(.A(G126), .B(G2105), .C1(new_n489), .C2(new_n461), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  OAI211_X1 g066(.A(G138), .B(new_n466), .C1(new_n489), .C2(new_n461), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(KEYINPUT4), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n470), .A2(new_n494), .A3(G138), .A4(new_n466), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n491), .B1(new_n493), .B2(new_n495), .ZN(G164));
  AND2_X1   g071(.A1(KEYINPUT5), .A2(G543), .ZN(new_n497));
  NOR2_X1   g072(.A1(KEYINPUT5), .A2(G543), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(G62), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(G75), .A2(G543), .ZN(new_n502));
  XNOR2_X1  g077(.A(new_n502), .B(KEYINPUT74), .ZN(new_n503));
  OAI21_X1  g078(.A(G651), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT75), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  OAI211_X1 g081(.A(KEYINPUT75), .B(G651), .C1(new_n501), .C2(new_n503), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AND2_X1   g083(.A1(KEYINPUT71), .A2(KEYINPUT6), .ZN(new_n509));
  NOR2_X1   g084(.A1(KEYINPUT71), .A2(KEYINPUT6), .ZN(new_n510));
  OAI21_X1  g085(.A(G651), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(KEYINPUT72), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT72), .ZN(new_n513));
  OAI211_X1 g088(.A(new_n513), .B(G651), .C1(new_n509), .C2(new_n510), .ZN(new_n514));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n512), .A2(new_n514), .B1(KEYINPUT6), .B2(new_n515), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n516), .A2(G50), .A3(G543), .ZN(new_n517));
  AND2_X1   g092(.A1(new_n508), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n512), .A2(new_n514), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n515), .A2(KEYINPUT6), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n520), .B1(new_n497), .B2(new_n498), .ZN(new_n521));
  INV_X1    g096(.A(new_n521), .ZN(new_n522));
  AOI21_X1  g097(.A(KEYINPUT73), .B1(new_n519), .B2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT73), .ZN(new_n524));
  AOI211_X1 g099(.A(new_n524), .B(new_n521), .C1(new_n512), .C2(new_n514), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G88), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n518), .A2(new_n527), .ZN(G303));
  INV_X1    g103(.A(G303), .ZN(G166));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n530), .B(KEYINPUT7), .ZN(new_n531));
  XNOR2_X1  g106(.A(KEYINPUT5), .B(G543), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n532), .A2(G63), .A3(G651), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  AND3_X1   g109(.A1(new_n519), .A2(G543), .A3(new_n520), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n534), .B1(new_n535), .B2(G51), .ZN(new_n536));
  INV_X1    g111(.A(G89), .ZN(new_n537));
  XNOR2_X1  g112(.A(KEYINPUT71), .B(KEYINPUT6), .ZN(new_n538));
  AOI21_X1  g113(.A(new_n513), .B1(new_n538), .B2(G651), .ZN(new_n539));
  INV_X1    g114(.A(new_n514), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n522), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(new_n524), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n519), .A2(KEYINPUT73), .A3(new_n522), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n536), .B1(new_n537), .B2(new_n544), .ZN(G286));
  INV_X1    g120(.A(G286), .ZN(G168));
  INV_X1    g121(.A(G90), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n519), .A2(G543), .A3(new_n520), .ZN(new_n549));
  INV_X1    g124(.A(G52), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n532), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n551));
  OAI22_X1  g126(.A1(new_n549), .A2(new_n550), .B1(new_n515), .B2(new_n551), .ZN(new_n552));
  OR2_X1    g127(.A1(new_n548), .A2(new_n552), .ZN(G301));
  INV_X1    g128(.A(G301), .ZN(G171));
  NAND2_X1  g129(.A1(new_n526), .A2(G81), .ZN(new_n555));
  NAND2_X1  g130(.A1(G68), .A2(G543), .ZN(new_n556));
  INV_X1    g131(.A(G56), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n556), .B1(new_n499), .B2(new_n557), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n535), .A2(G43), .B1(G651), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n555), .A2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G860), .ZN(G153));
  NAND4_X1  g137(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g138(.A1(G1), .A2(G3), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT8), .ZN(new_n565));
  NAND4_X1  g140(.A1(G319), .A2(G483), .A3(G661), .A4(new_n565), .ZN(G188));
  NAND3_X1  g141(.A1(new_n542), .A2(G91), .A3(new_n543), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n532), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n568));
  OR2_X1    g143(.A1(new_n568), .A2(new_n515), .ZN(new_n569));
  NAND4_X1  g144(.A1(new_n519), .A2(G53), .A3(G543), .A4(new_n520), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT9), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND4_X1  g147(.A1(new_n516), .A2(KEYINPUT9), .A3(G53), .A4(G543), .ZN(new_n573));
  NAND4_X1  g148(.A1(new_n567), .A2(new_n569), .A3(new_n572), .A4(new_n573), .ZN(G299));
  OAI21_X1  g149(.A(G651), .B1(new_n532), .B2(G74), .ZN(new_n575));
  INV_X1    g150(.A(G49), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n549), .B2(new_n576), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n577), .B1(G87), .B2(new_n526), .ZN(new_n578));
  INV_X1    g153(.A(new_n578), .ZN(G288));
  AND2_X1   g154(.A1(G48), .A2(G543), .ZN(new_n580));
  OAI211_X1 g155(.A(new_n520), .B(new_n580), .C1(new_n539), .C2(new_n540), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT76), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n516), .A2(KEYINPUT76), .A3(new_n580), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n526), .A2(G86), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(G73), .A2(G543), .ZN(new_n586));
  INV_X1    g161(.A(G61), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n499), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n588), .A2(G651), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n585), .A2(new_n589), .ZN(G305));
  NAND2_X1  g165(.A1(new_n526), .A2(G85), .ZN(new_n591));
  NAND2_X1  g166(.A1(G72), .A2(G543), .ZN(new_n592));
  INV_X1    g167(.A(G60), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n499), .B2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT77), .ZN(new_n595));
  OR2_X1    g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n515), .B1(new_n594), .B2(new_n595), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n535), .A2(G47), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n591), .A2(new_n598), .ZN(G290));
  NAND2_X1  g174(.A1(G301), .A2(G868), .ZN(new_n600));
  AND3_X1   g175(.A1(new_n516), .A2(G54), .A3(G543), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n532), .A2(G66), .ZN(new_n602));
  NAND2_X1  g177(.A1(G79), .A2(G543), .ZN(new_n603));
  XNOR2_X1  g178(.A(new_n603), .B(KEYINPUT78), .ZN(new_n604));
  AOI21_X1  g179(.A(new_n515), .B1(new_n602), .B2(new_n604), .ZN(new_n605));
  NOR2_X1   g180(.A1(new_n601), .A2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT10), .ZN(new_n608));
  INV_X1    g183(.A(G92), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n544), .B2(new_n609), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n526), .A2(KEYINPUT10), .A3(G92), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n607), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n600), .B1(new_n612), .B2(G868), .ZN(G284));
  XNOR2_X1  g188(.A(G284), .B(KEYINPUT79), .ZN(G321));
  NAND2_X1  g189(.A1(G286), .A2(G868), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n615), .A2(KEYINPUT80), .ZN(new_n616));
  AND2_X1   g191(.A1(new_n615), .A2(KEYINPUT80), .ZN(new_n617));
  INV_X1    g192(.A(G868), .ZN(new_n618));
  NAND2_X1  g193(.A1(G299), .A2(new_n618), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n616), .B1(new_n617), .B2(new_n619), .ZN(G297));
  AOI21_X1  g195(.A(new_n616), .B1(new_n617), .B2(new_n619), .ZN(G280));
  INV_X1    g196(.A(G559), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n612), .B1(new_n622), .B2(G860), .ZN(G148));
  NAND2_X1  g198(.A1(new_n560), .A2(new_n618), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n610), .A2(new_n611), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n625), .A2(new_n606), .ZN(new_n626));
  NOR2_X1   g201(.A1(new_n626), .A2(G559), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n624), .B1(new_n627), .B2(new_n618), .ZN(G323));
  XNOR2_X1  g203(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g204(.A1(new_n476), .A2(G123), .A3(new_n478), .ZN(new_n630));
  NOR2_X1   g205(.A1(new_n466), .A2(G111), .ZN(new_n631));
  OAI21_X1  g206(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n632));
  INV_X1    g207(.A(G135), .ZN(new_n633));
  OAI221_X1 g208(.A(new_n630), .B1(new_n631), .B2(new_n632), .C1(new_n482), .C2(new_n633), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(KEYINPUT82), .Z(new_n635));
  INV_X1    g210(.A(new_n635), .ZN(new_n636));
  INV_X1    g211(.A(G2096), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n635), .A2(G2096), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n470), .A2(new_n467), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT12), .ZN(new_n641));
  XOR2_X1   g216(.A(KEYINPUT81), .B(G2100), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT13), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n641), .B(new_n643), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n638), .A2(new_n639), .A3(new_n644), .ZN(G156));
  XNOR2_X1  g220(.A(KEYINPUT15), .B(G2435), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(G2438), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2427), .B(G2430), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n649), .A2(KEYINPUT14), .ZN(new_n650));
  AND2_X1   g225(.A1(new_n650), .A2(KEYINPUT83), .ZN(new_n651));
  NOR2_X1   g226(.A1(new_n650), .A2(KEYINPUT83), .ZN(new_n652));
  OAI22_X1  g227(.A1(new_n651), .A2(new_n652), .B1(new_n647), .B2(new_n648), .ZN(new_n653));
  XOR2_X1   g228(.A(G2443), .B(G2446), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1341), .B(G1348), .ZN(new_n656));
  OR2_X1    g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n655), .A2(new_n656), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2451), .B(G2454), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT16), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n657), .A2(new_n658), .A3(new_n661), .ZN(new_n664));
  AND3_X1   g239(.A1(new_n663), .A2(G14), .A3(new_n664), .ZN(G401));
  XNOR2_X1  g240(.A(G2067), .B(G2678), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n666), .B(KEYINPUT85), .Z(new_n667));
  XNOR2_X1  g242(.A(G2084), .B(G2090), .ZN(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(new_n669));
  OAI21_X1  g244(.A(KEYINPUT17), .B1(new_n667), .B2(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(G2072), .B(G2078), .Z(new_n671));
  AOI22_X1  g246(.A1(new_n670), .A2(new_n671), .B1(new_n669), .B2(new_n667), .ZN(new_n672));
  OAI21_X1  g247(.A(new_n672), .B1(new_n671), .B2(new_n670), .ZN(new_n673));
  INV_X1    g248(.A(new_n671), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n674), .A2(new_n669), .A3(new_n666), .ZN(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT84), .B(KEYINPUT18), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n673), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(new_n637), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT86), .B(G2100), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(G227));
  XNOR2_X1  g257(.A(G1961), .B(G1966), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT87), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1956), .B(G2474), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1971), .B(G1976), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT19), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT90), .ZN(new_n690));
  OR2_X1    g265(.A1(new_n684), .A2(new_n685), .ZN(new_n691));
  AND2_X1   g266(.A1(new_n686), .A2(new_n688), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n690), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n691), .A2(new_n688), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT89), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT88), .B(KEYINPUT20), .ZN(new_n696));
  AND2_X1   g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n695), .A2(new_n696), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n693), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(KEYINPUT91), .ZN(new_n700));
  INV_X1    g275(.A(KEYINPUT91), .ZN(new_n701));
  OAI211_X1 g276(.A(new_n701), .B(new_n693), .C1(new_n697), .C2(new_n698), .ZN(new_n702));
  XNOR2_X1  g277(.A(G1991), .B(G1996), .ZN(new_n703));
  XNOR2_X1  g278(.A(G1981), .B(G1986), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  XOR2_X1   g280(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n706));
  XOR2_X1   g281(.A(new_n705), .B(new_n706), .Z(new_n707));
  NAND3_X1  g282(.A1(new_n700), .A2(new_n702), .A3(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n707), .B1(new_n700), .B2(new_n702), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(G229));
  INV_X1    g287(.A(G29), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G27), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(G164), .B2(new_n713), .ZN(new_n715));
  XOR2_X1   g290(.A(new_n715), .B(KEYINPUT99), .Z(new_n716));
  INV_X1    g291(.A(G2078), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(G160), .ZN(new_n719));
  INV_X1    g294(.A(KEYINPUT24), .ZN(new_n720));
  AND2_X1   g295(.A1(new_n720), .A2(G34), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n713), .B1(new_n720), .B2(G34), .ZN(new_n722));
  OAI22_X1  g297(.A1(new_n719), .A2(new_n713), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(G2084), .ZN(new_n724));
  OR2_X1    g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n723), .A2(new_n724), .ZN(new_n726));
  INV_X1    g301(.A(G28), .ZN(new_n727));
  OR2_X1    g302(.A1(new_n727), .A2(KEYINPUT30), .ZN(new_n728));
  AOI21_X1  g303(.A(G29), .B1(new_n727), .B2(KEYINPUT30), .ZN(new_n729));
  OR2_X1    g304(.A1(KEYINPUT31), .A2(G11), .ZN(new_n730));
  NAND2_X1  g305(.A1(KEYINPUT31), .A2(G11), .ZN(new_n731));
  AOI22_X1  g306(.A1(new_n728), .A2(new_n729), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n725), .A2(new_n726), .A3(new_n732), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(KEYINPUT25), .Z(new_n735));
  AOI22_X1  g310(.A1(new_n470), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n736));
  INV_X1    g311(.A(G139), .ZN(new_n737));
  OAI221_X1 g312(.A(new_n735), .B1(new_n466), .B2(new_n736), .C1(new_n482), .C2(new_n737), .ZN(new_n738));
  MUX2_X1   g313(.A(G33), .B(new_n738), .S(G29), .Z(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(G2072), .ZN(new_n740));
  AOI211_X1 g315(.A(new_n733), .B(new_n740), .C1(G29), .C2(new_n636), .ZN(new_n741));
  NAND3_X1  g316(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n742));
  INV_X1    g317(.A(KEYINPUT26), .ZN(new_n743));
  OR2_X1    g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n742), .A2(new_n743), .ZN(new_n745));
  AOI22_X1  g320(.A1(new_n744), .A2(new_n745), .B1(G105), .B2(new_n467), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n476), .A2(new_n478), .ZN(new_n747));
  INV_X1    g322(.A(G129), .ZN(new_n748));
  INV_X1    g323(.A(G141), .ZN(new_n749));
  OAI221_X1 g324(.A(new_n746), .B1(new_n747), .B2(new_n748), .C1(new_n482), .C2(new_n749), .ZN(new_n750));
  MUX2_X1   g325(.A(G32), .B(new_n750), .S(G29), .Z(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT27), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(G1996), .ZN(new_n753));
  OR2_X1    g328(.A1(G104), .A2(G2105), .ZN(new_n754));
  OAI211_X1 g329(.A(new_n754), .B(G2104), .C1(G116), .C2(new_n466), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT96), .ZN(new_n756));
  INV_X1    g331(.A(G128), .ZN(new_n757));
  INV_X1    g332(.A(G140), .ZN(new_n758));
  OAI221_X1 g333(.A(new_n756), .B1(new_n747), .B2(new_n757), .C1(new_n482), .C2(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n759), .A2(G29), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n713), .A2(G26), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT28), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(G2067), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  AND3_X1   g340(.A1(new_n741), .A2(new_n753), .A3(new_n765), .ZN(new_n766));
  INV_X1    g341(.A(G16), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n561), .A2(new_n767), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(new_n767), .B2(G19), .ZN(new_n769));
  INV_X1    g344(.A(new_n769), .ZN(new_n770));
  OR2_X1    g345(.A1(new_n770), .A2(G1341), .ZN(new_n771));
  INV_X1    g346(.A(G1966), .ZN(new_n772));
  NOR2_X1   g347(.A1(G168), .A2(new_n767), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(new_n767), .B2(G21), .ZN(new_n774));
  AOI22_X1  g349(.A1(new_n772), .A2(new_n774), .B1(new_n770), .B2(G1341), .ZN(new_n775));
  AND4_X1   g350(.A1(new_n718), .A2(new_n766), .A3(new_n771), .A4(new_n775), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n774), .A2(new_n772), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(KEYINPUT97), .Z(new_n778));
  NAND2_X1  g353(.A1(new_n767), .A2(G5), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G171), .B2(new_n767), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT98), .ZN(new_n781));
  INV_X1    g356(.A(G1961), .ZN(new_n782));
  AND2_X1   g357(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NOR2_X1   g358(.A1(G4), .A2(G16), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(new_n612), .B2(G16), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(G1348), .ZN(new_n786));
  NOR3_X1   g361(.A1(new_n778), .A2(new_n783), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n713), .A2(G35), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G162), .B2(new_n713), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT29), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n790), .A2(G2090), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT100), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n790), .A2(G2090), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n781), .A2(new_n782), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n767), .A2(G20), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(KEYINPUT23), .Z(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(G299), .B2(G16), .ZN(new_n798));
  XOR2_X1   g373(.A(new_n798), .B(G1956), .Z(new_n799));
  NOR3_X1   g374(.A1(new_n794), .A2(new_n795), .A3(new_n799), .ZN(new_n800));
  NAND4_X1  g375(.A1(new_n776), .A2(new_n787), .A3(new_n793), .A4(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n767), .A2(G23), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(new_n578), .B2(new_n767), .ZN(new_n803));
  XOR2_X1   g378(.A(KEYINPUT33), .B(G1976), .Z(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n767), .A2(G6), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n583), .A2(new_n584), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n542), .A2(G86), .A3(new_n543), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(new_n589), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n806), .B1(new_n811), .B2(new_n767), .ZN(new_n812));
  XOR2_X1   g387(.A(KEYINPUT32), .B(G1981), .Z(new_n813));
  INV_X1    g388(.A(new_n813), .ZN(new_n814));
  AND2_X1   g389(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n812), .A2(new_n814), .ZN(new_n816));
  NOR3_X1   g391(.A1(new_n805), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  AND2_X1   g392(.A1(new_n767), .A2(G22), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n818), .B1(G303), .B2(G16), .ZN(new_n819));
  INV_X1    g394(.A(KEYINPUT93), .ZN(new_n820));
  AND2_X1   g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n819), .A2(new_n820), .ZN(new_n822));
  INV_X1    g397(.A(G1971), .ZN(new_n823));
  OR3_X1    g398(.A1(new_n821), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n823), .B1(new_n821), .B2(new_n822), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n817), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n826), .A2(KEYINPUT34), .ZN(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT34), .ZN(new_n829));
  NAND4_X1  g404(.A1(new_n817), .A2(new_n824), .A3(new_n829), .A4(new_n825), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n767), .A2(G24), .ZN(new_n831));
  INV_X1    g406(.A(G290), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n831), .B1(new_n832), .B2(new_n767), .ZN(new_n833));
  AND2_X1   g408(.A1(new_n833), .A2(G1986), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n476), .A2(G119), .A3(new_n478), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n466), .A2(G107), .ZN(new_n836));
  OAI21_X1  g411(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n837));
  INV_X1    g412(.A(G131), .ZN(new_n838));
  OAI221_X1 g413(.A(new_n835), .B1(new_n836), .B2(new_n837), .C1(new_n482), .C2(new_n838), .ZN(new_n839));
  MUX2_X1   g414(.A(G25), .B(new_n839), .S(G29), .Z(new_n840));
  XOR2_X1   g415(.A(KEYINPUT35), .B(G1991), .Z(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT92), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n840), .B(new_n842), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n833), .A2(G1986), .ZN(new_n844));
  NOR3_X1   g419(.A1(new_n834), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n830), .A2(new_n845), .ZN(new_n846));
  OAI21_X1  g421(.A(KEYINPUT95), .B1(new_n828), .B2(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(new_n846), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT95), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n848), .A2(new_n849), .A3(new_n827), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n847), .A2(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT94), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n852), .A2(KEYINPUT36), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(new_n853), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n847), .A2(new_n850), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n801), .B1(new_n854), .B2(new_n856), .ZN(G311));
  AND4_X1   g432(.A1(new_n776), .A2(new_n793), .A3(new_n787), .A4(new_n800), .ZN(new_n858));
  INV_X1    g433(.A(new_n856), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n855), .B1(new_n847), .B2(new_n850), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n858), .B1(new_n859), .B2(new_n860), .ZN(G150));
  AOI22_X1  g436(.A1(new_n532), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n862), .A2(new_n515), .ZN(new_n863));
  OR2_X1    g438(.A1(new_n863), .A2(KEYINPUT101), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(KEYINPUT101), .ZN(new_n865));
  AOI22_X1  g440(.A1(new_n864), .A2(new_n865), .B1(new_n535), .B2(G55), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n526), .A2(G93), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n868), .A2(G860), .ZN(new_n869));
  XOR2_X1   g444(.A(new_n869), .B(KEYINPUT37), .Z(new_n870));
  NOR2_X1   g445(.A1(new_n626), .A2(new_n622), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT38), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n868), .A2(new_n560), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  NAND4_X1  g449(.A1(new_n866), .A2(new_n867), .A3(new_n555), .A4(new_n559), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n872), .B(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT39), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(KEYINPUT102), .ZN(new_n881));
  INV_X1    g456(.A(G860), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n882), .B1(new_n878), .B2(new_n879), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n870), .B1(new_n881), .B2(new_n883), .ZN(G145));
  XNOR2_X1  g459(.A(new_n635), .B(new_n719), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(new_n485), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n750), .B(new_n738), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n476), .A2(G130), .A3(new_n478), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n466), .A2(G118), .ZN(new_n889));
  OAI21_X1  g464(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n890));
  INV_X1    g465(.A(G142), .ZN(new_n891));
  OAI221_X1 g466(.A(new_n888), .B1(new_n889), .B2(new_n890), .C1(new_n482), .C2(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(new_n641), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n887), .B(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n493), .A2(new_n495), .ZN(new_n895));
  AND2_X1   g470(.A1(new_n488), .A2(new_n490), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n759), .B(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n898), .B(new_n839), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n894), .B(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(G37), .B1(new_n886), .B2(new_n900), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n901), .B1(new_n886), .B2(new_n900), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n902), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g478(.A1(G166), .A2(G290), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n832), .A2(G303), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(G305), .A2(new_n578), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n811), .A2(G288), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n906), .A2(new_n909), .ZN(new_n910));
  NAND4_X1  g485(.A1(new_n904), .A2(new_n905), .A3(new_n907), .A4(new_n908), .ZN(new_n911));
  AOI21_X1  g486(.A(KEYINPUT42), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  AND3_X1   g487(.A1(new_n910), .A2(KEYINPUT104), .A3(new_n911), .ZN(new_n913));
  AOI21_X1  g488(.A(KEYINPUT104), .B1(new_n910), .B2(new_n911), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n912), .B1(new_n916), .B2(KEYINPUT42), .ZN(new_n917));
  XOR2_X1   g492(.A(new_n877), .B(new_n627), .Z(new_n918));
  INV_X1    g493(.A(KEYINPUT103), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n626), .A2(new_n919), .A3(G299), .ZN(new_n920));
  AND2_X1   g495(.A1(new_n567), .A2(new_n569), .ZN(new_n921));
  AND2_X1   g496(.A1(new_n572), .A2(new_n573), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n921), .A2(KEYINPUT103), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(G299), .A2(new_n919), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n612), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT41), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n920), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n920), .A2(new_n925), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(KEYINPUT41), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n918), .A2(new_n927), .A3(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n928), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n930), .B1(new_n918), .B2(new_n931), .ZN(new_n932));
  AND2_X1   g507(.A1(new_n917), .A2(new_n932), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n917), .A2(new_n932), .ZN(new_n934));
  OAI21_X1  g509(.A(G868), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n868), .A2(new_n618), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(G295));
  NAND2_X1  g512(.A1(new_n935), .A2(new_n936), .ZN(G331));
  INV_X1    g513(.A(G37), .ZN(new_n939));
  OAI21_X1  g514(.A(G171), .B1(new_n874), .B2(new_n876), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n873), .A2(G301), .A3(new_n875), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n940), .A2(G168), .A3(new_n941), .ZN(new_n942));
  AND3_X1   g517(.A1(new_n873), .A2(G301), .A3(new_n875), .ZN(new_n943));
  AOI21_X1  g518(.A(G301), .B1(new_n873), .B2(new_n875), .ZN(new_n944));
  OAI21_X1  g519(.A(G286), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  AND2_X1   g520(.A1(new_n942), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n929), .A2(new_n927), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n928), .B1(new_n942), .B2(new_n945), .ZN(new_n949));
  INV_X1    g524(.A(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n939), .B1(new_n951), .B2(new_n916), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n928), .A2(KEYINPUT105), .A3(KEYINPUT41), .ZN(new_n953));
  OAI211_X1 g528(.A(new_n946), .B(new_n953), .C1(KEYINPUT105), .C2(new_n947), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n915), .B1(new_n954), .B2(new_n950), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT43), .ZN(new_n956));
  NOR3_X1   g531(.A1(new_n952), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n949), .B1(new_n947), .B2(new_n946), .ZN(new_n958));
  AOI21_X1  g533(.A(G37), .B1(new_n958), .B2(new_n915), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n951), .A2(new_n916), .ZN(new_n960));
  AOI21_X1  g535(.A(KEYINPUT43), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  OAI21_X1  g536(.A(KEYINPUT44), .B1(new_n957), .B2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT44), .ZN(new_n963));
  NOR3_X1   g538(.A1(new_n952), .A2(new_n955), .A3(KEYINPUT43), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n956), .B1(new_n959), .B2(new_n960), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n963), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n962), .A2(new_n966), .ZN(G397));
  INV_X1    g542(.A(KEYINPUT61), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT57), .ZN(new_n969));
  NAND2_X1  g544(.A1(G299), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(KEYINPUT116), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT116), .ZN(new_n972));
  NAND3_X1  g547(.A1(G299), .A2(new_n972), .A3(new_n969), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n921), .A2(KEYINPUT117), .A3(new_n922), .A4(KEYINPUT57), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT117), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n976), .B1(G299), .B2(new_n969), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  AOI22_X1  g553(.A1(new_n464), .A2(G137), .B1(G101), .B2(new_n467), .ZN(new_n979));
  AND2_X1   g554(.A1(new_n471), .A2(new_n472), .ZN(new_n980));
  OAI211_X1 g555(.A(G40), .B(new_n979), .C1(new_n980), .C2(new_n466), .ZN(new_n981));
  INV_X1    g556(.A(G1384), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n897), .A2(new_n982), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n981), .B1(new_n983), .B2(KEYINPUT50), .ZN(new_n984));
  AOI21_X1  g559(.A(G1384), .B1(new_n895), .B2(new_n896), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT50), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n984), .A2(new_n987), .ZN(new_n988));
  XOR2_X1   g563(.A(KEYINPUT115), .B(G1956), .Z(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n985), .A2(KEYINPUT45), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT45), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n992), .B1(G164), .B2(G1384), .ZN(new_n993));
  INV_X1    g568(.A(G40), .ZN(new_n994));
  NOR3_X1   g569(.A1(new_n469), .A2(new_n473), .A3(new_n994), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n991), .A2(new_n993), .A3(new_n995), .ZN(new_n996));
  XNOR2_X1  g571(.A(KEYINPUT118), .B(KEYINPUT56), .ZN(new_n997));
  XNOR2_X1  g572(.A(new_n997), .B(G2072), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n990), .B1(new_n996), .B2(new_n999), .ZN(new_n1000));
  AND3_X1   g575(.A1(new_n974), .A2(new_n978), .A3(new_n1000), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n1000), .B1(new_n974), .B2(new_n978), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n968), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT60), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n983), .A2(new_n981), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(new_n764), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n995), .B1(new_n985), .B2(new_n986), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT108), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n987), .A2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n985), .A2(KEYINPUT108), .A3(new_n986), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1007), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1006), .B1(new_n1011), .B2(G1348), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(new_n612), .ZN(new_n1013));
  AOI21_X1  g588(.A(KEYINPUT108), .B1(new_n985), .B2(new_n986), .ZN(new_n1014));
  NOR4_X1   g589(.A1(G164), .A2(new_n1008), .A3(KEYINPUT50), .A4(G1384), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n984), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(G1348), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n626), .A2(new_n1018), .A3(new_n1006), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1004), .B1(new_n1013), .B2(new_n1019), .ZN(new_n1020));
  XNOR2_X1  g595(.A(KEYINPUT58), .B(G1341), .ZN(new_n1021));
  OAI22_X1  g596(.A1(new_n996), .A2(G1996), .B1(new_n1005), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(KEYINPUT119), .A2(KEYINPUT59), .ZN(new_n1023));
  AND3_X1   g598(.A1(new_n1022), .A2(new_n561), .A3(new_n1023), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1023), .B1(new_n1022), .B2(new_n561), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n612), .A2(new_n1004), .ZN(new_n1026));
  OAI22_X1  g601(.A1(new_n1024), .A2(new_n1025), .B1(new_n1026), .B2(new_n1012), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1020), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1000), .ZN(new_n1029));
  AND2_X1   g604(.A1(new_n975), .A2(new_n977), .ZN(new_n1030));
  AND3_X1   g605(.A1(G299), .A2(new_n972), .A3(new_n969), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n972), .B1(G299), .B2(new_n969), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1029), .B1(new_n1030), .B2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n974), .A2(new_n978), .A3(new_n1000), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1034), .A2(new_n1035), .A3(KEYINPUT61), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1003), .A2(new_n1028), .A3(new_n1036), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1002), .A2(new_n1013), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1038), .A2(new_n1001), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT120), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  XOR2_X1   g617(.A(KEYINPUT109), .B(G8), .Z(new_n1043));
  NOR2_X1   g618(.A1(new_n1005), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(G1976), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1044), .B1(G288), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(KEYINPUT52), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT52), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1048), .B1(new_n578), .B2(G1976), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1047), .B1(new_n1046), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1044), .ZN(new_n1051));
  XOR2_X1   g626(.A(KEYINPUT110), .B(G1981), .Z(new_n1052));
  NAND4_X1  g627(.A1(new_n585), .A2(KEYINPUT111), .A3(new_n589), .A4(new_n1052), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n807), .A2(new_n808), .A3(new_n589), .A4(new_n1052), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT111), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1053), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT112), .ZN(new_n1058));
  AND3_X1   g633(.A1(new_n807), .A2(new_n808), .A3(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1058), .B1(new_n807), .B2(new_n808), .ZN(new_n1060));
  NOR3_X1   g635(.A1(new_n1059), .A2(new_n1060), .A3(new_n810), .ZN(new_n1061));
  INV_X1    g636(.A(G1981), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1057), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT49), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1051), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  OAI211_X1 g640(.A(new_n1057), .B(KEYINPUT49), .C1(new_n1061), .C2(new_n1062), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1050), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n508), .A2(new_n517), .ZN(new_n1068));
  INV_X1    g643(.A(G88), .ZN(new_n1069));
  NOR3_X1   g644(.A1(new_n523), .A2(new_n525), .A3(new_n1069), .ZN(new_n1070));
  OAI21_X1  g645(.A(G8), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT55), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1074));
  INV_X1    g649(.A(new_n987), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1007), .A2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(G2090), .ZN(new_n1077));
  AOI22_X1  g652(.A1(new_n1076), .A2(new_n1077), .B1(new_n823), .B2(new_n996), .ZN(new_n1078));
  OAI211_X1 g653(.A(new_n1073), .B(new_n1074), .C1(new_n1078), .C2(new_n1043), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1074), .A2(new_n1073), .ZN(new_n1080));
  INV_X1    g655(.A(G8), .ZN(new_n1081));
  OAI211_X1 g656(.A(new_n984), .B(new_n1077), .C1(new_n1014), .C2(new_n1015), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n996), .A2(new_n823), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1081), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1080), .A2(new_n1084), .ZN(new_n1085));
  AND2_X1   g660(.A1(new_n1079), .A2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT121), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1043), .ZN(new_n1088));
  AOI21_X1  g663(.A(KEYINPUT51), .B1(G286), .B2(new_n1088), .ZN(new_n1089));
  AOI22_X1  g664(.A1(new_n1011), .A2(new_n724), .B1(new_n772), .B2(new_n996), .ZN(new_n1090));
  OAI211_X1 g665(.A(new_n1087), .B(new_n1089), .C1(new_n1090), .C2(new_n1043), .ZN(new_n1091));
  OAI211_X1 g666(.A(new_n984), .B(new_n724), .C1(new_n1014), .C2(new_n1015), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n996), .A2(new_n772), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1081), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(G286), .A2(new_n1088), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1095), .ZN(new_n1096));
  OAI21_X1  g671(.A(KEYINPUT51), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1043), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT51), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1095), .A2(new_n1099), .ZN(new_n1100));
  OAI21_X1  g675(.A(KEYINPUT121), .B1(new_n1098), .B2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1091), .A2(new_n1097), .A3(new_n1101), .ZN(new_n1102));
  OR2_X1    g677(.A1(new_n1090), .A2(new_n1095), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n991), .A2(new_n993), .A3(new_n717), .A4(new_n995), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT53), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT123), .ZN(new_n1108));
  AOI22_X1  g683(.A1(new_n1107), .A2(new_n1108), .B1(new_n1016), .B2(new_n782), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1105), .A2(KEYINPUT123), .A3(new_n1106), .ZN(new_n1110));
  AND2_X1   g685(.A1(new_n991), .A2(new_n993), .ZN(new_n1111));
  AOI211_X1 g686(.A(new_n1106), .B(G2078), .C1(new_n981), .C2(KEYINPUT125), .ZN(new_n1112));
  OAI211_X1 g687(.A(new_n1111), .B(new_n1112), .C1(KEYINPUT125), .C2(new_n981), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1109), .A2(new_n1110), .A3(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(G171), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1111), .A2(KEYINPUT53), .A3(new_n717), .A4(new_n995), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1109), .A2(G301), .A3(new_n1110), .A4(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1115), .A2(KEYINPUT54), .A3(new_n1117), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1067), .A2(new_n1086), .A3(new_n1104), .A4(new_n1118), .ZN(new_n1119));
  XNOR2_X1  g694(.A(KEYINPUT122), .B(KEYINPUT54), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1016), .A2(new_n782), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1121), .A2(new_n1122), .A3(new_n1110), .A4(new_n1116), .ZN(new_n1123));
  AND3_X1   g698(.A1(new_n1123), .A2(KEYINPUT124), .A3(G171), .ZN(new_n1124));
  AOI21_X1  g699(.A(KEYINPUT124), .B1(new_n1123), .B2(G171), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  OR2_X1    g701(.A1(new_n1114), .A2(G171), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1120), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1119), .A2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1037), .A2(KEYINPUT120), .A3(new_n1039), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1042), .A2(new_n1129), .A3(new_n1130), .ZN(new_n1131));
  XNOR2_X1  g706(.A(new_n1054), .B(KEYINPUT111), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n810), .B1(new_n809), .B2(KEYINPUT112), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n585), .A2(new_n1058), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1062), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1064), .B1(new_n1132), .B2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1136), .A2(new_n1066), .A3(new_n1044), .ZN(new_n1137));
  NOR2_X1   g712(.A1(G288), .A2(G1976), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1139), .A2(new_n1057), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1085), .ZN(new_n1141));
  AOI22_X1  g716(.A1(new_n1140), .A2(new_n1044), .B1(new_n1067), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1050), .ZN(new_n1143));
  AND2_X1   g718(.A1(new_n1098), .A2(G168), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1137), .A2(new_n1086), .A3(new_n1143), .A4(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT63), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT113), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1074), .A2(new_n1073), .A3(new_n1148), .ZN(new_n1149));
  AND2_X1   g724(.A1(new_n1149), .A2(new_n1084), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1149), .A2(new_n1084), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1098), .A2(KEYINPUT63), .A3(G168), .ZN(new_n1152));
  NOR3_X1   g727(.A1(new_n1150), .A2(new_n1151), .A3(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1067), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1147), .A2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT114), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1142), .A2(new_n1155), .A3(new_n1156), .ZN(new_n1157));
  AOI22_X1  g732(.A1(new_n1145), .A2(new_n1146), .B1(new_n1067), .B2(new_n1153), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1132), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1137), .A2(new_n1143), .ZN(new_n1160));
  OAI22_X1  g735(.A1(new_n1159), .A2(new_n1051), .B1(new_n1160), .B2(new_n1085), .ZN(new_n1161));
  OAI21_X1  g736(.A(KEYINPUT114), .B1(new_n1158), .B2(new_n1161), .ZN(new_n1162));
  AND2_X1   g737(.A1(new_n1067), .A2(new_n1086), .ZN(new_n1163));
  OR2_X1    g738(.A1(new_n1104), .A2(KEYINPUT62), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1104), .A2(KEYINPUT62), .ZN(new_n1165));
  INV_X1    g740(.A(new_n1126), .ZN(new_n1166));
  NAND4_X1  g741(.A1(new_n1163), .A2(new_n1164), .A3(new_n1165), .A4(new_n1166), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1131), .A2(new_n1157), .A3(new_n1162), .A4(new_n1167), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n993), .A2(new_n981), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1169), .A2(G1996), .A3(new_n750), .ZN(new_n1170));
  XNOR2_X1  g745(.A(new_n1170), .B(KEYINPUT107), .ZN(new_n1171));
  INV_X1    g746(.A(new_n1169), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1172), .A2(G1996), .ZN(new_n1173));
  XNOR2_X1  g748(.A(new_n1173), .B(KEYINPUT106), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n1174), .A2(new_n750), .ZN(new_n1175));
  XNOR2_X1  g750(.A(new_n759), .B(new_n764), .ZN(new_n1176));
  INV_X1    g751(.A(new_n1176), .ZN(new_n1177));
  AOI211_X1 g752(.A(new_n1171), .B(new_n1175), .C1(new_n1169), .C2(new_n1177), .ZN(new_n1178));
  AND2_X1   g753(.A1(new_n839), .A2(new_n842), .ZN(new_n1179));
  NOR2_X1   g754(.A1(new_n839), .A2(new_n842), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1169), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1178), .A2(new_n1181), .ZN(new_n1182));
  XNOR2_X1  g757(.A(G290), .B(G1986), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1182), .B1(new_n1169), .B2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1168), .A2(new_n1184), .ZN(new_n1185));
  AND2_X1   g760(.A1(new_n1178), .A2(new_n1180), .ZN(new_n1186));
  NOR2_X1   g761(.A1(new_n759), .A2(G2067), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1169), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n1169), .B1(new_n1177), .B2(new_n750), .ZN(new_n1189));
  AND2_X1   g764(.A1(new_n1174), .A2(KEYINPUT46), .ZN(new_n1190));
  NOR2_X1   g765(.A1(new_n1174), .A2(KEYINPUT46), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1189), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  XNOR2_X1  g767(.A(new_n1192), .B(KEYINPUT47), .ZN(new_n1193));
  NOR3_X1   g768(.A1(G290), .A2(new_n1172), .A3(G1986), .ZN(new_n1194));
  XNOR2_X1  g769(.A(KEYINPUT126), .B(KEYINPUT48), .ZN(new_n1195));
  XNOR2_X1  g770(.A(new_n1194), .B(new_n1195), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1178), .A2(new_n1181), .A3(new_n1196), .ZN(new_n1197));
  AND3_X1   g772(.A1(new_n1188), .A2(new_n1193), .A3(new_n1197), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1185), .A2(new_n1198), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g774(.A(KEYINPUT127), .ZN(new_n1201));
  INV_X1    g775(.A(new_n710), .ZN(new_n1202));
  NAND4_X1  g776(.A1(new_n1202), .A2(G319), .A3(new_n681), .A4(new_n708), .ZN(new_n1203));
  OAI21_X1  g777(.A(new_n1201), .B1(new_n1203), .B2(G401), .ZN(new_n1204));
  AND2_X1   g778(.A1(new_n681), .A2(G319), .ZN(new_n1205));
  NAND3_X1  g779(.A1(new_n663), .A2(G14), .A3(new_n664), .ZN(new_n1206));
  NAND4_X1  g780(.A1(new_n711), .A2(new_n1205), .A3(new_n1206), .A4(KEYINPUT127), .ZN(new_n1207));
  NAND2_X1  g781(.A1(new_n1204), .A2(new_n1207), .ZN(new_n1208));
  OAI211_X1 g782(.A(new_n1208), .B(new_n902), .C1(new_n964), .C2(new_n965), .ZN(G225));
  INV_X1    g783(.A(G225), .ZN(G308));
endmodule


