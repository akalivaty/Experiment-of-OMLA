//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 1 0 1 0 0 0 1 1 1 1 1 1 1 0 0 0 0 1 0 0 0 0 1 0 0 0 1 1 0 0 0 1 1 0 1 0 0 0 0 1 1 1 0 0 1 0 0 1 1 0 1 0 0 1 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n708, new_n709, new_n710, new_n711, new_n713, new_n714, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n754, new_n755, new_n756, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n801, new_n802, new_n803, new_n804, new_n806, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n837, new_n838,
    new_n839, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n886, new_n887, new_n889, new_n890, new_n891,
    new_n892, new_n894, new_n895, new_n896, new_n897, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n939, new_n940, new_n941, new_n943, new_n944, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n965, new_n966, new_n967, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n985, new_n986, new_n987,
    new_n988, new_n990, new_n991;
  NOR2_X1   g000(.A1(G71gat), .A2(G78gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT98), .ZN(new_n203));
  INV_X1    g002(.A(G57gat), .ZN(new_n204));
  INV_X1    g003(.A(G64gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(G57gat), .A2(G64gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n206), .A2(KEYINPUT9), .A3(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G71gat), .ZN(new_n209));
  INV_X1    g008(.A(G78gat), .ZN(new_n210));
  OAI211_X1 g009(.A(new_n203), .B(new_n208), .C1(new_n209), .C2(new_n210), .ZN(new_n211));
  XOR2_X1   g010(.A(new_n211), .B(KEYINPUT99), .Z(new_n212));
  NOR2_X1   g011(.A1(new_n209), .A2(new_n210), .ZN(new_n213));
  AOI21_X1  g012(.A(new_n213), .B1(KEYINPUT9), .B2(new_n202), .ZN(new_n214));
  NAND2_X1  g013(.A1(KEYINPUT100), .A2(G57gat), .ZN(new_n215));
  XNOR2_X1  g014(.A(new_n215), .B(new_n205), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n212), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(KEYINPUT21), .ZN(new_n219));
  XNOR2_X1  g018(.A(G15gat), .B(G22gat), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT95), .ZN(new_n221));
  XNOR2_X1  g020(.A(new_n220), .B(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT16), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n223), .A2(G1gat), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(G1gat), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n225), .B1(new_n226), .B2(new_n222), .ZN(new_n227));
  XNOR2_X1  g026(.A(new_n227), .B(G8gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n219), .A2(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n229), .B(G183gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(G231gat), .A2(G233gat), .ZN(new_n231));
  XNOR2_X1  g030(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(G127gat), .B(G155gat), .ZN(new_n233));
  INV_X1    g032(.A(G211gat), .ZN(new_n234));
  XNOR2_X1  g033(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(new_n232), .B(new_n235), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n218), .A2(KEYINPUT21), .ZN(new_n237));
  XNOR2_X1  g036(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g038(.A(new_n236), .B(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT105), .ZN(new_n241));
  NAND2_X1  g040(.A1(G85gat), .A2(G92gat), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n242), .B(KEYINPUT102), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n243), .B(KEYINPUT7), .ZN(new_n244));
  NAND2_X1  g043(.A1(G99gat), .A2(G106gat), .ZN(new_n245));
  INV_X1    g044(.A(G85gat), .ZN(new_n246));
  INV_X1    g045(.A(G92gat), .ZN(new_n247));
  AOI22_X1  g046(.A1(KEYINPUT8), .A2(new_n245), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n244), .A2(new_n248), .ZN(new_n249));
  XOR2_X1   g048(.A(G99gat), .B(G106gat), .Z(new_n250));
  OR2_X1    g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT103), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n249), .A2(new_n250), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n251), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n249), .A2(KEYINPUT103), .A3(new_n250), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT14), .ZN(new_n257));
  INV_X1    g056(.A(G29gat), .ZN(new_n258));
  INV_X1    g057(.A(G36gat), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n257), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  OAI21_X1  g059(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n261));
  AOI22_X1  g060(.A1(new_n260), .A2(new_n261), .B1(G29gat), .B2(G36gat), .ZN(new_n262));
  XNOR2_X1  g061(.A(G43gat), .B(G50gat), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n262), .B1(KEYINPUT15), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(KEYINPUT15), .ZN(new_n265));
  XOR2_X1   g064(.A(new_n264), .B(new_n265), .Z(new_n266));
  NAND2_X1  g065(.A1(new_n256), .A2(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(new_n266), .B(KEYINPUT17), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n268), .A2(new_n255), .A3(new_n254), .ZN(new_n269));
  NAND3_X1  g068(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n267), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(KEYINPUT104), .ZN(new_n272));
  XOR2_X1   g071(.A(G190gat), .B(G218gat), .Z(new_n273));
  INV_X1    g072(.A(KEYINPUT104), .ZN(new_n274));
  NAND4_X1  g073(.A1(new_n267), .A2(new_n269), .A3(new_n274), .A4(new_n270), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n272), .A2(new_n273), .A3(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n273), .B1(new_n272), .B2(new_n275), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n241), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(new_n278), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n280), .A2(KEYINPUT105), .A3(new_n276), .ZN(new_n281));
  AOI21_X1  g080(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n282), .B(KEYINPUT101), .ZN(new_n283));
  XNOR2_X1  g082(.A(G134gat), .B(G162gat), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n283), .B(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n279), .A2(new_n281), .A3(new_n286), .ZN(new_n287));
  OAI211_X1 g086(.A(new_n241), .B(new_n285), .C1(new_n277), .C2(new_n278), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT33), .ZN(new_n291));
  AND2_X1   g090(.A1(KEYINPUT71), .A2(G113gat), .ZN(new_n292));
  NOR2_X1   g091(.A1(KEYINPUT71), .A2(G113gat), .ZN(new_n293));
  OAI21_X1  g092(.A(G120gat), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(G113gat), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n295), .A2(G120gat), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(G127gat), .ZN(new_n298));
  AOI22_X1  g097(.A1(new_n294), .A2(new_n297), .B1(new_n298), .B2(G134gat), .ZN(new_n299));
  INV_X1    g098(.A(G134gat), .ZN(new_n300));
  AOI21_X1  g099(.A(KEYINPUT1), .B1(new_n300), .B2(G127gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n298), .A2(G134gat), .ZN(new_n302));
  XNOR2_X1  g101(.A(KEYINPUT70), .B(G134gat), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n302), .B1(new_n303), .B2(new_n298), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT1), .ZN(new_n305));
  INV_X1    g104(.A(G120gat), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n306), .A2(G113gat), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n305), .B1(new_n296), .B2(new_n307), .ZN(new_n308));
  AOI22_X1  g107(.A1(new_n299), .A2(new_n301), .B1(new_n304), .B2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(G183gat), .A2(G190gat), .ZN(new_n311));
  OR3_X1    g110(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n312));
  OAI21_X1  g111(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n313));
  INV_X1    g112(.A(G169gat), .ZN(new_n314));
  INV_X1    g113(.A(G176gat), .ZN(new_n315));
  OAI211_X1 g114(.A(new_n312), .B(new_n313), .C1(new_n314), .C2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT28), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(KEYINPUT68), .ZN(new_n318));
  XNOR2_X1  g117(.A(KEYINPUT27), .B(G183gat), .ZN(new_n319));
  INV_X1    g118(.A(G190gat), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n318), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  AND2_X1   g120(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n322));
  NOR2_X1   g121(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n323));
  OAI211_X1 g122(.A(new_n318), .B(new_n320), .C1(new_n322), .C2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  OAI211_X1 g124(.A(new_n311), .B(new_n316), .C1(new_n321), .C2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT69), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n320), .B1(new_n322), .B2(new_n323), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n329), .A2(KEYINPUT68), .A3(new_n317), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(new_n324), .ZN(new_n331));
  NAND4_X1  g130(.A1(new_n331), .A2(KEYINPUT69), .A3(new_n311), .A4(new_n316), .ZN(new_n332));
  AND2_X1   g131(.A1(new_n328), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT24), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n311), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n336));
  AND2_X1   g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(G183gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(new_n320), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(KEYINPUT67), .ZN(new_n340));
  OR3_X1    g139(.A1(KEYINPUT67), .A2(G183gat), .A3(G190gat), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n337), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  OAI21_X1  g141(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  NOR3_X1   g143(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n345));
  OAI22_X1  g144(.A1(new_n344), .A2(new_n345), .B1(new_n314), .B2(new_n315), .ZN(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  AND3_X1   g146(.A1(new_n342), .A2(new_n347), .A3(KEYINPUT25), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT25), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT66), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n346), .A2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT65), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n337), .A2(new_n352), .A3(new_n339), .ZN(new_n353));
  OAI221_X1 g152(.A(KEYINPUT66), .B1(new_n314), .B2(new_n315), .C1(new_n344), .C2(new_n345), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n335), .A2(new_n339), .A3(new_n336), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(KEYINPUT65), .ZN(new_n356));
  NAND4_X1  g155(.A1(new_n351), .A2(new_n353), .A3(new_n354), .A4(new_n356), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n348), .B1(new_n349), .B2(new_n357), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n310), .B1(new_n333), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n357), .A2(new_n349), .ZN(new_n360));
  INV_X1    g159(.A(new_n348), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n328), .A2(new_n332), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n362), .A2(new_n309), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n359), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(G227gat), .A2(G233gat), .ZN(new_n366));
  XOR2_X1   g165(.A(new_n366), .B(KEYINPUT64), .Z(new_n367));
  AOI21_X1  g166(.A(KEYINPUT72), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT72), .ZN(new_n369));
  INV_X1    g168(.A(new_n367), .ZN(new_n370));
  AOI211_X1 g169(.A(new_n369), .B(new_n370), .C1(new_n359), .C2(new_n364), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n291), .B1(new_n368), .B2(new_n371), .ZN(new_n372));
  XNOR2_X1  g171(.A(G15gat), .B(G43gat), .ZN(new_n373));
  XNOR2_X1  g172(.A(KEYINPUT73), .B(KEYINPUT74), .ZN(new_n374));
  XNOR2_X1  g173(.A(new_n373), .B(new_n374), .ZN(new_n375));
  XOR2_X1   g174(.A(G71gat), .B(G99gat), .Z(new_n376));
  XOR2_X1   g175(.A(new_n375), .B(new_n376), .Z(new_n377));
  NAND2_X1  g176(.A1(new_n372), .A2(new_n377), .ZN(new_n378));
  OAI21_X1  g177(.A(KEYINPUT32), .B1(new_n368), .B2(new_n371), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n359), .A2(new_n370), .A3(new_n364), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(KEYINPUT34), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT34), .ZN(new_n382));
  NAND4_X1  g181(.A1(new_n359), .A2(new_n382), .A3(new_n364), .A4(new_n370), .ZN(new_n383));
  AND2_X1   g182(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n379), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n381), .A2(new_n383), .ZN(new_n386));
  AND3_X1   g185(.A1(new_n362), .A2(new_n309), .A3(new_n363), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n309), .B1(new_n362), .B2(new_n363), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n367), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(new_n369), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n365), .A2(KEYINPUT72), .A3(new_n367), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n386), .B1(new_n392), .B2(KEYINPUT32), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n378), .B1(new_n385), .B2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(new_n377), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n395), .B1(new_n392), .B2(new_n291), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n379), .A2(new_n384), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n392), .A2(KEYINPUT32), .A3(new_n386), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n396), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  AND3_X1   g198(.A1(new_n394), .A2(KEYINPUT93), .A3(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(KEYINPUT93), .B1(new_n394), .B2(new_n399), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT85), .ZN(new_n403));
  NAND2_X1  g202(.A1(G225gat), .A2(G233gat), .ZN(new_n404));
  NOR2_X1   g203(.A1(G155gat), .A2(G162gat), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT79), .ZN(new_n407));
  NAND2_X1  g206(.A1(G155gat), .A2(G162gat), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  AND2_X1   g208(.A1(G155gat), .A2(G162gat), .ZN(new_n410));
  OAI21_X1  g209(.A(KEYINPUT79), .B1(new_n410), .B2(new_n405), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(G148gat), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(G141gat), .ZN(new_n414));
  INV_X1    g213(.A(G141gat), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(G148gat), .ZN(new_n416));
  AOI22_X1  g215(.A1(new_n414), .A2(new_n416), .B1(KEYINPUT2), .B2(new_n408), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n412), .A2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT81), .ZN(new_n420));
  INV_X1    g219(.A(G155gat), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(KEYINPUT81), .A2(G155gat), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n422), .A2(G162gat), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(KEYINPUT2), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n406), .A2(new_n408), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT80), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n427), .B1(new_n413), .B2(G141gat), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n415), .A2(KEYINPUT80), .A3(G148gat), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n428), .A2(new_n414), .A3(new_n429), .ZN(new_n430));
  AND4_X1   g229(.A1(KEYINPUT82), .A2(new_n425), .A3(new_n426), .A4(new_n430), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n410), .A2(new_n405), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n432), .B1(new_n424), .B2(KEYINPUT2), .ZN(new_n433));
  AOI21_X1  g232(.A(KEYINPUT82), .B1(new_n433), .B2(new_n430), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n419), .B1(new_n431), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(new_n310), .ZN(new_n436));
  OAI211_X1 g235(.A(new_n309), .B(new_n419), .C1(new_n431), .C2(new_n434), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n404), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT4), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  AND2_X1   g239(.A1(KEYINPUT81), .A2(G155gat), .ZN(new_n441));
  NOR2_X1   g240(.A1(KEYINPUT81), .A2(G155gat), .ZN(new_n442));
  INV_X1    g241(.A(G162gat), .ZN(new_n443));
  NOR3_X1   g242(.A1(new_n441), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT2), .ZN(new_n445));
  OAI211_X1 g244(.A(new_n430), .B(new_n426), .C1(new_n444), .C2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT82), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n433), .A2(KEYINPUT82), .A3(new_n430), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n418), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n450), .A2(KEYINPUT4), .A3(new_n309), .ZN(new_n451));
  AND3_X1   g250(.A1(new_n440), .A2(new_n451), .A3(new_n404), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT83), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n435), .A2(new_n453), .A3(KEYINPUT3), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT3), .ZN(new_n455));
  AOI21_X1  g254(.A(KEYINPUT83), .B1(new_n450), .B2(new_n455), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n450), .A2(new_n455), .ZN(new_n457));
  OAI211_X1 g256(.A(new_n310), .B(new_n454), .C1(new_n456), .C2(new_n457), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n438), .B1(new_n452), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(KEYINPUT5), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n440), .A2(new_n451), .A3(new_n404), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n435), .A2(KEYINPUT3), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n435), .A2(KEYINPUT3), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n462), .B1(new_n463), .B2(KEYINPUT83), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n309), .B1(new_n457), .B2(new_n453), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n461), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT5), .ZN(new_n467));
  AOI21_X1  g266(.A(KEYINPUT84), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n452), .A2(new_n458), .A3(KEYINPUT84), .A4(new_n467), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n460), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  XNOR2_X1  g270(.A(KEYINPUT0), .B(G57gat), .ZN(new_n472));
  XNOR2_X1  g271(.A(new_n472), .B(G85gat), .ZN(new_n473));
  XNOR2_X1  g272(.A(G1gat), .B(G29gat), .ZN(new_n474));
  XOR2_X1   g273(.A(new_n473), .B(new_n474), .Z(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n471), .A2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT6), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n403), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n452), .A2(new_n458), .A3(new_n467), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT84), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(new_n469), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n475), .B1(new_n483), .B2(new_n460), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n484), .A2(KEYINPUT85), .A3(KEYINPUT6), .ZN(new_n485));
  AOI22_X1  g284(.A1(new_n482), .A2(new_n469), .B1(KEYINPUT5), .B2(new_n459), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(new_n475), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n477), .A2(new_n487), .A3(new_n478), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n479), .A2(new_n485), .A3(new_n488), .ZN(new_n489));
  XOR2_X1   g288(.A(G78gat), .B(G106gat), .Z(new_n490));
  INV_X1    g289(.A(new_n490), .ZN(new_n491));
  XNOR2_X1  g290(.A(KEYINPUT90), .B(KEYINPUT31), .ZN(new_n492));
  INV_X1    g291(.A(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(G228gat), .ZN(new_n494));
  INV_X1    g293(.A(G233gat), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  XNOR2_X1  g296(.A(G211gat), .B(G218gat), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(G197gat), .A2(G204gat), .ZN(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  NOR2_X1   g300(.A1(G197gat), .A2(G204gat), .ZN(new_n502));
  OAI21_X1  g301(.A(KEYINPUT22), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(G218gat), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n234), .A2(new_n504), .A3(KEYINPUT22), .ZN(new_n505));
  NAND2_X1  g304(.A1(G211gat), .A2(G218gat), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  OR2_X1    g306(.A1(G197gat), .A2(G204gat), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(new_n500), .ZN(new_n509));
  AOI22_X1  g308(.A1(new_n499), .A2(new_n503), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  OAI21_X1  g309(.A(KEYINPUT88), .B1(new_n510), .B2(KEYINPUT29), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT88), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT29), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n498), .B1(new_n509), .B2(KEYINPUT22), .ZN(new_n514));
  AOI22_X1  g313(.A1(new_n505), .A2(new_n506), .B1(new_n508), .B2(new_n500), .ZN(new_n515));
  OAI211_X1 g314(.A(new_n512), .B(new_n513), .C1(new_n514), .C2(new_n515), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n511), .A2(new_n455), .A3(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT89), .ZN(new_n518));
  AND3_X1   g317(.A1(new_n517), .A2(new_n435), .A3(new_n518), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n518), .B1(new_n517), .B2(new_n435), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n510), .B1(new_n463), .B2(KEYINPUT29), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n497), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT86), .ZN(new_n524));
  OR2_X1    g323(.A1(new_n515), .A2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT87), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n514), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n499), .A2(new_n503), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(KEYINPUT87), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n515), .A2(new_n524), .ZN(new_n530));
  NAND4_X1  g329(.A1(new_n525), .A2(new_n527), .A3(new_n529), .A4(new_n530), .ZN(new_n531));
  AOI21_X1  g330(.A(KEYINPUT3), .B1(new_n531), .B2(new_n513), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n497), .B1(new_n532), .B2(new_n450), .ZN(new_n533));
  INV_X1    g332(.A(new_n510), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n450), .A2(new_n455), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n534), .B1(new_n535), .B2(new_n513), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n533), .A2(new_n536), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n493), .B1(new_n523), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n517), .A2(new_n435), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(KEYINPUT89), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n517), .A2(new_n435), .A3(new_n518), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n496), .B1(new_n542), .B2(new_n536), .ZN(new_n543));
  INV_X1    g342(.A(new_n537), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n543), .A2(new_n544), .A3(new_n492), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n491), .B1(new_n538), .B2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(G22gat), .B(G50gat), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n538), .A2(new_n491), .A3(new_n545), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(new_n548), .ZN(new_n551));
  AND3_X1   g350(.A1(new_n538), .A2(new_n491), .A3(new_n545), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n551), .B1(new_n552), .B2(new_n546), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(G8gat), .B(G36gat), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n556), .B(new_n205), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n557), .B(new_n247), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(G226gat), .A2(G233gat), .ZN(new_n560));
  XOR2_X1   g359(.A(new_n560), .B(KEYINPUT75), .Z(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n326), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n358), .A2(new_n563), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n562), .B1(new_n564), .B2(KEYINPUT29), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n562), .B1(new_n362), .B2(new_n363), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n510), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n564), .A2(new_n561), .ZN(new_n569));
  OAI211_X1 g368(.A(new_n513), .B(new_n562), .C1(new_n333), .C2(new_n358), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n534), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  OAI211_X1 g370(.A(KEYINPUT30), .B(new_n559), .C1(new_n568), .C2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT76), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  XOR2_X1   g373(.A(KEYINPUT78), .B(KEYINPUT30), .Z(new_n575));
  NOR2_X1   g374(.A1(new_n568), .A2(new_n571), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n575), .B1(new_n576), .B2(new_n558), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n558), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n569), .A2(new_n570), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(new_n510), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n362), .A2(new_n326), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n561), .B1(new_n581), .B2(new_n513), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n534), .B1(new_n582), .B2(new_n566), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  NAND4_X1  g383(.A1(new_n584), .A2(KEYINPUT76), .A3(KEYINPUT30), .A4(new_n559), .ZN(new_n585));
  NAND4_X1  g384(.A1(new_n574), .A2(new_n577), .A3(new_n578), .A4(new_n585), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n586), .A2(KEYINPUT35), .ZN(new_n587));
  NAND4_X1  g386(.A1(new_n402), .A2(new_n489), .A3(new_n555), .A4(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT94), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n574), .A2(new_n578), .A3(new_n585), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT77), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND4_X1  g391(.A1(new_n574), .A2(new_n585), .A3(KEYINPUT77), .A4(new_n578), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n489), .A2(new_n594), .A3(new_n577), .ZN(new_n595));
  NAND4_X1  g394(.A1(new_n550), .A2(new_n553), .A3(new_n394), .A4(new_n399), .ZN(new_n596));
  OAI211_X1 g395(.A(new_n589), .B(KEYINPUT35), .C1(new_n595), .C2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  AND4_X1   g397(.A1(new_n550), .A2(new_n553), .A3(new_n394), .A4(new_n399), .ZN(new_n599));
  NAND4_X1  g398(.A1(new_n599), .A2(new_n489), .A3(new_n577), .A4(new_n594), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n589), .B1(new_n600), .B2(KEYINPUT35), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n588), .B1(new_n598), .B2(new_n601), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n565), .A2(new_n510), .A3(new_n567), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n569), .A2(new_n534), .A3(new_n570), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n603), .A2(KEYINPUT37), .A3(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT38), .ZN(new_n606));
  AND3_X1   g405(.A1(new_n605), .A2(new_n606), .A3(new_n558), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT37), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n584), .A2(new_n608), .ZN(new_n609));
  AOI22_X1  g408(.A1(new_n607), .A2(new_n609), .B1(new_n584), .B2(new_n559), .ZN(new_n610));
  NAND4_X1  g409(.A1(new_n479), .A2(new_n488), .A3(new_n485), .A4(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT91), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  AOI21_X1  g412(.A(KEYINPUT85), .B1(new_n484), .B2(KEYINPUT6), .ZN(new_n614));
  NOR4_X1   g413(.A1(new_n486), .A2(new_n403), .A3(new_n478), .A4(new_n475), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND4_X1  g415(.A1(new_n616), .A2(KEYINPUT91), .A3(new_n488), .A4(new_n610), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n559), .B1(new_n576), .B2(KEYINPUT37), .ZN(new_n618));
  OR2_X1    g417(.A1(new_n618), .A2(KEYINPUT92), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(KEYINPUT92), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n619), .A2(new_n620), .A3(new_n609), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n621), .A2(KEYINPUT38), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n613), .A2(new_n617), .A3(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT39), .ZN(new_n624));
  AND2_X1   g423(.A1(new_n440), .A2(new_n451), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n404), .B1(new_n458), .B2(new_n625), .ZN(new_n626));
  AND2_X1   g425(.A1(new_n436), .A2(new_n437), .ZN(new_n627));
  AOI211_X1 g426(.A(new_n624), .B(new_n626), .C1(new_n404), .C2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT40), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n626), .A2(new_n624), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n630), .A2(new_n475), .ZN(new_n631));
  OR3_X1    g430(.A1(new_n628), .A2(new_n629), .A3(new_n631), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n629), .B1(new_n628), .B2(new_n631), .ZN(new_n633));
  NAND4_X1  g432(.A1(new_n632), .A2(new_n477), .A3(new_n633), .A4(new_n586), .ZN(new_n634));
  AND2_X1   g433(.A1(new_n555), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n623), .A2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT36), .ZN(new_n637));
  INV_X1    g436(.A(new_n394), .ZN(new_n638));
  INV_X1    g437(.A(new_n399), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n637), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n394), .A2(KEYINPUT36), .A3(new_n399), .ZN(new_n641));
  AOI22_X1  g440(.A1(new_n595), .A2(new_n554), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n636), .A2(new_n642), .ZN(new_n643));
  AOI211_X1 g442(.A(new_n240), .B(new_n290), .C1(new_n602), .C2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n266), .ZN(new_n645));
  AOI21_X1  g444(.A(KEYINPUT96), .B1(new_n228), .B2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(G8gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n227), .B(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n648), .A2(new_n266), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(G229gat), .A2(G233gat), .ZN(new_n651));
  XOR2_X1   g450(.A(new_n651), .B(KEYINPUT13), .Z(new_n652));
  NAND3_X1  g451(.A1(new_n648), .A2(KEYINPUT96), .A3(new_n266), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n650), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n268), .A2(new_n228), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n655), .A2(new_n649), .A3(new_n651), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT18), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND4_X1  g457(.A1(new_n655), .A2(new_n649), .A3(KEYINPUT18), .A4(new_n651), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n654), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  XNOR2_X1  g459(.A(KEYINPUT11), .B(G169gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(G197gat), .ZN(new_n662));
  XOR2_X1   g461(.A(G113gat), .B(G141gat), .Z(new_n663));
  XNOR2_X1  g462(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(KEYINPUT12), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n660), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT97), .ZN(new_n668));
  NAND4_X1  g467(.A1(new_n654), .A2(new_n658), .A3(new_n665), .A4(new_n659), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n667), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n660), .A2(KEYINPUT97), .A3(new_n666), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(G230gat), .A2(G233gat), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT10), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT106), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n251), .A2(new_n676), .A3(new_n253), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n249), .A2(KEYINPUT106), .A3(new_n250), .ZN(new_n678));
  AND3_X1   g477(.A1(new_n677), .A2(new_n218), .A3(new_n678), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n218), .B1(new_n254), .B2(new_n255), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n675), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n256), .A2(KEYINPUT10), .A3(new_n218), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n674), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  OR3_X1    g483(.A1(new_n679), .A2(new_n680), .A3(new_n673), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g485(.A(G120gat), .B(G148gat), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(new_n315), .ZN(new_n688));
  INV_X1    g487(.A(G204gat), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n688), .B(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n686), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n690), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n684), .A2(new_n685), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n672), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n644), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n696), .A2(new_n489), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n697), .B(new_n226), .ZN(G1324gat));
  INV_X1    g497(.A(new_n586), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n223), .A2(new_n647), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n700), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT42), .ZN(new_n704));
  OR2_X1    g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n703), .A2(new_n704), .ZN(new_n706));
  OAI211_X1 g505(.A(new_n705), .B(new_n706), .C1(new_n647), .C2(new_n700), .ZN(G1325gat));
  INV_X1    g506(.A(G15gat), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n640), .A2(new_n641), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n696), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n644), .A2(new_n402), .A3(new_n695), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n710), .B1(new_n708), .B2(new_n711), .ZN(G1326gat));
  NOR2_X1   g511(.A1(new_n696), .A2(new_n555), .ZN(new_n713));
  XOR2_X1   g512(.A(KEYINPUT43), .B(G22gat), .Z(new_n714));
  XNOR2_X1  g513(.A(new_n713), .B(new_n714), .ZN(G1327gat));
  AOI21_X1  g514(.A(new_n289), .B1(new_n602), .B2(new_n643), .ZN(new_n716));
  AND3_X1   g515(.A1(new_n716), .A2(new_n240), .A3(new_n695), .ZN(new_n717));
  INV_X1    g516(.A(new_n489), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n717), .A2(new_n258), .A3(new_n718), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n719), .B(KEYINPUT107), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(KEYINPUT45), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT110), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT109), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n643), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n636), .A2(KEYINPUT109), .A3(new_n642), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n724), .A2(new_n602), .A3(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT44), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n726), .A2(new_n727), .A3(new_n290), .ZN(new_n728));
  INV_X1    g527(.A(new_n588), .ZN(new_n729));
  OAI21_X1  g528(.A(KEYINPUT35), .B1(new_n595), .B2(new_n596), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(KEYINPUT94), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n729), .B1(new_n731), .B2(new_n597), .ZN(new_n732));
  AND2_X1   g531(.A1(new_n636), .A2(new_n642), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n290), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(KEYINPUT44), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n728), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n694), .B(KEYINPUT108), .ZN(new_n737));
  INV_X1    g536(.A(new_n737), .ZN(new_n738));
  AND2_X1   g537(.A1(new_n670), .A2(new_n671), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n240), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(new_n740), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n722), .B1(new_n736), .B2(new_n741), .ZN(new_n742));
  AOI211_X1 g541(.A(KEYINPUT110), .B(new_n740), .C1(new_n728), .C2(new_n735), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  OAI21_X1  g543(.A(KEYINPUT111), .B1(new_n744), .B2(new_n489), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n736), .A2(new_n741), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(KEYINPUT110), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n736), .A2(new_n722), .A3(new_n741), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT111), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n749), .A2(new_n750), .A3(new_n718), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n745), .A2(new_n751), .A3(G29gat), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n721), .A2(new_n752), .ZN(G1328gat));
  OAI21_X1  g552(.A(G36gat), .B1(new_n744), .B2(new_n699), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n717), .A2(new_n259), .A3(new_n586), .ZN(new_n755));
  XOR2_X1   g554(.A(KEYINPUT112), .B(KEYINPUT46), .Z(new_n756));
  XNOR2_X1  g555(.A(new_n755), .B(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n754), .A2(new_n757), .ZN(G1329gat));
  INV_X1    g557(.A(KEYINPUT113), .ZN(new_n759));
  OAI21_X1  g558(.A(G43gat), .B1(new_n746), .B2(new_n709), .ZN(new_n760));
  INV_X1    g559(.A(G43gat), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n717), .A2(new_n761), .A3(new_n402), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(KEYINPUT47), .ZN(new_n764));
  INV_X1    g563(.A(new_n709), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n761), .B1(new_n749), .B2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT47), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n762), .A2(new_n767), .ZN(new_n768));
  OAI211_X1 g567(.A(new_n759), .B(new_n764), .C1(new_n766), .C2(new_n768), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n765), .B1(new_n742), .B2(new_n743), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n768), .B1(new_n770), .B2(G43gat), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n767), .B1(new_n760), .B2(new_n762), .ZN(new_n772));
  OAI21_X1  g571(.A(KEYINPUT113), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n769), .A2(new_n773), .ZN(G1330gat));
  INV_X1    g573(.A(new_n717), .ZN(new_n775));
  NOR3_X1   g574(.A1(new_n775), .A2(G50gat), .A3(new_n555), .ZN(new_n776));
  INV_X1    g575(.A(new_n776), .ZN(new_n777));
  OAI21_X1  g576(.A(G50gat), .B1(new_n746), .B2(new_n555), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n777), .A2(KEYINPUT48), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n749), .A2(new_n554), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n776), .B1(new_n780), .B2(G50gat), .ZN(new_n781));
  XOR2_X1   g580(.A(KEYINPUT114), .B(KEYINPUT48), .Z(new_n782));
  OAI21_X1  g581(.A(new_n779), .B1(new_n781), .B2(new_n782), .ZN(G1331gat));
  NOR3_X1   g582(.A1(new_n240), .A2(new_n290), .A3(new_n739), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n726), .A2(new_n737), .A3(new_n784), .ZN(new_n785));
  OR2_X1    g584(.A1(new_n785), .A2(KEYINPUT115), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(KEYINPUT115), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n788), .A2(new_n489), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n789), .B(new_n204), .ZN(G1332gat));
  INV_X1    g589(.A(KEYINPUT49), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n791), .A2(new_n205), .ZN(new_n792));
  INV_X1    g591(.A(new_n792), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n786), .A2(new_n586), .A3(new_n787), .A4(new_n793), .ZN(new_n794));
  AND2_X1   g593(.A1(new_n794), .A2(KEYINPUT116), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n794), .A2(KEYINPUT116), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n791), .A2(new_n205), .ZN(new_n797));
  OR3_X1    g596(.A1(new_n795), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n797), .B1(new_n795), .B2(new_n796), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(new_n799), .ZN(G1333gat));
  INV_X1    g599(.A(new_n402), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n209), .B1(new_n788), .B2(new_n801), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n786), .A2(G71gat), .A3(new_n765), .A4(new_n787), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  XNOR2_X1  g603(.A(new_n804), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g604(.A1(new_n788), .A2(new_n555), .ZN(new_n806));
  XNOR2_X1  g605(.A(new_n806), .B(new_n210), .ZN(G1335gat));
  NAND2_X1  g606(.A1(new_n240), .A2(new_n672), .ZN(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n736), .A2(new_n694), .A3(new_n809), .ZN(new_n810));
  OAI21_X1  g609(.A(KEYINPUT117), .B1(new_n810), .B2(new_n489), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n808), .B1(new_n728), .B2(new_n735), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT117), .ZN(new_n813));
  NAND4_X1  g612(.A1(new_n812), .A2(new_n813), .A3(new_n718), .A4(new_n694), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n811), .A2(G85gat), .A3(new_n814), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n489), .A2(G85gat), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n726), .A2(new_n290), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n808), .B1(new_n817), .B2(KEYINPUT118), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT118), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n726), .A2(new_n819), .A3(new_n290), .ZN(new_n820));
  AND3_X1   g619(.A1(new_n818), .A2(KEYINPUT51), .A3(new_n820), .ZN(new_n821));
  AOI21_X1  g620(.A(KEYINPUT51), .B1(new_n818), .B2(new_n820), .ZN(new_n822));
  OAI211_X1 g621(.A(new_n694), .B(new_n816), .C1(new_n821), .C2(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n815), .A2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT119), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n815), .A2(KEYINPUT119), .A3(new_n823), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(G1336gat));
  NOR2_X1   g627(.A1(new_n699), .A2(G92gat), .ZN(new_n829));
  OAI211_X1 g628(.A(new_n737), .B(new_n829), .C1(new_n821), .C2(new_n822), .ZN(new_n830));
  OAI21_X1  g629(.A(G92gat), .B1(new_n810), .B2(new_n699), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(KEYINPUT52), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT52), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n830), .A2(new_n834), .A3(new_n831), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n833), .A2(new_n835), .ZN(G1337gat));
  OAI21_X1  g635(.A(G99gat), .B1(new_n810), .B2(new_n709), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n694), .B1(new_n821), .B2(new_n822), .ZN(new_n838));
  OR2_X1    g637(.A1(new_n801), .A2(G99gat), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n837), .B1(new_n838), .B2(new_n839), .ZN(G1338gat));
  NOR2_X1   g639(.A1(new_n555), .A2(G106gat), .ZN(new_n841));
  OAI211_X1 g640(.A(new_n737), .B(new_n841), .C1(new_n821), .C2(new_n822), .ZN(new_n842));
  OAI21_X1  g641(.A(G106gat), .B1(new_n810), .B2(new_n555), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(KEYINPUT53), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT53), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n842), .A2(new_n846), .A3(new_n843), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n845), .A2(new_n847), .ZN(G1339gat));
  NOR4_X1   g647(.A1(new_n240), .A2(new_n290), .A3(new_n694), .A4(new_n739), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n681), .A2(new_n674), .A3(new_n682), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n684), .A2(KEYINPUT54), .A3(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT54), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n692), .B1(new_n683), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT55), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(new_n669), .ZN(new_n857));
  AND2_X1   g656(.A1(new_n650), .A2(new_n653), .ZN(new_n858));
  AND2_X1   g657(.A1(new_n655), .A2(new_n649), .ZN(new_n859));
  OAI22_X1  g658(.A1(new_n858), .A2(new_n652), .B1(new_n651), .B2(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n857), .B1(new_n664), .B2(new_n860), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n851), .A2(KEYINPUT55), .A3(new_n853), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n856), .A2(new_n861), .A3(new_n693), .A4(new_n862), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n863), .A2(new_n289), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT120), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n694), .A2(new_n861), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n856), .A2(new_n693), .A3(new_n862), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n867), .B1(new_n868), .B2(new_n672), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(new_n289), .ZN(new_n870));
  OAI21_X1  g669(.A(KEYINPUT120), .B1(new_n863), .B2(new_n289), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n866), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n849), .B1(new_n240), .B2(new_n872), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n489), .A2(new_n586), .ZN(new_n874));
  INV_X1    g673(.A(new_n874), .ZN(new_n875));
  NOR3_X1   g674(.A1(new_n873), .A2(new_n596), .A3(new_n875), .ZN(new_n876));
  OAI211_X1 g675(.A(new_n876), .B(new_n739), .C1(new_n293), .C2(new_n292), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n872), .A2(new_n240), .ZN(new_n878));
  INV_X1    g677(.A(new_n694), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n784), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n801), .A2(new_n554), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NOR3_X1   g682(.A1(new_n883), .A2(new_n672), .A3(new_n875), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n877), .B1(new_n884), .B2(new_n295), .ZN(G1340gat));
  NAND3_X1  g684(.A1(new_n876), .A2(new_n306), .A3(new_n694), .ZN(new_n886));
  NOR3_X1   g685(.A1(new_n883), .A2(new_n738), .A3(new_n875), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n886), .B1(new_n887), .B2(new_n306), .ZN(G1341gat));
  INV_X1    g687(.A(new_n240), .ZN(new_n889));
  AOI21_X1  g688(.A(G127gat), .B1(new_n876), .B2(new_n889), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n883), .A2(new_n875), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n240), .A2(new_n298), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n890), .B1(new_n891), .B2(new_n892), .ZN(G1342gat));
  INV_X1    g692(.A(new_n303), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n876), .A2(new_n894), .A3(new_n290), .ZN(new_n895));
  XNOR2_X1  g694(.A(new_n895), .B(KEYINPUT56), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n300), .B1(new_n891), .B2(new_n290), .ZN(new_n897));
  OR2_X1    g696(.A1(new_n896), .A2(new_n897), .ZN(G1343gat));
  AOI21_X1  g697(.A(new_n555), .B1(new_n878), .B2(new_n880), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n765), .A2(new_n875), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n415), .B1(new_n901), .B2(new_n672), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n854), .A2(KEYINPUT121), .A3(new_n855), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n739), .A2(new_n903), .A3(new_n693), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n854), .B1(KEYINPUT121), .B2(new_n855), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n867), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(new_n289), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n907), .A2(new_n871), .A3(new_n866), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n849), .B1(new_n908), .B2(new_n240), .ZN(new_n909));
  OAI21_X1  g708(.A(KEYINPUT57), .B1(new_n909), .B2(new_n555), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT57), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n899), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n910), .A2(new_n912), .A3(new_n900), .ZN(new_n913));
  OR2_X1    g712(.A1(new_n913), .A2(new_n415), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n902), .B1(new_n914), .B2(new_n672), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT58), .ZN(new_n916));
  XNOR2_X1  g715(.A(new_n915), .B(new_n916), .ZN(G1344gat));
  OR2_X1    g716(.A1(new_n863), .A2(new_n289), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n889), .B1(new_n907), .B2(new_n918), .ZN(new_n919));
  OAI211_X1 g718(.A(new_n911), .B(new_n554), .C1(new_n919), .C2(new_n849), .ZN(new_n920));
  NOR3_X1   g719(.A1(new_n765), .A2(new_n875), .A3(new_n879), .ZN(new_n921));
  OAI211_X1 g720(.A(new_n920), .B(new_n921), .C1(new_n899), .C2(new_n911), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(KEYINPUT123), .ZN(new_n923));
  OAI21_X1  g722(.A(KEYINPUT57), .B1(new_n873), .B2(new_n555), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT123), .ZN(new_n925));
  NAND4_X1  g724(.A1(new_n924), .A2(new_n925), .A3(new_n920), .A4(new_n921), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n923), .A2(G148gat), .A3(new_n926), .ZN(new_n927));
  AND3_X1   g726(.A1(new_n927), .A2(KEYINPUT124), .A3(KEYINPUT59), .ZN(new_n928));
  AOI21_X1  g727(.A(KEYINPUT124), .B1(new_n927), .B2(KEYINPUT59), .ZN(new_n929));
  NAND4_X1  g728(.A1(new_n910), .A2(new_n912), .A3(new_n694), .A4(new_n900), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT59), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n930), .A2(new_n931), .A3(G148gat), .ZN(new_n932));
  AND2_X1   g731(.A1(new_n932), .A2(KEYINPUT122), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n932), .A2(KEYINPUT122), .ZN(new_n934));
  OAI22_X1  g733(.A1(new_n928), .A2(new_n929), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g734(.A(new_n901), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n936), .A2(new_n413), .A3(new_n694), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n935), .A2(new_n937), .ZN(G1345gat));
  NOR2_X1   g737(.A1(new_n441), .A2(new_n442), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n939), .B1(new_n936), .B2(new_n889), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n913), .A2(new_n240), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n940), .B1(new_n941), .B2(new_n939), .ZN(G1346gat));
  AOI21_X1  g741(.A(G162gat), .B1(new_n936), .B2(new_n290), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n913), .A2(new_n443), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n943), .B1(new_n944), .B2(new_n290), .ZN(G1347gat));
  NOR2_X1   g744(.A1(new_n718), .A2(new_n699), .ZN(new_n946));
  INV_X1    g745(.A(new_n946), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n883), .A2(new_n947), .ZN(new_n948));
  INV_X1    g747(.A(new_n948), .ZN(new_n949));
  OAI21_X1  g748(.A(G169gat), .B1(new_n949), .B2(new_n672), .ZN(new_n950));
  NOR3_X1   g749(.A1(new_n873), .A2(new_n596), .A3(new_n947), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n951), .A2(new_n314), .A3(new_n739), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n950), .A2(new_n952), .ZN(G1348gat));
  AOI21_X1  g752(.A(G176gat), .B1(new_n951), .B2(new_n694), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n949), .A2(new_n315), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n954), .B1(new_n955), .B2(new_n737), .ZN(G1349gat));
  NAND3_X1  g755(.A1(new_n951), .A2(new_n889), .A3(new_n319), .ZN(new_n957));
  NOR3_X1   g756(.A1(new_n883), .A2(new_n240), .A3(new_n947), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n957), .B1(new_n958), .B2(new_n338), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n959), .A2(KEYINPUT125), .ZN(new_n960));
  INV_X1    g759(.A(KEYINPUT125), .ZN(new_n961));
  OAI211_X1 g760(.A(new_n957), .B(new_n961), .C1(new_n958), .C2(new_n338), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  XNOR2_X1  g762(.A(new_n963), .B(KEYINPUT60), .ZN(G1350gat));
  AOI21_X1  g763(.A(new_n320), .B1(new_n948), .B2(new_n290), .ZN(new_n965));
  XOR2_X1   g764(.A(new_n965), .B(KEYINPUT61), .Z(new_n966));
  NAND3_X1  g765(.A1(new_n951), .A2(new_n320), .A3(new_n290), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n966), .A2(new_n967), .ZN(G1351gat));
  XOR2_X1   g767(.A(KEYINPUT126), .B(G197gat), .Z(new_n969));
  AND2_X1   g768(.A1(new_n924), .A2(new_n920), .ZN(new_n970));
  NOR2_X1   g769(.A1(new_n947), .A2(new_n765), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n969), .B1(new_n972), .B2(new_n672), .ZN(new_n973));
  AND2_X1   g772(.A1(new_n899), .A2(new_n971), .ZN(new_n974));
  INV_X1    g773(.A(new_n969), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n974), .A2(new_n739), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n973), .A2(new_n976), .ZN(G1352gat));
  NAND3_X1  g776(.A1(new_n974), .A2(new_n689), .A3(new_n694), .ZN(new_n978));
  NOR2_X1   g777(.A1(new_n978), .A2(KEYINPUT62), .ZN(new_n979));
  OR2_X1    g778(.A1(new_n979), .A2(KEYINPUT127), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n978), .A2(KEYINPUT62), .ZN(new_n981));
  OAI21_X1  g780(.A(G204gat), .B1(new_n972), .B2(new_n738), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n979), .A2(KEYINPUT127), .ZN(new_n983));
  NAND4_X1  g782(.A1(new_n980), .A2(new_n981), .A3(new_n982), .A4(new_n983), .ZN(G1353gat));
  NAND3_X1  g783(.A1(new_n974), .A2(new_n234), .A3(new_n889), .ZN(new_n985));
  NAND3_X1  g784(.A1(new_n970), .A2(new_n889), .A3(new_n971), .ZN(new_n986));
  AND3_X1   g785(.A1(new_n986), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n987));
  AOI21_X1  g786(.A(KEYINPUT63), .B1(new_n986), .B2(G211gat), .ZN(new_n988));
  OAI21_X1  g787(.A(new_n985), .B1(new_n987), .B2(new_n988), .ZN(G1354gat));
  OAI21_X1  g788(.A(G218gat), .B1(new_n972), .B2(new_n289), .ZN(new_n990));
  NAND3_X1  g789(.A1(new_n974), .A2(new_n504), .A3(new_n290), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n990), .A2(new_n991), .ZN(G1355gat));
endmodule


