//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 1 0 1 1 1 1 1 0 1 0 0 0 0 0 1 1 0 0 0 0 0 0 1 0 1 1 0 1 0 0 0 0 0 0 0 0 0 0 0 0 1 0 1 1 0 1 1 0 1 0 0 0 0 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:21 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1272, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355, new_n1356, new_n1357, new_n1358, new_n1359;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G68), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n206), .B(KEYINPUT64), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G68), .A2(G238), .B1(G107), .B2(G264), .ZN(new_n208));
  INV_X1    g0008(.A(G226), .ZN(new_n209));
  INV_X1    g0009(.A(G87), .ZN(new_n210));
  INV_X1    g0010(.A(G250), .ZN(new_n211));
  OAI221_X1 g0011(.A(new_n208), .B1(new_n201), .B2(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n207), .B1(new_n212), .B2(new_n215), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT1), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n207), .A2(G13), .ZN(new_n218));
  OAI211_X1 g0018(.A(new_n218), .B(G250), .C1(G257), .C2(G264), .ZN(new_n219));
  XOR2_X1   g0019(.A(new_n219), .B(KEYINPUT0), .Z(new_n220));
  NAND2_X1  g0020(.A1(G1), .A2(G13), .ZN(new_n221));
  INV_X1    g0021(.A(G20), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(G68), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n202), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n225), .A2(G50), .ZN(new_n226));
  INV_X1    g0026(.A(new_n226), .ZN(new_n227));
  AOI211_X1 g0027(.A(new_n217), .B(new_n220), .C1(new_n223), .C2(new_n227), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  INV_X1    g0029(.A(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(KEYINPUT2), .B(G226), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XOR2_X1   g0037(.A(G87), .B(G97), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT66), .ZN(new_n239));
  XOR2_X1   g0039(.A(G107), .B(G116), .Z(new_n240));
  XOR2_X1   g0040(.A(new_n239), .B(new_n240), .Z(new_n241));
  XNOR2_X1  g0041(.A(G68), .B(G77), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT65), .ZN(new_n243));
  XOR2_X1   g0043(.A(G50), .B(G58), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n241), .B(new_n245), .ZN(G351));
  INV_X1    g0046(.A(G41), .ZN(new_n247));
  INV_X1    g0047(.A(G45), .ZN(new_n248));
  AOI21_X1  g0048(.A(G1), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g0049(.A1(G33), .A2(G41), .ZN(new_n250));
  NAND3_X1  g0050(.A1(new_n250), .A2(G1), .A3(G13), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n249), .A2(new_n251), .A3(G274), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G1), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n254), .B1(G41), .B2(G45), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n251), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n253), .B1(G226), .B2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  XNOR2_X1  g0059(.A(KEYINPUT3), .B(G33), .ZN(new_n260));
  INV_X1    g0060(.A(G1698), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G222), .ZN(new_n263));
  OAI21_X1  g0063(.A(KEYINPUT67), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT67), .ZN(new_n265));
  NAND4_X1  g0065(.A1(new_n260), .A2(new_n265), .A3(G222), .A4(new_n261), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n260), .A2(G1698), .ZN(new_n268));
  INV_X1    g0068(.A(G223), .ZN(new_n269));
  INV_X1    g0069(.A(G77), .ZN(new_n270));
  OAI22_X1  g0070(.A1(new_n268), .A2(new_n269), .B1(new_n270), .B2(new_n260), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n267), .A2(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n221), .B1(G33), .B2(G41), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n259), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G179), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n271), .B1(new_n266), .B2(new_n264), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n258), .B1(new_n278), .B2(new_n251), .ZN(new_n279));
  INV_X1    g0079(.A(G169), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(new_n221), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n202), .A2(KEYINPUT8), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT8), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(G58), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n222), .A2(G33), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  NOR2_X1   g0090(.A1(G20), .A2(G33), .ZN(new_n291));
  AOI22_X1  g0091(.A1(new_n288), .A2(new_n290), .B1(G150), .B2(new_n291), .ZN(new_n292));
  OAI21_X1  g0092(.A(G20), .B1(new_n203), .B2(G68), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n284), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n254), .A2(G13), .A3(G20), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n284), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n254), .A2(G20), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(G50), .ZN(new_n298));
  OAI22_X1  g0098(.A1(new_n296), .A2(new_n298), .B1(G50), .B2(new_n295), .ZN(new_n299));
  OR2_X1    g0099(.A1(new_n294), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n277), .A2(new_n281), .A3(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT70), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n251), .B1(new_n267), .B2(new_n272), .ZN(new_n304));
  OAI211_X1 g0104(.A(new_n303), .B(G200), .C1(new_n304), .C2(new_n259), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n303), .B1(new_n279), .B2(G200), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT10), .ZN(new_n309));
  OAI211_X1 g0109(.A(G190), .B(new_n258), .C1(new_n278), .C2(new_n251), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT9), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n300), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT69), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n294), .A2(new_n299), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n313), .B1(new_n314), .B2(KEYINPUT9), .ZN(new_n315));
  NOR4_X1   g0115(.A1(new_n294), .A2(new_n299), .A3(KEYINPUT69), .A4(new_n311), .ZN(new_n316));
  OAI211_X1 g0116(.A(new_n310), .B(new_n312), .C1(new_n315), .C2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n308), .A2(new_n309), .A3(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(G200), .ZN(new_n320));
  OAI21_X1  g0120(.A(KEYINPUT70), .B1(new_n275), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(new_n305), .ZN(new_n322));
  OAI21_X1  g0122(.A(KEYINPUT10), .B1(new_n322), .B2(new_n317), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n302), .B1(new_n319), .B2(new_n323), .ZN(new_n324));
  AOI22_X1  g0124(.A1(new_n291), .A2(G50), .B1(G20), .B2(new_n224), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n325), .B1(new_n270), .B2(new_n289), .ZN(new_n326));
  AND2_X1   g0126(.A1(new_n326), .A2(new_n283), .ZN(new_n327));
  OR2_X1    g0127(.A1(new_n327), .A2(KEYINPUT11), .ZN(new_n328));
  INV_X1    g0128(.A(new_n295), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(new_n224), .ZN(new_n330));
  XNOR2_X1  g0130(.A(new_n330), .B(KEYINPUT12), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n327), .A2(KEYINPUT11), .ZN(new_n332));
  INV_X1    g0132(.A(new_n296), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n333), .A2(G68), .A3(new_n297), .ZN(new_n334));
  NAND4_X1  g0134(.A1(new_n328), .A2(new_n331), .A3(new_n332), .A4(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n256), .A2(KEYINPUT71), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT71), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n251), .A2(new_n337), .A3(new_n255), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n336), .A2(G238), .A3(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  NOR2_X1   g0140(.A1(G226), .A2(G1698), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n341), .B1(new_n230), .B2(G1698), .ZN(new_n342));
  AOI22_X1  g0142(.A1(new_n342), .A2(new_n260), .B1(G33), .B2(G97), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n252), .B1(new_n343), .B2(new_n251), .ZN(new_n344));
  OAI21_X1  g0144(.A(KEYINPUT13), .B1(new_n340), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n342), .A2(new_n260), .ZN(new_n346));
  NAND2_X1  g0146(.A1(G33), .A2(G97), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n253), .B1(new_n348), .B2(new_n274), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT13), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n349), .A2(new_n350), .A3(new_n339), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n345), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n335), .B1(new_n352), .B2(G200), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT72), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n345), .A2(new_n354), .ZN(new_n355));
  OAI211_X1 g0155(.A(KEYINPUT72), .B(KEYINPUT13), .C1(new_n340), .C2(new_n344), .ZN(new_n356));
  NAND4_X1  g0156(.A1(new_n355), .A2(G190), .A3(new_n356), .A4(new_n351), .ZN(new_n357));
  AND2_X1   g0157(.A1(new_n353), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n352), .A2(G169), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(KEYINPUT14), .ZN(new_n360));
  NAND4_X1  g0160(.A1(new_n355), .A2(G179), .A3(new_n356), .A4(new_n351), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT14), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n352), .A2(new_n362), .A3(G169), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n360), .A2(new_n361), .A3(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n358), .B1(new_n335), .B2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT73), .ZN(new_n366));
  NAND2_X1  g0166(.A1(G58), .A2(G68), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n222), .B1(new_n225), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n291), .A2(G159), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n366), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  AND2_X1   g0171(.A1(G58), .A2(G68), .ZN(new_n372));
  NOR2_X1   g0172(.A1(G58), .A2(G68), .ZN(new_n373));
  OAI21_X1  g0173(.A(G20), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n374), .A2(KEYINPUT73), .A3(new_n369), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n371), .A2(new_n375), .ZN(new_n376));
  AND2_X1   g0176(.A1(KEYINPUT3), .A2(G33), .ZN(new_n377));
  NOR2_X1   g0177(.A1(KEYINPUT3), .A2(G33), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(KEYINPUT7), .B1(new_n379), .B2(new_n222), .ZN(new_n380));
  OR2_X1    g0180(.A1(KEYINPUT3), .A2(G33), .ZN(new_n381));
  NAND2_X1  g0181(.A1(KEYINPUT3), .A2(G33), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n381), .A2(KEYINPUT7), .A3(new_n222), .A4(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(new_n383), .ZN(new_n384));
  OAI21_X1  g0184(.A(G68), .B1(new_n380), .B2(new_n384), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n376), .A2(new_n385), .A3(KEYINPUT16), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT16), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n381), .A2(new_n222), .A3(new_n382), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT7), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n224), .B1(new_n390), .B2(new_n383), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n374), .A2(new_n369), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n387), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n386), .A2(new_n393), .A3(new_n283), .ZN(new_n394));
  AND2_X1   g0194(.A1(new_n288), .A2(new_n297), .ZN(new_n395));
  INV_X1    g0195(.A(new_n288), .ZN(new_n396));
  AOI22_X1  g0196(.A1(new_n333), .A2(new_n395), .B1(new_n396), .B2(new_n329), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n394), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n209), .A2(G1698), .ZN(new_n399));
  OAI221_X1 g0199(.A(new_n399), .B1(G223), .B2(G1698), .C1(new_n377), .C2(new_n378), .ZN(new_n400));
  NAND2_X1  g0200(.A1(G33), .A2(G87), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(new_n274), .ZN(new_n403));
  INV_X1    g0203(.A(G274), .ZN(new_n404));
  INV_X1    g0204(.A(new_n221), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n404), .B1(new_n405), .B2(new_n250), .ZN(new_n406));
  AOI22_X1  g0206(.A1(new_n257), .A2(G232), .B1(new_n406), .B2(new_n249), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n403), .A2(new_n276), .A3(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n251), .B1(new_n400), .B2(new_n401), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n252), .B1(new_n230), .B2(new_n256), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n280), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n408), .A2(KEYINPUT74), .A3(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT74), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n403), .A2(new_n407), .A3(new_n413), .A4(new_n276), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n398), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(KEYINPUT18), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT18), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n398), .A2(new_n415), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(G190), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n403), .A2(new_n421), .A3(new_n407), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n320), .B1(new_n409), .B2(new_n410), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n394), .A2(new_n397), .A3(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT75), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n426), .A2(KEYINPUT17), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  XNOR2_X1  g0228(.A(KEYINPUT75), .B(KEYINPUT17), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n394), .A2(new_n424), .A3(new_n397), .A4(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n420), .A2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(G33), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n222), .A2(new_n433), .ZN(new_n434));
  OAI22_X1  g0234(.A1(new_n396), .A2(new_n434), .B1(new_n222), .B2(new_n270), .ZN(new_n435));
  XNOR2_X1  g0235(.A(KEYINPUT15), .B(G87), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n436), .A2(new_n289), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n283), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n329), .A2(new_n270), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n297), .A2(G77), .ZN(new_n440));
  OAI211_X1 g0240(.A(new_n438), .B(new_n439), .C1(new_n296), .C2(new_n440), .ZN(new_n441));
  OAI211_X1 g0241(.A(G238), .B(G1698), .C1(new_n377), .C2(new_n378), .ZN(new_n442));
  OAI211_X1 g0242(.A(G232), .B(new_n261), .C1(new_n377), .C2(new_n378), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n381), .A2(G107), .A3(new_n382), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n442), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(new_n274), .ZN(new_n446));
  AOI22_X1  g0246(.A1(new_n257), .A2(G244), .B1(new_n406), .B2(new_n249), .ZN(new_n447));
  AND3_X1   g0247(.A1(new_n446), .A2(new_n447), .A3(KEYINPUT68), .ZN(new_n448));
  AOI21_X1  g0248(.A(KEYINPUT68), .B1(new_n446), .B2(new_n447), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n441), .B1(new_n450), .B2(G200), .ZN(new_n451));
  OAI21_X1  g0251(.A(G190), .B1(new_n448), .B2(new_n449), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n450), .A2(new_n280), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n276), .B1(new_n448), .B2(new_n449), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n454), .A2(new_n441), .A3(new_n455), .ZN(new_n456));
  AND2_X1   g0256(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  AND4_X1   g0257(.A1(new_n324), .A2(new_n365), .A3(new_n432), .A4(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n248), .A2(G1), .ZN(new_n460));
  AND2_X1   g0260(.A1(KEYINPUT5), .A2(G41), .ZN(new_n461));
  NOR2_X1   g0261(.A1(KEYINPUT5), .A2(G41), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n460), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n463), .A2(G270), .A3(new_n251), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(KEYINPUT79), .ZN(new_n465));
  INV_X1    g0265(.A(G303), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n251), .B1(new_n379), .B2(new_n466), .ZN(new_n467));
  NOR2_X1   g0267(.A1(G257), .A2(G1698), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n261), .A2(G264), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n260), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n406), .B(new_n460), .C1(new_n462), .C2(new_n461), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT79), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n463), .A2(new_n473), .A3(G270), .A4(new_n251), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n465), .A2(new_n471), .A3(new_n472), .A4(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n254), .A2(G33), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n295), .A2(new_n477), .A3(new_n221), .A4(new_n282), .ZN(new_n478));
  AND2_X1   g0278(.A1(new_n478), .A2(G116), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n329), .A2(G116), .ZN(new_n480));
  INV_X1    g0280(.A(G116), .ZN(new_n481));
  AOI22_X1  g0281(.A1(new_n282), .A2(new_n221), .B1(G20), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(G33), .A2(G283), .ZN(new_n483));
  INV_X1    g0283(.A(G97), .ZN(new_n484));
  OAI211_X1 g0284(.A(new_n483), .B(new_n222), .C1(G33), .C2(new_n484), .ZN(new_n485));
  AND3_X1   g0285(.A1(new_n482), .A2(KEYINPUT20), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(KEYINPUT20), .B1(new_n482), .B2(new_n485), .ZN(new_n487));
  OAI22_X1  g0287(.A1(new_n479), .A2(new_n480), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n476), .A2(G179), .A3(new_n488), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n475), .A2(new_n488), .A3(KEYINPUT21), .A4(G169), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n475), .A2(new_n488), .A3(G169), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT21), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT80), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n492), .A2(KEYINPUT80), .A3(new_n493), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n491), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n488), .B1(new_n475), .B2(G200), .ZN(new_n499));
  AOI22_X1  g0299(.A1(new_n499), .A2(KEYINPUT81), .B1(G190), .B2(new_n476), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n500), .B1(KEYINPUT81), .B2(new_n499), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n498), .A2(new_n501), .ZN(new_n502));
  AND3_X1   g0302(.A1(new_n463), .A2(G264), .A3(new_n251), .ZN(new_n503));
  OAI211_X1 g0303(.A(G257), .B(G1698), .C1(new_n377), .C2(new_n378), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(KEYINPUT86), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT86), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n260), .A2(new_n506), .A3(G257), .A4(G1698), .ZN(new_n507));
  INV_X1    g0307(.A(G294), .ZN(new_n508));
  AND2_X1   g0308(.A1(new_n508), .A2(KEYINPUT87), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n508), .A2(KEYINPUT87), .ZN(new_n510));
  OAI21_X1  g0310(.A(G33), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n260), .A2(G250), .A3(new_n261), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n505), .A2(new_n507), .A3(new_n511), .A4(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n503), .B1(new_n513), .B2(new_n274), .ZN(new_n514));
  AOI21_X1  g0314(.A(G169), .B1(new_n514), .B2(new_n472), .ZN(new_n515));
  NOR3_X1   g0315(.A1(new_n463), .A2(new_n274), .A3(new_n404), .ZN(new_n516));
  AOI211_X1 g0316(.A(new_n516), .B(new_n503), .C1(new_n513), .C2(new_n274), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n515), .B1(new_n276), .B2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(G13), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n519), .A2(G1), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n222), .A2(G107), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT85), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n522), .A2(new_n523), .A3(KEYINPUT25), .ZN(new_n524));
  OR2_X1    g0324(.A1(new_n523), .A2(KEYINPUT25), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n523), .A2(KEYINPUT25), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n525), .A2(new_n520), .A3(new_n521), .A4(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(G107), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n524), .B(new_n527), .C1(new_n528), .C2(new_n478), .ZN(new_n529));
  INV_X1    g0329(.A(new_n529), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n222), .B(G87), .C1(new_n377), .C2(new_n378), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(KEYINPUT22), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT22), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n260), .A2(new_n533), .A3(new_n222), .A4(G87), .ZN(new_n534));
  AND2_X1   g0334(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT82), .ZN(new_n536));
  NAND2_X1  g0336(.A1(G33), .A2(G116), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n536), .B1(new_n537), .B2(G20), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n222), .A2(KEYINPUT82), .A3(G33), .A4(G116), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT23), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n538), .A2(new_n539), .B1(new_n540), .B2(new_n521), .ZN(new_n541));
  OAI21_X1  g0341(.A(KEYINPUT23), .B1(new_n222), .B2(G107), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(KEYINPUT83), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT83), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n544), .B(KEYINPUT23), .C1(new_n222), .C2(G107), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n541), .A2(new_n546), .ZN(new_n547));
  OAI21_X1  g0347(.A(KEYINPUT24), .B1(new_n535), .B2(new_n547), .ZN(new_n548));
  AND2_X1   g0348(.A1(new_n541), .A2(new_n546), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT24), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n532), .A2(new_n534), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n284), .B1(new_n548), .B2(new_n552), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n530), .B1(new_n553), .B2(KEYINPUT84), .ZN(new_n554));
  NOR3_X1   g0354(.A1(new_n535), .A2(KEYINPUT24), .A3(new_n547), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n550), .B1(new_n549), .B2(new_n551), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n283), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT84), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n518), .B1(new_n554), .B2(new_n559), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n295), .A2(G97), .ZN(new_n561));
  INV_X1    g0361(.A(new_n478), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n561), .B1(new_n562), .B2(G97), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  OAI21_X1  g0364(.A(G107), .B1(new_n380), .B2(new_n384), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT6), .ZN(new_n566));
  AND2_X1   g0366(.A1(G97), .A2(G107), .ZN(new_n567));
  NOR2_X1   g0367(.A1(G97), .A2(G107), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n566), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n528), .A2(KEYINPUT6), .A3(G97), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  AOI22_X1  g0371(.A1(new_n571), .A2(G20), .B1(G77), .B2(new_n291), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n565), .A2(new_n572), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n564), .B1(new_n573), .B2(new_n283), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n463), .A2(G257), .A3(new_n251), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT76), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n463), .A2(KEYINPUT76), .A3(G257), .A4(new_n251), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n516), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  OAI211_X1 g0379(.A(G244), .B(new_n261), .C1(new_n377), .C2(new_n378), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT4), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n260), .A2(KEYINPUT4), .A3(G244), .A4(new_n261), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n260), .A2(G250), .A3(G1698), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n582), .A2(new_n583), .A3(new_n483), .A4(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(new_n274), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n579), .A2(new_n586), .A3(G190), .ZN(new_n587));
  AND2_X1   g0387(.A1(new_n579), .A2(new_n586), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n574), .B(new_n587), .C1(new_n588), .C2(new_n320), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n579), .A2(new_n586), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n280), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n579), .A2(new_n586), .A3(new_n276), .ZN(new_n592));
  AND2_X1   g0392(.A1(new_n569), .A2(new_n570), .ZN(new_n593));
  OAI22_X1  g0393(.A1(new_n593), .A2(new_n222), .B1(new_n270), .B2(new_n434), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n528), .B1(new_n390), .B2(new_n383), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n283), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(new_n563), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n591), .A2(new_n592), .A3(new_n597), .ZN(new_n598));
  AND2_X1   g0398(.A1(new_n589), .A2(new_n598), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n529), .B1(new_n557), .B2(new_n558), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n553), .A2(KEYINPUT84), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n514), .A2(new_n421), .A3(new_n472), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n602), .B1(new_n517), .B2(G200), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n600), .A2(new_n601), .A3(new_n603), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n211), .B1(new_n248), .B2(G1), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n254), .A2(new_n404), .A3(G45), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n251), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(KEYINPUT77), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT77), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n251), .A2(new_n605), .A3(new_n606), .A4(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(G244), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(G1698), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n613), .B1(G238), .B2(G1698), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n537), .B1(new_n614), .B2(new_n379), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n274), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n611), .A2(new_n616), .A3(G190), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(KEYINPUT78), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n611), .A2(new_n616), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(G200), .ZN(new_n620));
  NAND3_X1  g0420(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(new_n222), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n568), .A2(new_n210), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n222), .B(G68), .C1(new_n377), .C2(new_n378), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT19), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n626), .B1(new_n289), .B2(new_n484), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n624), .A2(new_n625), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(new_n283), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n436), .A2(new_n329), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n562), .A2(G87), .ZN(new_n631));
  AND3_X1   g0431(.A1(new_n629), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT78), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n611), .A2(new_n616), .A3(new_n633), .A4(G190), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n618), .A2(new_n620), .A3(new_n632), .A4(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n619), .A2(new_n280), .ZN(new_n636));
  OAI211_X1 g0436(.A(new_n629), .B(new_n630), .C1(new_n436), .C2(new_n478), .ZN(new_n637));
  OAI211_X1 g0437(.A(new_n636), .B(new_n637), .C1(G179), .C2(new_n619), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n635), .A2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n560), .A2(new_n599), .A3(new_n604), .A4(new_n640), .ZN(new_n641));
  NOR3_X1   g0441(.A1(new_n459), .A2(new_n502), .A3(new_n641), .ZN(G372));
  AND3_X1   g0442(.A1(new_n611), .A2(new_n616), .A3(new_n276), .ZN(new_n643));
  AOI21_X1  g0443(.A(G169), .B1(new_n611), .B2(new_n616), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n320), .B1(new_n611), .B2(new_n616), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n629), .A2(new_n630), .A3(new_n631), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  AOI22_X1  g0448(.A1(new_n637), .A2(new_n645), .B1(new_n648), .B2(new_n617), .ZN(new_n649));
  AND3_X1   g0449(.A1(new_n649), .A2(new_n598), .A3(new_n589), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n517), .A2(new_n276), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n651), .B1(new_n517), .B2(G169), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n652), .B1(new_n600), .B2(new_n601), .ZN(new_n653));
  INV_X1    g0453(.A(new_n497), .ZN(new_n654));
  AOI21_X1  g0454(.A(KEYINPUT80), .B1(new_n492), .B2(new_n493), .ZN(new_n655));
  OAI211_X1 g0455(.A(new_n490), .B(new_n489), .C1(new_n654), .C2(new_n655), .ZN(new_n656));
  OAI211_X1 g0456(.A(new_n650), .B(new_n604), .C1(new_n653), .C2(new_n656), .ZN(new_n657));
  OAI21_X1  g0457(.A(KEYINPUT26), .B1(new_n639), .B2(new_n598), .ZN(new_n658));
  AND3_X1   g0458(.A1(new_n579), .A2(new_n586), .A3(new_n276), .ZN(new_n659));
  AOI21_X1  g0459(.A(G169), .B1(new_n579), .B2(new_n586), .ZN(new_n660));
  NOR3_X1   g0460(.A1(new_n659), .A2(new_n660), .A3(new_n574), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT26), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n661), .A2(new_n649), .A3(new_n662), .ZN(new_n663));
  AND3_X1   g0463(.A1(new_n658), .A2(new_n663), .A3(new_n638), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n657), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n458), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g0466(.A(new_n666), .B(KEYINPUT88), .Z(new_n667));
  AND3_X1   g0467(.A1(new_n398), .A2(new_n415), .A3(new_n418), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n418), .B1(new_n398), .B2(new_n415), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n353), .A2(new_n357), .ZN(new_n671));
  AND3_X1   g0471(.A1(new_n454), .A2(new_n441), .A3(new_n455), .ZN(new_n672));
  AOI22_X1  g0472(.A1(new_n364), .A2(new_n335), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n670), .B1(new_n673), .B2(new_n431), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n319), .A2(new_n323), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n302), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n667), .A2(new_n676), .ZN(G369));
  NAND2_X1  g0477(.A1(new_n520), .A2(new_n222), .ZN(new_n678));
  OR2_X1    g0478(.A1(new_n678), .A2(KEYINPUT27), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(KEYINPUT27), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n679), .A2(G213), .A3(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(G343), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  AND2_X1   g0483(.A1(new_n683), .A2(new_n488), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n656), .A2(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n685), .B1(new_n502), .B2(new_n684), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(G330), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  AND2_X1   g0488(.A1(new_n560), .A2(new_n604), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n683), .B1(new_n554), .B2(new_n559), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n653), .A2(new_n683), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n688), .A2(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n498), .A2(new_n683), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n689), .A2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT89), .ZN(new_n697));
  INV_X1    g0497(.A(new_n683), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n653), .A2(new_n698), .ZN(new_n699));
  AND3_X1   g0499(.A1(new_n696), .A2(new_n697), .A3(new_n699), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n697), .B1(new_n696), .B2(new_n699), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n694), .B1(new_n700), .B2(new_n701), .ZN(G399));
  INV_X1    g0502(.A(KEYINPUT90), .ZN(new_n703));
  INV_X1    g0503(.A(new_n218), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n703), .B1(new_n704), .B2(G41), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n218), .A2(KEYINPUT90), .A3(new_n247), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n623), .A2(G116), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n707), .A2(G1), .A3(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n709), .B1(new_n226), .B2(new_n707), .ZN(new_n710));
  XNOR2_X1  g0510(.A(new_n710), .B(KEYINPUT28), .ZN(new_n711));
  INV_X1    g0511(.A(G330), .ZN(new_n712));
  AND3_X1   g0512(.A1(new_n498), .A2(new_n501), .A3(new_n698), .ZN(new_n713));
  AND2_X1   g0513(.A1(new_n599), .A2(new_n640), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n689), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT30), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n276), .B1(new_n467), .B2(new_n470), .ZN(new_n717));
  AND3_X1   g0517(.A1(new_n717), .A2(new_n616), .A3(new_n611), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n465), .A2(new_n472), .A3(new_n474), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n718), .A2(new_n720), .A3(new_n514), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n716), .B1(new_n721), .B2(new_n590), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n717), .A2(new_n611), .A3(new_n616), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n723), .A2(new_n719), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n588), .A2(new_n724), .A3(KEYINPUT30), .A4(new_n514), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n514), .A2(new_n472), .ZN(new_n726));
  AOI21_X1  g0526(.A(G179), .B1(new_n611), .B2(new_n616), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n726), .A2(new_n727), .A3(new_n475), .A4(new_n590), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n722), .A2(new_n725), .A3(new_n728), .ZN(new_n729));
  AND3_X1   g0529(.A1(new_n729), .A2(KEYINPUT31), .A3(new_n683), .ZN(new_n730));
  AOI21_X1  g0530(.A(KEYINPUT31), .B1(new_n729), .B2(new_n683), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n712), .B1(new_n715), .B2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT29), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n658), .A2(new_n663), .A3(new_n638), .ZN(new_n735));
  AND3_X1   g0535(.A1(new_n599), .A2(new_n604), .A3(new_n649), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n560), .A2(new_n498), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n735), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n734), .B1(new_n738), .B2(new_n683), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n660), .A2(new_n574), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n740), .A2(new_n592), .A3(new_n635), .A4(new_n638), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n638), .B1(new_n741), .B2(KEYINPUT26), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n662), .B1(new_n661), .B2(new_n649), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n657), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n745), .A2(KEYINPUT29), .A3(new_n698), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n733), .B1(new_n739), .B2(new_n746), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n711), .B1(new_n747), .B2(G1), .ZN(G364));
  INV_X1    g0548(.A(new_n707), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n519), .A2(G20), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n254), .B1(new_n750), .B2(G45), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  OR3_X1    g0552(.A1(new_n749), .A2(KEYINPUT91), .A3(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(KEYINPUT91), .B1(new_n749), .B2(new_n752), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n688), .A2(new_n756), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n757), .B1(G330), .B2(new_n686), .ZN(new_n758));
  INV_X1    g0558(.A(KEYINPUT92), .ZN(new_n759));
  OAI21_X1  g0559(.A(G20), .B1(new_n759), .B2(G169), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n280), .A2(KEYINPUT92), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n405), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(KEYINPUT93), .ZN(new_n763));
  OR2_X1    g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n762), .A2(new_n763), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n222), .A2(G179), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n768), .A2(G190), .A3(G200), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(G87), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n768), .A2(new_n421), .A3(G200), .ZN(new_n772));
  OAI211_X1 g0572(.A(new_n771), .B(new_n260), .C1(new_n528), .C2(new_n772), .ZN(new_n773));
  XOR2_X1   g0573(.A(new_n773), .B(KEYINPUT96), .Z(new_n774));
  NOR2_X1   g0574(.A1(new_n222), .A2(new_n276), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n775), .A2(new_n421), .A3(G200), .ZN(new_n776));
  NOR2_X1   g0576(.A1(G190), .A2(G200), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  OAI22_X1  g0578(.A1(new_n776), .A2(new_n224), .B1(new_n778), .B2(new_n270), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n775), .A2(G190), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(G200), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NOR3_X1   g0582(.A1(new_n421), .A2(G179), .A3(G200), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(new_n222), .ZN(new_n784));
  OAI22_X1  g0584(.A1(new_n782), .A2(new_n202), .B1(new_n484), .B2(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n780), .A2(new_n320), .ZN(new_n786));
  AOI211_X1 g0586(.A(new_n779), .B(new_n785), .C1(G50), .C2(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n768), .A2(new_n777), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  XNOR2_X1  g0589(.A(KEYINPUT94), .B(G159), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  XOR2_X1   g0591(.A(new_n791), .B(KEYINPUT95), .Z(new_n792));
  OR2_X1    g0592(.A1(new_n792), .A2(KEYINPUT32), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n792), .A2(KEYINPUT32), .ZN(new_n794));
  NAND4_X1  g0594(.A1(new_n774), .A2(new_n787), .A3(new_n793), .A4(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(G322), .ZN(new_n796));
  INV_X1    g0596(.A(G283), .ZN(new_n797));
  OAI22_X1  g0597(.A1(new_n782), .A2(new_n796), .B1(new_n797), .B2(new_n772), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n509), .A2(new_n510), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n784), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n798), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  XOR2_X1   g0602(.A(KEYINPUT33), .B(G317), .Z(new_n803));
  INV_X1    g0603(.A(G311), .ZN(new_n804));
  OAI22_X1  g0604(.A1(new_n776), .A2(new_n803), .B1(new_n778), .B2(new_n804), .ZN(new_n805));
  AOI211_X1 g0605(.A(new_n260), .B(new_n805), .C1(G329), .C2(new_n789), .ZN(new_n806));
  AOI22_X1  g0606(.A1(new_n786), .A2(G326), .B1(new_n770), .B2(G303), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n802), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n767), .B1(new_n795), .B2(new_n808), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n218), .A2(G355), .A3(new_n260), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n810), .B1(G116), .B2(new_n218), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n245), .A2(G45), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n218), .A2(new_n379), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n813), .B1(new_n248), .B2(new_n227), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n811), .B1(new_n812), .B2(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(G13), .A2(G33), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n817), .A2(G20), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n766), .A2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n815), .A2(new_n820), .ZN(new_n821));
  NOR3_X1   g0621(.A1(new_n809), .A2(new_n821), .A3(new_n755), .ZN(new_n822));
  XNOR2_X1  g0622(.A(new_n818), .B(KEYINPUT97), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n822), .B1(new_n686), .B2(new_n823), .ZN(new_n824));
  AND2_X1   g0624(.A1(new_n758), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(G396));
  AOI21_X1  g0626(.A(new_n683), .B1(new_n657), .B2(new_n664), .ZN(new_n827));
  NAND4_X1  g0627(.A1(new_n454), .A2(new_n441), .A3(new_n455), .A4(new_n698), .ZN(new_n828));
  AOI22_X1  g0628(.A1(new_n451), .A2(new_n452), .B1(new_n441), .B2(new_n683), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n828), .B1(new_n829), .B2(new_n672), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  XNOR2_X1  g0631(.A(new_n827), .B(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n733), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n756), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n834), .B1(new_n833), .B2(new_n832), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n766), .A2(new_n816), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n755), .B1(new_n270), .B2(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n260), .B1(new_n789), .B2(G311), .ZN(new_n838));
  OAI221_X1 g0638(.A(new_n838), .B1(new_n481), .B2(new_n778), .C1(new_n797), .C2(new_n776), .ZN(new_n839));
  INV_X1    g0639(.A(new_n786), .ZN(new_n840));
  OAI22_X1  g0640(.A1(new_n782), .A2(new_n508), .B1(new_n840), .B2(new_n466), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n772), .A2(new_n210), .ZN(new_n842));
  OAI22_X1  g0642(.A1(new_n784), .A2(new_n484), .B1(new_n769), .B2(new_n528), .ZN(new_n843));
  NOR4_X1   g0643(.A1(new_n839), .A2(new_n841), .A3(new_n842), .A4(new_n843), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n772), .A2(new_n224), .ZN(new_n845));
  INV_X1    g0645(.A(G132), .ZN(new_n846));
  OAI221_X1 g0646(.A(new_n260), .B1(new_n788), .B2(new_n846), .C1(new_n201), .C2(new_n769), .ZN(new_n847));
  AOI211_X1 g0647(.A(new_n845), .B(new_n847), .C1(G58), .C2(new_n801), .ZN(new_n848));
  XOR2_X1   g0648(.A(new_n848), .B(KEYINPUT98), .Z(new_n849));
  INV_X1    g0649(.A(new_n776), .ZN(new_n850));
  INV_X1    g0650(.A(new_n778), .ZN(new_n851));
  AOI22_X1  g0651(.A1(new_n850), .A2(G150), .B1(new_n851), .B2(new_n790), .ZN(new_n852));
  INV_X1    g0652(.A(G143), .ZN(new_n853));
  INV_X1    g0653(.A(G137), .ZN(new_n854));
  OAI221_X1 g0654(.A(new_n852), .B1(new_n782), .B2(new_n853), .C1(new_n854), .C2(new_n840), .ZN(new_n855));
  XNOR2_X1  g0655(.A(new_n855), .B(KEYINPUT34), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n844), .B1(new_n849), .B2(new_n856), .ZN(new_n857));
  OAI221_X1 g0657(.A(new_n837), .B1(new_n857), .B2(new_n767), .C1(new_n831), .C2(new_n817), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n835), .A2(new_n858), .ZN(G384));
  INV_X1    g0659(.A(KEYINPUT40), .ZN(new_n860));
  INV_X1    g0660(.A(new_n397), .ZN(new_n861));
  AND3_X1   g0661(.A1(new_n374), .A2(KEYINPUT73), .A3(new_n369), .ZN(new_n862));
  AOI21_X1  g0662(.A(KEYINPUT73), .B1(new_n374), .B2(new_n369), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  OAI21_X1  g0664(.A(KEYINPUT102), .B1(new_n864), .B2(new_n391), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT102), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n376), .A2(new_n385), .A3(new_n866), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n865), .A2(new_n387), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n390), .A2(new_n383), .ZN(new_n869));
  AOI22_X1  g0669(.A1(new_n869), .A2(G68), .B1(new_n371), .B2(new_n375), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n284), .B1(new_n870), .B2(KEYINPUT16), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n861), .B1(new_n868), .B2(new_n871), .ZN(new_n872));
  AND2_X1   g0672(.A1(new_n412), .A2(new_n414), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n425), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n872), .A2(new_n681), .ZN(new_n875));
  OAI21_X1  g0675(.A(KEYINPUT37), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n416), .A2(KEYINPUT103), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT37), .ZN(new_n878));
  AND2_X1   g0678(.A1(new_n425), .A2(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n681), .B1(new_n394), .B2(new_n397), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT103), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n398), .A2(new_n415), .A3(new_n882), .ZN(new_n883));
  NAND4_X1  g0683(.A1(new_n877), .A2(new_n879), .A3(new_n881), .A4(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n876), .A2(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n875), .B1(new_n420), .B2(new_n431), .ZN(new_n886));
  AND3_X1   g0686(.A1(new_n885), .A2(KEYINPUT38), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(KEYINPUT38), .B1(new_n885), .B2(new_n886), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n364), .A2(new_n335), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n335), .A2(new_n683), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n890), .A2(new_n671), .A3(new_n891), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n335), .B(new_n683), .C1(new_n358), .C2(new_n364), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n830), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n729), .A2(new_n683), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT31), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n729), .A2(KEYINPUT31), .A3(new_n683), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n498), .A2(new_n501), .A3(new_n698), .ZN(new_n899));
  OAI211_X1 g0699(.A(new_n897), .B(new_n898), .C1(new_n641), .C2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n894), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n860), .B1(new_n889), .B2(new_n901), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n885), .A2(KEYINPUT38), .A3(new_n886), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT104), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n431), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n428), .A2(KEYINPUT104), .A3(new_n430), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n905), .A2(new_n670), .A3(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n881), .A2(new_n416), .A3(new_n425), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(KEYINPUT37), .ZN(new_n909));
  AOI22_X1  g0709(.A1(new_n907), .A2(new_n880), .B1(new_n884), .B2(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n903), .B1(new_n910), .B2(KEYINPUT38), .ZN(new_n911));
  NAND4_X1  g0711(.A1(new_n911), .A2(KEYINPUT40), .A3(new_n900), .A4(new_n894), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n902), .A2(new_n912), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n913), .B(KEYINPUT105), .ZN(new_n914));
  AND2_X1   g0714(.A1(new_n458), .A2(new_n900), .ZN(new_n915));
  AND2_X1   g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n914), .A2(new_n915), .ZN(new_n917));
  NOR3_X1   g0717(.A1(new_n916), .A2(new_n917), .A3(new_n712), .ZN(new_n918));
  AND2_X1   g0718(.A1(new_n892), .A2(new_n893), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n665), .A2(new_n698), .A3(new_n831), .ZN(new_n920));
  XOR2_X1   g0720(.A(new_n828), .B(KEYINPUT101), .Z(new_n921));
  AOI21_X1  g0721(.A(new_n919), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(new_n888), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n903), .ZN(new_n924));
  AOI22_X1  g0724(.A1(new_n922), .A2(new_n924), .B1(new_n420), .B2(new_n681), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT39), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n906), .A2(new_n417), .A3(new_n419), .ZN(new_n927));
  AOI21_X1  g0727(.A(KEYINPUT104), .B1(new_n428), .B2(new_n430), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n880), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n884), .A2(new_n909), .ZN(new_n930));
  AOI21_X1  g0730(.A(KEYINPUT38), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n926), .B1(new_n931), .B2(new_n887), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n923), .A2(KEYINPUT39), .A3(new_n903), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n890), .A2(new_n683), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  AND2_X1   g0735(.A1(new_n925), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n739), .A2(new_n458), .A3(new_n746), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(new_n676), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n936), .B(new_n938), .ZN(new_n939));
  OR2_X1    g0739(.A1(new_n918), .A2(new_n939), .ZN(new_n940));
  OR2_X1    g0740(.A1(new_n940), .A2(KEYINPUT106), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(KEYINPUT106), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n750), .A2(new_n254), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n943), .B1(new_n918), .B2(new_n939), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n941), .A2(new_n942), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n571), .A2(KEYINPUT35), .ZN(new_n946));
  OAI211_X1 g0746(.A(G116), .B(new_n223), .C1(new_n571), .C2(KEYINPUT35), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT99), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n946), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n949), .B1(new_n948), .B2(new_n947), .ZN(new_n950));
  XOR2_X1   g0750(.A(new_n950), .B(KEYINPUT36), .Z(new_n951));
  NAND2_X1  g0751(.A1(new_n367), .A2(G77), .ZN(new_n952));
  OAI22_X1  g0752(.A1(new_n226), .A2(new_n952), .B1(G50), .B2(new_n224), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n953), .A2(G1), .A3(new_n519), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n951), .A2(new_n954), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n955), .B(KEYINPUT100), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n945), .A2(new_n956), .ZN(G367));
  OAI22_X1  g0757(.A1(new_n813), .A2(new_n236), .B1(new_n218), .B2(new_n436), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n756), .B1(new_n820), .B2(new_n958), .ZN(new_n959));
  OAI22_X1  g0759(.A1(new_n840), .A2(new_n853), .B1(new_n769), .B2(new_n202), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n960), .B1(G150), .B2(new_n781), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n379), .B1(new_n850), .B2(new_n790), .ZN(new_n962));
  AOI22_X1  g0762(.A1(G50), .A2(new_n851), .B1(new_n789), .B2(G137), .ZN(new_n963));
  INV_X1    g0763(.A(new_n772), .ZN(new_n964));
  AOI22_X1  g0764(.A1(new_n801), .A2(G68), .B1(new_n964), .B2(G77), .ZN(new_n965));
  NAND4_X1  g0765(.A1(new_n961), .A2(new_n962), .A3(new_n963), .A4(new_n965), .ZN(new_n966));
  AOI22_X1  g0766(.A1(new_n781), .A2(G303), .B1(new_n964), .B2(G97), .ZN(new_n967));
  OAI221_X1 g0767(.A(new_n967), .B1(new_n528), .B2(new_n784), .C1(new_n804), .C2(new_n840), .ZN(new_n968));
  AOI22_X1  g0768(.A1(new_n800), .A2(new_n850), .B1(new_n789), .B2(G317), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n770), .A2(KEYINPUT46), .A3(G116), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT46), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n971), .B1(new_n769), .B2(new_n481), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n260), .B1(new_n851), .B2(G283), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n969), .A2(new_n970), .A3(new_n972), .A4(new_n973), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n966), .B1(new_n968), .B2(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT47), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n977), .A2(new_n767), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n975), .A2(new_n976), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n959), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n649), .B1(new_n632), .B2(new_n698), .ZN(new_n981));
  NAND4_X1  g0781(.A1(new_n645), .A2(new_n637), .A3(new_n647), .A4(new_n683), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  OR2_X1    g0783(.A1(new_n983), .A2(new_n823), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n980), .A2(new_n984), .ZN(new_n985));
  OAI211_X1 g0785(.A(new_n589), .B(new_n598), .C1(new_n574), .C2(new_n698), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n661), .A2(new_n683), .ZN(new_n987));
  AND2_X1   g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(new_n988), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n989), .B1(new_n700), .B2(new_n701), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT45), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  OAI211_X1 g0792(.A(KEYINPUT45), .B(new_n989), .C1(new_n700), .C2(new_n701), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n696), .A2(new_n699), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n995), .A2(KEYINPUT89), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n696), .A2(new_n697), .A3(new_n699), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n996), .A2(new_n997), .A3(new_n988), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT44), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND4_X1  g0800(.A1(new_n996), .A2(KEYINPUT44), .A3(new_n997), .A4(new_n988), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n994), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n694), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  OAI211_X1 g0805(.A(new_n691), .B(new_n692), .C1(new_n498), .C2(new_n683), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1006), .A2(new_n696), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1007), .A2(new_n688), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1006), .A2(new_n687), .A3(new_n696), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1010), .A2(new_n747), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n1011), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n994), .A2(new_n1002), .A3(new_n694), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1005), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1014), .A2(new_n747), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n707), .B(KEYINPUT41), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n752), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n989), .A2(new_n689), .A3(new_n695), .ZN(new_n1019));
  OR2_X1    g0819(.A1(new_n1019), .A2(KEYINPUT42), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n598), .B1(new_n560), .B2(new_n986), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n1019), .A2(KEYINPUT42), .B1(new_n698), .B2(new_n1021), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(new_n1020), .A2(new_n1022), .B1(KEYINPUT43), .B2(new_n983), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n983), .A2(KEYINPUT43), .ZN(new_n1024));
  XOR2_X1   g0824(.A(new_n1023), .B(new_n1024), .Z(new_n1025));
  NOR2_X1   g0825(.A1(new_n694), .A2(new_n988), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1025), .B(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n1027), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n985), .B1(new_n1018), .B2(new_n1028), .ZN(G387));
  OAI21_X1  g0829(.A(KEYINPUT108), .B1(new_n1010), .B2(new_n747), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n747), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT108), .ZN(new_n1032));
  NAND4_X1  g0832(.A1(new_n1031), .A2(new_n1032), .A3(new_n1008), .A4(new_n1009), .ZN(new_n1033));
  NAND4_X1  g0833(.A1(new_n1030), .A2(new_n1033), .A3(new_n749), .A4(new_n1011), .ZN(new_n1034));
  OR2_X1    g0834(.A1(new_n693), .A2(new_n823), .ZN(new_n1035));
  OR3_X1    g0835(.A1(new_n233), .A2(new_n248), .A3(new_n260), .ZN(new_n1036));
  XOR2_X1   g0836(.A(KEYINPUT107), .B(KEYINPUT50), .Z(new_n1037));
  OAI21_X1  g0837(.A(new_n1037), .B1(new_n396), .B2(G50), .ZN(new_n1038));
  OAI211_X1 g0838(.A(new_n1038), .B(new_n248), .C1(new_n224), .C2(new_n270), .ZN(new_n1039));
  NOR3_X1   g0839(.A1(new_n396), .A2(new_n1037), .A3(G50), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n379), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1041), .A2(new_n708), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n704), .B1(new_n1036), .B2(new_n1042), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n819), .B1(new_n528), .B2(new_n218), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n756), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g0845(.A(G150), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n778), .A2(new_n224), .B1(new_n788), .B2(new_n1046), .ZN(new_n1047));
  AOI211_X1 g0847(.A(new_n379), .B(new_n1047), .C1(new_n288), .C2(new_n850), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n769), .A2(new_n270), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n784), .A2(new_n436), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n1049), .B(new_n1050), .C1(G50), .C2(new_n781), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n786), .A2(G159), .B1(new_n964), .B2(G97), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1048), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n260), .B1(new_n789), .B2(G326), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n784), .A2(new_n797), .B1(new_n799), .B2(new_n769), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n850), .A2(G311), .B1(new_n851), .B2(G303), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n781), .A2(G317), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n1056), .B(new_n1057), .C1(new_n796), .C2(new_n840), .ZN(new_n1058));
  INV_X1    g0858(.A(KEYINPUT48), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1055), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1060), .B1(new_n1059), .B2(new_n1058), .ZN(new_n1061));
  INV_X1    g0861(.A(KEYINPUT49), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n1054), .B1(new_n481), .B2(new_n772), .C1(new_n1061), .C2(new_n1062), .ZN(new_n1063));
  AND2_X1   g0863(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1053), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1045), .B1(new_n1065), .B2(new_n766), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n1010), .A2(new_n752), .B1(new_n1035), .B2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1034), .A2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1068), .A2(KEYINPUT109), .ZN(new_n1069));
  INV_X1    g0869(.A(KEYINPUT109), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1034), .A2(new_n1070), .A3(new_n1067), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1069), .A2(new_n1071), .ZN(G393));
  INV_X1    g0872(.A(KEYINPUT110), .ZN(new_n1073));
  AND3_X1   g0873(.A1(new_n994), .A2(new_n1002), .A3(new_n694), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n694), .B1(new_n994), .B2(new_n1002), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1073), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1005), .A2(KEYINPUT110), .A3(new_n1013), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1076), .A2(new_n1077), .A3(new_n752), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1011), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1079), .A2(new_n1014), .A3(new_n749), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(G150), .A2(new_n786), .B1(new_n781), .B2(G159), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(new_n1081), .B(KEYINPUT111), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(KEYINPUT51), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n396), .A2(new_n778), .B1(new_n788), .B2(new_n853), .ZN(new_n1084));
  AOI211_X1 g0884(.A(new_n379), .B(new_n1084), .C1(G50), .C2(new_n850), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n784), .A2(new_n270), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n842), .B(new_n1086), .C1(G68), .C2(new_n770), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1083), .A2(new_n1085), .A3(new_n1087), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n1082), .A2(KEYINPUT51), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  OR2_X1    g0890(.A1(new_n1090), .A2(KEYINPUT112), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1090), .A2(KEYINPUT112), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(G311), .A2(new_n781), .B1(new_n786), .B2(G317), .ZN(new_n1093));
  XOR2_X1   g0893(.A(new_n1093), .B(KEYINPUT52), .Z(new_n1094));
  OAI22_X1  g0894(.A1(new_n778), .A2(new_n508), .B1(new_n788), .B2(new_n796), .ZN(new_n1095));
  AOI211_X1 g0895(.A(new_n260), .B(new_n1095), .C1(G303), .C2(new_n850), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n784), .A2(new_n481), .B1(new_n772), .B2(new_n528), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1097), .B1(G283), .B2(new_n770), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1094), .A2(new_n1096), .A3(new_n1098), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1091), .A2(new_n1092), .A3(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1100), .A2(new_n766), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n988), .A2(new_n818), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n241), .ZN(new_n1103));
  OAI221_X1 g0903(.A(new_n819), .B1(new_n484), .B2(new_n218), .C1(new_n1103), .C2(new_n813), .ZN(new_n1104));
  NAND4_X1  g0904(.A1(new_n1101), .A2(new_n756), .A3(new_n1102), .A4(new_n1104), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1078), .A2(new_n1080), .A3(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(KEYINPUT113), .ZN(new_n1107));
  XNOR2_X1  g0907(.A(new_n1106), .B(new_n1107), .ZN(G390));
  AND3_X1   g0908(.A1(new_n894), .A2(new_n900), .A3(G330), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n892), .A2(new_n893), .ZN(new_n1110));
  AOI211_X1 g0910(.A(new_n683), .B(new_n830), .C1(new_n657), .C2(new_n664), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n921), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1110), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n934), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n932), .A2(new_n933), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n911), .A2(new_n1114), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n683), .B1(new_n657), .B2(new_n744), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n829), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1118), .A2(new_n456), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1117), .A2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n919), .B1(new_n1120), .B2(new_n828), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n1116), .A2(new_n1121), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1109), .B1(new_n1115), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n733), .A2(new_n894), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n1117), .A2(new_n1119), .B1(new_n672), .B2(new_n698), .ZN(new_n1125));
  OAI211_X1 g0925(.A(new_n1114), .B(new_n911), .C1(new_n1125), .C2(new_n919), .ZN(new_n1126));
  AND2_X1   g0926(.A1(new_n932), .A2(new_n933), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n922), .A2(new_n934), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n1124), .B(new_n1126), .C1(new_n1127), .C2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1123), .A2(new_n1129), .A3(new_n752), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n379), .B1(new_n789), .B2(G125), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1131), .B1(new_n201), .B2(new_n772), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(new_n1132), .B(KEYINPUT114), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n770), .A2(G150), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(new_n1134), .B(KEYINPUT53), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(KEYINPUT54), .B(G143), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(new_n850), .A2(G137), .B1(new_n851), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(G128), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1138), .B1(new_n1139), .B2(new_n840), .ZN(new_n1140));
  INV_X1    g0940(.A(G159), .ZN(new_n1141));
  OAI22_X1  g0941(.A1(new_n782), .A2(new_n846), .B1(new_n1141), .B2(new_n784), .ZN(new_n1142));
  OR4_X1    g0942(.A1(new_n1133), .A2(new_n1135), .A3(new_n1140), .A4(new_n1142), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n840), .A2(new_n797), .ZN(new_n1144));
  AOI211_X1 g0944(.A(new_n1086), .B(new_n1144), .C1(G116), .C2(new_n781), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n845), .ZN(new_n1146));
  OAI22_X1  g0946(.A1(new_n778), .A2(new_n484), .B1(new_n788), .B2(new_n508), .ZN(new_n1147));
  AOI211_X1 g0947(.A(new_n260), .B(new_n1147), .C1(G107), .C2(new_n850), .ZN(new_n1148));
  NAND4_X1  g0948(.A1(new_n1145), .A2(new_n771), .A3(new_n1146), .A4(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n767), .B1(new_n1143), .B2(new_n1149), .ZN(new_n1150));
  AOI211_X1 g0950(.A(new_n755), .B(new_n1150), .C1(new_n396), .C2(new_n836), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1151), .B1(new_n1127), .B2(new_n817), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1130), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1123), .A2(new_n1129), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n733), .A2(new_n458), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n937), .A2(new_n676), .A3(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1112), .B1(new_n827), .B2(new_n831), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1110), .B1(new_n733), .B2(new_n831), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1158), .B1(new_n1159), .B2(new_n1109), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n900), .A2(G330), .A3(new_n831), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1161), .A2(new_n919), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1162), .A2(new_n1124), .A3(new_n1125), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1156), .B1(new_n1160), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n707), .B1(new_n1154), .B2(new_n1165), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1123), .A2(new_n1129), .A3(new_n1164), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1153), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(G378));
  NAND2_X1  g0969(.A1(new_n925), .A2(new_n935), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n309), .B1(new_n308), .B2(new_n318), .ZN(new_n1171));
  NOR3_X1   g0971(.A1(new_n322), .A2(KEYINPUT10), .A3(new_n317), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n301), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n314), .A2(new_n681), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(new_n1174), .B(KEYINPUT55), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1173), .A2(new_n1175), .ZN(new_n1176));
  XOR2_X1   g0976(.A(KEYINPUT115), .B(KEYINPUT56), .Z(new_n1177));
  INV_X1    g0977(.A(new_n1175), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n324), .A2(new_n1178), .ZN(new_n1179));
  AND3_X1   g0979(.A1(new_n1176), .A2(new_n1177), .A3(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1177), .B1(new_n1176), .B2(new_n1179), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  AND4_X1   g0982(.A1(G330), .A2(new_n902), .A3(new_n1182), .A4(new_n912), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n900), .B(new_n894), .C1(new_n887), .C2(new_n888), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n712), .B1(new_n1184), .B2(new_n860), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1182), .B1(new_n1185), .B2(new_n912), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1170), .B1(new_n1183), .B2(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(KEYINPUT116), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n902), .A2(G330), .A3(new_n912), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1182), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1185), .A2(new_n912), .A3(new_n1182), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1191), .A2(new_n936), .A3(new_n1192), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1187), .A2(new_n1188), .A3(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1156), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1167), .A2(new_n1195), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n1170), .B(KEYINPUT116), .C1(new_n1183), .C2(new_n1186), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1194), .A2(new_n1196), .A3(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(KEYINPUT57), .ZN(new_n1199));
  AND2_X1   g0999(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1187), .A2(KEYINPUT117), .A3(new_n1193), .ZN(new_n1201));
  INV_X1    g1001(.A(KEYINPUT117), .ZN(new_n1202));
  OAI211_X1 g1002(.A(new_n1170), .B(new_n1202), .C1(new_n1183), .C2(new_n1186), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1201), .A2(new_n1196), .A3(KEYINPUT57), .A4(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1204), .A2(new_n749), .ZN(new_n1205));
  OR2_X1    g1005(.A1(new_n1200), .A2(new_n1205), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1194), .A2(new_n752), .A3(new_n1197), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n836), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n756), .B1(G50), .B2(new_n1208), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n776), .A2(new_n846), .B1(new_n778), .B2(new_n854), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(G150), .A2(new_n801), .B1(new_n786), .B2(G125), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1211), .B1(new_n1139), .B2(new_n782), .ZN(new_n1212));
  AOI211_X1 g1012(.A(new_n1210), .B(new_n1212), .C1(new_n770), .C2(new_n1137), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT59), .ZN(new_n1214));
  OR2_X1    g1014(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n964), .A2(new_n790), .ZN(new_n1217));
  AOI211_X1 g1017(.A(G33), .B(G41), .C1(new_n789), .C2(G124), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1215), .A2(new_n1216), .A3(new_n1217), .A4(new_n1218), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n201), .B1(G33), .B2(G41), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1220), .B1(new_n379), .B2(new_n247), .ZN(new_n1221));
  OAI22_X1  g1021(.A1(new_n782), .A2(new_n528), .B1(new_n202), .B2(new_n772), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1222), .B1(G116), .B2(new_n786), .ZN(new_n1223));
  AOI211_X1 g1023(.A(G41), .B(new_n260), .C1(new_n850), .C2(G97), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n436), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(new_n1225), .A2(new_n851), .B1(new_n789), .B2(G283), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1049), .B1(G68), .B2(new_n801), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1223), .A2(new_n1224), .A3(new_n1226), .A4(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT58), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1221), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1230));
  OAI211_X1 g1030(.A(new_n1219), .B(new_n1230), .C1(new_n1229), .C2(new_n1228), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1209), .B1(new_n1231), .B2(new_n766), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1232), .B1(new_n1182), .B2(new_n817), .ZN(new_n1233));
  AND2_X1   g1033(.A1(new_n1207), .A2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1206), .A2(new_n1234), .ZN(G375));
  NAND3_X1  g1035(.A1(new_n1160), .A2(new_n1156), .A3(new_n1163), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1165), .A2(new_n1017), .A3(new_n1236), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n919), .A2(new_n1161), .B1(new_n733), .B2(new_n894), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1163), .B1(new_n1238), .B2(new_n1157), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n919), .A2(new_n816), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n756), .B1(G68), .B2(new_n1208), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n840), .A2(new_n508), .B1(new_n769), .B2(new_n484), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1242), .B1(G283), .B2(new_n781), .ZN(new_n1243));
  OAI22_X1  g1043(.A1(new_n778), .A2(new_n528), .B1(new_n788), .B2(new_n466), .ZN(new_n1244));
  AOI211_X1 g1044(.A(new_n260), .B(new_n1244), .C1(G116), .C2(new_n850), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1050), .B1(G77), .B2(new_n964), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1243), .A2(new_n1245), .A3(new_n1246), .ZN(new_n1247));
  OR2_X1    g1047(.A1(new_n1247), .A2(KEYINPUT118), .ZN(new_n1248));
  OAI22_X1  g1048(.A1(new_n782), .A2(new_n854), .B1(new_n769), .B2(new_n1141), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1249), .B1(G132), .B2(new_n786), .ZN(new_n1250));
  OAI22_X1  g1050(.A1(new_n776), .A2(new_n1136), .B1(new_n788), .B2(new_n1139), .ZN(new_n1251));
  AOI211_X1 g1051(.A(new_n379), .B(new_n1251), .C1(G150), .C2(new_n851), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(new_n801), .A2(G50), .B1(new_n964), .B2(G58), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1250), .A2(new_n1252), .A3(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1247), .A2(KEYINPUT118), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1248), .A2(new_n1254), .A3(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1241), .B1(new_n766), .B2(new_n1256), .ZN(new_n1257));
  AOI22_X1  g1057(.A1(new_n1239), .A2(new_n752), .B1(new_n1240), .B2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1237), .A2(new_n1258), .ZN(G381));
  XNOR2_X1  g1059(.A(new_n1106), .B(KEYINPUT113), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n985), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1031), .B1(new_n1262), .B2(new_n1010), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n751), .B1(new_n1263), .B2(new_n1016), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1261), .B1(new_n1264), .B2(new_n1027), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1069), .A2(new_n825), .A3(new_n1071), .ZN(new_n1266));
  NOR3_X1   g1066(.A1(new_n1266), .A2(G384), .A3(G381), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1260), .A2(new_n1265), .A3(new_n1267), .ZN(new_n1268));
  XNOR2_X1  g1068(.A(new_n1268), .B(KEYINPUT119), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(G375), .A2(G378), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(new_n1270), .ZN(G407));
  INV_X1    g1071(.A(new_n1270), .ZN(new_n1272));
  OAI211_X1 g1072(.A(G407), .B(G213), .C1(G343), .C2(new_n1272), .ZN(G409));
  INV_X1    g1073(.A(new_n1071), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1070), .B1(new_n1034), .B2(new_n1067), .ZN(new_n1275));
  OAI21_X1  g1075(.A(G396), .B1(new_n1274), .B2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(new_n1266), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT125), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1277), .B1(new_n1265), .B2(new_n1278), .ZN(new_n1279));
  AND2_X1   g1079(.A1(new_n1276), .A2(new_n1266), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1280), .A2(G387), .ZN(new_n1281));
  AND3_X1   g1081(.A1(new_n1279), .A2(G390), .A3(new_n1281), .ZN(new_n1282));
  AOI21_X1  g1082(.A(G390), .B1(new_n1279), .B2(new_n1281), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  NAND4_X1  g1084(.A1(new_n1194), .A2(new_n1196), .A3(new_n1017), .A4(new_n1197), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1201), .A2(new_n752), .A3(new_n1203), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1285), .A2(new_n1233), .A3(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1287), .A2(new_n1168), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1288), .A2(KEYINPUT120), .ZN(new_n1289));
  OAI211_X1 g1089(.A(G378), .B(new_n1234), .C1(new_n1200), .C2(new_n1205), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT120), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1287), .A2(new_n1291), .A3(new_n1168), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1289), .A2(new_n1290), .A3(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n682), .A2(G213), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT122), .ZN(new_n1295));
  AND3_X1   g1095(.A1(new_n1162), .A2(new_n1124), .A3(new_n1125), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1157), .B1(new_n1162), .B2(new_n1124), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT121), .ZN(new_n1299));
  NAND4_X1  g1099(.A1(new_n1298), .A2(new_n1299), .A3(KEYINPUT60), .A4(new_n1156), .ZN(new_n1300));
  NAND4_X1  g1100(.A1(new_n1160), .A2(new_n1156), .A3(KEYINPUT60), .A4(new_n1163), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(KEYINPUT121), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT60), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1236), .A2(new_n1303), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n707), .B1(new_n1239), .B2(new_n1195), .ZN(new_n1305));
  NAND4_X1  g1105(.A1(new_n1300), .A2(new_n1302), .A3(new_n1304), .A4(new_n1305), .ZN(new_n1306));
  AND3_X1   g1106(.A1(new_n1306), .A2(G384), .A3(new_n1258), .ZN(new_n1307));
  AOI21_X1  g1107(.A(G384), .B1(new_n1306), .B2(new_n1258), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1295), .B1(new_n1307), .B2(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1306), .A2(new_n1258), .ZN(new_n1310));
  INV_X1    g1110(.A(G384), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1306), .A2(G384), .A3(new_n1258), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1312), .A2(KEYINPUT122), .A3(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1309), .A2(new_n1314), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1293), .A2(new_n1294), .A3(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1316), .A2(KEYINPUT62), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT62), .ZN(new_n1318));
  NAND4_X1  g1118(.A1(new_n1293), .A2(new_n1318), .A3(new_n1294), .A4(new_n1315), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n682), .A2(G213), .A3(G2897), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1321), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1322), .B1(new_n1309), .B2(new_n1314), .ZN(new_n1323));
  NOR2_X1   g1123(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1324));
  NOR2_X1   g1124(.A1(new_n1324), .A2(new_n1321), .ZN(new_n1325));
  NOR2_X1   g1125(.A1(new_n1323), .A2(new_n1325), .ZN(new_n1326));
  AOI21_X1  g1126(.A(KEYINPUT61), .B1(new_n1320), .B2(new_n1326), .ZN(new_n1327));
  OAI211_X1 g1127(.A(new_n1317), .B(new_n1319), .C1(new_n1327), .C2(KEYINPUT127), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT127), .ZN(new_n1329));
  AOI211_X1 g1129(.A(new_n1329), .B(KEYINPUT61), .C1(new_n1320), .C2(new_n1326), .ZN(new_n1330));
  OAI21_X1  g1130(.A(new_n1284), .B1(new_n1328), .B2(new_n1330), .ZN(new_n1331));
  NOR3_X1   g1131(.A1(new_n1307), .A2(new_n1308), .A3(new_n1295), .ZN(new_n1332));
  AOI21_X1  g1132(.A(KEYINPUT122), .B1(new_n1312), .B2(new_n1313), .ZN(new_n1333));
  OAI21_X1  g1133(.A(new_n1321), .B1(new_n1332), .B2(new_n1333), .ZN(new_n1334));
  INV_X1    g1134(.A(new_n1325), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1334), .A2(new_n1335), .A3(KEYINPUT123), .ZN(new_n1336));
  INV_X1    g1136(.A(KEYINPUT123), .ZN(new_n1337));
  OAI21_X1  g1137(.A(new_n1337), .B1(new_n1323), .B2(new_n1325), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1336), .A2(new_n1338), .ZN(new_n1339));
  AND3_X1   g1139(.A1(new_n1339), .A2(KEYINPUT124), .A3(new_n1320), .ZN(new_n1340));
  AOI21_X1  g1140(.A(KEYINPUT124), .B1(new_n1339), .B2(new_n1320), .ZN(new_n1341));
  NOR2_X1   g1141(.A1(new_n1340), .A2(new_n1341), .ZN(new_n1342));
  INV_X1    g1142(.A(KEYINPUT61), .ZN(new_n1343));
  OAI21_X1  g1143(.A(new_n1343), .B1(new_n1282), .B2(new_n1283), .ZN(new_n1344));
  INV_X1    g1144(.A(KEYINPUT63), .ZN(new_n1345));
  AOI21_X1  g1145(.A(new_n1344), .B1(new_n1345), .B2(new_n1316), .ZN(new_n1346));
  NAND4_X1  g1146(.A1(new_n1293), .A2(KEYINPUT63), .A3(new_n1294), .A4(new_n1315), .ZN(new_n1347));
  XNOR2_X1  g1147(.A(new_n1347), .B(KEYINPUT126), .ZN(new_n1348));
  NAND3_X1  g1148(.A1(new_n1342), .A2(new_n1346), .A3(new_n1348), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1331), .A2(new_n1349), .ZN(G405));
  NAND2_X1  g1150(.A1(G375), .A2(G378), .ZN(new_n1351));
  INV_X1    g1151(.A(new_n1351), .ZN(new_n1352));
  NOR2_X1   g1152(.A1(new_n1352), .A2(new_n1270), .ZN(new_n1353));
  NOR2_X1   g1153(.A1(new_n1353), .A2(new_n1324), .ZN(new_n1354));
  AND3_X1   g1154(.A1(new_n1272), .A2(new_n1315), .A3(new_n1351), .ZN(new_n1355));
  OAI21_X1  g1155(.A(new_n1284), .B1(new_n1354), .B2(new_n1355), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1353), .A2(new_n1315), .ZN(new_n1357));
  INV_X1    g1157(.A(new_n1284), .ZN(new_n1358));
  OAI211_X1 g1158(.A(new_n1357), .B(new_n1358), .C1(new_n1324), .C2(new_n1353), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1356), .A2(new_n1359), .ZN(G402));
endmodule


