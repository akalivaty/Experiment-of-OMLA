//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 1 0 0 1 0 0 0 0 0 1 0 0 1 0 0 1 0 0 1 1 1 0 1 1 1 0 0 0 1 1 1 0 1 1 1 0 1 1 0 1 0 1 0 1 1 1 1 0 0 1 0 0 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:26 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n450, new_n451, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n531, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n550,
    new_n551, new_n552, new_n553, new_n555, new_n557, new_n558, new_n559,
    new_n561, new_n562, new_n563, new_n564, new_n566, new_n567, new_n568,
    new_n569, new_n571, new_n572, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n580, new_n581, new_n582, new_n583, new_n584, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n601, new_n602,
    new_n605, new_n606, new_n608, new_n609, new_n610, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1118,
    new_n1119;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT64), .B(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  INV_X1    g024(.A(G2106), .ZN(new_n450));
  NOR2_X1   g025(.A1(new_n447), .A2(new_n450), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT65), .Z(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  NOR4_X1   g029(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT66), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  XNOR2_X1  g032(.A(new_n457), .B(KEYINPUT67), .ZN(G261));
  INV_X1    g033(.A(G261), .ZN(G325));
  OR2_X1    g034(.A1(new_n454), .A2(new_n450), .ZN(new_n460));
  INV_X1    g035(.A(G567), .ZN(new_n461));
  OR2_X1    g036(.A1(new_n456), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n465), .A2(G2105), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G101), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT68), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT3), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n468), .B1(new_n469), .B2(G2104), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n465), .A2(KEYINPUT68), .A3(KEYINPUT3), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n469), .A2(G2104), .ZN(new_n473));
  NAND4_X1  g048(.A1(new_n470), .A2(new_n471), .A3(new_n472), .A4(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(G137), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n467), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(KEYINPUT69), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT69), .ZN(new_n478));
  OAI211_X1 g053(.A(new_n478), .B(new_n467), .C1(new_n474), .C2(new_n475), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(G113), .A2(G2104), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(new_n473), .ZN(new_n483));
  INV_X1    g058(.A(G125), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n481), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n480), .B1(G2105), .B2(new_n485), .ZN(G160));
  NAND4_X1  g061(.A1(new_n470), .A2(new_n471), .A3(G2105), .A4(new_n473), .ZN(new_n487));
  INV_X1    g062(.A(G124), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n472), .A2(G112), .ZN(new_n489));
  OAI21_X1  g064(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n490));
  OAI22_X1  g065(.A1(new_n487), .A2(new_n488), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n474), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n491), .B1(new_n492), .B2(G136), .ZN(G162));
  INV_X1    g068(.A(G138), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n494), .A2(G2105), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n470), .A2(new_n471), .A3(new_n495), .A4(new_n473), .ZN(new_n496));
  AND2_X1   g071(.A1(new_n482), .A2(new_n473), .ZN(new_n497));
  NOR3_X1   g072(.A1(new_n494), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n498));
  AOI22_X1  g073(.A1(new_n496), .A2(KEYINPUT4), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(G126), .ZN(new_n500));
  OR2_X1    g075(.A1(KEYINPUT70), .A2(G114), .ZN(new_n501));
  NAND2_X1  g076(.A1(KEYINPUT70), .A2(G114), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n472), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  OAI21_X1  g078(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n504));
  OAI22_X1  g079(.A1(new_n487), .A2(new_n500), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n499), .A2(new_n505), .ZN(G164));
  INV_X1    g081(.A(KEYINPUT5), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n507), .B1(new_n508), .B2(KEYINPUT71), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT71), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n510), .A2(KEYINPUT5), .A3(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n512), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  OR2_X1    g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  OR2_X1    g090(.A1(KEYINPUT6), .A2(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n509), .A2(new_n511), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  XNOR2_X1  g093(.A(KEYINPUT72), .B(G88), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n508), .B1(new_n516), .B2(new_n517), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n518), .A2(new_n519), .B1(new_n520), .B2(G50), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n515), .A2(new_n521), .ZN(G303));
  INV_X1    g097(.A(G303), .ZN(G166));
  NAND2_X1  g098(.A1(new_n518), .A2(G89), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n512), .A2(G63), .A3(G651), .ZN(new_n525));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  XNOR2_X1  g101(.A(new_n526), .B(KEYINPUT7), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n520), .A2(G51), .ZN(new_n528));
  NAND4_X1  g103(.A1(new_n524), .A2(new_n525), .A3(new_n527), .A4(new_n528), .ZN(G286));
  INV_X1    g104(.A(G286), .ZN(G168));
  AND3_X1   g105(.A1(new_n510), .A2(KEYINPUT5), .A3(G543), .ZN(new_n531));
  AOI21_X1  g106(.A(KEYINPUT5), .B1(new_n510), .B2(G543), .ZN(new_n532));
  OAI21_X1  g107(.A(G64), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(G77), .A2(G543), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n514), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  XNOR2_X1  g110(.A(KEYINPUT6), .B(G651), .ZN(new_n536));
  OAI211_X1 g111(.A(new_n536), .B(G90), .C1(new_n531), .C2(new_n532), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n536), .A2(G52), .A3(G543), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NOR3_X1   g114(.A1(new_n535), .A2(new_n539), .A3(KEYINPUT73), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT73), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n518), .A2(G90), .B1(new_n520), .B2(G52), .ZN(new_n542));
  INV_X1    g117(.A(G64), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n543), .B1(new_n509), .B2(new_n511), .ZN(new_n544));
  INV_X1    g119(.A(new_n534), .ZN(new_n545));
  OAI21_X1  g120(.A(G651), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  AOI21_X1  g121(.A(new_n541), .B1(new_n542), .B2(new_n546), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n540), .A2(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(new_n548), .ZN(G171));
  AOI22_X1  g124(.A1(new_n518), .A2(G81), .B1(new_n520), .B2(G43), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n512), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n550), .B1(new_n514), .B2(new_n551), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT74), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G860), .ZN(G153));
  NAND4_X1  g129(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n555));
  XOR2_X1   g130(.A(new_n555), .B(KEYINPUT75), .Z(G176));
  XOR2_X1   g131(.A(KEYINPUT76), .B(KEYINPUT8), .Z(new_n557));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n557), .B(new_n558), .ZN(new_n559));
  NAND4_X1  g134(.A1(G319), .A2(G483), .A3(G661), .A4(new_n559), .ZN(G188));
  NAND2_X1  g135(.A1(new_n520), .A2(G53), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT9), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n518), .A2(G91), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n512), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n564));
  OAI211_X1 g139(.A(new_n562), .B(new_n563), .C1(new_n514), .C2(new_n564), .ZN(G299));
  OAI21_X1  g140(.A(KEYINPUT73), .B1(new_n535), .B2(new_n539), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n542), .A2(new_n541), .A3(new_n546), .ZN(new_n567));
  AND3_X1   g142(.A1(new_n566), .A2(KEYINPUT77), .A3(new_n567), .ZN(new_n568));
  AOI21_X1  g143(.A(KEYINPUT77), .B1(new_n566), .B2(new_n567), .ZN(new_n569));
  NOR2_X1   g144(.A1(new_n568), .A2(new_n569), .ZN(G301));
  AOI22_X1  g145(.A1(new_n518), .A2(G87), .B1(new_n520), .B2(G49), .ZN(new_n571));
  OAI21_X1  g146(.A(G651), .B1(new_n512), .B2(G74), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n571), .A2(new_n572), .ZN(G288));
  AND2_X1   g148(.A1(new_n512), .A2(G61), .ZN(new_n574));
  NAND2_X1  g149(.A1(G73), .A2(G543), .ZN(new_n575));
  XOR2_X1   g150(.A(new_n575), .B(KEYINPUT78), .Z(new_n576));
  OAI21_X1  g151(.A(G651), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n518), .A2(G86), .B1(new_n520), .B2(G48), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(G305));
  AOI22_X1  g154(.A1(new_n518), .A2(G85), .B1(new_n520), .B2(G47), .ZN(new_n580));
  XOR2_X1   g155(.A(new_n580), .B(KEYINPUT80), .Z(new_n581));
  AOI22_X1  g156(.A1(new_n512), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n582), .A2(new_n514), .ZN(new_n583));
  XNOR2_X1  g158(.A(new_n583), .B(KEYINPUT79), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n581), .A2(new_n584), .ZN(G290));
  NAND2_X1  g160(.A1(new_n512), .A2(G66), .ZN(new_n586));
  INV_X1    g161(.A(G79), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n587), .B2(new_n508), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n588), .A2(G651), .B1(G54), .B2(new_n520), .ZN(new_n589));
  XOR2_X1   g164(.A(KEYINPUT81), .B(KEYINPUT10), .Z(new_n590));
  NAND3_X1  g165(.A1(new_n518), .A2(G92), .A3(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n590), .ZN(new_n592));
  INV_X1    g167(.A(new_n518), .ZN(new_n593));
  INV_X1    g168(.A(G92), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n592), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n589), .A2(new_n591), .A3(new_n595), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n596), .A2(G868), .ZN(new_n597));
  INV_X1    g172(.A(G301), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n597), .B1(new_n598), .B2(G868), .ZN(G321));
  XOR2_X1   g174(.A(G321), .B(KEYINPUT82), .Z(G284));
  INV_X1    g175(.A(G868), .ZN(new_n601));
  NAND2_X1  g176(.A1(G299), .A2(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n602), .B1(new_n601), .B2(G168), .ZN(G297));
  OAI21_X1  g178(.A(new_n602), .B1(new_n601), .B2(G168), .ZN(G280));
  INV_X1    g179(.A(new_n596), .ZN(new_n605));
  INV_X1    g180(.A(G559), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n606), .B2(G860), .ZN(G148));
  INV_X1    g182(.A(new_n553), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(new_n601), .ZN(new_n609));
  NOR2_X1   g184(.A1(new_n596), .A2(G559), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n601), .B2(new_n610), .ZN(G323));
  XNOR2_X1  g186(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g187(.A1(new_n497), .A2(new_n466), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT12), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT13), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(G2100), .ZN(new_n616));
  INV_X1    g191(.A(G123), .ZN(new_n617));
  OAI21_X1  g192(.A(KEYINPUT83), .B1(new_n472), .B2(G111), .ZN(new_n618));
  OR2_X1    g193(.A1(G99), .A2(G2105), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n618), .A2(G2104), .A3(new_n619), .ZN(new_n620));
  NOR3_X1   g195(.A1(new_n472), .A2(KEYINPUT83), .A3(G111), .ZN(new_n621));
  OAI22_X1  g196(.A1(new_n487), .A2(new_n617), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  AOI21_X1  g197(.A(new_n622), .B1(new_n492), .B2(G135), .ZN(new_n623));
  INV_X1    g198(.A(new_n623), .ZN(new_n624));
  OR2_X1    g199(.A1(new_n624), .A2(G2096), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n624), .A2(G2096), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n616), .A2(new_n625), .A3(new_n626), .ZN(G156));
  XNOR2_X1  g202(.A(G2427), .B(G2438), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(G2430), .ZN(new_n629));
  XNOR2_X1  g204(.A(KEYINPUT15), .B(G2435), .ZN(new_n630));
  OR2_X1    g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n629), .A2(new_n630), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n631), .A2(KEYINPUT14), .A3(new_n632), .ZN(new_n633));
  XOR2_X1   g208(.A(G1341), .B(G1348), .Z(new_n634));
  XNOR2_X1  g209(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n633), .B(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(G2451), .B(G2454), .Z(new_n638));
  XNOR2_X1  g213(.A(G2443), .B(G2446), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n637), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n637), .A2(new_n640), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n641), .A2(G14), .A3(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT85), .ZN(G401));
  XOR2_X1   g219(.A(G2084), .B(G2090), .Z(new_n645));
  XNOR2_X1  g220(.A(G2067), .B(G2678), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NOR2_X1   g222(.A1(G2072), .A2(G2078), .ZN(new_n648));
  NOR2_X1   g223(.A1(new_n442), .A2(new_n648), .ZN(new_n649));
  NOR2_X1   g224(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(KEYINPUT86), .B(KEYINPUT18), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  OR2_X1    g227(.A1(new_n645), .A2(new_n646), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n649), .B(KEYINPUT88), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  INV_X1    g230(.A(KEYINPUT17), .ZN(new_n656));
  OAI21_X1  g231(.A(new_n653), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  AOI21_X1  g232(.A(new_n657), .B1(new_n656), .B2(new_n655), .ZN(new_n658));
  INV_X1    g233(.A(KEYINPUT87), .ZN(new_n659));
  AOI21_X1  g234(.A(new_n653), .B1(new_n659), .B2(new_n649), .ZN(new_n660));
  OAI21_X1  g235(.A(new_n660), .B1(new_n659), .B2(new_n649), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n661), .A2(new_n647), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n652), .B1(new_n658), .B2(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(G2096), .B(G2100), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(G227));
  XNOR2_X1  g240(.A(G1971), .B(G1976), .ZN(new_n666));
  INV_X1    g241(.A(KEYINPUT19), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(G1956), .B(G2474), .Z(new_n669));
  XOR2_X1   g244(.A(G1961), .B(G1966), .Z(new_n670));
  AND2_X1   g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT20), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n669), .A2(new_n670), .ZN(new_n674));
  NOR3_X1   g249(.A1(new_n668), .A2(new_n671), .A3(new_n674), .ZN(new_n675));
  AOI21_X1  g250(.A(new_n675), .B1(new_n668), .B2(new_n674), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1991), .B(G1996), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1981), .B(G1986), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(G229));
  MUX2_X1   g258(.A(G23), .B(G288), .S(G16), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT33), .ZN(new_n685));
  INV_X1    g260(.A(G1976), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(G16), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n688), .A2(G6), .ZN(new_n689));
  INV_X1    g264(.A(G305), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n689), .B1(new_n690), .B2(new_n688), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT32), .B(G1981), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT92), .ZN(new_n693));
  XOR2_X1   g268(.A(new_n691), .B(new_n693), .Z(new_n694));
  XOR2_X1   g269(.A(KEYINPUT91), .B(G16), .Z(new_n695));
  NAND2_X1  g270(.A1(new_n695), .A2(G22), .ZN(new_n696));
  XOR2_X1   g271(.A(new_n696), .B(KEYINPUT93), .Z(new_n697));
  INV_X1    g272(.A(new_n695), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n697), .B1(G303), .B2(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(G1971), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  NOR3_X1   g276(.A1(new_n687), .A2(new_n694), .A3(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(KEYINPUT34), .ZN(new_n703));
  OR2_X1    g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n702), .A2(new_n703), .ZN(new_n705));
  MUX2_X1   g280(.A(G24), .B(G290), .S(new_n698), .Z(new_n706));
  XOR2_X1   g281(.A(new_n706), .B(G1986), .Z(new_n707));
  INV_X1    g282(.A(G29), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(G25), .ZN(new_n709));
  OAI21_X1  g284(.A(KEYINPUT89), .B1(G95), .B2(G2105), .ZN(new_n710));
  INV_X1    g285(.A(new_n710), .ZN(new_n711));
  NOR3_X1   g286(.A1(KEYINPUT89), .A2(G95), .A3(G2105), .ZN(new_n712));
  OAI221_X1 g287(.A(G2104), .B1(G107), .B2(new_n472), .C1(new_n711), .C2(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(G119), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n713), .B1(new_n714), .B2(new_n487), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n715), .B1(G131), .B2(new_n492), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n709), .B1(new_n716), .B2(new_n708), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT90), .ZN(new_n718));
  XOR2_X1   g293(.A(KEYINPUT35), .B(G1991), .Z(new_n719));
  XOR2_X1   g294(.A(new_n718), .B(new_n719), .Z(new_n720));
  NAND4_X1  g295(.A1(new_n704), .A2(new_n705), .A3(new_n707), .A4(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(KEYINPUT36), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n722), .A2(KEYINPUT94), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n721), .B(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n605), .A2(G16), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(G4), .B2(G16), .ZN(new_n726));
  XNOR2_X1  g301(.A(KEYINPUT95), .B(G1348), .ZN(new_n727));
  OR2_X1    g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n708), .A2(G32), .ZN(new_n729));
  NAND3_X1  g304(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT100), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(KEYINPUT26), .ZN(new_n732));
  AOI22_X1  g307(.A1(new_n492), .A2(G141), .B1(G105), .B2(new_n466), .ZN(new_n733));
  INV_X1    g308(.A(G129), .ZN(new_n734));
  OR2_X1    g309(.A1(new_n487), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n732), .A2(new_n733), .A3(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(new_n736), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n729), .B1(new_n737), .B2(new_n708), .ZN(new_n738));
  XOR2_X1   g313(.A(KEYINPUT27), .B(G1996), .Z(new_n739));
  NAND2_X1  g314(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n726), .A2(new_n727), .ZN(new_n741));
  NOR2_X1   g316(.A1(G286), .A2(new_n688), .ZN(new_n742));
  INV_X1    g317(.A(KEYINPUT101), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  OAI21_X1  g319(.A(KEYINPUT101), .B1(G16), .B2(G21), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n744), .B1(new_n742), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n746), .A2(G1966), .ZN(new_n747));
  NAND4_X1  g322(.A1(new_n728), .A2(new_n740), .A3(new_n741), .A4(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n695), .A2(G20), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT23), .Z(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(G299), .B2(G16), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(G1956), .ZN(new_n752));
  NOR2_X1   g327(.A1(G29), .A2(G35), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(G162), .B2(G29), .ZN(new_n754));
  XNOR2_X1  g329(.A(KEYINPUT105), .B(KEYINPUT29), .ZN(new_n755));
  INV_X1    g330(.A(G2090), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n754), .B(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n708), .A2(G26), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT98), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT28), .ZN(new_n761));
  OR2_X1    g336(.A1(G104), .A2(G2105), .ZN(new_n762));
  OAI211_X1 g337(.A(new_n762), .B(G2104), .C1(G116), .C2(new_n472), .ZN(new_n763));
  INV_X1    g338(.A(G128), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n763), .B1(new_n487), .B2(new_n764), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(new_n492), .B2(G140), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n761), .B1(new_n766), .B2(new_n708), .ZN(new_n767));
  XOR2_X1   g342(.A(KEYINPUT99), .B(G2067), .Z(new_n768));
  XNOR2_X1  g343(.A(new_n767), .B(new_n768), .ZN(new_n769));
  NAND3_X1  g344(.A1(new_n752), .A2(new_n758), .A3(new_n769), .ZN(new_n770));
  OR2_X1    g345(.A1(G29), .A2(G33), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n492), .A2(G139), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n472), .A2(G103), .A3(G2104), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(KEYINPUT25), .Z(new_n774));
  AOI22_X1  g349(.A1(new_n497), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n775));
  OAI211_X1 g350(.A(new_n772), .B(new_n774), .C1(new_n472), .C2(new_n775), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n771), .B1(new_n776), .B2(new_n708), .ZN(new_n777));
  INV_X1    g352(.A(G2072), .ZN(new_n778));
  AND2_X1   g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g354(.A(KEYINPUT30), .B(G28), .ZN(new_n780));
  OR2_X1    g355(.A1(KEYINPUT31), .A2(G11), .ZN(new_n781));
  NAND2_X1  g356(.A1(KEYINPUT31), .A2(G11), .ZN(new_n782));
  AOI22_X1  g357(.A1(new_n780), .A2(new_n708), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(new_n624), .B2(new_n708), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n777), .A2(new_n778), .ZN(new_n785));
  NOR3_X1   g360(.A1(new_n779), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  OAI221_X1 g361(.A(new_n786), .B1(G1966), .B2(new_n746), .C1(new_n738), .C2(new_n739), .ZN(new_n787));
  NOR3_X1   g362(.A1(new_n748), .A2(new_n770), .A3(new_n787), .ZN(new_n788));
  NOR2_X1   g363(.A1(G5), .A2(G16), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(G171), .B2(G16), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT102), .ZN(new_n791));
  INV_X1    g366(.A(G1961), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n698), .A2(G19), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(new_n553), .B2(new_n698), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT97), .ZN(new_n796));
  XNOR2_X1  g371(.A(KEYINPUT96), .B(G1341), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  NOR2_X1   g373(.A1(G27), .A2(G29), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n799), .B1(G164), .B2(G29), .ZN(new_n800));
  XNOR2_X1  g375(.A(KEYINPUT103), .B(G2078), .ZN(new_n801));
  XOR2_X1   g376(.A(new_n800), .B(new_n801), .Z(new_n802));
  AND2_X1   g377(.A1(new_n802), .A2(KEYINPUT104), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n802), .A2(KEYINPUT104), .ZN(new_n804));
  INV_X1    g379(.A(KEYINPUT24), .ZN(new_n805));
  INV_X1    g380(.A(G34), .ZN(new_n806));
  AOI21_X1  g381(.A(G29), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(new_n805), .B2(new_n806), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(G160), .B2(new_n708), .ZN(new_n809));
  AND2_X1   g384(.A1(new_n809), .A2(G2084), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n809), .A2(G2084), .ZN(new_n811));
  NOR4_X1   g386(.A1(new_n803), .A2(new_n804), .A3(new_n810), .A4(new_n811), .ZN(new_n812));
  AND4_X1   g387(.A1(new_n788), .A2(new_n793), .A3(new_n798), .A4(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n724), .A2(new_n813), .ZN(G150));
  INV_X1    g389(.A(G150), .ZN(G311));
  NAND2_X1  g390(.A1(new_n520), .A2(G55), .ZN(new_n816));
  XOR2_X1   g391(.A(KEYINPUT106), .B(G93), .Z(new_n817));
  AOI22_X1  g392(.A1(new_n512), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n818));
  OAI221_X1 g393(.A(new_n816), .B1(new_n593), .B2(new_n817), .C1(new_n818), .C2(new_n514), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n819), .A2(new_n552), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n820), .B1(new_n608), .B2(new_n819), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT38), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n596), .A2(new_n606), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT39), .ZN(new_n825));
  AOI21_X1  g400(.A(G860), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(new_n825), .B2(new_n824), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n819), .A2(G860), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(KEYINPUT107), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT37), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n827), .A2(new_n830), .ZN(G145));
  NAND2_X1  g406(.A1(new_n776), .A2(KEYINPUT108), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n737), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n736), .A2(KEYINPUT108), .A3(new_n776), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n835), .A2(G164), .ZN(new_n836));
  OR2_X1    g411(.A1(new_n499), .A2(new_n505), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n833), .A2(new_n837), .A3(new_n834), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(new_n766), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n836), .A2(new_n766), .A3(new_n838), .ZN(new_n842));
  INV_X1    g417(.A(G130), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n472), .A2(G118), .ZN(new_n844));
  OAI21_X1  g419(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n845));
  OAI22_X1  g420(.A1(new_n487), .A2(new_n843), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n846), .B1(new_n492), .B2(G142), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(new_n614), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(new_n716), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n841), .A2(new_n842), .A3(new_n849), .ZN(new_n850));
  OR2_X1    g425(.A1(new_n850), .A2(KEYINPUT109), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n841), .A2(new_n842), .ZN(new_n852));
  INV_X1    g427(.A(new_n849), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n850), .A2(KEYINPUT109), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n851), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(G160), .B(new_n624), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(G162), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  XOR2_X1   g434(.A(KEYINPUT110), .B(G37), .Z(new_n860));
  AOI21_X1  g435(.A(new_n858), .B1(new_n852), .B2(new_n853), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT111), .ZN(new_n862));
  NAND4_X1  g437(.A1(new_n841), .A2(new_n849), .A3(new_n862), .A4(new_n842), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n850), .A2(KEYINPUT111), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n861), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  AND2_X1   g440(.A1(new_n865), .A2(KEYINPUT112), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n865), .A2(KEYINPUT112), .ZN(new_n867));
  OAI211_X1 g442(.A(new_n859), .B(new_n860), .C1(new_n866), .C2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(KEYINPUT113), .B(KEYINPUT40), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n868), .B(new_n869), .ZN(G395));
  NAND2_X1  g445(.A1(new_n608), .A2(new_n819), .ZN(new_n871));
  INV_X1    g446(.A(new_n820), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(new_n610), .ZN(new_n874));
  XNOR2_X1  g449(.A(G299), .B(new_n596), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(KEYINPUT41), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  AND2_X1   g452(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n875), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n874), .A2(new_n879), .ZN(new_n880));
  OR3_X1    g455(.A1(new_n878), .A2(new_n880), .A3(KEYINPUT42), .ZN(new_n881));
  XNOR2_X1  g456(.A(G290), .B(G305), .ZN(new_n882));
  XOR2_X1   g457(.A(G303), .B(G288), .Z(new_n883));
  XNOR2_X1  g458(.A(new_n882), .B(new_n883), .ZN(new_n884));
  OAI21_X1  g459(.A(KEYINPUT42), .B1(new_n878), .B2(new_n880), .ZN(new_n885));
  AND3_X1   g460(.A1(new_n881), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n884), .B1(new_n881), .B2(new_n885), .ZN(new_n887));
  OAI21_X1  g462(.A(G868), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n819), .A2(new_n601), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(G295));
  NAND2_X1  g465(.A1(new_n888), .A2(new_n889), .ZN(G331));
  INV_X1    g466(.A(new_n884), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT77), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n893), .B1(new_n540), .B2(new_n547), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n566), .A2(KEYINPUT77), .A3(new_n567), .ZN(new_n895));
  AOI21_X1  g470(.A(G286), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NOR3_X1   g471(.A1(new_n540), .A2(G168), .A3(new_n547), .ZN(new_n897));
  NOR3_X1   g472(.A1(new_n896), .A2(KEYINPUT114), .A3(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT114), .ZN(new_n899));
  OAI21_X1  g474(.A(G168), .B1(new_n568), .B2(new_n569), .ZN(new_n900));
  INV_X1    g475(.A(new_n897), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n899), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n873), .B1(new_n898), .B2(new_n902), .ZN(new_n903));
  OAI21_X1  g478(.A(KEYINPUT114), .B1(new_n896), .B2(new_n897), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n900), .A2(new_n899), .A3(new_n901), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n904), .A2(new_n905), .A3(new_n821), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n903), .A2(new_n879), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(KEYINPUT116), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT116), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n903), .A2(new_n909), .A3(new_n879), .A4(new_n906), .ZN(new_n910));
  AND2_X1   g485(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT115), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n903), .A2(new_n912), .ZN(new_n913));
  OAI211_X1 g488(.A(KEYINPUT115), .B(new_n873), .C1(new_n898), .C2(new_n902), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n913), .A2(new_n906), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(new_n876), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n892), .B1(new_n911), .B2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT43), .ZN(new_n918));
  NAND4_X1  g493(.A1(new_n913), .A2(new_n914), .A3(new_n879), .A4(new_n906), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n903), .A2(new_n906), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(new_n876), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n919), .A2(new_n892), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(new_n860), .ZN(new_n923));
  NOR3_X1   g498(.A1(new_n917), .A2(new_n918), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n919), .A2(new_n921), .ZN(new_n925));
  AOI21_X1  g500(.A(G37), .B1(new_n925), .B2(new_n884), .ZN(new_n926));
  AOI21_X1  g501(.A(KEYINPUT43), .B1(new_n926), .B2(new_n922), .ZN(new_n927));
  OAI21_X1  g502(.A(KEYINPUT44), .B1(new_n924), .B2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT44), .ZN(new_n929));
  NOR3_X1   g504(.A1(new_n917), .A2(KEYINPUT43), .A3(new_n923), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n918), .B1(new_n926), .B2(new_n922), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n929), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n928), .A2(new_n932), .ZN(G397));
  NAND2_X1  g508(.A1(G303), .A2(G8), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n934), .B(KEYINPUT55), .ZN(new_n935));
  XNOR2_X1  g510(.A(KEYINPUT117), .B(G40), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n936), .B1(new_n485), .B2(G2105), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n477), .A2(new_n479), .A3(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(G1384), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n939), .B1(new_n499), .B2(new_n505), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n938), .B1(KEYINPUT50), .B2(new_n940), .ZN(new_n941));
  NOR2_X1   g516(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n942), .B1(new_n499), .B2(new_n505), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n944), .A2(G2090), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n837), .A2(KEYINPUT45), .A3(new_n939), .ZN(new_n946));
  AND3_X1   g521(.A1(new_n477), .A2(new_n479), .A3(new_n937), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT45), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n940), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n946), .A2(new_n947), .A3(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT118), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n946), .A2(KEYINPUT118), .A3(new_n947), .A4(new_n949), .ZN(new_n953));
  AND2_X1   g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n945), .B1(new_n954), .B2(new_n700), .ZN(new_n955));
  INV_X1    g530(.A(G8), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n935), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(new_n940), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n947), .A2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT120), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n959), .A2(new_n960), .A3(G8), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n938), .A2(new_n940), .ZN(new_n962));
  OAI21_X1  g537(.A(KEYINPUT120), .B1(new_n962), .B2(new_n956), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(G305), .A2(G1981), .ZN(new_n965));
  INV_X1    g540(.A(G1981), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n577), .A2(new_n966), .A3(new_n578), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(KEYINPUT49), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT49), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n965), .A2(new_n970), .A3(new_n967), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n964), .A2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT121), .ZN(new_n974));
  XNOR2_X1  g549(.A(new_n973), .B(new_n974), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n571), .A2(G1976), .A3(new_n572), .ZN(new_n976));
  AOI21_X1  g551(.A(KEYINPUT52), .B1(G288), .B2(new_n686), .ZN(new_n977));
  AND3_X1   g552(.A1(new_n964), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n964), .A2(new_n976), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n978), .B1(KEYINPUT52), .B2(new_n979), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n952), .A2(new_n700), .A3(new_n953), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n837), .A2(KEYINPUT119), .A3(new_n942), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT119), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n943), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(new_n941), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n981), .B1(G2090), .B2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(new_n935), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n987), .A2(G8), .A3(new_n988), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n957), .A2(new_n975), .A3(new_n980), .A4(new_n989), .ZN(new_n990));
  XNOR2_X1  g565(.A(G299), .B(KEYINPUT57), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(KEYINPUT123), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT57), .ZN(new_n993));
  XNOR2_X1  g568(.A(G299), .B(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT123), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(G1956), .B1(new_n941), .B2(new_n943), .ZN(new_n997));
  XNOR2_X1  g572(.A(KEYINPUT56), .B(G2072), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n950), .A2(new_n999), .ZN(new_n1000));
  OAI211_X1 g575(.A(new_n992), .B(new_n996), .C1(new_n997), .C2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT61), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n1000), .A2(new_n997), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n1002), .B1(new_n1003), .B2(new_n994), .ZN(new_n1004));
  INV_X1    g579(.A(G1348), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n959), .A2(G2067), .ZN(new_n1006));
  AOI22_X1  g581(.A1(new_n986), .A2(new_n1005), .B1(new_n1006), .B2(KEYINPUT122), .ZN(new_n1007));
  OR2_X1    g582(.A1(new_n1006), .A2(KEYINPUT122), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT60), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n596), .A2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1007), .A2(new_n1008), .A3(new_n1010), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n596), .A2(new_n1009), .ZN(new_n1012));
  AOI22_X1  g587(.A1(new_n1001), .A2(new_n1004), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(G1956), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n944), .A2(new_n1014), .ZN(new_n1015));
  OAI211_X1 g590(.A(new_n1015), .B(new_n994), .C1(new_n950), .C2(new_n999), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n991), .B1(new_n1000), .B2(new_n997), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  XNOR2_X1  g593(.A(KEYINPUT58), .B(G1341), .ZN(new_n1019));
  OAI22_X1  g594(.A1(new_n950), .A2(G1996), .B1(new_n962), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(new_n553), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(KEYINPUT59), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT59), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1020), .A2(new_n1023), .A3(new_n553), .ZN(new_n1024));
  AOI22_X1  g599(.A1(new_n1018), .A2(new_n1002), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1025));
  OR2_X1    g600(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1013), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1028), .A2(new_n605), .A3(new_n1016), .ZN(new_n1029));
  AND2_X1   g604(.A1(new_n1029), .A2(new_n1001), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n990), .B1(new_n1027), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(G1966), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n950), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(G2084), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n985), .A2(new_n1034), .A3(new_n941), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1033), .A2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(G8), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT125), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT51), .ZN(new_n1039));
  NOR2_X1   g614(.A1(G168), .A2(new_n956), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1040), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n1037), .A2(new_n1038), .A3(new_n1039), .A4(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1039), .B1(new_n1037), .B2(new_n1041), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT124), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1042), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n956), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1046));
  OAI211_X1 g621(.A(new_n1044), .B(KEYINPUT51), .C1(new_n1046), .C2(new_n1040), .ZN(new_n1047));
  NOR3_X1   g622(.A1(new_n1046), .A2(KEYINPUT51), .A3(new_n1040), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1047), .B1(new_n1048), .B2(new_n1038), .ZN(new_n1049));
  OAI22_X1  g624(.A1(new_n1045), .A2(new_n1049), .B1(G168), .B2(new_n1037), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT54), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT126), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT53), .ZN(new_n1053));
  OAI211_X1 g628(.A(new_n1052), .B(new_n1053), .C1(new_n954), .C2(G2078), .ZN(new_n1054));
  AOI21_X1  g629(.A(G2078), .B1(new_n952), .B2(new_n953), .ZN(new_n1055));
  OAI21_X1  g630(.A(KEYINPUT126), .B1(new_n1055), .B2(KEYINPUT53), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1054), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(new_n950), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1053), .A2(G2078), .ZN(new_n1059));
  AOI22_X1  g634(.A1(new_n1058), .A2(new_n1059), .B1(new_n986), .B2(new_n792), .ZN(new_n1060));
  AOI21_X1  g635(.A(G301), .B1(new_n1057), .B2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n986), .A2(new_n792), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n946), .A2(new_n949), .ZN(new_n1063));
  NAND3_X1  g638(.A1(G160), .A2(G40), .A3(new_n1059), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1062), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  AOI211_X1 g640(.A(new_n598), .B(new_n1065), .C1(new_n1054), .C2(new_n1056), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1051), .B1(new_n1061), .B2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1057), .A2(G301), .A3(new_n1060), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1065), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1069));
  OAI211_X1 g644(.A(new_n1068), .B(KEYINPUT54), .C1(new_n548), .C2(new_n1069), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1031), .A2(new_n1050), .A3(new_n1067), .A4(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(new_n989), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1072), .A2(new_n975), .A3(new_n980), .ZN(new_n1073));
  NOR2_X1   g648(.A1(G288), .A2(G1976), .ZN(new_n1074));
  AOI22_X1  g649(.A1(new_n975), .A2(new_n1074), .B1(new_n966), .B2(new_n690), .ZN(new_n1075));
  INV_X1    g650(.A(new_n964), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1073), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT63), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1046), .A2(G168), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1078), .B1(new_n990), .B2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n988), .B1(new_n987), .B2(G8), .ZN(new_n1081));
  NOR3_X1   g656(.A1(new_n1081), .A2(new_n1078), .A3(new_n1079), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1082), .A2(new_n989), .A3(new_n975), .A4(new_n980), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1077), .B1(new_n1080), .B2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1050), .A2(KEYINPUT62), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1057), .A2(new_n1060), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(new_n598), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1087), .A2(new_n990), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT62), .ZN(new_n1089));
  OAI221_X1 g664(.A(new_n1089), .B1(G168), .B2(new_n1037), .C1(new_n1045), .C2(new_n1049), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1085), .A2(new_n1088), .A3(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1071), .A2(new_n1084), .A3(new_n1091), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n949), .A2(new_n938), .ZN(new_n1093));
  XOR2_X1   g668(.A(new_n716), .B(new_n719), .Z(new_n1094));
  XOR2_X1   g669(.A(new_n736), .B(G1996), .Z(new_n1095));
  XNOR2_X1  g670(.A(new_n766), .B(G2067), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1094), .A2(new_n1095), .A3(new_n1096), .ZN(new_n1097));
  XNOR2_X1  g672(.A(G290), .B(G1986), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1093), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1092), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1093), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1101), .B1(new_n737), .B2(new_n1096), .ZN(new_n1102));
  OR3_X1    g677(.A1(new_n1101), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1103));
  OAI21_X1  g678(.A(KEYINPUT46), .B1(new_n1101), .B2(G1996), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1102), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  XOR2_X1   g680(.A(new_n1105), .B(KEYINPUT47), .Z(new_n1106));
  NAND4_X1  g681(.A1(new_n1095), .A2(new_n719), .A3(new_n716), .A4(new_n1096), .ZN(new_n1107));
  OR2_X1    g682(.A1(new_n840), .A2(G2067), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1101), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  NOR3_X1   g684(.A1(new_n1101), .A2(G290), .A3(G1986), .ZN(new_n1110));
  OR2_X1    g685(.A1(new_n1110), .A2(KEYINPUT48), .ZN(new_n1111));
  AOI22_X1  g686(.A1(new_n1097), .A2(new_n1093), .B1(new_n1110), .B2(KEYINPUT48), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1109), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1106), .A2(new_n1113), .ZN(new_n1114));
  XOR2_X1   g689(.A(new_n1114), .B(KEYINPUT127), .Z(new_n1115));
  NAND2_X1  g690(.A1(new_n1100), .A2(new_n1115), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g691(.A(new_n643), .ZN(new_n1118));
  NOR4_X1   g692(.A1(G229), .A2(new_n463), .A3(new_n1118), .A4(G227), .ZN(new_n1119));
  OAI211_X1 g693(.A(new_n868), .B(new_n1119), .C1(new_n930), .C2(new_n931), .ZN(G225));
  INV_X1    g694(.A(G225), .ZN(G308));
endmodule


