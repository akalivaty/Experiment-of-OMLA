//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 0 1 1 0 1 0 0 1 0 0 0 0 0 1 1 1 1 1 0 0 1 0 0 0 1 0 1 1 0 0 0 0 0 1 1 1 0 0 1 0 0 1 0 1 0 0 1 0 1 1 1 1 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:46 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n591, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n599, new_n600, new_n601, new_n602,
    new_n603, new_n604, new_n605, new_n606, new_n608, new_n609, new_n610,
    new_n611, new_n612, new_n613, new_n614, new_n615, new_n616, new_n617,
    new_n618, new_n619, new_n620, new_n621, new_n622, new_n623, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n667, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n707, new_n708, new_n709, new_n710,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962;
  OAI21_X1  g000(.A(G210), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(G104), .ZN(new_n188));
  NOR3_X1   g002(.A1(new_n188), .A2(KEYINPUT3), .A3(G107), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT75), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(KEYINPUT74), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT74), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G104), .ZN(new_n193));
  AOI21_X1  g007(.A(G107), .B1(new_n191), .B2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT3), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n190), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  XNOR2_X1  g010(.A(KEYINPUT74), .B(G104), .ZN(new_n197));
  OAI211_X1 g011(.A(KEYINPUT75), .B(KEYINPUT3), .C1(new_n197), .C2(G107), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n189), .B1(new_n196), .B2(new_n198), .ZN(new_n199));
  AOI21_X1  g013(.A(G101), .B1(new_n197), .B2(G107), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT76), .ZN(new_n201));
  INV_X1    g015(.A(G107), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n201), .B1(new_n202), .B2(G104), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n188), .A2(KEYINPUT76), .A3(G107), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  OAI21_X1  g019(.A(G101), .B1(new_n194), .B2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT77), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  OAI211_X1 g022(.A(KEYINPUT77), .B(G101), .C1(new_n194), .C2(new_n205), .ZN(new_n209));
  AOI22_X1  g023(.A1(new_n199), .A2(new_n200), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  XOR2_X1   g024(.A(KEYINPUT2), .B(G113), .Z(new_n211));
  XNOR2_X1  g025(.A(G116), .B(G119), .ZN(new_n212));
  AND2_X1   g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(KEYINPUT5), .ZN(new_n214));
  INV_X1    g028(.A(G116), .ZN(new_n215));
  NOR3_X1   g029(.A1(new_n215), .A2(KEYINPUT5), .A3(G119), .ZN(new_n216));
  INV_X1    g030(.A(G113), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n213), .B1(new_n214), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n210), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(new_n189), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n192), .A2(G104), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n188), .A2(KEYINPUT74), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n202), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  AOI21_X1  g038(.A(KEYINPUT75), .B1(new_n224), .B2(KEYINPUT3), .ZN(new_n225));
  NOR3_X1   g039(.A1(new_n194), .A2(new_n190), .A3(new_n195), .ZN(new_n226));
  OAI211_X1 g040(.A(new_n221), .B(new_n200), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(KEYINPUT4), .ZN(new_n228));
  INV_X1    g042(.A(G101), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n197), .A2(G107), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n229), .B1(new_n199), .B2(new_n230), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n228), .A2(new_n231), .ZN(new_n232));
  OAI211_X1 g046(.A(new_n230), .B(new_n221), .C1(new_n225), .C2(new_n226), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n229), .A2(KEYINPUT4), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n211), .A2(new_n212), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n213), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n235), .A2(new_n238), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n220), .B1(new_n232), .B2(new_n239), .ZN(new_n240));
  XNOR2_X1  g054(.A(G110), .B(G122), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  OAI211_X1 g057(.A(new_n220), .B(new_n241), .C1(new_n232), .C2(new_n239), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n243), .A2(KEYINPUT6), .A3(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(G146), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G143), .ZN(new_n247));
  INV_X1    g061(.A(G143), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(G146), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n247), .A2(new_n249), .A3(KEYINPUT0), .A4(G128), .ZN(new_n250));
  AND2_X1   g064(.A1(new_n247), .A2(new_n249), .ZN(new_n251));
  XNOR2_X1  g065(.A(KEYINPUT0), .B(G128), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n250), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G125), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n247), .A2(new_n249), .ZN(new_n255));
  OAI21_X1  g069(.A(KEYINPUT1), .B1(new_n248), .B2(G146), .ZN(new_n256));
  AND2_X1   g070(.A1(new_n256), .A2(KEYINPUT64), .ZN(new_n257));
  OAI21_X1  g071(.A(G128), .B1(new_n256), .B2(KEYINPUT64), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n255), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(G128), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n260), .A2(KEYINPUT1), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n261), .A2(new_n247), .A3(new_n249), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n259), .A2(new_n262), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n254), .B1(new_n263), .B2(G125), .ZN(new_n264));
  INV_X1    g078(.A(G224), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n265), .A2(G953), .ZN(new_n266));
  XNOR2_X1  g080(.A(new_n264), .B(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT6), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n240), .A2(new_n268), .A3(new_n242), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n245), .A2(new_n267), .A3(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT80), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND4_X1  g086(.A1(new_n245), .A2(KEYINPUT80), .A3(new_n267), .A4(new_n269), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(G902), .ZN(new_n275));
  OAI21_X1  g089(.A(KEYINPUT7), .B1(new_n265), .B2(G953), .ZN(new_n276));
  XOR2_X1   g090(.A(new_n264), .B(new_n276), .Z(new_n277));
  NAND2_X1  g091(.A1(new_n208), .A2(new_n209), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n227), .A2(new_n278), .ZN(new_n279));
  XNOR2_X1  g093(.A(new_n279), .B(new_n219), .ZN(new_n280));
  XOR2_X1   g094(.A(new_n241), .B(KEYINPUT8), .Z(new_n281));
  OAI21_X1  g095(.A(new_n277), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(new_n244), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n275), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n187), .B1(new_n274), .B2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(new_n187), .ZN(new_n287));
  AOI211_X1 g101(.A(new_n287), .B(new_n284), .C1(new_n272), .C2(new_n273), .ZN(new_n288));
  NOR3_X1   g102(.A1(new_n286), .A2(new_n288), .A3(KEYINPUT81), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(KEYINPUT81), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(G214), .B1(G237), .B2(G902), .ZN(new_n293));
  INV_X1    g107(.A(G475), .ZN(new_n294));
  INV_X1    g108(.A(G953), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(KEYINPUT67), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT67), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(G953), .ZN(new_n298));
  AND2_X1   g112(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  XOR2_X1   g113(.A(KEYINPUT66), .B(G237), .Z(new_n300));
  NAND3_X1  g114(.A1(new_n299), .A2(new_n300), .A3(G214), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(new_n248), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n299), .A2(new_n300), .A3(G143), .A4(G214), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT18), .ZN(new_n304));
  INV_X1    g118(.A(G131), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n302), .A2(new_n303), .A3(new_n307), .ZN(new_n308));
  XNOR2_X1  g122(.A(G125), .B(G140), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(new_n246), .ZN(new_n310));
  XNOR2_X1  g124(.A(new_n309), .B(KEYINPUT83), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n310), .B1(new_n311), .B2(new_n246), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n308), .A2(new_n312), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n307), .B1(new_n302), .B2(new_n303), .ZN(new_n314));
  OAI21_X1  g128(.A(KEYINPUT84), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n302), .A2(new_n303), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(new_n306), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT84), .ZN(new_n318));
  NAND4_X1  g132(.A1(new_n317), .A2(new_n318), .A3(new_n312), .A4(new_n308), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n305), .B1(new_n302), .B2(new_n303), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT17), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n302), .A2(new_n305), .A3(new_n303), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n321), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n309), .A2(KEYINPUT16), .ZN(new_n325));
  INV_X1    g139(.A(G140), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(G125), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n325), .B1(KEYINPUT16), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(new_n246), .ZN(new_n329));
  OAI211_X1 g143(.A(new_n325), .B(G146), .C1(KEYINPUT16), .C2(new_n327), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n331), .B1(new_n320), .B2(KEYINPUT17), .ZN(new_n332));
  AOI22_X1  g146(.A1(new_n315), .A2(new_n319), .B1(new_n324), .B2(new_n332), .ZN(new_n333));
  XNOR2_X1  g147(.A(G113), .B(G122), .ZN(new_n334));
  XNOR2_X1  g148(.A(new_n334), .B(new_n188), .ZN(new_n335));
  XNOR2_X1  g149(.A(new_n333), .B(new_n335), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n294), .B1(new_n336), .B2(new_n275), .ZN(new_n337));
  XOR2_X1   g151(.A(KEYINPUT82), .B(KEYINPUT20), .Z(new_n338));
  NAND2_X1  g152(.A1(new_n315), .A2(new_n319), .ZN(new_n339));
  INV_X1    g153(.A(new_n330), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n311), .A2(KEYINPUT19), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n341), .B1(KEYINPUT19), .B2(new_n309), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n340), .B1(new_n342), .B2(new_n246), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n321), .A2(new_n323), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n335), .B1(new_n339), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(KEYINPUT85), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT85), .ZN(new_n348));
  AOI22_X1  g162(.A1(new_n315), .A2(new_n319), .B1(new_n343), .B2(new_n344), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n348), .B1(new_n349), .B2(new_n335), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n333), .A2(new_n335), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n347), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  NOR2_X1   g166(.A1(G475), .A2(G902), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n338), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT20), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n352), .A2(new_n356), .A3(new_n353), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n337), .B1(new_n355), .B2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(G952), .ZN(new_n359));
  AOI211_X1 g173(.A(G953), .B(new_n359), .C1(G234), .C2(G237), .ZN(new_n360));
  INV_X1    g174(.A(new_n299), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n275), .B1(G234), .B2(G237), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  XNOR2_X1  g177(.A(new_n363), .B(KEYINPUT91), .ZN(new_n364));
  XNOR2_X1  g178(.A(KEYINPUT21), .B(G898), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n360), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  XNOR2_X1  g181(.A(KEYINPUT9), .B(G234), .ZN(new_n368));
  INV_X1    g182(.A(G217), .ZN(new_n369));
  NOR3_X1   g183(.A1(new_n368), .A2(new_n369), .A3(G953), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n260), .A2(G143), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n248), .A2(G128), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT88), .ZN(new_n375));
  XNOR2_X1  g189(.A(new_n374), .B(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(G134), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  XNOR2_X1  g192(.A(G116), .B(G122), .ZN(new_n379));
  XNOR2_X1  g193(.A(new_n379), .B(new_n202), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT86), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n382), .B1(new_n372), .B2(KEYINPUT13), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT13), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n373), .A2(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n383), .B1(new_n385), .B2(new_n372), .ZN(new_n386));
  INV_X1    g200(.A(new_n372), .ZN(new_n387));
  OAI211_X1 g201(.A(new_n387), .B(new_n382), .C1(new_n384), .C2(new_n373), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n386), .A2(G134), .A3(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT87), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  OR2_X1    g205(.A1(new_n389), .A2(new_n390), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n381), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT14), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n379), .A2(new_n394), .ZN(new_n395));
  AND2_X1   g209(.A1(new_n215), .A2(G122), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n202), .B1(new_n396), .B2(KEYINPUT14), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n379), .A2(new_n202), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT89), .ZN(new_n399));
  AOI22_X1  g213(.A1(new_n395), .A2(new_n397), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n400), .B1(new_n399), .B2(new_n398), .ZN(new_n401));
  XNOR2_X1  g215(.A(new_n374), .B(KEYINPUT88), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(G134), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n401), .B1(new_n378), .B2(new_n403), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n371), .B1(new_n393), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n392), .A2(new_n391), .ZN(new_n406));
  INV_X1    g220(.A(new_n381), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n404), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n408), .A2(new_n409), .A3(new_n370), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n405), .A2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT90), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n411), .A2(new_n412), .A3(new_n275), .ZN(new_n413));
  INV_X1    g227(.A(G478), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n414), .A2(KEYINPUT15), .ZN(new_n415));
  AND2_X1   g229(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n413), .A2(new_n415), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n358), .A2(new_n367), .A3(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(G469), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n299), .A2(G227), .ZN(new_n421));
  XOR2_X1   g235(.A(G110), .B(G140), .Z(new_n422));
  XNOR2_X1  g236(.A(new_n421), .B(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n263), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n279), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n256), .A2(G128), .ZN(new_n426));
  AOI22_X1  g240(.A1(new_n255), .A2(new_n426), .B1(new_n262), .B2(KEYINPUT78), .ZN(new_n427));
  OR2_X1    g241(.A1(new_n262), .A2(KEYINPUT78), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n227), .A2(new_n278), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n425), .A2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT11), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n432), .B1(new_n377), .B2(G137), .ZN(new_n433));
  INV_X1    g247(.A(G137), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n434), .A2(KEYINPUT11), .A3(G134), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n377), .A2(G137), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n433), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(G131), .ZN(new_n438));
  NAND4_X1  g252(.A1(new_n433), .A2(new_n435), .A3(new_n305), .A4(new_n436), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n431), .A2(KEYINPUT12), .A3(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT12), .ZN(new_n442));
  AOI22_X1  g256(.A1(new_n208), .A2(new_n209), .B1(new_n428), .B2(new_n427), .ZN(new_n443));
  AOI22_X1  g257(.A1(new_n279), .A2(new_n424), .B1(new_n443), .B2(new_n227), .ZN(new_n444));
  INV_X1    g258(.A(new_n440), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n442), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT10), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n447), .B1(new_n259), .B2(new_n262), .ZN(new_n448));
  AOI22_X1  g262(.A1(new_n430), .A2(new_n447), .B1(new_n210), .B2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(new_n253), .ZN(new_n450));
  OAI211_X1 g264(.A(new_n450), .B(new_n235), .C1(new_n228), .C2(new_n231), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n449), .A2(new_n451), .A3(new_n445), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT79), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n449), .A2(new_n451), .A3(KEYINPUT79), .A4(new_n445), .ZN(new_n455));
  AOI221_X4 g269(.A(new_n423), .B1(new_n441), .B2(new_n446), .C1(new_n454), .C2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(new_n423), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n454), .A2(new_n455), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n449), .A2(new_n451), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(new_n440), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n457), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  OAI211_X1 g275(.A(new_n420), .B(new_n275), .C1(new_n456), .C2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(G469), .A2(G902), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n458), .A2(new_n460), .A3(new_n457), .ZN(new_n464));
  AOI22_X1  g278(.A1(new_n454), .A2(new_n455), .B1(new_n441), .B2(new_n446), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n464), .B(G469), .C1(new_n457), .C2(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n462), .A2(new_n463), .A3(new_n466), .ZN(new_n467));
  OAI21_X1  g281(.A(G221), .B1(new_n368), .B2(G902), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n419), .A2(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n369), .B1(G234), .B2(new_n275), .ZN(new_n471));
  INV_X1    g285(.A(G119), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n472), .A2(G128), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n472), .A2(G128), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  XNOR2_X1  g290(.A(KEYINPUT24), .B(G110), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n260), .A2(KEYINPUT23), .A3(G119), .ZN(new_n479));
  OAI211_X1 g293(.A(new_n479), .B(new_n475), .C1(new_n473), .C2(KEYINPUT23), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n478), .B1(new_n480), .B2(G110), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n481), .A2(new_n310), .A3(new_n330), .ZN(new_n482));
  XNOR2_X1  g296(.A(new_n482), .B(KEYINPUT71), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n480), .A2(G110), .ZN(new_n484));
  XOR2_X1   g298(.A(new_n484), .B(KEYINPUT69), .Z(new_n485));
  INV_X1    g299(.A(KEYINPUT70), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n476), .A2(new_n477), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n487), .B1(new_n329), .B2(new_n330), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n485), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n486), .B1(new_n485), .B2(new_n488), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n483), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n299), .A2(G221), .A3(G234), .ZN(new_n493));
  XNOR2_X1  g307(.A(new_n493), .B(KEYINPUT72), .ZN(new_n494));
  XNOR2_X1  g308(.A(KEYINPUT22), .B(G137), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n494), .B(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n492), .A2(new_n497), .ZN(new_n498));
  OAI211_X1 g312(.A(new_n496), .B(new_n483), .C1(new_n490), .C2(new_n491), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g314(.A(KEYINPUT25), .B1(new_n500), .B2(new_n275), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT25), .ZN(new_n502));
  AOI211_X1 g316(.A(new_n502), .B(G902), .C1(new_n498), .C2(new_n499), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n471), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n471), .A2(G902), .ZN(new_n505));
  XNOR2_X1  g319(.A(new_n505), .B(KEYINPUT73), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n500), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT29), .ZN(new_n510));
  INV_X1    g324(.A(new_n436), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n377), .A2(G137), .ZN(new_n512));
  OAI21_X1  g326(.A(G131), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(new_n439), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n514), .B1(new_n259), .B2(new_n262), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n253), .B1(new_n438), .B2(new_n439), .ZN(new_n516));
  NOR3_X1   g330(.A1(new_n515), .A2(new_n516), .A3(KEYINPUT30), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  OAI21_X1  g332(.A(KEYINPUT30), .B1(new_n515), .B2(new_n516), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n237), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(new_n514), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n263), .A2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(new_n516), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n522), .A2(new_n523), .A3(new_n237), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(KEYINPUT65), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n515), .A2(new_n516), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT65), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n526), .A2(new_n527), .A3(new_n237), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n525), .A2(new_n528), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n520), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n299), .A2(new_n300), .A3(G210), .ZN(new_n531));
  XNOR2_X1  g345(.A(new_n531), .B(KEYINPUT27), .ZN(new_n532));
  XNOR2_X1  g346(.A(KEYINPUT26), .B(G101), .ZN(new_n533));
  XNOR2_X1  g347(.A(new_n532), .B(new_n533), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n510), .B1(new_n530), .B2(new_n534), .ZN(new_n535));
  AOI21_X1  g349(.A(KEYINPUT28), .B1(new_n526), .B2(new_n237), .ZN(new_n536));
  INV_X1    g350(.A(new_n534), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n238), .B1(new_n515), .B2(new_n516), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n525), .A2(new_n538), .A3(new_n528), .ZN(new_n539));
  AOI211_X1 g353(.A(new_n536), .B(new_n537), .C1(new_n539), .C2(KEYINPUT28), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n535), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n536), .B1(new_n539), .B2(KEYINPUT28), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n542), .A2(KEYINPUT29), .A3(new_n534), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(new_n275), .ZN(new_n544));
  OAI21_X1  g358(.A(G472), .B1(new_n541), .B2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT30), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n546), .B1(new_n522), .B2(new_n523), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n238), .B1(new_n547), .B2(new_n517), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n548), .A2(new_n525), .A3(new_n528), .A4(new_n534), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(KEYINPUT31), .ZN(new_n550));
  AND2_X1   g364(.A1(new_n525), .A2(new_n528), .ZN(new_n551));
  XNOR2_X1  g365(.A(KEYINPUT68), .B(KEYINPUT31), .ZN(new_n552));
  NAND4_X1  g366(.A1(new_n551), .A2(new_n534), .A3(new_n548), .A4(new_n552), .ZN(new_n553));
  OAI211_X1 g367(.A(new_n550), .B(new_n553), .C1(new_n542), .C2(new_n534), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT32), .ZN(new_n555));
  NOR2_X1   g369(.A1(G472), .A2(G902), .ZN(new_n556));
  AND3_X1   g370(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n555), .B1(new_n554), .B2(new_n556), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n545), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n509), .A2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  NAND4_X1  g375(.A1(new_n292), .A2(new_n293), .A3(new_n470), .A4(new_n561), .ZN(new_n562));
  XNOR2_X1  g376(.A(new_n562), .B(G101), .ZN(G3));
  INV_X1    g377(.A(G472), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n564), .B1(new_n554), .B2(new_n275), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(KEYINPUT92), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n554), .A2(new_n556), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT92), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n565), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n567), .A2(new_n568), .A3(new_n570), .ZN(new_n571));
  NOR3_X1   g385(.A1(new_n571), .A2(new_n469), .A3(new_n508), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n293), .B1(new_n286), .B2(new_n288), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n337), .ZN(new_n575));
  INV_X1    g389(.A(new_n357), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n575), .B1(new_n576), .B2(new_n354), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n411), .A2(new_n414), .A3(new_n275), .ZN(new_n578));
  NAND2_X1  g392(.A1(G478), .A2(G902), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  OAI21_X1  g394(.A(KEYINPUT33), .B1(new_n370), .B2(KEYINPUT93), .ZN(new_n581));
  OR2_X1    g395(.A1(new_n411), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n411), .A2(new_n581), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n580), .B1(new_n584), .B2(G478), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n577), .A2(new_n585), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n586), .A2(new_n366), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n572), .A2(new_n574), .A3(new_n587), .ZN(new_n588));
  XOR2_X1   g402(.A(KEYINPUT34), .B(G104), .Z(new_n589));
  XNOR2_X1  g403(.A(new_n588), .B(new_n589), .ZN(G6));
  XNOR2_X1  g404(.A(new_n413), .B(new_n415), .ZN(new_n591));
  AND3_X1   g405(.A1(new_n352), .A2(new_n338), .A3(new_n353), .ZN(new_n592));
  OAI211_X1 g406(.A(new_n591), .B(new_n575), .C1(new_n592), .C2(new_n354), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n593), .A2(new_n366), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n572), .A2(new_n574), .A3(new_n594), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n595), .B(KEYINPUT94), .ZN(new_n596));
  XNOR2_X1  g410(.A(KEYINPUT35), .B(G107), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n596), .B(new_n597), .ZN(G9));
  NOR2_X1   g412(.A1(new_n496), .A2(KEYINPUT36), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n492), .B(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(new_n506), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n504), .A2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n571), .A2(new_n603), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n292), .A2(new_n293), .A3(new_n470), .A4(new_n604), .ZN(new_n605));
  XOR2_X1   g419(.A(KEYINPUT37), .B(G110), .Z(new_n606));
  XNOR2_X1  g420(.A(new_n605), .B(new_n606), .ZN(G12));
  INV_X1    g421(.A(new_n353), .ZN(new_n608));
  AOI22_X1  g422(.A1(new_n346), .A2(KEYINPUT85), .B1(new_n333), .B2(new_n335), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n608), .B1(new_n609), .B2(new_n350), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(new_n338), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n337), .B1(new_n355), .B2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT96), .ZN(new_n613));
  INV_X1    g427(.A(G900), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n360), .B1(new_n364), .B2(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(KEYINPUT95), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n612), .A2(new_n613), .A3(new_n591), .A4(new_n617), .ZN(new_n618));
  OAI21_X1  g432(.A(KEYINPUT96), .B1(new_n593), .B2(new_n616), .ZN(new_n619));
  AND2_X1   g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n467), .A2(new_n559), .A3(new_n468), .A4(new_n602), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n621), .A2(new_n573), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n623), .B(G128), .ZN(G30));
  NAND2_X1  g438(.A1(new_n274), .A2(new_n285), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n625), .A2(new_n287), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT81), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n274), .A2(new_n187), .A3(new_n285), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n626), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(new_n290), .ZN(new_n630));
  XOR2_X1   g444(.A(KEYINPUT97), .B(KEYINPUT38), .Z(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XOR2_X1   g446(.A(new_n616), .B(KEYINPUT39), .Z(new_n633));
  NAND3_X1  g447(.A1(new_n467), .A2(new_n468), .A3(new_n633), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n634), .A2(KEYINPUT40), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n634), .A2(KEYINPUT40), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n568), .A2(KEYINPUT32), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n530), .A2(new_n537), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n275), .B1(new_n539), .B2(new_n534), .ZN(new_n641));
  OAI21_X1  g455(.A(G472), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n639), .A2(new_n642), .ZN(new_n643));
  OAI21_X1  g457(.A(new_n357), .B1(new_n338), .B2(new_n610), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n418), .B1(new_n644), .B2(new_n575), .ZN(new_n645));
  INV_X1    g459(.A(new_n293), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n602), .A2(new_n646), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n636), .A2(new_n643), .A3(new_n645), .A4(new_n647), .ZN(new_n648));
  OR3_X1    g462(.A1(new_n632), .A2(new_n635), .A3(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(G143), .ZN(G45));
  INV_X1    g464(.A(new_n621), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n577), .A2(new_n585), .A3(new_n617), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n651), .A2(new_n574), .A3(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT98), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n622), .A2(KEYINPUT98), .A3(new_n653), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(G146), .ZN(G48));
  NOR2_X1   g473(.A1(new_n456), .A2(new_n461), .ZN(new_n660));
  OAI21_X1  g474(.A(G469), .B1(new_n660), .B2(G902), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n661), .A2(new_n468), .A3(new_n462), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n560), .A2(new_n662), .ZN(new_n663));
  AND3_X1   g477(.A1(new_n663), .A2(new_n574), .A3(new_n587), .ZN(new_n664));
  XOR2_X1   g478(.A(KEYINPUT41), .B(G113), .Z(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G15));
  AND3_X1   g480(.A1(new_n663), .A2(new_n574), .A3(new_n594), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(new_n215), .ZN(G18));
  NOR2_X1   g482(.A1(new_n573), .A2(new_n662), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n559), .A2(new_n602), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n419), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G119), .ZN(G21));
  OAI211_X1 g487(.A(new_n645), .B(new_n293), .C1(new_n288), .C2(new_n286), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n550), .B1(new_n542), .B2(new_n534), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT99), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  OAI211_X1 g492(.A(new_n550), .B(KEYINPUT99), .C1(new_n542), .C2(new_n534), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n678), .A2(new_n679), .A3(new_n553), .ZN(new_n680));
  AND2_X1   g494(.A1(new_n680), .A2(new_n556), .ZN(new_n681));
  NOR3_X1   g495(.A1(new_n681), .A2(new_n508), .A3(new_n565), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n662), .A2(new_n366), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n675), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G122), .ZN(G24));
  NAND2_X1  g499(.A1(new_n680), .A2(new_n556), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n686), .A2(new_n602), .A3(new_n566), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n652), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n669), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G125), .ZN(G27));
  NAND2_X1  g504(.A1(new_n467), .A2(KEYINPUT100), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT100), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n462), .A2(new_n692), .A3(new_n463), .A4(new_n466), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n691), .A2(new_n468), .A3(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT101), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n646), .B1(new_n629), .B2(new_n290), .ZN(new_n697));
  INV_X1    g511(.A(new_n468), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n698), .B1(new_n467), .B2(KEYINPUT100), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n699), .A2(KEYINPUT101), .A3(new_n693), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n696), .A2(new_n697), .A3(new_n561), .A4(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT42), .ZN(new_n702));
  OR3_X1    g516(.A1(new_n701), .A2(new_n702), .A3(new_n652), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n702), .B1(new_n701), .B2(new_n652), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G131), .ZN(G33));
  OAI21_X1  g520(.A(new_n293), .B1(new_n289), .B2(new_n291), .ZN(new_n707));
  AOI21_X1  g521(.A(KEYINPUT101), .B1(new_n699), .B2(new_n693), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n709), .A2(new_n561), .A3(new_n620), .A4(new_n700), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G134), .ZN(G36));
  NAND2_X1  g525(.A1(new_n358), .A2(new_n585), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(KEYINPUT43), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT43), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n358), .A2(new_n714), .A3(new_n585), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(new_n716), .ZN(new_n717));
  AND2_X1   g531(.A1(new_n571), .A2(new_n602), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n717), .A2(KEYINPUT44), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(new_n697), .ZN(new_n720));
  AOI21_X1  g534(.A(KEYINPUT44), .B1(new_n717), .B2(new_n718), .ZN(new_n721));
  INV_X1    g535(.A(new_n633), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n464), .B1(new_n457), .B2(new_n465), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT45), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n420), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n725), .B1(new_n724), .B2(new_n723), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(new_n463), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT46), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n726), .A2(KEYINPUT46), .A3(new_n463), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n729), .A2(new_n462), .A3(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(new_n468), .ZN(new_n732));
  NOR4_X1   g546(.A1(new_n720), .A2(new_n721), .A3(new_n722), .A4(new_n732), .ZN(new_n733));
  XOR2_X1   g547(.A(KEYINPUT102), .B(G137), .Z(new_n734));
  XNOR2_X1  g548(.A(new_n733), .B(new_n734), .ZN(G39));
  INV_X1    g549(.A(KEYINPUT47), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n732), .B(new_n736), .ZN(new_n737));
  NOR3_X1   g551(.A1(new_n652), .A2(new_n509), .A3(new_n559), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n697), .A2(new_n738), .ZN(new_n739));
  XOR2_X1   g553(.A(new_n739), .B(KEYINPUT103), .Z(new_n740));
  NAND2_X1  g554(.A1(new_n737), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G140), .ZN(G42));
  NAND2_X1  g556(.A1(new_n682), .A2(new_n360), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n716), .A2(new_n743), .ZN(new_n744));
  AOI211_X1 g558(.A(new_n359), .B(G953), .C1(new_n744), .C2(new_n669), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n509), .A2(new_n639), .A3(new_n642), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n661), .A2(new_n468), .A3(new_n462), .A4(new_n360), .ZN(new_n747));
  NOR3_X1   g561(.A1(new_n707), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(new_n586), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n745), .A2(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT48), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n707), .A2(new_n747), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n753), .A2(new_n561), .A3(new_n717), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n751), .B1(new_n752), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n661), .A2(new_n462), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(KEYINPUT104), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT109), .ZN(new_n758));
  AND2_X1   g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n757), .A2(new_n758), .ZN(new_n760));
  NOR3_X1   g574(.A1(new_n759), .A2(new_n760), .A3(new_n468), .ZN(new_n761));
  OAI211_X1 g575(.A(new_n697), .B(new_n744), .C1(new_n737), .C2(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(KEYINPUT51), .ZN(new_n763));
  NOR4_X1   g577(.A1(new_n716), .A2(new_n743), .A3(new_n293), .A4(new_n662), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n764), .A2(new_n632), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT50), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n662), .A2(new_n293), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n632), .A2(KEYINPUT50), .A3(new_n744), .A4(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(new_n687), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n753), .A2(new_n771), .A3(new_n717), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(KEYINPUT110), .ZN(new_n773));
  OR2_X1    g587(.A1(new_n577), .A2(new_n585), .ZN(new_n774));
  INV_X1    g588(.A(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n748), .A2(new_n775), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n770), .A2(new_n773), .A3(new_n776), .ZN(new_n777));
  OAI221_X1 g591(.A(new_n755), .B1(new_n752), .B2(new_n754), .C1(new_n763), .C2(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT111), .ZN(new_n779));
  INV_X1    g593(.A(new_n769), .ZN(new_n780));
  AOI21_X1  g594(.A(KEYINPUT50), .B1(new_n764), .B2(new_n632), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n776), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT110), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n772), .B(new_n783), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n779), .B1(new_n782), .B2(new_n784), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n770), .A2(new_n773), .A3(KEYINPUT111), .A4(new_n776), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n785), .A2(new_n786), .A3(new_n762), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT51), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n789), .A2(KEYINPUT112), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT112), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n787), .A2(new_n791), .A3(new_n788), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n778), .B1(new_n790), .B2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(new_n620), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n701), .A2(new_n794), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n696), .A2(new_n697), .A3(new_n688), .A4(new_n700), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n591), .A2(new_n616), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n697), .A2(new_n612), .A3(new_n651), .A4(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  OAI21_X1  g613(.A(KEYINPUT106), .B1(new_n795), .B2(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT106), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n710), .A2(new_n801), .A3(new_n798), .A4(new_n796), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  AOI22_X1  g617(.A1(new_n620), .A2(new_n622), .B1(new_n669), .B2(new_n688), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n643), .A2(new_n603), .A3(new_n617), .ZN(new_n805));
  OR3_X1    g619(.A1(new_n694), .A2(new_n674), .A3(new_n805), .ZN(new_n806));
  AOI21_X1  g620(.A(KEYINPUT98), .B1(new_n622), .B2(new_n653), .ZN(new_n807));
  NOR4_X1   g621(.A1(new_n621), .A2(new_n573), .A3(new_n652), .A4(new_n655), .ZN(new_n808));
  OAI211_X1 g622(.A(new_n804), .B(new_n806), .C1(new_n807), .C2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT52), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n658), .A2(KEYINPUT52), .A3(new_n804), .A4(new_n806), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n577), .A2(new_n366), .A3(new_n418), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n629), .A2(new_n814), .A3(new_n293), .A4(new_n290), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT105), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n817), .A2(new_n572), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n815), .A2(new_n816), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n572), .A2(new_n292), .A3(new_n293), .A4(new_n587), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n821), .A2(new_n562), .A3(new_n605), .ZN(new_n822));
  OAI211_X1 g636(.A(new_n663), .B(new_n574), .C1(new_n587), .C2(new_n594), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n823), .A2(new_n684), .A3(new_n672), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n820), .A2(new_n822), .A3(new_n824), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n803), .A2(new_n813), .A3(new_n705), .A4(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT53), .ZN(new_n827));
  OR2_X1    g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n826), .A2(new_n827), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n828), .A2(KEYINPUT107), .A3(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT107), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n826), .A2(new_n831), .A3(new_n827), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n830), .A2(KEYINPUT54), .A3(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT108), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n824), .A2(new_n834), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n823), .A2(new_n684), .A3(KEYINPUT108), .A4(new_n672), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n835), .A2(KEYINPUT53), .A3(new_n836), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n837), .A2(new_n820), .A3(new_n822), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n838), .A2(new_n705), .A3(new_n803), .A4(new_n813), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT54), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n829), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n793), .A2(new_n833), .A3(new_n841), .ZN(new_n842));
  NOR2_X1   g656(.A1(G952), .A2(G953), .ZN(new_n843));
  XNOR2_X1  g657(.A(new_n843), .B(KEYINPUT113), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n358), .A2(new_n293), .A3(new_n468), .A4(new_n585), .ZN(new_n846));
  AOI211_X1 g660(.A(new_n746), .B(new_n846), .C1(new_n757), .C2(KEYINPUT49), .ZN(new_n847));
  OAI211_X1 g661(.A(new_n847), .B(new_n632), .C1(KEYINPUT49), .C2(new_n757), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n845), .A2(new_n848), .ZN(G75));
  NOR2_X1   g663(.A1(new_n299), .A2(G952), .ZN(new_n850));
  INV_X1    g664(.A(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT56), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n829), .A2(new_n839), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(G902), .ZN(new_n854));
  INV_X1    g668(.A(G210), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n852), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n245), .A2(new_n269), .ZN(new_n857));
  XNOR2_X1  g671(.A(new_n857), .B(new_n267), .ZN(new_n858));
  XOR2_X1   g672(.A(new_n858), .B(KEYINPUT55), .Z(new_n859));
  OAI21_X1  g673(.A(new_n851), .B1(new_n856), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n856), .A2(new_n859), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT114), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n856), .A2(KEYINPUT114), .A3(new_n859), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n860), .B1(new_n863), .B2(new_n864), .ZN(G51));
  INV_X1    g679(.A(KEYINPUT115), .ZN(new_n866));
  AOI211_X1 g680(.A(new_n275), .B(new_n726), .C1(new_n829), .C2(new_n839), .ZN(new_n867));
  XOR2_X1   g681(.A(new_n463), .B(KEYINPUT57), .Z(new_n868));
  AND3_X1   g682(.A1(new_n829), .A2(new_n840), .A3(new_n839), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n840), .B1(new_n829), .B2(new_n839), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n868), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(new_n660), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n867), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n866), .B1(new_n873), .B2(new_n850), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n853), .A2(KEYINPUT54), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(new_n841), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n660), .B1(new_n876), .B2(new_n868), .ZN(new_n877));
  OAI211_X1 g691(.A(KEYINPUT115), .B(new_n851), .C1(new_n877), .C2(new_n867), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n874), .A2(new_n878), .ZN(G54));
  INV_X1    g693(.A(new_n352), .ZN(new_n880));
  NAND2_X1  g694(.A1(KEYINPUT58), .A2(G475), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n880), .B1(new_n854), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(KEYINPUT117), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT117), .ZN(new_n884));
  OAI211_X1 g698(.A(new_n884), .B(new_n880), .C1(new_n854), .C2(new_n881), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(new_n881), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n853), .A2(G902), .A3(new_n352), .A4(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT116), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n888), .B(new_n889), .ZN(new_n890));
  AND3_X1   g704(.A1(new_n886), .A2(new_n851), .A3(new_n890), .ZN(G60));
  INV_X1    g705(.A(new_n876), .ZN(new_n892));
  XOR2_X1   g706(.A(new_n579), .B(KEYINPUT59), .Z(new_n893));
  INV_X1    g707(.A(new_n893), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n582), .A2(new_n583), .A3(new_n894), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n851), .B1(new_n892), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n833), .A2(new_n841), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(new_n894), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n896), .B1(new_n898), .B2(new_n584), .ZN(G63));
  XOR2_X1   g713(.A(KEYINPUT118), .B(KEYINPUT61), .Z(new_n900));
  NAND2_X1  g714(.A1(G217), .A2(G902), .ZN(new_n901));
  XOR2_X1   g715(.A(new_n901), .B(KEYINPUT60), .Z(new_n902));
  AOI21_X1  g716(.A(new_n500), .B1(new_n853), .B2(new_n902), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n903), .A2(new_n850), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n853), .A2(new_n600), .A3(new_n902), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT119), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n904), .A2(new_n907), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n905), .A2(new_n906), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n900), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n904), .A2(KEYINPUT61), .A3(new_n905), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(G66));
  OAI21_X1  g726(.A(G953), .B1(new_n365), .B2(new_n265), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n913), .B1(new_n825), .B2(new_n361), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n857), .B1(G898), .B2(new_n299), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n915), .B(KEYINPUT120), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n914), .B(new_n916), .ZN(G69));
  AOI21_X1  g731(.A(new_n749), .B1(new_n358), .B2(new_n591), .ZN(new_n918));
  NOR4_X1   g732(.A1(new_n918), .A2(new_n707), .A3(new_n560), .A4(new_n634), .ZN(new_n919));
  AOI211_X1 g733(.A(new_n919), .B(new_n733), .C1(new_n737), .C2(new_n740), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n649), .A2(new_n658), .A3(new_n804), .ZN(new_n921));
  OR2_X1    g735(.A1(new_n921), .A2(KEYINPUT62), .ZN(new_n922));
  AOI21_X1  g736(.A(KEYINPUT121), .B1(new_n921), .B2(KEYINPUT62), .ZN(new_n923));
  AND3_X1   g737(.A1(new_n921), .A2(KEYINPUT121), .A3(KEYINPUT62), .ZN(new_n924));
  OAI211_X1 g738(.A(new_n920), .B(new_n922), .C1(new_n923), .C2(new_n924), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n547), .A2(new_n517), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n926), .B(new_n342), .Z(new_n927));
  INV_X1    g741(.A(new_n927), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n925), .A2(new_n299), .A3(new_n928), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n733), .B1(new_n737), .B2(new_n740), .ZN(new_n930));
  NOR4_X1   g744(.A1(new_n732), .A2(new_n560), .A3(new_n722), .A4(new_n674), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT123), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n931), .B(new_n932), .ZN(new_n933));
  AND3_X1   g747(.A1(new_n710), .A2(new_n658), .A3(new_n804), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n930), .A2(new_n933), .A3(new_n705), .A4(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n935), .A2(new_n299), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n299), .A2(G900), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n937), .B(KEYINPUT122), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n936), .A2(new_n927), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n299), .B1(G227), .B2(G900), .ZN(new_n940));
  OAI211_X1 g754(.A(new_n929), .B(new_n939), .C1(KEYINPUT124), .C2(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n940), .A2(KEYINPUT124), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n941), .B(new_n942), .ZN(G72));
  NAND2_X1  g757(.A1(G472), .A2(G902), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n944), .B(KEYINPUT63), .Z(new_n945));
  XNOR2_X1  g759(.A(new_n945), .B(KEYINPUT125), .ZN(new_n946));
  INV_X1    g760(.A(new_n825), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n946), .B1(new_n925), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n948), .A2(KEYINPUT126), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT126), .ZN(new_n950));
  OAI211_X1 g764(.A(new_n950), .B(new_n946), .C1(new_n925), .C2(new_n947), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n949), .A2(new_n640), .A3(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(new_n945), .ZN(new_n953));
  NOR3_X1   g767(.A1(new_n520), .A2(new_n529), .A3(new_n534), .ZN(new_n954));
  NOR3_X1   g768(.A1(new_n640), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n830), .A2(new_n832), .A3(new_n955), .ZN(new_n956));
  OAI211_X1 g770(.A(KEYINPUT127), .B(new_n946), .C1(new_n935), .C2(new_n947), .ZN(new_n957));
  AND2_X1   g771(.A1(new_n957), .A2(new_n954), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n946), .B1(new_n935), .B2(new_n947), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT127), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n850), .B1(new_n958), .B2(new_n961), .ZN(new_n962));
  AND3_X1   g776(.A1(new_n952), .A2(new_n956), .A3(new_n962), .ZN(G57));
endmodule


