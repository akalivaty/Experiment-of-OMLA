//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 1 0 1 1 0 0 1 0 0 0 0 0 1 1 0 1 1 1 1 0 0 1 0 0 1 0 1 0 0 1 0 1 1 1 1 1 1 0 1 1 1 1 0 0 1 1 1 0 1 0 1 1 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:00 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n651, new_n652,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n716, new_n717, new_n718, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n726, new_n727, new_n728, new_n730,
    new_n731, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n835, new_n836, new_n838, new_n839, new_n840, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n912, new_n913, new_n914, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n945, new_n946, new_n947, new_n948,
    new_n950, new_n951, new_n952, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n962, new_n963, new_n964, new_n965,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981;
  XNOR2_X1  g000(.A(G155gat), .B(G162gat), .ZN(new_n202));
  NOR2_X1   g001(.A1(new_n202), .A2(KEYINPUT75), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT2), .ZN(new_n204));
  AOI21_X1  g003(.A(new_n204), .B1(G155gat), .B2(G162gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(G141gat), .B(G148gat), .ZN(new_n206));
  NOR3_X1   g005(.A1(new_n203), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n202), .A2(KEYINPUT75), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  OAI211_X1 g008(.A(KEYINPUT75), .B(new_n202), .C1(new_n206), .C2(new_n205), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(G113gat), .B(G120gat), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT70), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT1), .ZN(new_n216));
  XNOR2_X1  g015(.A(G127gat), .B(G134gat), .ZN(new_n217));
  INV_X1    g016(.A(G120gat), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n218), .A2(KEYINPUT70), .A3(G113gat), .ZN(new_n219));
  NAND4_X1  g018(.A1(new_n215), .A2(new_n216), .A3(new_n217), .A4(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(new_n217), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n221), .B1(KEYINPUT1), .B2(new_n213), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n212), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(G225gat), .A2(G233gat), .ZN(new_n225));
  INV_X1    g024(.A(new_n223), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n211), .A2(new_n226), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n224), .A2(new_n225), .A3(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(KEYINPUT39), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT4), .ZN(new_n230));
  XNOR2_X1  g029(.A(new_n223), .B(KEYINPUT71), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n230), .B1(new_n231), .B2(new_n212), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT3), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n211), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n209), .A2(KEYINPUT3), .A3(new_n210), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n234), .A2(new_n223), .A3(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n211), .A2(KEYINPUT4), .A3(new_n226), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n232), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(new_n225), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n229), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  XNOR2_X1  g040(.A(G1gat), .B(G29gat), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n242), .B(KEYINPUT0), .ZN(new_n243));
  XNOR2_X1  g042(.A(G57gat), .B(G85gat), .ZN(new_n244));
  XOR2_X1   g043(.A(new_n243), .B(new_n244), .Z(new_n245));
  INV_X1    g044(.A(KEYINPUT39), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n238), .A2(new_n246), .A3(new_n239), .ZN(new_n247));
  NAND4_X1  g046(.A1(new_n241), .A2(KEYINPUT40), .A3(new_n245), .A4(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT40), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n247), .A2(new_n245), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n249), .B1(new_n250), .B2(new_n240), .ZN(new_n251));
  AND2_X1   g050(.A1(new_n248), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT76), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT71), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n223), .B(new_n254), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n255), .A2(KEYINPUT4), .A3(new_n211), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n227), .A2(new_n230), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n236), .A2(new_n225), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n253), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  AND2_X1   g059(.A1(new_n235), .A2(new_n223), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n239), .B1(new_n261), .B2(new_n234), .ZN(new_n262));
  NAND4_X1  g061(.A1(new_n262), .A2(KEYINPUT76), .A3(new_n256), .A4(new_n257), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n260), .A2(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(KEYINPUT77), .B(KEYINPUT5), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  AND2_X1   g065(.A1(new_n224), .A2(new_n227), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n266), .B1(new_n267), .B2(new_n225), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT78), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n232), .A2(new_n237), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n235), .A2(new_n223), .ZN(new_n272));
  AOI21_X1  g071(.A(KEYINPUT3), .B1(new_n209), .B2(new_n210), .ZN(new_n273));
  OAI211_X1 g072(.A(new_n225), .B(new_n265), .C1(new_n272), .C2(new_n273), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n270), .B1(new_n271), .B2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n274), .ZN(new_n276));
  NAND4_X1  g075(.A1(new_n276), .A2(KEYINPUT78), .A3(new_n232), .A4(new_n237), .ZN(new_n277));
  AOI22_X1  g076(.A1(new_n264), .A2(new_n269), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  OAI21_X1  g077(.A(KEYINPUT83), .B1(new_n278), .B2(new_n245), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT83), .ZN(new_n280));
  INV_X1    g079(.A(new_n245), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n277), .A2(new_n275), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n268), .B1(new_n260), .B2(new_n263), .ZN(new_n284));
  OAI211_X1 g083(.A(new_n280), .B(new_n281), .C1(new_n283), .C2(new_n284), .ZN(new_n285));
  AND3_X1   g084(.A1(new_n252), .A2(new_n279), .A3(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(G8gat), .B(G36gat), .ZN(new_n287));
  XNOR2_X1  g086(.A(G64gat), .B(G92gat), .ZN(new_n288));
  XOR2_X1   g087(.A(new_n287), .B(new_n288), .Z(new_n289));
  XNOR2_X1  g088(.A(G197gat), .B(G204gat), .ZN(new_n290));
  INV_X1    g089(.A(G211gat), .ZN(new_n291));
  INV_X1    g090(.A(G218gat), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n290), .B1(KEYINPUT22), .B2(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(G211gat), .B(G218gat), .ZN(new_n295));
  XNOR2_X1  g094(.A(new_n294), .B(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(G226gat), .ZN(new_n298));
  INV_X1    g097(.A(G233gat), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n300), .A2(KEYINPUT29), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT25), .ZN(new_n303));
  NAND3_X1  g102(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n304), .B1(G183gat), .B2(G190gat), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT64), .ZN(new_n306));
  AOI21_X1  g105(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n307));
  OR3_X1    g106(.A1(new_n305), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  NOR2_X1   g107(.A1(G169gat), .A2(G176gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(G169gat), .A2(G176gat), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n309), .B1(KEYINPUT23), .B2(new_n310), .ZN(new_n311));
  XOR2_X1   g110(.A(KEYINPUT65), .B(G169gat), .Z(new_n312));
  INV_X1    g111(.A(G176gat), .ZN(new_n313));
  AND2_X1   g112(.A1(new_n313), .A2(KEYINPUT23), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n311), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n306), .B1(new_n305), .B2(new_n307), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n308), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(G169gat), .ZN(new_n318));
  AOI211_X1 g117(.A(new_n303), .B(new_n311), .C1(new_n318), .C2(new_n314), .ZN(new_n319));
  XNOR2_X1  g118(.A(new_n307), .B(KEYINPUT66), .ZN(new_n320));
  OR2_X1    g119(.A1(new_n320), .A2(new_n305), .ZN(new_n321));
  AOI22_X1  g120(.A1(new_n303), .A2(new_n317), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  AOI22_X1  g121(.A1(new_n309), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n323));
  OR2_X1    g122(.A1(new_n309), .A2(KEYINPUT26), .ZN(new_n324));
  INV_X1    g123(.A(new_n310), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n323), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(KEYINPUT27), .B(G183gat), .ZN(new_n327));
  INV_X1    g126(.A(G190gat), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n327), .A2(KEYINPUT28), .A3(new_n328), .ZN(new_n329));
  XNOR2_X1  g128(.A(new_n329), .B(KEYINPUT69), .ZN(new_n330));
  NAND2_X1  g129(.A1(KEYINPUT67), .A2(G183gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(KEYINPUT27), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT27), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n333), .A2(KEYINPUT67), .A3(G183gat), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n332), .A2(new_n334), .A3(new_n328), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT68), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT28), .ZN(new_n338));
  NAND4_X1  g137(.A1(new_n332), .A2(new_n334), .A3(KEYINPUT68), .A4(new_n328), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n337), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n326), .B1(new_n330), .B2(new_n340), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n322), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(KEYINPUT73), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT73), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n344), .B1(new_n322), .B2(new_n341), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n302), .B1(new_n343), .B2(new_n345), .ZN(new_n346));
  AND2_X1   g145(.A1(new_n342), .A2(new_n300), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n297), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n343), .A2(new_n300), .A3(new_n345), .ZN(new_n349));
  OR2_X1    g148(.A1(new_n322), .A2(new_n341), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(new_n301), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n349), .A2(new_n296), .A3(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n289), .B1(new_n348), .B2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  NAND4_X1  g153(.A1(new_n348), .A2(new_n352), .A3(KEYINPUT30), .A4(new_n289), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT74), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n348), .A2(new_n352), .A3(new_n289), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT30), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n357), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n356), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n358), .A2(new_n357), .A3(new_n359), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n286), .A2(new_n363), .A3(KEYINPUT84), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT84), .ZN(new_n365));
  INV_X1    g164(.A(new_n362), .ZN(new_n366));
  NOR3_X1   g165(.A1(new_n366), .A2(new_n356), .A3(new_n360), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n252), .A2(new_n279), .A3(new_n285), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n365), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n296), .B1(new_n273), .B2(KEYINPUT29), .ZN(new_n370));
  NAND2_X1  g169(.A1(G228gat), .A2(G233gat), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT81), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n233), .B1(new_n296), .B2(KEYINPUT29), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n212), .A2(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n370), .A2(new_n373), .A3(new_n375), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n371), .A2(new_n372), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n377), .ZN(new_n379));
  NAND4_X1  g178(.A1(new_n370), .A2(new_n375), .A3(new_n379), .A4(new_n373), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n378), .A2(G22gat), .A3(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT82), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  XNOR2_X1  g182(.A(G78gat), .B(G106gat), .ZN(new_n384));
  XNOR2_X1  g183(.A(KEYINPUT31), .B(G50gat), .ZN(new_n385));
  XNOR2_X1  g184(.A(new_n384), .B(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n383), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n378), .A2(new_n380), .ZN(new_n388));
  INV_X1    g187(.A(G22gat), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(new_n381), .ZN(new_n391));
  AND2_X1   g190(.A1(new_n387), .A2(new_n391), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n387), .A2(new_n391), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n358), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT37), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n289), .A2(new_n397), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n353), .A2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  AND2_X1   g199(.A1(new_n349), .A2(new_n351), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n397), .B1(new_n401), .B2(new_n297), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n296), .B1(new_n346), .B2(new_n347), .ZN(new_n403));
  AOI21_X1  g202(.A(KEYINPUT38), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n396), .B1(new_n400), .B2(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(KEYINPUT6), .B1(new_n278), .B2(new_n245), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n279), .A2(new_n406), .A3(new_n285), .ZN(new_n407));
  OAI211_X1 g206(.A(KEYINPUT6), .B(new_n281), .C1(new_n283), .C2(new_n284), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n397), .B1(new_n348), .B2(new_n352), .ZN(new_n409));
  OAI21_X1  g208(.A(KEYINPUT38), .B1(new_n399), .B2(new_n409), .ZN(new_n410));
  NAND4_X1  g209(.A1(new_n405), .A2(new_n407), .A3(new_n408), .A4(new_n410), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n364), .A2(new_n369), .A3(new_n395), .A4(new_n411), .ZN(new_n412));
  XNOR2_X1  g211(.A(G15gat), .B(G43gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(G71gat), .B(G99gat), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n413), .B(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n350), .A2(new_n255), .ZN(new_n416));
  INV_X1    g215(.A(G227gat), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n417), .A2(new_n299), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n342), .A2(new_n231), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n416), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT33), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n415), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n420), .A2(KEYINPUT32), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  OAI211_X1 g223(.A(new_n420), .B(KEYINPUT32), .C1(new_n421), .C2(new_n415), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n416), .A2(new_n419), .ZN(new_n427));
  INV_X1    g226(.A(new_n418), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(KEYINPUT34), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT34), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n427), .A2(new_n431), .A3(new_n428), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n426), .A2(new_n433), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n424), .A2(new_n430), .A3(new_n425), .A4(new_n432), .ZN(new_n435));
  AOI21_X1  g234(.A(KEYINPUT36), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n434), .A2(KEYINPUT72), .A3(new_n435), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT72), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n426), .A2(new_n438), .A3(new_n433), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n436), .B1(new_n440), .B2(KEYINPUT36), .ZN(new_n441));
  OAI21_X1  g240(.A(KEYINPUT80), .B1(new_n278), .B2(new_n245), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT80), .ZN(new_n443));
  OAI211_X1 g242(.A(new_n443), .B(new_n281), .C1(new_n283), .C2(new_n284), .ZN(new_n444));
  OAI211_X1 g243(.A(new_n442), .B(new_n444), .C1(new_n406), .C2(KEYINPUT79), .ZN(new_n445));
  NOR3_X1   g244(.A1(new_n283), .A2(new_n284), .A3(new_n281), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT79), .ZN(new_n447));
  NOR3_X1   g246(.A1(new_n446), .A2(new_n447), .A3(KEYINPUT6), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n408), .B1(new_n445), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(new_n367), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n441), .B1(new_n450), .B2(new_n394), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n394), .B1(new_n439), .B2(new_n437), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n449), .A2(new_n452), .A3(new_n367), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(KEYINPUT35), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n434), .A2(new_n435), .ZN(new_n455));
  NOR3_X1   g254(.A1(new_n394), .A2(new_n455), .A3(KEYINPUT35), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n407), .A2(new_n408), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n456), .A2(new_n367), .A3(new_n457), .ZN(new_n458));
  AOI22_X1  g257(.A1(new_n412), .A2(new_n451), .B1(new_n454), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(G29gat), .A2(G36gat), .ZN(new_n460));
  OAI21_X1  g259(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n461));
  NOR3_X1   g260(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n461), .B1(new_n462), .B2(KEYINPUT87), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT14), .ZN(new_n464));
  INV_X1    g263(.A(G29gat), .ZN(new_n465));
  INV_X1    g264(.A(G36gat), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n464), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT87), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n460), .B1(new_n463), .B2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT86), .ZN(new_n471));
  AND2_X1   g270(.A1(G43gat), .A2(G50gat), .ZN(new_n472));
  NOR2_X1   g271(.A1(G43gat), .A2(G50gat), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n471), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(G43gat), .ZN(new_n475));
  INV_X1    g274(.A(G50gat), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(G43gat), .A2(G50gat), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n477), .A2(KEYINPUT86), .A3(new_n478), .ZN(new_n479));
  AND3_X1   g278(.A1(new_n474), .A2(new_n479), .A3(KEYINPUT15), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n470), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n474), .A2(new_n479), .A3(KEYINPUT15), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n472), .A2(new_n473), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT15), .ZN(new_n484));
  AOI22_X1  g283(.A1(new_n483), .A2(new_n484), .B1(G29gat), .B2(G36gat), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n467), .A2(new_n461), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n482), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n481), .A2(KEYINPUT17), .A3(new_n487), .ZN(new_n488));
  XNOR2_X1  g287(.A(G15gat), .B(G22gat), .ZN(new_n489));
  INV_X1    g288(.A(G1gat), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(KEYINPUT16), .ZN(new_n491));
  AND2_X1   g290(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n489), .A2(G1gat), .ZN(new_n493));
  NOR3_X1   g292(.A1(new_n492), .A2(new_n493), .A3(G8gat), .ZN(new_n494));
  INV_X1    g293(.A(G8gat), .ZN(new_n495));
  XOR2_X1   g294(.A(G15gat), .B(G22gat), .Z(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(new_n490), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n489), .A2(new_n491), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n495), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n494), .A2(new_n499), .ZN(new_n500));
  AND2_X1   g299(.A1(new_n488), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n481), .A2(new_n487), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT17), .ZN(new_n503));
  AOI21_X1  g302(.A(KEYINPUT88), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT88), .ZN(new_n505));
  AOI211_X1 g304(.A(new_n505), .B(KEYINPUT17), .C1(new_n481), .C2(new_n487), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n501), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(G229gat), .A2(G233gat), .ZN(new_n508));
  OAI21_X1  g307(.A(G8gat), .B1(new_n492), .B2(new_n493), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n497), .A2(new_n495), .A3(new_n498), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n502), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n507), .A2(new_n508), .A3(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT18), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(KEYINPUT89), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n507), .A2(KEYINPUT18), .A3(new_n508), .A4(new_n512), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n481), .A2(new_n487), .A3(new_n509), .A4(new_n510), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n512), .A2(new_n518), .ZN(new_n519));
  XOR2_X1   g318(.A(new_n508), .B(KEYINPUT13), .Z(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  AND2_X1   g320(.A1(new_n517), .A2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT89), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n513), .A2(new_n523), .A3(new_n514), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n516), .A2(new_n522), .A3(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(G113gat), .B(G141gat), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n526), .B(G197gat), .ZN(new_n527));
  XOR2_X1   g326(.A(KEYINPUT11), .B(G169gat), .Z(new_n528));
  XNOR2_X1  g327(.A(new_n527), .B(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(KEYINPUT85), .B(KEYINPUT12), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n529), .B(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n525), .A2(new_n532), .ZN(new_n533));
  AND3_X1   g332(.A1(new_n517), .A2(new_n531), .A3(new_n521), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT90), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n515), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n513), .A2(KEYINPUT90), .A3(new_n514), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n534), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n533), .A2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n459), .A2(new_n540), .ZN(new_n541));
  AND2_X1   g340(.A1(G71gat), .A2(G78gat), .ZN(new_n542));
  NOR2_X1   g341(.A1(G71gat), .A2(G78gat), .ZN(new_n543));
  NOR2_X1   g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(G57gat), .B(G64gat), .ZN(new_n545));
  AOI21_X1  g344(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(G57gat), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(G64gat), .ZN(new_n549));
  INV_X1    g348(.A(G64gat), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(G57gat), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  XNOR2_X1  g351(.A(G71gat), .B(G78gat), .ZN(new_n553));
  INV_X1    g352(.A(new_n546), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n547), .A2(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(KEYINPUT91), .B(KEYINPUT21), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(G231gat), .A2(G233gat), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n558), .B(new_n559), .ZN(new_n560));
  XOR2_X1   g359(.A(G127gat), .B(G155gat), .Z(new_n561));
  XNOR2_X1  g360(.A(new_n561), .B(KEYINPUT20), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n560), .B(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(G183gat), .B(G211gat), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n563), .B(new_n564), .ZN(new_n565));
  AND2_X1   g364(.A1(new_n547), .A2(new_n555), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n511), .B1(KEYINPUT21), .B2(new_n566), .ZN(new_n567));
  XOR2_X1   g366(.A(KEYINPUT92), .B(KEYINPUT19), .Z(new_n568));
  XNOR2_X1  g367(.A(new_n567), .B(new_n568), .ZN(new_n569));
  OR2_X1    g368(.A1(new_n565), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n565), .A2(new_n569), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  XOR2_X1   g371(.A(G134gat), .B(G162gat), .Z(new_n573));
  AND2_X1   g372(.A1(G232gat), .A2(G233gat), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n574), .A2(KEYINPUT41), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n573), .B(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(KEYINPUT95), .ZN(new_n577));
  NAND3_X1  g376(.A1(KEYINPUT93), .A2(G85gat), .A3(G92gat), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  OR2_X1    g378(.A1(KEYINPUT94), .A2(KEYINPUT7), .ZN(new_n580));
  NAND2_X1  g379(.A1(KEYINPUT94), .A2(KEYINPUT7), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  AND2_X1   g381(.A1(KEYINPUT94), .A2(KEYINPUT7), .ZN(new_n583));
  NOR2_X1   g382(.A1(KEYINPUT94), .A2(KEYINPUT7), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n578), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(G99gat), .A2(G106gat), .ZN(new_n586));
  INV_X1    g385(.A(G85gat), .ZN(new_n587));
  INV_X1    g386(.A(G92gat), .ZN(new_n588));
  AOI22_X1  g387(.A1(KEYINPUT8), .A2(new_n586), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n582), .A2(new_n585), .A3(new_n589), .ZN(new_n590));
  XOR2_X1   g389(.A(G99gat), .B(G106gat), .Z(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n582), .A2(new_n591), .A3(new_n585), .A4(new_n589), .ZN(new_n594));
  AND2_X1   g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  OAI211_X1 g394(.A(new_n488), .B(new_n595), .C1(new_n504), .C2(new_n506), .ZN(new_n596));
  XOR2_X1   g395(.A(G190gat), .B(G218gat), .Z(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n593), .A2(new_n594), .ZN(new_n599));
  AOI22_X1  g398(.A1(new_n502), .A2(new_n599), .B1(KEYINPUT41), .B2(new_n574), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n596), .A2(new_n598), .A3(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n598), .B1(new_n596), .B2(new_n600), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n577), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n596), .A2(new_n600), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n605), .A2(new_n597), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n576), .B(KEYINPUT95), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n606), .A2(new_n601), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n604), .A2(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(G120gat), .B(G148gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(G176gat), .B(G204gat), .ZN(new_n611));
  XOR2_X1   g410(.A(new_n610), .B(new_n611), .Z(new_n612));
  NAND2_X1  g411(.A1(G230gat), .A2(G233gat), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n590), .A2(KEYINPUT96), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n566), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n615), .A2(new_n599), .ZN(new_n616));
  NAND4_X1  g415(.A1(new_n566), .A2(new_n593), .A3(new_n614), .A4(new_n594), .ZN(new_n617));
  AOI21_X1  g416(.A(KEYINPUT10), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n599), .A2(KEYINPUT10), .A3(new_n566), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n613), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n613), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n616), .A2(new_n622), .A3(new_n617), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT97), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n612), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n612), .ZN(new_n627));
  AOI211_X1 g426(.A(KEYINPUT97), .B(new_n627), .C1(new_n621), .C2(new_n623), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  NOR3_X1   g428(.A1(new_n572), .A2(new_n609), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n541), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n631), .A2(new_n449), .ZN(new_n632));
  XOR2_X1   g431(.A(KEYINPUT98), .B(G1gat), .Z(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(G1324gat));
  NAND3_X1  g433(.A1(new_n541), .A2(new_n363), .A3(new_n630), .ZN(new_n635));
  XOR2_X1   g434(.A(KEYINPUT16), .B(G8gat), .Z(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  OR3_X1    g436(.A1(new_n635), .A2(KEYINPUT42), .A3(new_n637), .ZN(new_n638));
  OAI21_X1  g437(.A(KEYINPUT42), .B1(new_n635), .B2(new_n637), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n635), .A2(G8gat), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n641), .A2(KEYINPUT99), .ZN(new_n642));
  OR2_X1    g441(.A1(new_n641), .A2(KEYINPUT99), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n640), .A2(new_n642), .A3(new_n643), .ZN(G1325gat));
  NAND2_X1  g443(.A1(new_n440), .A2(KEYINPUT36), .ZN(new_n645));
  INV_X1    g444(.A(new_n436), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  OAI21_X1  g446(.A(G15gat), .B1(new_n631), .B2(new_n647), .ZN(new_n648));
  OR2_X1    g447(.A1(new_n455), .A2(G15gat), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n648), .B1(new_n631), .B2(new_n649), .ZN(G1326gat));
  NOR2_X1   g449(.A1(new_n631), .A2(new_n395), .ZN(new_n651));
  XOR2_X1   g450(.A(KEYINPUT43), .B(G22gat), .Z(new_n652));
  XNOR2_X1  g451(.A(new_n651), .B(new_n652), .ZN(G1327gat));
  AND4_X1   g452(.A1(new_n395), .A2(new_n364), .A3(new_n369), .A4(new_n411), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n447), .B1(new_n446), .B2(KEYINPUT6), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n278), .A2(new_n245), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT6), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n656), .A2(KEYINPUT79), .A3(new_n657), .ZN(new_n658));
  NAND4_X1  g457(.A1(new_n655), .A2(new_n658), .A3(new_n442), .A4(new_n444), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n363), .B1(new_n659), .B2(new_n408), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n647), .B1(new_n660), .B2(new_n395), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT35), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n662), .B1(new_n660), .B2(new_n452), .ZN(new_n663));
  INV_X1    g462(.A(new_n458), .ZN(new_n664));
  OAI22_X1  g463(.A1(new_n654), .A2(new_n661), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n572), .ZN(new_n666));
  INV_X1    g465(.A(new_n609), .ZN(new_n667));
  NOR3_X1   g466(.A1(new_n666), .A2(new_n667), .A3(new_n629), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n665), .A2(new_n539), .A3(new_n668), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n449), .A2(G29gat), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  OR3_X1    g470(.A1(new_n669), .A2(KEYINPUT100), .A3(new_n671), .ZN(new_n672));
  OAI21_X1  g471(.A(KEYINPUT100), .B1(new_n669), .B2(new_n671), .ZN(new_n673));
  AND3_X1   g472(.A1(new_n672), .A2(KEYINPUT45), .A3(new_n673), .ZN(new_n674));
  AOI21_X1  g473(.A(KEYINPUT45), .B1(new_n672), .B2(new_n673), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT44), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n677), .B1(new_n459), .B2(new_n667), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n665), .A2(KEYINPUT44), .A3(new_n609), .ZN(new_n679));
  INV_X1    g478(.A(new_n449), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT101), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n572), .B(new_n681), .ZN(new_n682));
  NOR3_X1   g481(.A1(new_n682), .A2(new_n540), .A3(new_n629), .ZN(new_n683));
  NAND4_X1  g482(.A1(new_n678), .A2(new_n679), .A3(new_n680), .A4(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT102), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n465), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n686), .B1(new_n685), .B2(new_n684), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n676), .A2(new_n687), .ZN(G1328gat));
  NOR3_X1   g487(.A1(new_n669), .A2(G36gat), .A3(new_n367), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(KEYINPUT46), .ZN(new_n690));
  NOR3_X1   g489(.A1(new_n459), .A2(new_n677), .A3(new_n667), .ZN(new_n691));
  AOI21_X1  g490(.A(KEYINPUT44), .B1(new_n665), .B2(new_n609), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  AND3_X1   g492(.A1(new_n693), .A2(new_n363), .A3(new_n683), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n690), .B1(new_n466), .B2(new_n694), .ZN(G1329gat));
  NOR2_X1   g494(.A1(new_n647), .A2(new_n475), .ZN(new_n696));
  NAND4_X1  g495(.A1(new_n678), .A2(new_n679), .A3(new_n683), .A4(new_n696), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n475), .B1(new_n669), .B2(new_n455), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g499(.A1(new_n678), .A2(new_n679), .A3(new_n394), .A4(new_n683), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(G50gat), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n669), .A2(KEYINPUT103), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT103), .ZN(new_n704));
  NAND4_X1  g503(.A1(new_n665), .A2(new_n704), .A3(new_n539), .A4(new_n668), .ZN(new_n705));
  NAND4_X1  g504(.A1(new_n703), .A2(new_n476), .A3(new_n394), .A4(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n702), .A2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT48), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT104), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n476), .B1(new_n701), .B2(new_n710), .ZN(new_n711));
  NAND4_X1  g510(.A1(new_n693), .A2(KEYINPUT104), .A3(new_n394), .A4(new_n683), .ZN(new_n712));
  AND2_X1   g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n706), .A2(KEYINPUT48), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n709), .B1(new_n713), .B2(new_n714), .ZN(G1331gat));
  NAND4_X1  g514(.A1(new_n666), .A2(new_n540), .A3(new_n667), .A4(new_n629), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n459), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(new_n680), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g518(.A(new_n367), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n717), .A2(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT105), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n721), .B(new_n722), .ZN(new_n723));
  NOR2_X1   g522(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n723), .B(new_n724), .ZN(G1333gat));
  NAND2_X1  g524(.A1(new_n717), .A2(new_n441), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n455), .A2(G71gat), .ZN(new_n727));
  AOI22_X1  g526(.A1(new_n726), .A2(G71gat), .B1(new_n717), .B2(new_n727), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g528(.A1(new_n717), .A2(new_n394), .ZN(new_n730));
  XOR2_X1   g529(.A(KEYINPUT106), .B(G78gat), .Z(new_n731));
  XNOR2_X1  g530(.A(new_n730), .B(new_n731), .ZN(G1335gat));
  NAND2_X1  g531(.A1(new_n540), .A2(new_n572), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(KEYINPUT107), .ZN(new_n734));
  INV_X1    g533(.A(new_n629), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  AND3_X1   g535(.A1(new_n693), .A2(new_n680), .A3(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(new_n734), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n665), .A2(new_n609), .A3(new_n738), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n735), .B1(new_n739), .B2(KEYINPUT51), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n740), .B1(KEYINPUT51), .B2(new_n739), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n680), .A2(new_n587), .ZN(new_n742));
  OAI22_X1  g541(.A1(new_n737), .A2(new_n587), .B1(new_n741), .B2(new_n742), .ZN(G1336gat));
  NAND4_X1  g542(.A1(new_n678), .A2(new_n679), .A3(new_n363), .A4(new_n736), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(G92gat), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n363), .A2(new_n588), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n745), .B1(new_n741), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(KEYINPUT52), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT52), .ZN(new_n749));
  OAI211_X1 g548(.A(new_n745), .B(new_n749), .C1(new_n741), .C2(new_n746), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n748), .A2(new_n750), .ZN(G1337gat));
  NAND4_X1  g550(.A1(new_n678), .A2(new_n679), .A3(new_n441), .A4(new_n736), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(G99gat), .ZN(new_n753));
  OR2_X1    g552(.A1(new_n455), .A2(G99gat), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n753), .B1(new_n741), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(KEYINPUT108), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT108), .ZN(new_n757));
  OAI211_X1 g556(.A(new_n753), .B(new_n757), .C1(new_n741), .C2(new_n754), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n756), .A2(new_n758), .ZN(G1338gat));
  NAND4_X1  g558(.A1(new_n678), .A2(new_n679), .A3(new_n394), .A4(new_n736), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(G106gat), .ZN(new_n761));
  OR2_X1    g560(.A1(new_n395), .A2(G106gat), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n761), .B1(new_n741), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(KEYINPUT53), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT53), .ZN(new_n765));
  OAI211_X1 g564(.A(new_n761), .B(new_n765), .C1(new_n741), .C2(new_n762), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n764), .A2(new_n766), .ZN(G1339gat));
  NAND2_X1  g566(.A1(new_n630), .A2(new_n540), .ZN(new_n768));
  INV_X1    g567(.A(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT55), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT10), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n615), .A2(new_n599), .ZN(new_n772));
  AOI22_X1  g571(.A1(new_n566), .A2(new_n614), .B1(new_n593), .B2(new_n594), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n771), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n774), .A2(new_n622), .A3(new_n619), .ZN(new_n775));
  AND3_X1   g574(.A1(new_n775), .A2(new_n621), .A3(KEYINPUT54), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT54), .ZN(new_n777));
  OAI211_X1 g576(.A(new_n777), .B(new_n613), .C1(new_n618), .C2(new_n620), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(new_n627), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n770), .B1(new_n776), .B2(new_n779), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n621), .A2(new_n623), .A3(new_n612), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n775), .A2(new_n621), .A3(KEYINPUT54), .ZN(new_n782));
  NAND4_X1  g581(.A1(new_n782), .A2(KEYINPUT55), .A3(new_n627), .A4(new_n778), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n780), .A2(new_n781), .A3(new_n783), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n784), .B1(new_n533), .B2(new_n538), .ZN(new_n785));
  INV_X1    g584(.A(new_n520), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n512), .A2(new_n518), .A3(new_n786), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n787), .B(KEYINPUT110), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n508), .B1(new_n507), .B2(new_n512), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n788), .B1(new_n789), .B2(KEYINPUT109), .ZN(new_n790));
  INV_X1    g589(.A(new_n512), .ZN(new_n791));
  INV_X1    g590(.A(new_n487), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n467), .A2(new_n468), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n462), .A2(KEYINPUT87), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n793), .A2(new_n794), .A3(new_n461), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n482), .B1(new_n460), .B2(new_n795), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n503), .B1(new_n792), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(new_n505), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n502), .A2(KEYINPUT88), .A3(new_n503), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n791), .B1(new_n800), .B2(new_n501), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT109), .ZN(new_n802));
  NOR3_X1   g601(.A1(new_n801), .A2(new_n802), .A3(new_n508), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n529), .B1(new_n790), .B2(new_n803), .ZN(new_n804));
  AND3_X1   g603(.A1(new_n804), .A2(new_n538), .A3(new_n629), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n667), .B1(new_n785), .B2(new_n805), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n609), .A2(new_n781), .A3(new_n783), .A4(new_n780), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n804), .A2(new_n538), .ZN(new_n808));
  OAI21_X1  g607(.A(KEYINPUT111), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  AND3_X1   g608(.A1(new_n513), .A2(KEYINPUT90), .A3(new_n514), .ZN(new_n810));
  AOI21_X1  g609(.A(KEYINPUT90), .B1(new_n513), .B2(new_n514), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n802), .B1(new_n801), .B2(new_n508), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n789), .A2(KEYINPUT109), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n813), .A2(new_n814), .A3(new_n788), .ZN(new_n815));
  AOI22_X1  g614(.A1(new_n812), .A2(new_n534), .B1(new_n815), .B2(new_n529), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT111), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n783), .A2(new_n781), .ZN(new_n818));
  INV_X1    g617(.A(new_n779), .ZN(new_n819));
  AOI21_X1  g618(.A(KEYINPUT55), .B1(new_n819), .B2(new_n782), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n816), .A2(new_n817), .A3(new_n821), .A4(new_n609), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n806), .A2(new_n809), .A3(new_n822), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n682), .B1(new_n823), .B2(KEYINPUT112), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT112), .ZN(new_n825));
  NAND4_X1  g624(.A1(new_n806), .A2(new_n825), .A3(new_n809), .A4(new_n822), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n769), .B1(new_n824), .B2(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(new_n452), .ZN(new_n828));
  NOR4_X1   g627(.A1(new_n827), .A2(new_n449), .A3(new_n363), .A4(new_n828), .ZN(new_n829));
  AOI21_X1  g628(.A(G113gat), .B1(new_n829), .B2(new_n539), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n680), .A2(new_n367), .ZN(new_n831));
  NOR4_X1   g630(.A1(new_n827), .A2(new_n394), .A3(new_n455), .A4(new_n831), .ZN(new_n832));
  AND2_X1   g631(.A1(new_n539), .A2(G113gat), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n830), .B1(new_n832), .B2(new_n833), .ZN(G1340gat));
  AOI21_X1  g633(.A(G120gat), .B1(new_n829), .B2(new_n629), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n735), .A2(new_n218), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n835), .B1(new_n832), .B2(new_n836), .ZN(G1341gat));
  INV_X1    g636(.A(G127gat), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n829), .A2(new_n838), .A3(new_n666), .ZN(new_n839));
  AND2_X1   g638(.A1(new_n832), .A2(new_n682), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n839), .B1(new_n840), .B2(new_n838), .ZN(G1342gat));
  AND2_X1   g640(.A1(new_n832), .A2(new_n609), .ZN(new_n842));
  INV_X1    g641(.A(G134gat), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n829), .A2(new_n843), .A3(new_n609), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n844), .B1(KEYINPUT56), .B2(new_n845), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n846), .B1(KEYINPUT56), .B2(new_n845), .ZN(G1343gat));
  INV_X1    g646(.A(KEYINPUT57), .ZN(new_n848));
  OAI211_X1 g647(.A(KEYINPUT113), .B(new_n848), .C1(new_n827), .C2(new_n395), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT113), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n809), .A2(new_n822), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n523), .B1(new_n513), .B2(new_n514), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n517), .A2(new_n521), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n531), .B1(new_n854), .B2(new_n524), .ZN(new_n855));
  AND3_X1   g654(.A1(new_n534), .A2(new_n536), .A3(new_n537), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n821), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n804), .A2(new_n538), .A3(new_n629), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n609), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  OAI21_X1  g658(.A(KEYINPUT112), .B1(new_n851), .B2(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(new_n682), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n860), .A2(new_n826), .A3(new_n861), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n395), .B1(new_n862), .B2(new_n768), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n850), .B1(new_n863), .B2(KEYINPUT57), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT114), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n865), .B1(new_n776), .B2(new_n779), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n819), .A2(KEYINPUT114), .A3(new_n782), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n866), .A2(new_n867), .A3(new_n770), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n539), .A2(new_n781), .A3(new_n783), .A4(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n609), .B1(new_n869), .B2(new_n858), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n870), .A2(new_n851), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n768), .B1(new_n871), .B2(new_n666), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n872), .A2(KEYINPUT57), .A3(new_n394), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n849), .A2(new_n864), .A3(new_n873), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n831), .A2(new_n441), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n874), .A2(new_n539), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(G141gat), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT115), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n827), .A2(new_n449), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n441), .A2(new_n395), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(new_n367), .ZN(new_n882));
  INV_X1    g681(.A(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  OR3_X1    g683(.A1(new_n884), .A2(G141gat), .A3(new_n540), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n877), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n879), .A2(new_n886), .A3(KEYINPUT58), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT58), .ZN(new_n888));
  OAI211_X1 g687(.A(new_n877), .B(new_n885), .C1(new_n878), .C2(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n887), .A2(new_n889), .ZN(G1344gat));
  OR3_X1    g689(.A1(new_n831), .A2(KEYINPUT117), .A3(new_n441), .ZN(new_n891));
  OAI21_X1  g690(.A(KEYINPUT117), .B1(new_n831), .B2(new_n441), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n891), .A2(new_n629), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n862), .A2(new_n768), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(new_n394), .ZN(new_n895));
  OR3_X1    g694(.A1(new_n895), .A2(KEYINPUT118), .A3(new_n848), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n807), .A2(new_n808), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n572), .B1(new_n870), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(new_n768), .ZN(new_n899));
  AOI21_X1  g698(.A(KEYINPUT57), .B1(new_n899), .B2(new_n394), .ZN(new_n900));
  OAI22_X1  g699(.A1(KEYINPUT118), .A2(new_n900), .B1(new_n895), .B2(new_n848), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n893), .B1(new_n896), .B2(new_n901), .ZN(new_n902));
  INV_X1    g701(.A(G148gat), .ZN(new_n903));
  OAI21_X1  g702(.A(KEYINPUT59), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n874), .A2(new_n629), .A3(new_n875), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n903), .A2(KEYINPUT59), .ZN(new_n906));
  AND3_X1   g705(.A1(new_n905), .A2(KEYINPUT116), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g706(.A(KEYINPUT116), .B1(new_n905), .B2(new_n906), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n904), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND4_X1  g708(.A1(new_n880), .A2(new_n903), .A3(new_n629), .A4(new_n883), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(G1345gat));
  NAND2_X1  g710(.A1(new_n874), .A2(new_n875), .ZN(new_n912));
  OAI21_X1  g711(.A(G155gat), .B1(new_n912), .B2(new_n861), .ZN(new_n913));
  OR2_X1    g712(.A1(new_n572), .A2(G155gat), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n913), .B1(new_n884), .B2(new_n914), .ZN(G1346gat));
  OR3_X1    g714(.A1(new_n884), .A2(G162gat), .A3(new_n667), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT119), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n917), .B1(new_n912), .B2(new_n667), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(G162gat), .ZN(new_n919));
  NOR3_X1   g718(.A1(new_n912), .A2(new_n917), .A3(new_n667), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n916), .B1(new_n919), .B2(new_n920), .ZN(G1347gat));
  NOR2_X1   g720(.A1(new_n394), .A2(new_n455), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n680), .A2(new_n367), .ZN(new_n923));
  NAND4_X1  g722(.A1(new_n894), .A2(new_n539), .A3(new_n922), .A4(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(G169gat), .ZN(new_n925));
  XOR2_X1   g724(.A(new_n925), .B(KEYINPUT122), .Z(new_n926));
  NOR2_X1   g725(.A1(new_n828), .A2(new_n367), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n894), .A2(new_n449), .A3(new_n927), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT120), .ZN(new_n929));
  XNOR2_X1  g728(.A(new_n928), .B(new_n929), .ZN(new_n930));
  AND2_X1   g729(.A1(new_n539), .A2(new_n312), .ZN(new_n931));
  AOI21_X1  g730(.A(KEYINPUT121), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  OR2_X1    g731(.A1(new_n928), .A2(KEYINPUT120), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n928), .A2(KEYINPUT120), .ZN(new_n934));
  AND4_X1   g733(.A1(KEYINPUT121), .A2(new_n933), .A3(new_n934), .A4(new_n931), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n926), .B1(new_n932), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n936), .A2(KEYINPUT123), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT123), .ZN(new_n938));
  OAI211_X1 g737(.A(new_n926), .B(new_n938), .C1(new_n932), .C2(new_n935), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n937), .A2(new_n939), .ZN(G1348gat));
  NAND3_X1  g739(.A1(new_n930), .A2(new_n313), .A3(new_n629), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n894), .A2(new_n922), .A3(new_n923), .ZN(new_n942));
  OAI21_X1  g741(.A(G176gat), .B1(new_n942), .B2(new_n735), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n941), .A2(new_n943), .ZN(G1349gat));
  OAI21_X1  g743(.A(G183gat), .B1(new_n942), .B2(new_n861), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT124), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n666), .A2(new_n327), .ZN(new_n947));
  OAI211_X1 g746(.A(new_n945), .B(new_n946), .C1(new_n928), .C2(new_n947), .ZN(new_n948));
  XNOR2_X1  g747(.A(new_n948), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g748(.A(G190gat), .B1(new_n942), .B2(new_n667), .ZN(new_n950));
  XNOR2_X1  g749(.A(new_n950), .B(KEYINPUT61), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n930), .A2(new_n328), .A3(new_n609), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n951), .A2(new_n952), .ZN(G1351gat));
  AND4_X1   g752(.A1(new_n449), .A2(new_n894), .A3(new_n363), .A4(new_n881), .ZN(new_n954));
  AOI21_X1  g753(.A(G197gat), .B1(new_n954), .B2(new_n539), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n896), .A2(new_n901), .ZN(new_n956));
  NOR3_X1   g755(.A1(new_n680), .A2(new_n441), .A3(new_n367), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  INV_X1    g757(.A(new_n958), .ZN(new_n959));
  AND2_X1   g758(.A1(new_n539), .A2(G197gat), .ZN(new_n960));
  AOI21_X1  g759(.A(new_n955), .B1(new_n959), .B2(new_n960), .ZN(G1352gat));
  OAI21_X1  g760(.A(G204gat), .B1(new_n958), .B2(new_n735), .ZN(new_n962));
  INV_X1    g761(.A(G204gat), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n954), .A2(new_n963), .A3(new_n629), .ZN(new_n964));
  XOR2_X1   g763(.A(new_n964), .B(KEYINPUT62), .Z(new_n965));
  NAND2_X1  g764(.A1(new_n962), .A2(new_n965), .ZN(G1353gat));
  OAI21_X1  g765(.A(G211gat), .B1(new_n958), .B2(new_n572), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n967), .A2(KEYINPUT63), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT63), .ZN(new_n969));
  OAI211_X1 g768(.A(new_n969), .B(G211gat), .C1(new_n958), .C2(new_n572), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n954), .A2(new_n291), .A3(new_n666), .ZN(new_n971));
  XOR2_X1   g770(.A(new_n971), .B(KEYINPUT125), .Z(new_n972));
  NAND3_X1  g771(.A1(new_n968), .A2(new_n970), .A3(new_n972), .ZN(G1354gat));
  NAND2_X1  g772(.A1(new_n954), .A2(new_n609), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n974), .A2(new_n292), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n609), .A2(G218gat), .ZN(new_n976));
  XOR2_X1   g775(.A(new_n976), .B(KEYINPUT126), .Z(new_n977));
  OAI21_X1  g776(.A(new_n975), .B1(new_n958), .B2(new_n977), .ZN(new_n978));
  INV_X1    g777(.A(KEYINPUT127), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  OAI211_X1 g779(.A(KEYINPUT127), .B(new_n975), .C1(new_n958), .C2(new_n977), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n980), .A2(new_n981), .ZN(G1355gat));
endmodule


