//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 0 1 1 1 1 0 0 1 0 1 1 0 0 1 1 0 0 1 0 0 0 1 0 1 1 1 1 1 1 1 1 1 1 1 1 0 1 0 1 0 0 1 0 0 0 1 1 1 0 0 1 1 1 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n773, new_n774, new_n775, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n784, new_n785, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n870, new_n871, new_n872, new_n874, new_n875, new_n876, new_n878,
    new_n879, new_n880, new_n881, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n931, new_n932, new_n933, new_n934, new_n936, new_n937, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n946, new_n947,
    new_n949, new_n950, new_n951, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n987, new_n988;
  XNOR2_X1  g000(.A(KEYINPUT89), .B(G29gat), .ZN(new_n202));
  INV_X1    g001(.A(G36gat), .ZN(new_n203));
  OAI21_X1  g002(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  NOR3_X1   g004(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n206));
  OAI22_X1  g005(.A1(new_n202), .A2(new_n203), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT90), .ZN(new_n209));
  XNOR2_X1  g008(.A(G43gat), .B(G50gat), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT15), .ZN(new_n212));
  AOI21_X1  g011(.A(new_n209), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n210), .A2(KEYINPUT15), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n208), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  OAI211_X1 g014(.A(KEYINPUT15), .B(new_n210), .C1(new_n207), .C2(new_n209), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  XNOR2_X1  g016(.A(KEYINPUT91), .B(KEYINPUT17), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n215), .A2(new_n216), .A3(KEYINPUT17), .ZN(new_n220));
  INV_X1    g019(.A(G22gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(G15gat), .ZN(new_n222));
  INV_X1    g021(.A(G15gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(G22gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(G1gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(KEYINPUT16), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n228), .A2(new_n222), .A3(new_n224), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(G8gat), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT92), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n229), .A2(new_n232), .ZN(new_n233));
  NAND4_X1  g032(.A1(new_n228), .A2(new_n222), .A3(new_n224), .A4(KEYINPUT92), .ZN(new_n234));
  XOR2_X1   g033(.A(KEYINPUT93), .B(G8gat), .Z(new_n235));
  NAND4_X1  g034(.A1(new_n233), .A2(new_n227), .A3(new_n234), .A4(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n231), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(KEYINPUT94), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT94), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n231), .A2(new_n236), .A3(new_n239), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n219), .A2(new_n220), .A3(new_n238), .A4(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(G229gat), .A2(G233gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n217), .A2(new_n237), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n241), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT18), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n217), .B(new_n237), .ZN(new_n247));
  XOR2_X1   g046(.A(new_n242), .B(KEYINPUT13), .Z(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n241), .A2(KEYINPUT18), .A3(new_n242), .A4(new_n243), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n246), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  XNOR2_X1  g050(.A(G113gat), .B(G141gat), .ZN(new_n252));
  XNOR2_X1  g051(.A(new_n252), .B(G197gat), .ZN(new_n253));
  XOR2_X1   g052(.A(KEYINPUT11), .B(G169gat), .Z(new_n254));
  XNOR2_X1  g053(.A(new_n253), .B(new_n254), .ZN(new_n255));
  XOR2_X1   g054(.A(new_n255), .B(KEYINPUT12), .Z(new_n256));
  NAND2_X1  g055(.A1(new_n251), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(new_n256), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n246), .A2(new_n258), .A3(new_n249), .A4(new_n250), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  XNOR2_X1  g060(.A(G78gat), .B(G106gat), .ZN(new_n262));
  XNOR2_X1  g061(.A(KEYINPUT31), .B(G50gat), .ZN(new_n263));
  XOR2_X1   g062(.A(new_n262), .B(new_n263), .Z(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(G228gat), .ZN(new_n266));
  INV_X1    g065(.A(G233gat), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT29), .ZN(new_n269));
  XNOR2_X1  g068(.A(G155gat), .B(G162gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(KEYINPUT79), .ZN(new_n271));
  NAND2_X1  g070(.A1(G155gat), .A2(G162gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(KEYINPUT2), .ZN(new_n273));
  INV_X1    g072(.A(G141gat), .ZN(new_n274));
  INV_X1    g073(.A(G148gat), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(G141gat), .A2(G148gat), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n273), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT79), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n272), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n271), .A2(new_n278), .A3(new_n280), .ZN(new_n281));
  XOR2_X1   g080(.A(G141gat), .B(G148gat), .Z(new_n282));
  NAND2_X1  g081(.A1(new_n273), .A2(KEYINPUT80), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT80), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n272), .A2(new_n284), .A3(KEYINPUT2), .ZN(new_n285));
  NAND4_X1  g084(.A1(new_n282), .A2(new_n283), .A3(new_n270), .A4(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n281), .A2(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(KEYINPUT81), .B(KEYINPUT3), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n269), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  XOR2_X1   g089(.A(G211gat), .B(G218gat), .Z(new_n291));
  AOI21_X1  g090(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n292));
  AND2_X1   g091(.A1(G197gat), .A2(G204gat), .ZN(new_n293));
  NOR2_X1   g092(.A1(G197gat), .A2(G204gat), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n291), .B1(new_n292), .B2(new_n295), .ZN(new_n296));
  XNOR2_X1  g095(.A(G211gat), .B(G218gat), .ZN(new_n297));
  XNOR2_X1  g096(.A(G197gat), .B(G204gat), .ZN(new_n298));
  INV_X1    g097(.A(new_n292), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n297), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n296), .A2(KEYINPUT76), .A3(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT76), .ZN(new_n302));
  OAI211_X1 g101(.A(new_n291), .B(new_n302), .C1(new_n292), .C2(new_n295), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n290), .A2(new_n304), .ZN(new_n305));
  AOI21_X1  g104(.A(KEYINPUT29), .B1(new_n296), .B2(new_n300), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n287), .B1(new_n306), .B2(new_n289), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n268), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n301), .A2(new_n269), .A3(new_n303), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT3), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(new_n287), .ZN(new_n313));
  INV_X1    g112(.A(new_n268), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n314), .B1(new_n290), .B2(new_n304), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT83), .ZN(new_n316));
  AND3_X1   g115(.A1(new_n313), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n316), .B1(new_n313), .B2(new_n315), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n309), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n265), .B1(new_n319), .B2(new_n221), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n305), .A2(new_n268), .ZN(new_n321));
  AND2_X1   g120(.A1(new_n281), .A2(new_n286), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n322), .B1(new_n310), .B2(new_n311), .ZN(new_n323));
  OAI21_X1  g122(.A(KEYINPUT83), .B1(new_n321), .B2(new_n323), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n313), .A2(new_n315), .A3(new_n316), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n308), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(G22gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n320), .A2(new_n327), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n221), .A2(KEYINPUT84), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n265), .B1(new_n326), .B2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT85), .ZN(new_n332));
  AOI211_X1 g131(.A(new_n308), .B(new_n329), .C1(new_n324), .C2(new_n325), .ZN(new_n333));
  NOR3_X1   g132(.A1(new_n331), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n264), .B1(new_n319), .B2(new_n329), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n326), .A2(new_n330), .ZN(new_n336));
  AOI21_X1  g135(.A(KEYINPUT85), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n328), .B1(new_n334), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(G169gat), .A2(G176gat), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(G169gat), .ZN(new_n341));
  INV_X1    g140(.A(G176gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n340), .B1(KEYINPUT26), .B2(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n341), .A2(new_n342), .A3(KEYINPUT65), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT65), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n346), .B1(G169gat), .B2(G176gat), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT26), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n345), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n344), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(G183gat), .A2(G190gat), .ZN(new_n351));
  AND2_X1   g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT27), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n353), .A2(G183gat), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  AOI21_X1  g154(.A(G190gat), .B1(new_n353), .B2(G183gat), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n355), .A2(KEYINPUT28), .A3(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(G183gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(KEYINPUT66), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT66), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(G183gat), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n359), .A2(new_n361), .A3(KEYINPUT27), .ZN(new_n362));
  AOI21_X1  g161(.A(KEYINPUT28), .B1(new_n362), .B2(new_n356), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT68), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n357), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  AOI211_X1 g164(.A(KEYINPUT68), .B(KEYINPUT28), .C1(new_n362), .C2(new_n356), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n352), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT25), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n339), .A2(KEYINPUT23), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n368), .B1(new_n369), .B2(new_n343), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n345), .A2(new_n347), .A3(KEYINPUT23), .ZN(new_n371));
  AND2_X1   g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(G190gat), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n359), .A2(new_n361), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n351), .A2(KEYINPUT24), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT24), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n376), .A2(G183gat), .A3(G190gat), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  AND3_X1   g177(.A1(new_n374), .A2(new_n378), .A3(KEYINPUT67), .ZN(new_n379));
  AOI21_X1  g178(.A(KEYINPUT67), .B1(new_n374), .B2(new_n378), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n372), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  AND2_X1   g180(.A1(KEYINPUT64), .A2(G176gat), .ZN(new_n382));
  NOR2_X1   g181(.A1(KEYINPUT64), .A2(G176gat), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  AND2_X1   g183(.A1(new_n341), .A2(KEYINPUT23), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n369), .A2(new_n343), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n358), .A2(new_n373), .ZN(new_n389));
  AND2_X1   g188(.A1(new_n378), .A2(new_n389), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n368), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n381), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(G226gat), .A2(G233gat), .ZN(new_n393));
  AND3_X1   g192(.A1(new_n367), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  AOI21_X1  g193(.A(KEYINPUT29), .B1(G226gat), .B2(G233gat), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n395), .B1(new_n367), .B2(new_n392), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n304), .B1(new_n394), .B2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT77), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n367), .A2(new_n392), .A3(new_n393), .ZN(new_n399));
  INV_X1    g198(.A(new_n304), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n353), .A2(G183gat), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(new_n373), .ZN(new_n402));
  XNOR2_X1  g201(.A(KEYINPUT66), .B(G183gat), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n402), .B1(new_n403), .B2(KEYINPUT27), .ZN(new_n404));
  OAI21_X1  g203(.A(KEYINPUT68), .B1(new_n404), .B2(KEYINPUT28), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n363), .A2(new_n364), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n405), .A2(new_n406), .A3(new_n357), .ZN(new_n407));
  AOI22_X1  g206(.A1(new_n407), .A2(new_n352), .B1(new_n381), .B2(new_n391), .ZN(new_n408));
  OAI211_X1 g207(.A(new_n399), .B(new_n400), .C1(new_n408), .C2(new_n395), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n397), .A2(new_n398), .A3(new_n409), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n394), .A2(new_n396), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n411), .A2(KEYINPUT77), .A3(new_n400), .ZN(new_n412));
  XNOR2_X1  g211(.A(G8gat), .B(G36gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(G64gat), .B(G92gat), .ZN(new_n414));
  XOR2_X1   g213(.A(new_n413), .B(new_n414), .Z(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n410), .A2(new_n412), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n410), .A2(new_n412), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(new_n415), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT30), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n417), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(KEYINPUT78), .B1(new_n418), .B2(new_n415), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT78), .ZN(new_n423));
  AOI211_X1 g222(.A(new_n423), .B(new_n416), .C1(new_n410), .C2(new_n412), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n421), .B1(new_n425), .B2(new_n420), .ZN(new_n426));
  XOR2_X1   g225(.A(G1gat), .B(G29gat), .Z(new_n427));
  XNOR2_X1  g226(.A(KEYINPUT82), .B(KEYINPUT0), .ZN(new_n428));
  XNOR2_X1  g227(.A(new_n427), .B(new_n428), .ZN(new_n429));
  XNOR2_X1  g228(.A(G57gat), .B(G85gat), .ZN(new_n430));
  XNOR2_X1  g229(.A(new_n429), .B(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT5), .ZN(new_n432));
  XOR2_X1   g231(.A(G113gat), .B(G120gat), .Z(new_n433));
  INV_X1    g232(.A(KEYINPUT1), .ZN(new_n434));
  XNOR2_X1  g233(.A(G127gat), .B(G134gat), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  XNOR2_X1  g235(.A(KEYINPUT69), .B(G134gat), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(G127gat), .ZN(new_n438));
  OR2_X1    g237(.A1(KEYINPUT70), .A2(G127gat), .ZN(new_n439));
  NAND2_X1  g238(.A1(KEYINPUT70), .A2(G127gat), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n439), .A2(G134gat), .A3(new_n440), .ZN(new_n441));
  AND2_X1   g240(.A1(new_n438), .A2(new_n441), .ZN(new_n442));
  AND2_X1   g241(.A1(new_n433), .A2(new_n434), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n436), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(new_n287), .ZN(new_n445));
  AOI22_X1  g244(.A1(new_n438), .A2(new_n441), .B1(new_n433), .B2(new_n434), .ZN(new_n446));
  INV_X1    g245(.A(new_n436), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(new_n322), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n445), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(G225gat), .A2(G233gat), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n432), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT4), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n449), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n287), .A2(KEYINPUT3), .ZN(new_n456));
  OAI211_X1 g255(.A(new_n456), .B(new_n444), .C1(new_n287), .C2(new_n289), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n448), .A2(new_n322), .A3(KEYINPUT4), .ZN(new_n458));
  AND3_X1   g257(.A1(new_n455), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n453), .B1(new_n459), .B2(new_n451), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n455), .A2(new_n457), .A3(new_n451), .A4(new_n458), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n461), .A2(new_n432), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n431), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT6), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n459), .A2(KEYINPUT5), .A3(new_n451), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n450), .A2(new_n452), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(KEYINPUT5), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(new_n461), .ZN(new_n468));
  INV_X1    g267(.A(new_n431), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n465), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n463), .A2(new_n464), .A3(new_n470), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n465), .A2(new_n468), .A3(KEYINPUT6), .A4(new_n469), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n338), .B1(new_n426), .B2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n350), .A2(new_n351), .ZN(new_n476));
  INV_X1    g275(.A(new_n357), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n362), .A2(new_n356), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT28), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n477), .B1(new_n480), .B2(KEYINPUT68), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n476), .B1(new_n481), .B2(new_n406), .ZN(new_n482));
  AOI22_X1  g281(.A1(new_n384), .A2(new_n385), .B1(new_n343), .B2(new_n369), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n378), .A2(new_n389), .ZN(new_n484));
  AOI21_X1  g283(.A(KEYINPUT25), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n374), .A2(new_n378), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT67), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n374), .A2(new_n378), .A3(KEYINPUT67), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n485), .B1(new_n490), .B2(new_n372), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n448), .B1(new_n482), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(G227gat), .A2(G233gat), .ZN(new_n493));
  INV_X1    g292(.A(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n367), .A2(new_n392), .A3(new_n444), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n492), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT33), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n496), .A2(KEYINPUT32), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT72), .ZN(new_n500));
  XNOR2_X1  g299(.A(G15gat), .B(G43gat), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT71), .ZN(new_n502));
  XNOR2_X1  g301(.A(new_n501), .B(new_n502), .ZN(new_n503));
  XNOR2_X1  g302(.A(G71gat), .B(G99gat), .ZN(new_n504));
  XNOR2_X1  g303(.A(new_n503), .B(new_n504), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n498), .A2(new_n499), .A3(new_n500), .A4(new_n505), .ZN(new_n506));
  AND3_X1   g305(.A1(new_n498), .A2(new_n499), .A3(new_n505), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT73), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n497), .B1(new_n505), .B2(new_n508), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n509), .B1(new_n508), .B2(new_n505), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n496), .A2(new_n510), .A3(KEYINPUT32), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(KEYINPUT72), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n506), .B1(new_n507), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n492), .A2(new_n495), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT34), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n514), .A2(new_n515), .A3(new_n493), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(KEYINPUT74), .ZN(new_n517));
  INV_X1    g316(.A(new_n514), .ZN(new_n518));
  OAI21_X1  g317(.A(KEYINPUT34), .B1(new_n518), .B2(new_n494), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT74), .ZN(new_n520));
  NAND4_X1  g319(.A1(new_n514), .A2(new_n520), .A3(new_n515), .A4(new_n493), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n517), .A2(new_n519), .A3(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n513), .A2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT75), .ZN(new_n525));
  OAI211_X1 g324(.A(new_n522), .B(new_n506), .C1(new_n507), .C2(new_n512), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n524), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT36), .ZN(new_n528));
  INV_X1    g327(.A(new_n513), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n529), .A2(KEYINPUT75), .A3(new_n522), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n527), .A2(new_n528), .A3(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n524), .A2(KEYINPUT36), .A3(new_n526), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT86), .ZN(new_n534));
  NOR3_X1   g333(.A1(new_n422), .A2(new_n424), .A3(KEYINPUT30), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n534), .B1(new_n535), .B2(new_n421), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n419), .A2(new_n423), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n418), .A2(KEYINPUT78), .A3(new_n415), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n537), .A2(new_n420), .A3(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(new_n421), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n539), .A2(new_n540), .A3(KEYINPUT86), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT40), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n450), .A2(new_n452), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n543), .B(KEYINPUT87), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n455), .A2(new_n457), .A3(new_n458), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(new_n452), .ZN(new_n546));
  AND3_X1   g345(.A1(new_n544), .A2(KEYINPUT39), .A3(new_n546), .ZN(new_n547));
  OR2_X1    g346(.A1(new_n546), .A2(KEYINPUT39), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(new_n431), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n542), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n544), .A2(KEYINPUT39), .A3(new_n546), .ZN(new_n551));
  NAND4_X1  g350(.A1(new_n551), .A2(KEYINPUT40), .A3(new_n431), .A4(new_n548), .ZN(new_n552));
  AND3_X1   g351(.A1(new_n550), .A2(new_n470), .A3(new_n552), .ZN(new_n553));
  AND3_X1   g352(.A1(new_n536), .A2(new_n541), .A3(new_n553), .ZN(new_n554));
  AND2_X1   g353(.A1(new_n471), .A2(new_n472), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT88), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n416), .A2(KEYINPUT37), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n417), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n397), .A2(new_n409), .ZN(new_n559));
  AOI21_X1  g358(.A(KEYINPUT38), .B1(new_n559), .B2(KEYINPUT37), .ZN(new_n560));
  AND2_X1   g359(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  OAI211_X1 g360(.A(new_n555), .B(new_n425), .C1(new_n556), .C2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT37), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n558), .B1(new_n563), .B2(new_n418), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n564), .A2(KEYINPUT38), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n558), .A2(new_n556), .A3(new_n560), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n338), .B1(new_n562), .B2(new_n567), .ZN(new_n568));
  OAI211_X1 g367(.A(new_n475), .B(new_n533), .C1(new_n554), .C2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n536), .A2(new_n541), .ZN(new_n570));
  AOI21_X1  g369(.A(KEYINPUT35), .B1(new_n471), .B2(new_n472), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n338), .A2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n527), .A2(new_n530), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n570), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  AND2_X1   g374(.A1(new_n524), .A2(new_n526), .ZN(new_n576));
  NAND4_X1  g375(.A1(new_n576), .A2(new_n473), .A3(new_n426), .A4(new_n338), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n577), .A2(KEYINPUT35), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n575), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n261), .B1(new_n569), .B2(new_n579), .ZN(new_n580));
  XOR2_X1   g379(.A(G57gat), .B(G64gat), .Z(new_n581));
  AND2_X1   g380(.A1(G71gat), .A2(G78gat), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n581), .B1(KEYINPUT9), .B2(new_n582), .ZN(new_n583));
  XOR2_X1   g382(.A(G71gat), .B(G78gat), .Z(new_n584));
  XNOR2_X1  g383(.A(new_n583), .B(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT21), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(G231gat), .A2(G233gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n587), .B(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(G127gat), .ZN(new_n590));
  OR2_X1    g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n589), .A2(new_n590), .ZN(new_n592));
  XNOR2_X1  g391(.A(G183gat), .B(G211gat), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  AND3_X1   g393(.A1(new_n591), .A2(new_n592), .A3(new_n594), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n594), .B1(new_n591), .B2(new_n592), .ZN(new_n596));
  OAI211_X1 g395(.A(new_n231), .B(new_n236), .C1(new_n585), .C2(new_n586), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n597), .B(KEYINPUT96), .ZN(new_n598));
  XNOR2_X1  g397(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(KEYINPUT95), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n600), .B(G155gat), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  AND2_X1   g401(.A1(new_n598), .A2(new_n601), .ZN(new_n603));
  OAI22_X1  g402(.A1(new_n595), .A2(new_n596), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n591), .A2(new_n592), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n605), .A2(new_n593), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n603), .A2(new_n602), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n591), .A2(new_n592), .A3(new_n594), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n604), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(G99gat), .A2(G106gat), .ZN(new_n611));
  INV_X1    g410(.A(G85gat), .ZN(new_n612));
  INV_X1    g411(.A(G92gat), .ZN(new_n613));
  AOI22_X1  g412(.A1(KEYINPUT8), .A2(new_n611), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND4_X1  g413(.A1(KEYINPUT98), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n615));
  NAND3_X1  g414(.A1(KEYINPUT98), .A2(G85gat), .A3(G92gat), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT7), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n614), .A2(new_n615), .A3(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT99), .ZN(new_n620));
  XNOR2_X1  g419(.A(G99gat), .B(G106gat), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n619), .A2(new_n620), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n619), .A2(new_n622), .ZN(new_n624));
  NAND4_X1  g423(.A1(new_n614), .A2(new_n621), .A3(new_n615), .A4(new_n618), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n624), .A2(KEYINPUT99), .A3(new_n625), .ZN(new_n626));
  NAND4_X1  g425(.A1(new_n219), .A2(new_n220), .A3(new_n623), .A4(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n623), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n628), .A2(new_n217), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT41), .ZN(new_n630));
  NAND2_X1  g429(.A1(G232gat), .A2(G233gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n631), .B(KEYINPUT97), .ZN(new_n632));
  OAI211_X1 g431(.A(new_n627), .B(new_n629), .C1(new_n630), .C2(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(G190gat), .B(G218gat), .ZN(new_n634));
  OR2_X1    g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n633), .A2(new_n634), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  AOI21_X1  g436(.A(KEYINPUT100), .B1(new_n633), .B2(new_n634), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n632), .A2(new_n630), .ZN(new_n639));
  XOR2_X1   g438(.A(new_n639), .B(G134gat), .Z(new_n640));
  INV_X1    g439(.A(G162gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n640), .B(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n637), .B1(new_n638), .B2(new_n643), .ZN(new_n644));
  NAND4_X1  g443(.A1(new_n635), .A2(KEYINPUT100), .A3(new_n636), .A4(new_n642), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n610), .A2(new_n646), .ZN(new_n647));
  XOR2_X1   g446(.A(G120gat), .B(G148gat), .Z(new_n648));
  XNOR2_X1  g447(.A(new_n648), .B(KEYINPUT103), .ZN(new_n649));
  XNOR2_X1  g448(.A(G176gat), .B(G204gat), .ZN(new_n650));
  XOR2_X1   g449(.A(new_n649), .B(new_n650), .Z(new_n651));
  NAND2_X1  g450(.A1(G230gat), .A2(G233gat), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  XOR2_X1   g452(.A(new_n583), .B(new_n584), .Z(new_n654));
  INV_X1    g453(.A(KEYINPUT101), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n621), .B1(new_n619), .B2(new_n655), .ZN(new_n656));
  NAND4_X1  g455(.A1(new_n614), .A2(KEYINPUT101), .A3(new_n615), .A4(new_n618), .ZN(new_n657));
  AND3_X1   g456(.A1(new_n656), .A2(KEYINPUT102), .A3(new_n657), .ZN(new_n658));
  AOI22_X1  g457(.A1(new_n656), .A2(new_n657), .B1(KEYINPUT102), .B2(new_n625), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n654), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n628), .A2(new_n585), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT10), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n654), .A2(KEYINPUT10), .A3(new_n628), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n653), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n662), .A2(new_n652), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n651), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  AOI21_X1  g467(.A(KEYINPUT10), .B1(new_n660), .B2(new_n661), .ZN(new_n669));
  INV_X1    g468(.A(new_n665), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n652), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n651), .ZN(new_n672));
  OAI211_X1 g471(.A(new_n671), .B(new_n672), .C1(new_n662), .C2(new_n652), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n668), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n647), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n580), .A2(new_n675), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n676), .A2(new_n473), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(new_n226), .ZN(G1324gat));
  OAI21_X1  g477(.A(G8gat), .B1(new_n676), .B2(new_n570), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT42), .ZN(new_n680));
  INV_X1    g479(.A(new_n676), .ZN(new_n681));
  INV_X1    g480(.A(new_n570), .ZN(new_n682));
  XOR2_X1   g481(.A(KEYINPUT16), .B(G8gat), .Z(new_n683));
  NAND3_X1  g482(.A1(new_n681), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  AND3_X1   g483(.A1(new_n684), .A2(KEYINPUT104), .A3(new_n680), .ZN(new_n685));
  AOI21_X1  g484(.A(KEYINPUT104), .B1(new_n684), .B2(new_n680), .ZN(new_n686));
  OAI221_X1 g485(.A(new_n679), .B1(new_n680), .B2(new_n684), .C1(new_n685), .C2(new_n686), .ZN(G1325gat));
  NAND2_X1  g486(.A1(new_n533), .A2(KEYINPUT105), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT105), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n531), .A2(new_n689), .A3(new_n532), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  OAI21_X1  g490(.A(G15gat), .B1(new_n676), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n574), .A2(new_n223), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n692), .B1(new_n676), .B2(new_n693), .ZN(G1326gat));
  NOR2_X1   g493(.A1(new_n676), .A2(new_n338), .ZN(new_n695));
  XOR2_X1   g494(.A(KEYINPUT43), .B(G22gat), .Z(new_n696));
  XNOR2_X1  g495(.A(new_n695), .B(new_n696), .ZN(G1327gat));
  INV_X1    g496(.A(new_n610), .ZN(new_n698));
  INV_X1    g497(.A(new_n646), .ZN(new_n699));
  INV_X1    g498(.A(new_n674), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n698), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(KEYINPUT106), .ZN(new_n702));
  NAND4_X1  g501(.A1(new_n580), .A2(new_n555), .A3(new_n202), .A4(new_n702), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(KEYINPUT45), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT44), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n569), .A2(new_n579), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n705), .B1(new_n706), .B2(new_n699), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n705), .A2(KEYINPUT107), .ZN(new_n708));
  OR2_X1    g507(.A1(new_n705), .A2(KEYINPUT107), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n646), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(new_n337), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n335), .A2(KEYINPUT85), .A3(new_n336), .ZN(new_n713));
  AOI22_X1  g512(.A1(new_n712), .A2(new_n713), .B1(new_n327), .B2(new_n320), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n537), .A2(new_n538), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n556), .B1(new_n558), .B2(new_n560), .ZN(new_n716));
  NOR3_X1   g515(.A1(new_n715), .A2(new_n716), .A3(new_n473), .ZN(new_n717));
  AOI22_X1  g516(.A1(new_n556), .A2(new_n561), .B1(new_n564), .B2(KEYINPUT38), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n714), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n536), .A2(new_n541), .A3(new_n553), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n474), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(new_n690), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n689), .B1(new_n531), .B2(new_n532), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n721), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n711), .B1(new_n724), .B2(new_n579), .ZN(new_n725));
  OR2_X1    g524(.A1(new_n707), .A2(new_n725), .ZN(new_n726));
  NOR3_X1   g525(.A1(new_n610), .A2(new_n261), .A3(new_n674), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n726), .A2(new_n555), .A3(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(new_n728), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n704), .B1(new_n729), .B2(new_n202), .ZN(G1328gat));
  NAND3_X1  g529(.A1(new_n726), .A2(new_n682), .A3(new_n727), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(G36gat), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n580), .A2(new_n702), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n682), .A2(new_n203), .ZN(new_n734));
  OR3_X1    g533(.A1(new_n733), .A2(KEYINPUT108), .A3(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT46), .ZN(new_n736));
  OAI21_X1  g535(.A(KEYINPUT108), .B1(new_n733), .B2(new_n734), .ZN(new_n737));
  AND3_X1   g536(.A1(new_n735), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n736), .B1(new_n735), .B2(new_n737), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n732), .B1(new_n738), .B2(new_n739), .ZN(G1329gat));
  INV_X1    g539(.A(new_n691), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n726), .A2(G43gat), .A3(new_n741), .A4(new_n727), .ZN(new_n742));
  INV_X1    g541(.A(G43gat), .ZN(new_n743));
  INV_X1    g542(.A(new_n574), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n743), .B1(new_n733), .B2(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n742), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(KEYINPUT47), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT47), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n742), .A2(new_n748), .A3(new_n745), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n747), .A2(new_n749), .ZN(G1330gat));
  NAND4_X1  g549(.A1(new_n726), .A2(G50gat), .A3(new_n714), .A4(new_n727), .ZN(new_n751));
  INV_X1    g550(.A(G50gat), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n752), .B1(new_n733), .B2(new_n338), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(KEYINPUT48), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT48), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n751), .A2(new_n756), .A3(new_n753), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n755), .A2(new_n757), .ZN(G1331gat));
  INV_X1    g557(.A(KEYINPUT109), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n572), .B1(new_n530), .B2(new_n527), .ZN(new_n760));
  AOI22_X1  g559(.A1(new_n760), .A2(new_n570), .B1(KEYINPUT35), .B2(new_n577), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n761), .B1(new_n691), .B2(new_n721), .ZN(new_n762));
  NOR3_X1   g561(.A1(new_n647), .A2(new_n260), .A3(new_n700), .ZN(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n759), .B1(new_n762), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n724), .A2(new_n579), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n766), .A2(KEYINPUT109), .A3(new_n763), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n765), .A2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(new_n555), .ZN(new_n770));
  XNOR2_X1  g569(.A(KEYINPUT110), .B(G57gat), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n770), .B(new_n771), .ZN(G1332gat));
  XNOR2_X1  g571(.A(KEYINPUT49), .B(G64gat), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n769), .A2(new_n682), .A3(new_n773), .ZN(new_n774));
  OAI22_X1  g573(.A1(new_n768), .A2(new_n570), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(G1333gat));
  OAI21_X1  g575(.A(G71gat), .B1(new_n768), .B2(new_n691), .ZN(new_n777));
  OR2_X1    g576(.A1(new_n744), .A2(G71gat), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n777), .B1(new_n768), .B2(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT50), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  OAI211_X1 g580(.A(new_n777), .B(KEYINPUT50), .C1(new_n768), .C2(new_n778), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(G1334gat));
  NOR2_X1   g582(.A1(new_n768), .A2(new_n338), .ZN(new_n784));
  XNOR2_X1  g583(.A(KEYINPUT111), .B(G78gat), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n784), .B(new_n785), .ZN(G1335gat));
  INV_X1    g585(.A(KEYINPUT51), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n610), .A2(new_n260), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT112), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n788), .B(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(new_n699), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n787), .B1(new_n762), .B2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(new_n791), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n766), .A2(KEYINPUT51), .A3(new_n793), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n700), .B1(new_n792), .B2(new_n794), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n795), .A2(new_n612), .A3(new_n555), .ZN(new_n796));
  INV_X1    g595(.A(new_n790), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n797), .A2(new_n700), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n726), .A2(new_n555), .A3(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(new_n799), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n796), .B1(new_n800), .B2(new_n612), .ZN(G1336gat));
  NAND3_X1  g600(.A1(new_n795), .A2(new_n613), .A3(new_n682), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT113), .ZN(new_n803));
  OAI211_X1 g602(.A(new_n682), .B(new_n798), .C1(new_n707), .C2(new_n725), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(G92gat), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n802), .A2(new_n803), .A3(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(KEYINPUT52), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT52), .ZN(new_n808));
  NAND4_X1  g607(.A1(new_n802), .A2(new_n803), .A3(new_n808), .A4(new_n805), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n807), .A2(new_n809), .ZN(G1337gat));
  NOR2_X1   g609(.A1(new_n744), .A2(G99gat), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n811), .ZN(new_n812));
  OAI211_X1 g611(.A(new_n741), .B(new_n798), .C1(new_n707), .C2(new_n725), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(G99gat), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  XNOR2_X1  g614(.A(new_n815), .B(KEYINPUT114), .ZN(G1338gat));
  INV_X1    g615(.A(KEYINPUT116), .ZN(new_n817));
  OAI211_X1 g616(.A(new_n714), .B(new_n798), .C1(new_n707), .C2(new_n725), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(G106gat), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n338), .A2(G106gat), .ZN(new_n820));
  AOI21_X1  g619(.A(KEYINPUT51), .B1(new_n766), .B2(new_n793), .ZN(new_n821));
  AOI211_X1 g620(.A(new_n787), .B(new_n791), .C1(new_n724), .C2(new_n579), .ZN(new_n822));
  OAI211_X1 g621(.A(new_n674), .B(new_n820), .C1(new_n821), .C2(new_n822), .ZN(new_n823));
  XOR2_X1   g622(.A(KEYINPUT115), .B(KEYINPUT53), .Z(new_n824));
  AND4_X1   g623(.A1(new_n817), .A2(new_n819), .A3(new_n823), .A4(new_n824), .ZN(new_n825));
  AOI22_X1  g624(.A1(new_n795), .A2(new_n820), .B1(new_n818), .B2(G106gat), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n817), .B1(new_n826), .B2(new_n824), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n819), .A2(new_n823), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(KEYINPUT53), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n825), .B1(new_n827), .B2(new_n829), .ZN(G1339gat));
  AOI21_X1  g629(.A(new_n242), .B1(new_n241), .B2(new_n243), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n247), .A2(new_n248), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n255), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  AND2_X1   g632(.A1(new_n259), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(new_n674), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(KEYINPUT118), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT55), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n665), .A2(new_n653), .ZN(new_n838));
  OAI21_X1  g637(.A(KEYINPUT54), .B1(new_n669), .B2(new_n838), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n666), .A2(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT54), .ZN(new_n841));
  OAI211_X1 g640(.A(new_n841), .B(new_n652), .C1(new_n669), .C2(new_n670), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(new_n651), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n837), .B1(new_n840), .B2(new_n843), .ZN(new_n844));
  OAI211_X1 g643(.A(new_n671), .B(KEYINPUT54), .C1(new_n669), .C2(new_n838), .ZN(new_n845));
  NAND4_X1  g644(.A1(new_n845), .A2(KEYINPUT55), .A3(new_n651), .A4(new_n842), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n260), .A2(new_n844), .A3(new_n846), .A4(new_n673), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n836), .A2(new_n847), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n835), .A2(KEYINPUT118), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n646), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  AND4_X1   g649(.A1(new_n645), .A2(new_n644), .A3(new_n673), .A4(new_n846), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT117), .ZN(new_n852));
  XNOR2_X1  g651(.A(new_n834), .B(new_n852), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n851), .A2(new_n853), .A3(new_n844), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n610), .B1(new_n850), .B2(new_n854), .ZN(new_n855));
  NOR3_X1   g654(.A1(new_n647), .A2(new_n260), .A3(new_n674), .ZN(new_n856));
  OR2_X1    g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n744), .A2(new_n714), .ZN(new_n858));
  AND2_X1   g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n859), .A2(new_n555), .A3(new_n570), .ZN(new_n860));
  INV_X1    g659(.A(G113gat), .ZN(new_n861));
  NOR3_X1   g660(.A1(new_n860), .A2(new_n861), .A3(new_n261), .ZN(new_n862));
  AND2_X1   g661(.A1(new_n857), .A2(new_n555), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n576), .A2(new_n338), .ZN(new_n864));
  INV_X1    g663(.A(new_n864), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n863), .A2(new_n570), .A3(new_n865), .ZN(new_n866));
  INV_X1    g665(.A(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(new_n260), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n862), .B1(new_n868), .B2(new_n861), .ZN(G1340gat));
  INV_X1    g668(.A(G120gat), .ZN(new_n870));
  NOR3_X1   g669(.A1(new_n860), .A2(new_n870), .A3(new_n700), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n867), .A2(new_n674), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n871), .B1(new_n872), .B2(new_n870), .ZN(G1341gat));
  NAND2_X1  g672(.A1(new_n439), .A2(new_n440), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n874), .B1(new_n860), .B2(new_n698), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n610), .A2(new_n439), .A3(new_n440), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n875), .B1(new_n866), .B2(new_n876), .ZN(G1342gat));
  NAND3_X1  g676(.A1(new_n867), .A2(new_n437), .A3(new_n699), .ZN(new_n878));
  OR2_X1    g677(.A1(new_n878), .A2(KEYINPUT56), .ZN(new_n879));
  OAI21_X1  g678(.A(G134gat), .B1(new_n860), .B2(new_n646), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n878), .A2(KEYINPUT56), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(G1343gat));
  INV_X1    g681(.A(KEYINPUT57), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n857), .A2(new_n883), .A3(new_n714), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n847), .A2(KEYINPUT119), .A3(new_n835), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(new_n646), .ZN(new_n886));
  AOI21_X1  g685(.A(KEYINPUT119), .B1(new_n847), .B2(new_n835), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n854), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n856), .B1(new_n888), .B2(new_n698), .ZN(new_n889));
  OAI21_X1  g688(.A(KEYINPUT57), .B1(new_n889), .B2(new_n338), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n691), .A2(new_n555), .A3(new_n570), .ZN(new_n891));
  INV_X1    g690(.A(new_n891), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n884), .A2(new_n890), .A3(new_n892), .ZN(new_n893));
  OAI21_X1  g692(.A(G141gat), .B1(new_n893), .B2(new_n261), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT120), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n863), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n857), .A2(new_n555), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(KEYINPUT120), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n691), .A2(new_n570), .A3(new_n714), .ZN(new_n899));
  INV_X1    g698(.A(new_n899), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n896), .A2(new_n898), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n260), .A2(new_n274), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n894), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  XNOR2_X1  g702(.A(new_n903), .B(KEYINPUT58), .ZN(G1344gat));
  INV_X1    g703(.A(KEYINPUT59), .ZN(new_n905));
  OAI211_X1 g704(.A(new_n905), .B(G148gat), .C1(new_n893), .C2(new_n700), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT122), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT121), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n847), .A2(new_n835), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT119), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n911), .A2(new_n646), .A3(new_n885), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n610), .B1(new_n912), .B2(new_n854), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n908), .B1(new_n913), .B2(new_n856), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n888), .A2(new_n698), .ZN(new_n915));
  INV_X1    g714(.A(new_n856), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n915), .A2(KEYINPUT121), .A3(new_n916), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n338), .A2(KEYINPUT57), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n914), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n891), .A2(new_n700), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n714), .B1(new_n855), .B2(new_n856), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(KEYINPUT57), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n919), .A2(new_n920), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n923), .A2(G148gat), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n907), .B1(new_n924), .B2(KEYINPUT59), .ZN(new_n925));
  AOI211_X1 g724(.A(KEYINPUT122), .B(new_n905), .C1(new_n923), .C2(G148gat), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n906), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  INV_X1    g726(.A(new_n901), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n928), .A2(new_n275), .A3(new_n674), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n927), .A2(new_n929), .ZN(G1345gat));
  AOI21_X1  g729(.A(G155gat), .B1(new_n928), .B2(new_n610), .ZN(new_n931));
  INV_X1    g730(.A(new_n893), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n610), .A2(G155gat), .ZN(new_n933));
  XOR2_X1   g732(.A(new_n933), .B(KEYINPUT123), .Z(new_n934));
  AOI21_X1  g733(.A(new_n931), .B1(new_n932), .B2(new_n934), .ZN(G1346gat));
  OAI21_X1  g734(.A(G162gat), .B1(new_n893), .B2(new_n646), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n699), .A2(new_n641), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n936), .B1(new_n901), .B2(new_n937), .ZN(G1347gat));
  NOR2_X1   g737(.A1(new_n570), .A2(new_n555), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n859), .A2(new_n939), .ZN(new_n940));
  OAI21_X1  g739(.A(G169gat), .B1(new_n940), .B2(new_n261), .ZN(new_n941));
  AND3_X1   g740(.A1(new_n857), .A2(new_n865), .A3(new_n939), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n942), .A2(new_n341), .A3(new_n260), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  XNOR2_X1  g743(.A(new_n944), .B(KEYINPUT124), .ZN(G1348gat));
  NOR3_X1   g744(.A1(new_n940), .A2(new_n384), .A3(new_n700), .ZN(new_n946));
  AOI21_X1  g745(.A(G176gat), .B1(new_n942), .B2(new_n674), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n946), .A2(new_n947), .ZN(G1349gat));
  NAND4_X1  g747(.A1(new_n942), .A2(new_n401), .A3(new_n355), .A4(new_n610), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n940), .A2(new_n698), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n949), .B1(new_n950), .B2(new_n403), .ZN(new_n951));
  XNOR2_X1  g750(.A(new_n951), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g751(.A1(new_n942), .A2(new_n373), .A3(new_n699), .ZN(new_n953));
  NAND4_X1  g752(.A1(new_n857), .A2(new_n699), .A3(new_n858), .A4(new_n939), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n954), .A2(G190gat), .ZN(new_n955));
  OR2_X1    g754(.A1(new_n955), .A2(KEYINPUT125), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT61), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n955), .A2(KEYINPUT125), .ZN(new_n958));
  AND3_X1   g757(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n957), .B1(new_n956), .B2(new_n958), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n953), .B1(new_n959), .B2(new_n960), .ZN(G1351gat));
  NAND2_X1  g760(.A1(new_n691), .A2(new_n939), .ZN(new_n962));
  NOR2_X1   g761(.A1(new_n962), .A2(new_n921), .ZN(new_n963));
  AOI21_X1  g762(.A(G197gat), .B1(new_n963), .B2(new_n260), .ZN(new_n964));
  XOR2_X1   g763(.A(new_n962), .B(KEYINPUT126), .Z(new_n965));
  OAI21_X1  g764(.A(new_n918), .B1(new_n889), .B2(KEYINPUT121), .ZN(new_n966));
  NOR3_X1   g765(.A1(new_n913), .A2(new_n908), .A3(new_n856), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n922), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NOR2_X1   g767(.A1(new_n965), .A2(new_n968), .ZN(new_n969));
  AND2_X1   g768(.A1(new_n260), .A2(G197gat), .ZN(new_n970));
  AOI21_X1  g769(.A(new_n964), .B1(new_n969), .B2(new_n970), .ZN(G1352gat));
  NOR4_X1   g770(.A1(new_n962), .A2(new_n921), .A3(G204gat), .A4(new_n700), .ZN(new_n972));
  INV_X1    g771(.A(KEYINPUT62), .ZN(new_n973));
  OR2_X1    g772(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n972), .A2(new_n973), .ZN(new_n975));
  NOR3_X1   g774(.A1(new_n965), .A2(new_n700), .A3(new_n968), .ZN(new_n976));
  INV_X1    g775(.A(G204gat), .ZN(new_n977));
  OAI211_X1 g776(.A(new_n974), .B(new_n975), .C1(new_n976), .C2(new_n977), .ZN(G1353gat));
  NAND3_X1  g777(.A1(new_n691), .A2(new_n610), .A3(new_n939), .ZN(new_n979));
  OAI21_X1  g778(.A(G211gat), .B1(new_n968), .B2(new_n979), .ZN(new_n980));
  INV_X1    g779(.A(KEYINPUT63), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  OAI211_X1 g781(.A(KEYINPUT63), .B(G211gat), .C1(new_n968), .C2(new_n979), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n982), .A2(KEYINPUT127), .A3(new_n983), .ZN(new_n984));
  OR3_X1    g783(.A1(new_n979), .A2(new_n921), .A3(G211gat), .ZN(new_n985));
  OAI211_X1 g784(.A(new_n984), .B(new_n985), .C1(KEYINPUT127), .C2(new_n982), .ZN(G1354gat));
  AOI21_X1  g785(.A(G218gat), .B1(new_n963), .B2(new_n699), .ZN(new_n987));
  AND2_X1   g786(.A1(new_n699), .A2(G218gat), .ZN(new_n988));
  AOI21_X1  g787(.A(new_n987), .B1(new_n969), .B2(new_n988), .ZN(G1355gat));
endmodule


