

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U552 ( .A1(G2105), .A2(G2104), .ZN(n524) );
  NOR2_X2 U553 ( .A1(n998), .A2(n703), .ZN(n710) );
  XNOR2_X1 U554 ( .A(n689), .B(n688), .ZN(n691) );
  NOR2_X1 U555 ( .A1(n769), .A2(n768), .ZN(n516) );
  OR2_X1 U556 ( .A1(KEYINPUT33), .A2(n754), .ZN(n517) );
  OR2_X1 U557 ( .A1(G171), .A2(n724), .ZN(n518) );
  AND2_X1 U558 ( .A1(n697), .A2(G1996), .ZN(n699) );
  XNOR2_X1 U559 ( .A(KEYINPUT99), .B(KEYINPUT30), .ZN(n688) );
  INV_X1 U560 ( .A(G168), .ZN(n690) );
  AND2_X1 U561 ( .A1(n694), .A2(n518), .ZN(n696) );
  INV_X1 U562 ( .A(KEYINPUT101), .ZN(n728) );
  NOR2_X1 U563 ( .A1(n742), .A2(n741), .ZN(n745) );
  INV_X1 U564 ( .A(n1013), .ZN(n756) );
  NOR2_X1 U565 ( .A1(n757), .A2(n756), .ZN(n758) );
  INV_X1 U566 ( .A(KEYINPUT89), .ZN(n561) );
  XNOR2_X1 U567 ( .A(n562), .B(n561), .ZN(n563) );
  NOR2_X1 U568 ( .A1(G651), .A2(n652), .ZN(n646) );
  NOR2_X1 U569 ( .A1(n531), .A2(n530), .ZN(G160) );
  INV_X1 U570 ( .A(G2105), .ZN(n523) );
  INV_X1 U571 ( .A(G2104), .ZN(n519) );
  NOR2_X1 U572 ( .A1(n523), .A2(n519), .ZN(n879) );
  NAND2_X1 U573 ( .A1(n879), .A2(G113), .ZN(n522) );
  NOR2_X2 U574 ( .A1(G2105), .A2(n519), .ZN(n875) );
  NAND2_X1 U575 ( .A1(G101), .A2(n875), .ZN(n520) );
  XOR2_X1 U576 ( .A(KEYINPUT23), .B(n520), .Z(n521) );
  NAND2_X1 U577 ( .A1(n522), .A2(n521), .ZN(n531) );
  NOR2_X1 U578 ( .A1(G2104), .A2(n523), .ZN(n880) );
  NAND2_X1 U579 ( .A1(n880), .A2(G125), .ZN(n529) );
  XNOR2_X1 U580 ( .A(n524), .B(KEYINPUT66), .ZN(n526) );
  XNOR2_X1 U581 ( .A(KEYINPUT67), .B(KEYINPUT17), .ZN(n525) );
  XNOR2_X1 U582 ( .A(n526), .B(n525), .ZN(n560) );
  INV_X1 U583 ( .A(n560), .ZN(n527) );
  INV_X1 U584 ( .A(n527), .ZN(n876) );
  NAND2_X1 U585 ( .A1(G137), .A2(n876), .ZN(n528) );
  NAND2_X1 U586 ( .A1(n529), .A2(n528), .ZN(n530) );
  INV_X1 U587 ( .A(G651), .ZN(n536) );
  NOR2_X1 U588 ( .A1(G543), .A2(n536), .ZN(n532) );
  XOR2_X1 U589 ( .A(KEYINPUT1), .B(n532), .Z(n651) );
  NAND2_X1 U590 ( .A1(G63), .A2(n651), .ZN(n534) );
  XOR2_X1 U591 ( .A(KEYINPUT0), .B(G543), .Z(n652) );
  NAND2_X1 U592 ( .A1(G51), .A2(n646), .ZN(n533) );
  NAND2_X1 U593 ( .A1(n534), .A2(n533), .ZN(n535) );
  XOR2_X1 U594 ( .A(KEYINPUT6), .B(n535), .Z(n544) );
  NOR2_X1 U595 ( .A1(n652), .A2(n536), .ZN(n639) );
  NAND2_X1 U596 ( .A1(G76), .A2(n639), .ZN(n540) );
  XOR2_X1 U597 ( .A(KEYINPUT4), .B(KEYINPUT73), .Z(n538) );
  NOR2_X1 U598 ( .A1(G651), .A2(G543), .ZN(n636) );
  NAND2_X1 U599 ( .A1(G89), .A2(n636), .ZN(n537) );
  XNOR2_X1 U600 ( .A(n538), .B(n537), .ZN(n539) );
  NAND2_X1 U601 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U602 ( .A(n541), .B(KEYINPUT5), .ZN(n542) );
  XNOR2_X1 U603 ( .A(KEYINPUT74), .B(n542), .ZN(n543) );
  NAND2_X1 U604 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U605 ( .A(KEYINPUT7), .B(n545), .ZN(G168) );
  NAND2_X1 U606 ( .A1(G85), .A2(n636), .ZN(n547) );
  NAND2_X1 U607 ( .A1(G72), .A2(n639), .ZN(n546) );
  NAND2_X1 U608 ( .A1(n547), .A2(n546), .ZN(n551) );
  NAND2_X1 U609 ( .A1(G60), .A2(n651), .ZN(n549) );
  NAND2_X1 U610 ( .A1(G47), .A2(n646), .ZN(n548) );
  NAND2_X1 U611 ( .A1(n549), .A2(n548), .ZN(n550) );
  OR2_X1 U612 ( .A1(n551), .A2(n550), .ZN(G290) );
  NAND2_X1 U613 ( .A1(G64), .A2(n651), .ZN(n553) );
  NAND2_X1 U614 ( .A1(G52), .A2(n646), .ZN(n552) );
  NAND2_X1 U615 ( .A1(n553), .A2(n552), .ZN(n559) );
  NAND2_X1 U616 ( .A1(n639), .A2(G77), .ZN(n554) );
  XNOR2_X1 U617 ( .A(n554), .B(KEYINPUT68), .ZN(n556) );
  NAND2_X1 U618 ( .A1(G90), .A2(n636), .ZN(n555) );
  NAND2_X1 U619 ( .A1(n556), .A2(n555), .ZN(n557) );
  XOR2_X1 U620 ( .A(KEYINPUT9), .B(n557), .Z(n558) );
  NOR2_X1 U621 ( .A1(n559), .A2(n558), .ZN(G171) );
  INV_X1 U622 ( .A(G57), .ZN(G237) );
  INV_X1 U623 ( .A(G82), .ZN(G220) );
  NAND2_X1 U624 ( .A1(n879), .A2(G114), .ZN(n564) );
  NAND2_X1 U625 ( .A1(n560), .A2(G138), .ZN(n562) );
  NAND2_X1 U626 ( .A1(n564), .A2(n563), .ZN(n568) );
  NAND2_X1 U627 ( .A1(G102), .A2(n875), .ZN(n566) );
  NAND2_X1 U628 ( .A1(G126), .A2(n880), .ZN(n565) );
  NAND2_X1 U629 ( .A1(n566), .A2(n565), .ZN(n567) );
  NOR2_X1 U630 ( .A1(n568), .A2(n567), .ZN(n683) );
  BUF_X1 U631 ( .A(n683), .Z(G164) );
  NAND2_X1 U632 ( .A1(G94), .A2(G452), .ZN(n569) );
  XNOR2_X1 U633 ( .A(n569), .B(KEYINPUT69), .ZN(G173) );
  NAND2_X1 U634 ( .A1(G7), .A2(G661), .ZN(n570) );
  XNOR2_X1 U635 ( .A(n570), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U636 ( .A(G223), .ZN(n825) );
  NAND2_X1 U637 ( .A1(n825), .A2(G567), .ZN(n571) );
  XOR2_X1 U638 ( .A(KEYINPUT11), .B(n571), .Z(G234) );
  NAND2_X1 U639 ( .A1(G56), .A2(n651), .ZN(n572) );
  XOR2_X1 U640 ( .A(KEYINPUT14), .B(n572), .Z(n579) );
  NAND2_X1 U641 ( .A1(G81), .A2(n636), .ZN(n573) );
  XNOR2_X1 U642 ( .A(n573), .B(KEYINPUT72), .ZN(n574) );
  XNOR2_X1 U643 ( .A(n574), .B(KEYINPUT12), .ZN(n576) );
  NAND2_X1 U644 ( .A1(G68), .A2(n639), .ZN(n575) );
  NAND2_X1 U645 ( .A1(n576), .A2(n575), .ZN(n577) );
  XOR2_X1 U646 ( .A(KEYINPUT13), .B(n577), .Z(n578) );
  NOR2_X1 U647 ( .A1(n579), .A2(n578), .ZN(n581) );
  NAND2_X1 U648 ( .A1(n646), .A2(G43), .ZN(n580) );
  NAND2_X1 U649 ( .A1(n581), .A2(n580), .ZN(n998) );
  INV_X1 U650 ( .A(G860), .ZN(n620) );
  OR2_X1 U651 ( .A1(n998), .A2(n620), .ZN(G153) );
  INV_X1 U652 ( .A(G171), .ZN(G301) );
  NAND2_X1 U653 ( .A1(G868), .A2(G301), .ZN(n590) );
  NAND2_X1 U654 ( .A1(G66), .A2(n651), .ZN(n583) );
  NAND2_X1 U655 ( .A1(G92), .A2(n636), .ZN(n582) );
  NAND2_X1 U656 ( .A1(n583), .A2(n582), .ZN(n587) );
  NAND2_X1 U657 ( .A1(G79), .A2(n639), .ZN(n585) );
  NAND2_X1 U658 ( .A1(G54), .A2(n646), .ZN(n584) );
  NAND2_X1 U659 ( .A1(n585), .A2(n584), .ZN(n586) );
  NOR2_X1 U660 ( .A1(n587), .A2(n586), .ZN(n588) );
  XOR2_X1 U661 ( .A(KEYINPUT15), .B(n588), .Z(n1001) );
  OR2_X1 U662 ( .A1(n1001), .A2(G868), .ZN(n589) );
  NAND2_X1 U663 ( .A1(n590), .A2(n589), .ZN(G284) );
  XOR2_X1 U664 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U665 ( .A1(G65), .A2(n651), .ZN(n592) );
  NAND2_X1 U666 ( .A1(G91), .A2(n636), .ZN(n591) );
  NAND2_X1 U667 ( .A1(n592), .A2(n591), .ZN(n596) );
  NAND2_X1 U668 ( .A1(G78), .A2(n639), .ZN(n594) );
  NAND2_X1 U669 ( .A1(G53), .A2(n646), .ZN(n593) );
  NAND2_X1 U670 ( .A1(n594), .A2(n593), .ZN(n595) );
  NOR2_X1 U671 ( .A1(n596), .A2(n595), .ZN(n597) );
  XOR2_X1 U672 ( .A(KEYINPUT70), .B(n597), .Z(G299) );
  INV_X1 U673 ( .A(G868), .ZN(n665) );
  NOR2_X1 U674 ( .A1(G286), .A2(n665), .ZN(n598) );
  XOR2_X1 U675 ( .A(KEYINPUT75), .B(n598), .Z(n600) );
  NOR2_X1 U676 ( .A1(G299), .A2(G868), .ZN(n599) );
  NOR2_X1 U677 ( .A1(n600), .A2(n599), .ZN(G297) );
  NAND2_X1 U678 ( .A1(n620), .A2(G559), .ZN(n601) );
  NAND2_X1 U679 ( .A1(n601), .A2(n1001), .ZN(n602) );
  XNOR2_X1 U680 ( .A(n602), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U681 ( .A1(G868), .A2(n998), .ZN(n603) );
  XNOR2_X1 U682 ( .A(KEYINPUT76), .B(n603), .ZN(n606) );
  NAND2_X1 U683 ( .A1(G868), .A2(n1001), .ZN(n604) );
  NOR2_X1 U684 ( .A1(G559), .A2(n604), .ZN(n605) );
  NOR2_X1 U685 ( .A1(n606), .A2(n605), .ZN(n607) );
  XOR2_X1 U686 ( .A(KEYINPUT77), .B(n607), .Z(G282) );
  NAND2_X1 U687 ( .A1(n879), .A2(G111), .ZN(n608) );
  XNOR2_X1 U688 ( .A(n608), .B(KEYINPUT78), .ZN(n610) );
  NAND2_X1 U689 ( .A1(G99), .A2(n875), .ZN(n609) );
  NAND2_X1 U690 ( .A1(n610), .A2(n609), .ZN(n611) );
  XNOR2_X1 U691 ( .A(n611), .B(KEYINPUT79), .ZN(n613) );
  NAND2_X1 U692 ( .A1(G135), .A2(n876), .ZN(n612) );
  NAND2_X1 U693 ( .A1(n613), .A2(n612), .ZN(n616) );
  NAND2_X1 U694 ( .A1(n880), .A2(G123), .ZN(n614) );
  XOR2_X1 U695 ( .A(KEYINPUT18), .B(n614), .Z(n615) );
  NOR2_X1 U696 ( .A1(n616), .A2(n615), .ZN(n927) );
  XNOR2_X1 U697 ( .A(n927), .B(G2096), .ZN(n618) );
  INV_X1 U698 ( .A(G2100), .ZN(n617) );
  NAND2_X1 U699 ( .A1(n618), .A2(n617), .ZN(G156) );
  NAND2_X1 U700 ( .A1(G559), .A2(n1001), .ZN(n619) );
  XOR2_X1 U701 ( .A(n998), .B(n619), .Z(n662) );
  NAND2_X1 U702 ( .A1(n620), .A2(n662), .ZN(n627) );
  NAND2_X1 U703 ( .A1(G67), .A2(n651), .ZN(n622) );
  NAND2_X1 U704 ( .A1(G93), .A2(n636), .ZN(n621) );
  NAND2_X1 U705 ( .A1(n622), .A2(n621), .ZN(n626) );
  NAND2_X1 U706 ( .A1(G80), .A2(n639), .ZN(n624) );
  NAND2_X1 U707 ( .A1(G55), .A2(n646), .ZN(n623) );
  NAND2_X1 U708 ( .A1(n624), .A2(n623), .ZN(n625) );
  NOR2_X1 U709 ( .A1(n626), .A2(n625), .ZN(n664) );
  XOR2_X1 U710 ( .A(n627), .B(n664), .Z(G145) );
  NAND2_X1 U711 ( .A1(G88), .A2(n636), .ZN(n628) );
  XOR2_X1 U712 ( .A(KEYINPUT84), .B(n628), .Z(n633) );
  NAND2_X1 U713 ( .A1(G62), .A2(n651), .ZN(n630) );
  NAND2_X1 U714 ( .A1(G50), .A2(n646), .ZN(n629) );
  NAND2_X1 U715 ( .A1(n630), .A2(n629), .ZN(n631) );
  XOR2_X1 U716 ( .A(KEYINPUT83), .B(n631), .Z(n632) );
  NOR2_X1 U717 ( .A1(n633), .A2(n632), .ZN(n635) );
  NAND2_X1 U718 ( .A1(n639), .A2(G75), .ZN(n634) );
  NAND2_X1 U719 ( .A1(n635), .A2(n634), .ZN(G303) );
  INV_X1 U720 ( .A(G303), .ZN(G166) );
  NAND2_X1 U721 ( .A1(G61), .A2(n651), .ZN(n638) );
  NAND2_X1 U722 ( .A1(G86), .A2(n636), .ZN(n637) );
  NAND2_X1 U723 ( .A1(n638), .A2(n637), .ZN(n642) );
  NAND2_X1 U724 ( .A1(n639), .A2(G73), .ZN(n640) );
  XOR2_X1 U725 ( .A(KEYINPUT2), .B(n640), .Z(n641) );
  NOR2_X1 U726 ( .A1(n642), .A2(n641), .ZN(n643) );
  XNOR2_X1 U727 ( .A(n643), .B(KEYINPUT82), .ZN(n645) );
  NAND2_X1 U728 ( .A1(G48), .A2(n646), .ZN(n644) );
  NAND2_X1 U729 ( .A1(n645), .A2(n644), .ZN(G305) );
  NAND2_X1 U730 ( .A1(n646), .A2(G49), .ZN(n647) );
  XNOR2_X1 U731 ( .A(n647), .B(KEYINPUT80), .ZN(n649) );
  NAND2_X1 U732 ( .A1(G74), .A2(G651), .ZN(n648) );
  NAND2_X1 U733 ( .A1(n649), .A2(n648), .ZN(n650) );
  NOR2_X1 U734 ( .A1(n651), .A2(n650), .ZN(n655) );
  NAND2_X1 U735 ( .A1(G87), .A2(n652), .ZN(n653) );
  XOR2_X1 U736 ( .A(KEYINPUT81), .B(n653), .Z(n654) );
  NAND2_X1 U737 ( .A1(n655), .A2(n654), .ZN(G288) );
  XNOR2_X1 U738 ( .A(KEYINPUT85), .B(KEYINPUT19), .ZN(n657) );
  XNOR2_X1 U739 ( .A(G290), .B(G299), .ZN(n656) );
  XNOR2_X1 U740 ( .A(n657), .B(n656), .ZN(n659) );
  XNOR2_X1 U741 ( .A(G166), .B(G305), .ZN(n658) );
  XNOR2_X1 U742 ( .A(n659), .B(n658), .ZN(n661) );
  XNOR2_X1 U743 ( .A(G288), .B(n664), .ZN(n660) );
  XNOR2_X1 U744 ( .A(n661), .B(n660), .ZN(n897) );
  XOR2_X1 U745 ( .A(n897), .B(n662), .Z(n663) );
  NOR2_X1 U746 ( .A1(n665), .A2(n663), .ZN(n667) );
  AND2_X1 U747 ( .A1(n665), .A2(n664), .ZN(n666) );
  NOR2_X1 U748 ( .A1(n667), .A2(n666), .ZN(G295) );
  NAND2_X1 U749 ( .A1(G2078), .A2(G2084), .ZN(n668) );
  XOR2_X1 U750 ( .A(KEYINPUT20), .B(n668), .Z(n669) );
  NAND2_X1 U751 ( .A1(n669), .A2(G2090), .ZN(n670) );
  XNOR2_X1 U752 ( .A(n670), .B(KEYINPUT21), .ZN(n671) );
  XNOR2_X1 U753 ( .A(KEYINPUT86), .B(n671), .ZN(n672) );
  NAND2_X1 U754 ( .A1(G2072), .A2(n672), .ZN(G158) );
  XOR2_X1 U755 ( .A(KEYINPUT87), .B(G44), .Z(n673) );
  XNOR2_X1 U756 ( .A(KEYINPUT3), .B(n673), .ZN(G218) );
  XNOR2_X1 U757 ( .A(KEYINPUT71), .B(G132), .ZN(G219) );
  NOR2_X1 U758 ( .A1(G220), .A2(G219), .ZN(n674) );
  XOR2_X1 U759 ( .A(KEYINPUT22), .B(n674), .Z(n675) );
  XNOR2_X1 U760 ( .A(n675), .B(KEYINPUT88), .ZN(n676) );
  NOR2_X1 U761 ( .A1(G218), .A2(n676), .ZN(n677) );
  NAND2_X1 U762 ( .A1(G96), .A2(n677), .ZN(n831) );
  NAND2_X1 U763 ( .A1(n831), .A2(G2106), .ZN(n681) );
  NAND2_X1 U764 ( .A1(G120), .A2(G69), .ZN(n678) );
  NOR2_X1 U765 ( .A1(G237), .A2(n678), .ZN(n679) );
  NAND2_X1 U766 ( .A1(G108), .A2(n679), .ZN(n832) );
  NAND2_X1 U767 ( .A1(n832), .A2(G567), .ZN(n680) );
  NAND2_X1 U768 ( .A1(n681), .A2(n680), .ZN(n833) );
  NAND2_X1 U769 ( .A1(G483), .A2(G661), .ZN(n682) );
  NOR2_X1 U770 ( .A1(n833), .A2(n682), .ZN(n830) );
  NAND2_X1 U771 ( .A1(n830), .A2(G36), .ZN(G176) );
  NAND2_X1 U772 ( .A1(G160), .A2(G40), .ZN(n774) );
  NOR2_X1 U773 ( .A1(G1384), .A2(n683), .ZN(n684) );
  XNOR2_X1 U774 ( .A(n684), .B(KEYINPUT64), .ZN(n773) );
  INV_X1 U775 ( .A(n773), .ZN(n685) );
  NOR2_X2 U776 ( .A1(n774), .A2(n685), .ZN(n697) );
  INV_X1 U777 ( .A(n697), .ZN(n700) );
  NAND2_X1 U778 ( .A1(G8), .A2(n700), .ZN(n769) );
  NOR2_X1 U779 ( .A1(G1966), .A2(n769), .ZN(n742) );
  NOR2_X1 U780 ( .A1(G2084), .A2(n700), .ZN(n743) );
  NOR2_X1 U781 ( .A1(n742), .A2(n743), .ZN(n686) );
  XNOR2_X1 U782 ( .A(n686), .B(KEYINPUT98), .ZN(n687) );
  NAND2_X1 U783 ( .A1(n687), .A2(G8), .ZN(n689) );
  NAND2_X1 U784 ( .A1(n691), .A2(n690), .ZN(n694) );
  XNOR2_X1 U785 ( .A(KEYINPUT25), .B(G2078), .ZN(n977) );
  NOR2_X1 U786 ( .A1(n700), .A2(n977), .ZN(n693) );
  AND2_X1 U787 ( .A1(n700), .A2(G1961), .ZN(n692) );
  NOR2_X1 U788 ( .A1(n693), .A2(n692), .ZN(n724) );
  INV_X1 U789 ( .A(KEYINPUT31), .ZN(n695) );
  XNOR2_X1 U790 ( .A(n696), .B(n695), .ZN(n739) );
  XNOR2_X1 U791 ( .A(KEYINPUT65), .B(KEYINPUT26), .ZN(n698) );
  XNOR2_X1 U792 ( .A(n699), .B(n698), .ZN(n702) );
  NAND2_X1 U793 ( .A1(n700), .A2(G1341), .ZN(n701) );
  NAND2_X1 U794 ( .A1(n702), .A2(n701), .ZN(n703) );
  NAND2_X1 U795 ( .A1(n710), .A2(n1001), .ZN(n707) );
  NOR2_X1 U796 ( .A1(n697), .A2(G1348), .ZN(n705) );
  NOR2_X1 U797 ( .A1(G2067), .A2(n700), .ZN(n704) );
  NOR2_X1 U798 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND2_X1 U799 ( .A1(n707), .A2(n706), .ZN(n709) );
  INV_X1 U800 ( .A(KEYINPUT96), .ZN(n708) );
  XNOR2_X1 U801 ( .A(n709), .B(n708), .ZN(n712) );
  NOR2_X1 U802 ( .A1(n1001), .A2(n710), .ZN(n711) );
  NOR2_X1 U803 ( .A1(n712), .A2(n711), .ZN(n718) );
  NAND2_X1 U804 ( .A1(n697), .A2(G2072), .ZN(n713) );
  XOR2_X1 U805 ( .A(KEYINPUT27), .B(n713), .Z(n715) );
  NAND2_X1 U806 ( .A1(G1956), .A2(n700), .ZN(n714) );
  NAND2_X1 U807 ( .A1(n715), .A2(n714), .ZN(n719) );
  NOR2_X1 U808 ( .A1(G299), .A2(n719), .ZN(n716) );
  XOR2_X1 U809 ( .A(KEYINPUT97), .B(n716), .Z(n717) );
  NOR2_X1 U810 ( .A1(n718), .A2(n717), .ZN(n722) );
  NAND2_X1 U811 ( .A1(G299), .A2(n719), .ZN(n720) );
  XOR2_X1 U812 ( .A(KEYINPUT28), .B(n720), .Z(n721) );
  NOR2_X1 U813 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U814 ( .A(n723), .B(KEYINPUT29), .ZN(n726) );
  NAND2_X1 U815 ( .A1(n724), .A2(G171), .ZN(n725) );
  NAND2_X1 U816 ( .A1(n726), .A2(n725), .ZN(n740) );
  NAND2_X1 U817 ( .A1(n739), .A2(n740), .ZN(n727) );
  NAND2_X1 U818 ( .A1(n727), .A2(G286), .ZN(n729) );
  XNOR2_X1 U819 ( .A(n729), .B(n728), .ZN(n735) );
  NOR2_X1 U820 ( .A1(G1971), .A2(n769), .ZN(n731) );
  NOR2_X1 U821 ( .A1(G2090), .A2(n700), .ZN(n730) );
  NOR2_X1 U822 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U823 ( .A1(n732), .A2(G303), .ZN(n733) );
  XNOR2_X1 U824 ( .A(KEYINPUT102), .B(n733), .ZN(n734) );
  NAND2_X1 U825 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U826 ( .A1(n736), .A2(G8), .ZN(n738) );
  XOR2_X1 U827 ( .A(KEYINPUT32), .B(KEYINPUT103), .Z(n737) );
  XNOR2_X1 U828 ( .A(n738), .B(n737), .ZN(n759) );
  AND2_X1 U829 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U830 ( .A1(G8), .A2(n743), .ZN(n744) );
  NAND2_X1 U831 ( .A1(n745), .A2(n744), .ZN(n746) );
  XNOR2_X1 U832 ( .A(KEYINPUT100), .B(n746), .ZN(n760) );
  NAND2_X1 U833 ( .A1(G1976), .A2(G288), .ZN(n1003) );
  AND2_X1 U834 ( .A1(n760), .A2(n1003), .ZN(n747) );
  NAND2_X1 U835 ( .A1(n759), .A2(n747), .ZN(n752) );
  INV_X1 U836 ( .A(n1003), .ZN(n750) );
  NOR2_X1 U837 ( .A1(G1976), .A2(G288), .ZN(n1002) );
  NOR2_X1 U838 ( .A1(G1971), .A2(G303), .ZN(n748) );
  NOR2_X1 U839 ( .A1(n1002), .A2(n748), .ZN(n749) );
  OR2_X1 U840 ( .A1(n750), .A2(n749), .ZN(n751) );
  AND2_X1 U841 ( .A1(n752), .A2(n751), .ZN(n753) );
  NOR2_X1 U842 ( .A1(n769), .A2(n753), .ZN(n754) );
  NAND2_X1 U843 ( .A1(n1002), .A2(KEYINPUT33), .ZN(n755) );
  NOR2_X1 U844 ( .A1(n755), .A2(n769), .ZN(n757) );
  XOR2_X1 U845 ( .A(G1981), .B(G305), .Z(n1013) );
  NAND2_X1 U846 ( .A1(n517), .A2(n758), .ZN(n772) );
  NAND2_X1 U847 ( .A1(n760), .A2(n759), .ZN(n763) );
  NOR2_X1 U848 ( .A1(G2090), .A2(G303), .ZN(n761) );
  NAND2_X1 U849 ( .A1(G8), .A2(n761), .ZN(n762) );
  NAND2_X1 U850 ( .A1(n763), .A2(n762), .ZN(n764) );
  XNOR2_X1 U851 ( .A(n764), .B(KEYINPUT104), .ZN(n765) );
  AND2_X1 U852 ( .A1(n765), .A2(n769), .ZN(n770) );
  NOR2_X1 U853 ( .A1(G1981), .A2(G305), .ZN(n766) );
  XNOR2_X1 U854 ( .A(n766), .B(KEYINPUT24), .ZN(n767) );
  XNOR2_X1 U855 ( .A(KEYINPUT95), .B(n767), .ZN(n768) );
  NOR2_X1 U856 ( .A1(n770), .A2(n516), .ZN(n771) );
  NAND2_X1 U857 ( .A1(n772), .A2(n771), .ZN(n809) );
  XNOR2_X1 U858 ( .A(G1986), .B(G290), .ZN(n1010) );
  NOR2_X1 U859 ( .A1(n774), .A2(n773), .ZN(n820) );
  NAND2_X1 U860 ( .A1(n1010), .A2(n820), .ZN(n807) );
  XNOR2_X1 U861 ( .A(KEYINPUT90), .B(KEYINPUT34), .ZN(n778) );
  NAND2_X1 U862 ( .A1(G104), .A2(n875), .ZN(n776) );
  NAND2_X1 U863 ( .A1(G140), .A2(n876), .ZN(n775) );
  NAND2_X1 U864 ( .A1(n776), .A2(n775), .ZN(n777) );
  XNOR2_X1 U865 ( .A(n778), .B(n777), .ZN(n784) );
  XNOR2_X1 U866 ( .A(KEYINPUT35), .B(KEYINPUT91), .ZN(n782) );
  NAND2_X1 U867 ( .A1(G116), .A2(n879), .ZN(n780) );
  NAND2_X1 U868 ( .A1(G128), .A2(n880), .ZN(n779) );
  NAND2_X1 U869 ( .A1(n780), .A2(n779), .ZN(n781) );
  XNOR2_X1 U870 ( .A(n782), .B(n781), .ZN(n783) );
  NOR2_X1 U871 ( .A1(n784), .A2(n783), .ZN(n785) );
  XNOR2_X1 U872 ( .A(n785), .B(KEYINPUT36), .ZN(n786) );
  XNOR2_X1 U873 ( .A(n786), .B(KEYINPUT92), .ZN(n889) );
  XNOR2_X1 U874 ( .A(G2067), .B(KEYINPUT37), .ZN(n818) );
  NOR2_X1 U875 ( .A1(n889), .A2(n818), .ZN(n923) );
  NAND2_X1 U876 ( .A1(n820), .A2(n923), .ZN(n815) );
  NAND2_X1 U877 ( .A1(G107), .A2(n879), .ZN(n788) );
  NAND2_X1 U878 ( .A1(G119), .A2(n880), .ZN(n787) );
  NAND2_X1 U879 ( .A1(n788), .A2(n787), .ZN(n793) );
  NAND2_X1 U880 ( .A1(G95), .A2(n875), .ZN(n790) );
  NAND2_X1 U881 ( .A1(G131), .A2(n876), .ZN(n789) );
  NAND2_X1 U882 ( .A1(n790), .A2(n789), .ZN(n791) );
  XOR2_X1 U883 ( .A(KEYINPUT93), .B(n791), .Z(n792) );
  NOR2_X1 U884 ( .A1(n793), .A2(n792), .ZN(n888) );
  INV_X1 U885 ( .A(G1991), .ZN(n978) );
  NOR2_X1 U886 ( .A1(n888), .A2(n978), .ZN(n803) );
  XOR2_X1 U887 ( .A(KEYINPUT94), .B(KEYINPUT38), .Z(n795) );
  NAND2_X1 U888 ( .A1(G105), .A2(n875), .ZN(n794) );
  XNOR2_X1 U889 ( .A(n795), .B(n794), .ZN(n799) );
  NAND2_X1 U890 ( .A1(G117), .A2(n879), .ZN(n797) );
  NAND2_X1 U891 ( .A1(G141), .A2(n876), .ZN(n796) );
  NAND2_X1 U892 ( .A1(n797), .A2(n796), .ZN(n798) );
  NOR2_X1 U893 ( .A1(n799), .A2(n798), .ZN(n801) );
  NAND2_X1 U894 ( .A1(n880), .A2(G129), .ZN(n800) );
  NAND2_X1 U895 ( .A1(n801), .A2(n800), .ZN(n872) );
  AND2_X1 U896 ( .A1(n872), .A2(G1996), .ZN(n802) );
  NOR2_X1 U897 ( .A1(n803), .A2(n802), .ZN(n921) );
  INV_X1 U898 ( .A(n820), .ZN(n804) );
  NOR2_X1 U899 ( .A1(n921), .A2(n804), .ZN(n812) );
  INV_X1 U900 ( .A(n812), .ZN(n805) );
  AND2_X1 U901 ( .A1(n815), .A2(n805), .ZN(n806) );
  AND2_X1 U902 ( .A1(n807), .A2(n806), .ZN(n808) );
  NAND2_X1 U903 ( .A1(n809), .A2(n808), .ZN(n823) );
  NOR2_X1 U904 ( .A1(G1996), .A2(n872), .ZN(n918) );
  NOR2_X1 U905 ( .A1(G1986), .A2(G290), .ZN(n810) );
  AND2_X1 U906 ( .A1(n978), .A2(n888), .ZN(n922) );
  NOR2_X1 U907 ( .A1(n810), .A2(n922), .ZN(n811) );
  NOR2_X1 U908 ( .A1(n812), .A2(n811), .ZN(n813) );
  NOR2_X1 U909 ( .A1(n918), .A2(n813), .ZN(n814) );
  XNOR2_X1 U910 ( .A(n814), .B(KEYINPUT39), .ZN(n816) );
  NAND2_X1 U911 ( .A1(n816), .A2(n815), .ZN(n817) );
  XOR2_X1 U912 ( .A(KEYINPUT105), .B(n817), .Z(n819) );
  NAND2_X1 U913 ( .A1(n889), .A2(n818), .ZN(n931) );
  NAND2_X1 U914 ( .A1(n819), .A2(n931), .ZN(n821) );
  NAND2_X1 U915 ( .A1(n821), .A2(n820), .ZN(n822) );
  NAND2_X1 U916 ( .A1(n823), .A2(n822), .ZN(n824) );
  XNOR2_X1 U917 ( .A(KEYINPUT40), .B(n824), .ZN(G329) );
  NAND2_X1 U918 ( .A1(G2106), .A2(n825), .ZN(G217) );
  NAND2_X1 U919 ( .A1(G15), .A2(G2), .ZN(n827) );
  INV_X1 U920 ( .A(G661), .ZN(n826) );
  NOR2_X1 U921 ( .A1(n827), .A2(n826), .ZN(n828) );
  XNOR2_X1 U922 ( .A(n828), .B(KEYINPUT107), .ZN(G259) );
  NAND2_X1 U923 ( .A1(G3), .A2(G1), .ZN(n829) );
  NAND2_X1 U924 ( .A1(n830), .A2(n829), .ZN(G188) );
  XOR2_X1 U925 ( .A(G69), .B(KEYINPUT108), .Z(G235) );
  INV_X1 U927 ( .A(G120), .ZN(G236) );
  NOR2_X1 U928 ( .A1(n832), .A2(n831), .ZN(G325) );
  INV_X1 U929 ( .A(G325), .ZN(G261) );
  INV_X1 U930 ( .A(n833), .ZN(G319) );
  XOR2_X1 U931 ( .A(KEYINPUT42), .B(G2090), .Z(n835) );
  XNOR2_X1 U932 ( .A(G2072), .B(G2084), .ZN(n834) );
  XNOR2_X1 U933 ( .A(n835), .B(n834), .ZN(n836) );
  XOR2_X1 U934 ( .A(n836), .B(G2100), .Z(n838) );
  XNOR2_X1 U935 ( .A(G2067), .B(G2078), .ZN(n837) );
  XNOR2_X1 U936 ( .A(n838), .B(n837), .ZN(n842) );
  XOR2_X1 U937 ( .A(G2096), .B(KEYINPUT43), .Z(n840) );
  XNOR2_X1 U938 ( .A(KEYINPUT109), .B(G2678), .ZN(n839) );
  XNOR2_X1 U939 ( .A(n840), .B(n839), .ZN(n841) );
  XOR2_X1 U940 ( .A(n842), .B(n841), .Z(G227) );
  XNOR2_X1 U941 ( .A(G1991), .B(KEYINPUT41), .ZN(n852) );
  XOR2_X1 U942 ( .A(G1976), .B(G1956), .Z(n844) );
  XNOR2_X1 U943 ( .A(G1996), .B(G1961), .ZN(n843) );
  XNOR2_X1 U944 ( .A(n844), .B(n843), .ZN(n848) );
  XOR2_X1 U945 ( .A(G1981), .B(G1971), .Z(n846) );
  XNOR2_X1 U946 ( .A(G1986), .B(G1966), .ZN(n845) );
  XNOR2_X1 U947 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U948 ( .A(n848), .B(n847), .Z(n850) );
  XNOR2_X1 U949 ( .A(G2474), .B(KEYINPUT110), .ZN(n849) );
  XNOR2_X1 U950 ( .A(n850), .B(n849), .ZN(n851) );
  XNOR2_X1 U951 ( .A(n852), .B(n851), .ZN(G229) );
  NAND2_X1 U952 ( .A1(G124), .A2(n880), .ZN(n853) );
  XNOR2_X1 U953 ( .A(n853), .B(KEYINPUT44), .ZN(n855) );
  NAND2_X1 U954 ( .A1(n879), .A2(G112), .ZN(n854) );
  NAND2_X1 U955 ( .A1(n855), .A2(n854), .ZN(n859) );
  NAND2_X1 U956 ( .A1(G100), .A2(n875), .ZN(n857) );
  NAND2_X1 U957 ( .A1(G136), .A2(n876), .ZN(n856) );
  NAND2_X1 U958 ( .A1(n857), .A2(n856), .ZN(n858) );
  NOR2_X1 U959 ( .A1(n859), .A2(n858), .ZN(G162) );
  NAND2_X1 U960 ( .A1(G118), .A2(n879), .ZN(n861) );
  NAND2_X1 U961 ( .A1(G130), .A2(n880), .ZN(n860) );
  NAND2_X1 U962 ( .A1(n861), .A2(n860), .ZN(n868) );
  XNOR2_X1 U963 ( .A(KEYINPUT112), .B(KEYINPUT45), .ZN(n866) );
  NAND2_X1 U964 ( .A1(n875), .A2(G106), .ZN(n864) );
  NAND2_X1 U965 ( .A1(G142), .A2(n876), .ZN(n862) );
  XOR2_X1 U966 ( .A(KEYINPUT111), .B(n862), .Z(n863) );
  NAND2_X1 U967 ( .A1(n864), .A2(n863), .ZN(n865) );
  XOR2_X1 U968 ( .A(n866), .B(n865), .Z(n867) );
  NOR2_X1 U969 ( .A1(n868), .A2(n867), .ZN(n893) );
  XOR2_X1 U970 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n870) );
  XNOR2_X1 U971 ( .A(G160), .B(n927), .ZN(n869) );
  XNOR2_X1 U972 ( .A(n870), .B(n869), .ZN(n871) );
  XOR2_X1 U973 ( .A(n871), .B(G162), .Z(n874) );
  XOR2_X1 U974 ( .A(G164), .B(n872), .Z(n873) );
  XNOR2_X1 U975 ( .A(n874), .B(n873), .ZN(n887) );
  NAND2_X1 U976 ( .A1(G103), .A2(n875), .ZN(n878) );
  NAND2_X1 U977 ( .A1(G139), .A2(n876), .ZN(n877) );
  NAND2_X1 U978 ( .A1(n878), .A2(n877), .ZN(n885) );
  NAND2_X1 U979 ( .A1(G115), .A2(n879), .ZN(n882) );
  NAND2_X1 U980 ( .A1(G127), .A2(n880), .ZN(n881) );
  NAND2_X1 U981 ( .A1(n882), .A2(n881), .ZN(n883) );
  XOR2_X1 U982 ( .A(KEYINPUT47), .B(n883), .Z(n884) );
  NOR2_X1 U983 ( .A1(n885), .A2(n884), .ZN(n886) );
  XOR2_X1 U984 ( .A(KEYINPUT113), .B(n886), .Z(n933) );
  XOR2_X1 U985 ( .A(n887), .B(n933), .Z(n891) );
  XNOR2_X1 U986 ( .A(n889), .B(n888), .ZN(n890) );
  XNOR2_X1 U987 ( .A(n891), .B(n890), .ZN(n892) );
  XOR2_X1 U988 ( .A(n893), .B(n892), .Z(n894) );
  NOR2_X1 U989 ( .A1(G37), .A2(n894), .ZN(G395) );
  XNOR2_X1 U990 ( .A(n998), .B(KEYINPUT114), .ZN(n896) );
  XNOR2_X1 U991 ( .A(G171), .B(n1001), .ZN(n895) );
  XNOR2_X1 U992 ( .A(n896), .B(n895), .ZN(n899) );
  XOR2_X1 U993 ( .A(G286), .B(n897), .Z(n898) );
  XNOR2_X1 U994 ( .A(n899), .B(n898), .ZN(n900) );
  NOR2_X1 U995 ( .A1(G37), .A2(n900), .ZN(G397) );
  XOR2_X1 U996 ( .A(KEYINPUT106), .B(G2446), .Z(n902) );
  XNOR2_X1 U997 ( .A(G2443), .B(G2454), .ZN(n901) );
  XNOR2_X1 U998 ( .A(n902), .B(n901), .ZN(n903) );
  XOR2_X1 U999 ( .A(n903), .B(G2451), .Z(n905) );
  XNOR2_X1 U1000 ( .A(G1341), .B(G1348), .ZN(n904) );
  XNOR2_X1 U1001 ( .A(n905), .B(n904), .ZN(n909) );
  XOR2_X1 U1002 ( .A(G2435), .B(G2427), .Z(n907) );
  XNOR2_X1 U1003 ( .A(G2430), .B(G2438), .ZN(n906) );
  XNOR2_X1 U1004 ( .A(n907), .B(n906), .ZN(n908) );
  XOR2_X1 U1005 ( .A(n909), .B(n908), .Z(n910) );
  NAND2_X1 U1006 ( .A1(G14), .A2(n910), .ZN(n916) );
  NAND2_X1 U1007 ( .A1(G319), .A2(n916), .ZN(n913) );
  NOR2_X1 U1008 ( .A1(G227), .A2(G229), .ZN(n911) );
  XNOR2_X1 U1009 ( .A(KEYINPUT49), .B(n911), .ZN(n912) );
  NOR2_X1 U1010 ( .A1(n913), .A2(n912), .ZN(n915) );
  NOR2_X1 U1011 ( .A1(G395), .A2(G397), .ZN(n914) );
  NAND2_X1 U1012 ( .A1(n915), .A2(n914), .ZN(G225) );
  INV_X1 U1013 ( .A(G225), .ZN(G308) );
  INV_X1 U1014 ( .A(G96), .ZN(G221) );
  INV_X1 U1015 ( .A(G108), .ZN(G238) );
  INV_X1 U1016 ( .A(n916), .ZN(G401) );
  XOR2_X1 U1017 ( .A(G2090), .B(G162), .Z(n917) );
  NOR2_X1 U1018 ( .A1(n918), .A2(n917), .ZN(n919) );
  XOR2_X1 U1019 ( .A(KEYINPUT51), .B(n919), .Z(n920) );
  NAND2_X1 U1020 ( .A1(n921), .A2(n920), .ZN(n930) );
  XNOR2_X1 U1021 ( .A(G160), .B(G2084), .ZN(n925) );
  NOR2_X1 U1022 ( .A1(n923), .A2(n922), .ZN(n924) );
  NAND2_X1 U1023 ( .A1(n925), .A2(n924), .ZN(n926) );
  NOR2_X1 U1024 ( .A1(n927), .A2(n926), .ZN(n928) );
  XNOR2_X1 U1025 ( .A(KEYINPUT115), .B(n928), .ZN(n929) );
  NOR2_X1 U1026 ( .A1(n930), .A2(n929), .ZN(n932) );
  NAND2_X1 U1027 ( .A1(n932), .A2(n931), .ZN(n938) );
  XOR2_X1 U1028 ( .A(G2072), .B(n933), .Z(n935) );
  XOR2_X1 U1029 ( .A(G164), .B(G2078), .Z(n934) );
  NOR2_X1 U1030 ( .A1(n935), .A2(n934), .ZN(n936) );
  XOR2_X1 U1031 ( .A(KEYINPUT50), .B(n936), .Z(n937) );
  NOR2_X1 U1032 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1033 ( .A(KEYINPUT52), .B(n939), .ZN(n941) );
  INV_X1 U1034 ( .A(KEYINPUT55), .ZN(n940) );
  NAND2_X1 U1035 ( .A1(n941), .A2(n940), .ZN(n942) );
  NAND2_X1 U1036 ( .A1(n942), .A2(G29), .ZN(n943) );
  XNOR2_X1 U1037 ( .A(KEYINPUT116), .B(n943), .ZN(n996) );
  XNOR2_X1 U1038 ( .A(G1341), .B(KEYINPUT123), .ZN(n944) );
  XNOR2_X1 U1039 ( .A(n944), .B(G19), .ZN(n950) );
  XNOR2_X1 U1040 ( .A(G1956), .B(G20), .ZN(n945) );
  XNOR2_X1 U1041 ( .A(n945), .B(KEYINPUT122), .ZN(n948) );
  XNOR2_X1 U1042 ( .A(G1981), .B(KEYINPUT124), .ZN(n946) );
  XNOR2_X1 U1043 ( .A(n946), .B(G6), .ZN(n947) );
  NOR2_X1 U1044 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1045 ( .A1(n950), .A2(n949), .ZN(n953) );
  XOR2_X1 U1046 ( .A(KEYINPUT59), .B(G1348), .Z(n951) );
  XNOR2_X1 U1047 ( .A(G4), .B(n951), .ZN(n952) );
  NOR2_X1 U1048 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1049 ( .A(KEYINPUT60), .B(n954), .ZN(n956) );
  XOR2_X1 U1050 ( .A(G1961), .B(G5), .Z(n955) );
  NAND2_X1 U1051 ( .A1(n956), .A2(n955), .ZN(n967) );
  XOR2_X1 U1052 ( .A(G1966), .B(G21), .Z(n965) );
  XOR2_X1 U1053 ( .A(G1971), .B(G22), .Z(n959) );
  XOR2_X1 U1054 ( .A(G24), .B(KEYINPUT126), .Z(n957) );
  XNOR2_X1 U1055 ( .A(n957), .B(G1986), .ZN(n958) );
  NAND2_X1 U1056 ( .A1(n959), .A2(n958), .ZN(n962) );
  XOR2_X1 U1057 ( .A(KEYINPUT125), .B(G1976), .Z(n960) );
  XNOR2_X1 U1058 ( .A(G23), .B(n960), .ZN(n961) );
  NOR2_X1 U1059 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1060 ( .A(n963), .B(KEYINPUT58), .ZN(n964) );
  NAND2_X1 U1061 ( .A1(n965), .A2(n964), .ZN(n966) );
  NOR2_X1 U1062 ( .A1(n967), .A2(n966), .ZN(n968) );
  XOR2_X1 U1063 ( .A(KEYINPUT61), .B(n968), .Z(n969) );
  NOR2_X1 U1064 ( .A1(G16), .A2(n969), .ZN(n994) );
  XOR2_X1 U1065 ( .A(G2090), .B(G35), .Z(n973) );
  XOR2_X1 U1066 ( .A(G2084), .B(KEYINPUT118), .Z(n970) );
  XNOR2_X1 U1067 ( .A(G34), .B(n970), .ZN(n971) );
  XNOR2_X1 U1068 ( .A(n971), .B(KEYINPUT54), .ZN(n972) );
  NAND2_X1 U1069 ( .A1(n973), .A2(n972), .ZN(n988) );
  XOR2_X1 U1070 ( .A(G2067), .B(G26), .Z(n974) );
  NAND2_X1 U1071 ( .A1(n974), .A2(G28), .ZN(n984) );
  XNOR2_X1 U1072 ( .A(G1996), .B(G32), .ZN(n976) );
  XNOR2_X1 U1073 ( .A(G33), .B(G2072), .ZN(n975) );
  NOR2_X1 U1074 ( .A1(n976), .A2(n975), .ZN(n982) );
  XOR2_X1 U1075 ( .A(n977), .B(G27), .Z(n980) );
  XOR2_X1 U1076 ( .A(n978), .B(G25), .Z(n979) );
  NOR2_X1 U1077 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1078 ( .A1(n982), .A2(n981), .ZN(n983) );
  NOR2_X1 U1079 ( .A1(n984), .A2(n983), .ZN(n985) );
  XOR2_X1 U1080 ( .A(KEYINPUT53), .B(n985), .Z(n986) );
  XNOR2_X1 U1081 ( .A(n986), .B(KEYINPUT117), .ZN(n987) );
  NOR2_X1 U1082 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1083 ( .A(n989), .B(KEYINPUT55), .ZN(n991) );
  XNOR2_X1 U1084 ( .A(G29), .B(KEYINPUT119), .ZN(n990) );
  NAND2_X1 U1085 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1086 ( .A1(G11), .A2(n992), .ZN(n993) );
  NOR2_X1 U1087 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1088 ( .A1(n996), .A2(n995), .ZN(n1024) );
  XOR2_X1 U1089 ( .A(G16), .B(KEYINPUT56), .Z(n1022) );
  XNOR2_X1 U1090 ( .A(G1971), .B(KEYINPUT120), .ZN(n997) );
  XNOR2_X1 U1091 ( .A(n997), .B(G303), .ZN(n1000) );
  XNOR2_X1 U1092 ( .A(G1341), .B(n998), .ZN(n999) );
  NOR2_X1 U1093 ( .A1(n1000), .A2(n999), .ZN(n1012) );
  XNOR2_X1 U1094 ( .A(n1001), .B(G1348), .ZN(n1008) );
  INV_X1 U1095 ( .A(n1002), .ZN(n1004) );
  NAND2_X1 U1096 ( .A1(n1004), .A2(n1003), .ZN(n1006) );
  XNOR2_X1 U1097 ( .A(G1956), .B(G299), .ZN(n1005) );
  NOR2_X1 U1098 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1099 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NOR2_X1 U1100 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1101 ( .A1(n1012), .A2(n1011), .ZN(n1019) );
  XNOR2_X1 U1102 ( .A(G171), .B(G1961), .ZN(n1017) );
  XNOR2_X1 U1103 ( .A(G168), .B(G1966), .ZN(n1014) );
  NAND2_X1 U1104 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XNOR2_X1 U1105 ( .A(n1015), .B(KEYINPUT57), .ZN(n1016) );
  NAND2_X1 U1106 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NOR2_X1 U1107 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XOR2_X1 U1108 ( .A(KEYINPUT121), .B(n1020), .Z(n1021) );
  NOR2_X1 U1109 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NOR2_X1 U1110 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XNOR2_X1 U1111 ( .A(n1025), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1112 ( .A(G311), .ZN(G150) );
endmodule

