//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 0 1 1 1 1 1 1 0 1 0 1 1 1 1 0 1 1 0 1 0 0 1 0 0 1 1 1 1 1 0 1 0 1 1 1 0 1 1 0 1 1 1 0 0 0 1 0 0 0 0 0 1 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:04 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n444, new_n448, new_n449, new_n451, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n565, new_n567,
    new_n568, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n604, new_n605, new_n606, new_n607, new_n610, new_n611,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1146;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT65), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  XOR2_X1   g016(.A(KEYINPUT66), .B(G108), .Z(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XOR2_X1   g019(.A(new_n444), .B(KEYINPUT67), .Z(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g022(.A(KEYINPUT68), .B(KEYINPUT1), .ZN(new_n448));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n448), .B(new_n449), .ZN(G223));
  INV_X1    g025(.A(new_n449), .ZN(new_n451));
  NAND2_X1  g026(.A1(new_n451), .A2(G567), .ZN(G234));
  NAND2_X1  g027(.A1(new_n451), .A2(G2106), .ZN(G217));
  NAND4_X1  g028(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n454));
  XNOR2_X1  g029(.A(KEYINPUT69), .B(KEYINPUT2), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n454), .B(new_n455), .ZN(new_n456));
  NOR4_X1   g031(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n456), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  NAND2_X1  g035(.A1(new_n456), .A2(G2106), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n458), .A2(G567), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  INV_X1    g041(.A(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(KEYINPUT70), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT70), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n467), .B1(new_n472), .B2(KEYINPUT3), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G137), .ZN(new_n474));
  XNOR2_X1  g049(.A(KEYINPUT70), .B(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G101), .ZN(new_n476));
  AOI21_X1  g051(.A(G2105), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(G113), .A2(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n468), .A2(KEYINPUT3), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n466), .A2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(G125), .ZN(new_n481));
  OAI21_X1  g056(.A(new_n478), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G2105), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n477), .A2(new_n484), .ZN(G160));
  INV_X1    g060(.A(G2105), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n473), .A2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(G136), .ZN(new_n488));
  NOR2_X1   g063(.A1(G100), .A2(G2105), .ZN(new_n489));
  OAI21_X1  g064(.A(G2104), .B1(new_n486), .B2(G112), .ZN(new_n490));
  OAI22_X1  g065(.A1(new_n487), .A2(new_n488), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n473), .A2(G2105), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n491), .B1(G124), .B2(new_n493), .ZN(G162));
  OAI211_X1 g069(.A(G126), .B(new_n466), .C1(new_n475), .C2(new_n465), .ZN(new_n495));
  NAND2_X1  g070(.A1(G114), .A2(G2104), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(G2105), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n470), .A2(G2104), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n468), .A2(KEYINPUT70), .ZN(new_n500));
  OAI21_X1  g075(.A(KEYINPUT3), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  AND2_X1   g076(.A1(KEYINPUT4), .A2(G138), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n501), .A2(new_n486), .A3(new_n466), .A4(new_n502), .ZN(new_n503));
  AND3_X1   g078(.A1(new_n486), .A2(G102), .A3(G2104), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n466), .A2(new_n479), .A3(G138), .A4(new_n486), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT4), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND4_X1  g082(.A1(new_n498), .A2(KEYINPUT71), .A3(new_n503), .A4(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT71), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n503), .A2(new_n507), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n486), .B1(new_n495), .B2(new_n496), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n508), .A2(new_n512), .ZN(G164));
  NAND2_X1  g088(.A1(KEYINPUT73), .A2(G543), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT5), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n514), .A2(KEYINPUT72), .A3(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT72), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n517), .B1(KEYINPUT73), .B2(G543), .ZN(new_n518));
  INV_X1    g093(.A(G543), .ZN(new_n519));
  OAI21_X1  g094(.A(KEYINPUT5), .B1(new_n519), .B2(KEYINPUT72), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n516), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n521), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n522));
  INV_X1    g097(.A(G651), .ZN(new_n523));
  OR2_X1    g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  XNOR2_X1  g099(.A(KEYINPUT6), .B(G651), .ZN(new_n525));
  XNOR2_X1  g100(.A(KEYINPUT74), .B(G88), .ZN(new_n526));
  AND2_X1   g101(.A1(new_n521), .A2(new_n526), .ZN(new_n527));
  AND2_X1   g102(.A1(G50), .A2(G543), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n525), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n524), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(KEYINPUT75), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT75), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n524), .A2(new_n532), .A3(new_n529), .ZN(new_n533));
  AND2_X1   g108(.A1(new_n531), .A2(new_n533), .ZN(G303));
  INV_X1    g109(.A(G303), .ZN(G166));
  XOR2_X1   g110(.A(KEYINPUT6), .B(G651), .Z(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(KEYINPUT76), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT76), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n525), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n537), .A2(G543), .A3(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G51), .ZN(new_n542));
  INV_X1    g117(.A(new_n521), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n525), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n544));
  OR2_X1    g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g120(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT7), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n542), .A2(new_n545), .A3(new_n547), .ZN(G286));
  INV_X1    g123(.A(G286), .ZN(G168));
  INV_X1    g124(.A(G52), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n521), .A2(new_n525), .ZN(new_n551));
  INV_X1    g126(.A(G90), .ZN(new_n552));
  OAI22_X1  g127(.A1(new_n540), .A2(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  AOI22_X1  g128(.A1(new_n521), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n554), .A2(new_n523), .ZN(new_n555));
  OR2_X1    g130(.A1(new_n553), .A2(new_n555), .ZN(G301));
  INV_X1    g131(.A(G301), .ZN(G171));
  INV_X1    g132(.A(G43), .ZN(new_n558));
  INV_X1    g133(.A(G81), .ZN(new_n559));
  OAI22_X1  g134(.A1(new_n540), .A2(new_n558), .B1(new_n551), .B2(new_n559), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n521), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n561));
  NOR2_X1   g136(.A1(new_n561), .A2(new_n523), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G860), .ZN(G153));
  AND3_X1   g139(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G36), .ZN(G176));
  NAND2_X1  g141(.A1(G1), .A2(G3), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT8), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n565), .A2(new_n568), .ZN(G188));
  INV_X1    g144(.A(new_n551), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(G91), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n521), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n572));
  NAND4_X1  g147(.A1(new_n537), .A2(G53), .A3(G543), .A4(new_n539), .ZN(new_n573));
  AND2_X1   g148(.A1(new_n573), .A2(KEYINPUT9), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n573), .A2(KEYINPUT9), .ZN(new_n575));
  OAI221_X1 g150(.A(new_n571), .B1(new_n523), .B2(new_n572), .C1(new_n574), .C2(new_n575), .ZN(G299));
  NAND2_X1  g151(.A1(new_n541), .A2(G49), .ZN(new_n577));
  OAI21_X1  g152(.A(G651), .B1(new_n521), .B2(G74), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n570), .A2(G87), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(G288));
  AOI22_X1  g155(.A1(new_n521), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n521), .A2(G86), .B1(G48), .B2(G543), .ZN(new_n582));
  OAI22_X1  g157(.A1(new_n523), .A2(new_n581), .B1(new_n582), .B2(new_n536), .ZN(G305));
  INV_X1    g158(.A(G47), .ZN(new_n584));
  INV_X1    g159(.A(G85), .ZN(new_n585));
  OAI22_X1  g160(.A1(new_n540), .A2(new_n584), .B1(new_n551), .B2(new_n585), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n521), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n587), .A2(new_n523), .ZN(new_n588));
  OR2_X1    g163(.A1(new_n586), .A2(new_n588), .ZN(G290));
  NAND2_X1  g164(.A1(G301), .A2(G868), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n570), .A2(KEYINPUT10), .A3(G92), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT10), .ZN(new_n592));
  INV_X1    g167(.A(G92), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n551), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(G79), .A2(G543), .ZN(new_n595));
  INV_X1    g170(.A(G66), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n543), .B2(new_n596), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n591), .A2(new_n594), .B1(G651), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n541), .A2(G54), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n590), .B1(new_n601), .B2(G868), .ZN(G321));
  XOR2_X1   g177(.A(G321), .B(KEYINPUT77), .Z(G284));
  NAND2_X1  g178(.A1(G286), .A2(G868), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n574), .A2(new_n575), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n571), .B1(new_n572), .B2(new_n523), .ZN(new_n606));
  NOR2_X1   g181(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n604), .B1(new_n607), .B2(G868), .ZN(G297));
  OAI21_X1  g183(.A(new_n604), .B1(new_n607), .B2(G868), .ZN(G280));
  XOR2_X1   g184(.A(KEYINPUT78), .B(G559), .Z(new_n610));
  OAI21_X1  g185(.A(new_n601), .B1(G860), .B2(new_n610), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT79), .ZN(G148));
  OR2_X1    g187(.A1(new_n560), .A2(new_n562), .ZN(new_n613));
  NOR2_X1   g188(.A1(new_n613), .A2(G868), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n601), .A2(new_n610), .ZN(new_n615));
  XOR2_X1   g190(.A(new_n615), .B(KEYINPUT80), .Z(new_n616));
  AOI21_X1  g191(.A(new_n614), .B1(new_n616), .B2(G868), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT81), .ZN(G323));
  XNOR2_X1  g193(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR3_X1   g194(.A1(new_n480), .A2(new_n472), .A3(G2105), .ZN(new_n620));
  XOR2_X1   g195(.A(new_n620), .B(KEYINPUT12), .Z(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT13), .ZN(new_n622));
  NOR2_X1   g197(.A1(KEYINPUT82), .A2(G2100), .ZN(new_n623));
  AND2_X1   g198(.A1(KEYINPUT82), .A2(G2100), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n622), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n493), .A2(G123), .ZN(new_n626));
  INV_X1    g201(.A(new_n487), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n627), .A2(G135), .ZN(new_n628));
  NOR2_X1   g203(.A1(G99), .A2(G2105), .ZN(new_n629));
  OAI21_X1  g204(.A(G2104), .B1(new_n486), .B2(G111), .ZN(new_n630));
  OAI211_X1 g205(.A(new_n626), .B(new_n628), .C1(new_n629), .C2(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(G2096), .Z(new_n632));
  OAI211_X1 g207(.A(new_n625), .B(new_n632), .C1(new_n623), .C2(new_n622), .ZN(G156));
  XOR2_X1   g208(.A(KEYINPUT84), .B(G2438), .Z(new_n634));
  XNOR2_X1  g209(.A(G2427), .B(G2430), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(KEYINPUT15), .B(G2435), .Z(new_n637));
  INV_X1    g212(.A(KEYINPUT14), .ZN(new_n638));
  AOI22_X1  g213(.A1(new_n636), .A2(new_n637), .B1(KEYINPUT83), .B2(new_n638), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n638), .A2(KEYINPUT83), .ZN(new_n640));
  OAI211_X1 g215(.A(new_n639), .B(new_n640), .C1(new_n637), .C2(new_n636), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2451), .B(G2454), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT85), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT16), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n641), .B(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(G1341), .B(G1348), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2443), .B(G2446), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n647), .B(new_n648), .Z(new_n649));
  AND2_X1   g224(.A1(new_n649), .A2(G14), .ZN(G401));
  XOR2_X1   g225(.A(G2084), .B(G2090), .Z(new_n651));
  XNOR2_X1  g226(.A(G2067), .B(G2678), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2072), .B(G2078), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n651), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n654), .B(KEYINPUT18), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n652), .B(KEYINPUT86), .ZN(new_n656));
  OAI21_X1  g231(.A(KEYINPUT17), .B1(new_n656), .B2(new_n651), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n657), .B(new_n653), .Z(new_n658));
  AND2_X1   g233(.A1(new_n656), .A2(new_n651), .ZN(new_n659));
  OAI21_X1  g234(.A(new_n655), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(G2100), .ZN(new_n661));
  XNOR2_X1  g236(.A(KEYINPUT87), .B(G2096), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(G227));
  XNOR2_X1  g238(.A(G1961), .B(G1966), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(G1956), .B(G2474), .Z(new_n666));
  NAND2_X1  g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n667), .A2(KEYINPUT89), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n667), .A2(KEYINPUT89), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1971), .B(G1976), .ZN(new_n670));
  XNOR2_X1  g245(.A(KEYINPUT88), .B(KEYINPUT19), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n668), .A2(new_n669), .A3(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(KEYINPUT90), .B(KEYINPUT20), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n665), .A2(new_n666), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n672), .A2(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(new_n676), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n678), .A2(new_n667), .ZN(new_n679));
  OAI211_X1 g254(.A(new_n675), .B(new_n677), .C1(new_n672), .C2(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(G1986), .B(G1996), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n683));
  INV_X1    g258(.A(G1981), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(G1991), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n682), .B(new_n686), .ZN(G229));
  INV_X1    g262(.A(G16), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n688), .A2(G24), .ZN(new_n689));
  INV_X1    g264(.A(G290), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n689), .B1(new_n690), .B2(new_n688), .ZN(new_n691));
  MUX2_X1   g266(.A(new_n689), .B(new_n691), .S(KEYINPUT92), .Z(new_n692));
  AND2_X1   g267(.A1(new_n692), .A2(G1986), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n627), .A2(KEYINPUT91), .A3(G131), .ZN(new_n694));
  INV_X1    g269(.A(KEYINPUT91), .ZN(new_n695));
  INV_X1    g270(.A(G131), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n695), .B1(new_n487), .B2(new_n696), .ZN(new_n697));
  AOI22_X1  g272(.A1(new_n694), .A2(new_n697), .B1(G119), .B2(new_n493), .ZN(new_n698));
  OR2_X1    g273(.A1(G95), .A2(G2105), .ZN(new_n699));
  OAI211_X1 g274(.A(new_n699), .B(G2104), .C1(G107), .C2(new_n486), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  MUX2_X1   g276(.A(G25), .B(new_n701), .S(G29), .Z(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT35), .B(G1991), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n688), .A2(G23), .ZN(new_n705));
  INV_X1    g280(.A(G288), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n705), .B1(new_n706), .B2(new_n688), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT33), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(G1976), .ZN(new_n709));
  NOR2_X1   g284(.A1(G16), .A2(G22), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n710), .B1(G166), .B2(G16), .ZN(new_n711));
  INV_X1    g286(.A(G1971), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n688), .A2(G6), .ZN(new_n714));
  INV_X1    g289(.A(G305), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n714), .B1(new_n715), .B2(new_n688), .ZN(new_n716));
  XOR2_X1   g291(.A(KEYINPUT32), .B(G1981), .Z(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT93), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n716), .B(new_n718), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n709), .A2(new_n713), .A3(new_n719), .ZN(new_n720));
  AOI211_X1 g295(.A(new_n693), .B(new_n704), .C1(new_n720), .C2(KEYINPUT34), .ZN(new_n721));
  OAI221_X1 g296(.A(new_n721), .B1(KEYINPUT34), .B2(new_n720), .C1(G1986), .C2(new_n692), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT36), .ZN(new_n723));
  XNOR2_X1  g298(.A(KEYINPUT31), .B(G11), .ZN(new_n724));
  NOR2_X1   g299(.A1(G27), .A2(G29), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n725), .B1(G164), .B2(G29), .ZN(new_n726));
  XNOR2_X1  g301(.A(KEYINPUT101), .B(G2078), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n627), .A2(G141), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n493), .A2(G129), .ZN(new_n730));
  NAND3_X1  g305(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(KEYINPUT26), .Z(new_n732));
  NAND3_X1  g307(.A1(new_n475), .A2(G105), .A3(new_n486), .ZN(new_n733));
  NAND4_X1  g308(.A1(new_n729), .A2(new_n730), .A3(new_n732), .A4(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n735), .A2(G29), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(G29), .B2(G32), .ZN(new_n737));
  XNOR2_X1  g312(.A(KEYINPUT27), .B(G1996), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g314(.A1(G5), .A2(G16), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(G171), .B2(G16), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n741), .A2(G1961), .ZN(new_n742));
  AND2_X1   g317(.A1(new_n739), .A2(new_n742), .ZN(new_n743));
  OR2_X1    g318(.A1(KEYINPUT24), .A2(G34), .ZN(new_n744));
  INV_X1    g319(.A(G29), .ZN(new_n745));
  NAND2_X1  g320(.A1(KEYINPUT24), .A2(G34), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n744), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(G160), .B2(new_n745), .ZN(new_n748));
  OAI221_X1 g323(.A(new_n743), .B1(G2084), .B2(new_n748), .C1(new_n737), .C2(new_n738), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n748), .A2(G2084), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(new_n741), .B2(G1961), .ZN(new_n751));
  NAND2_X1  g326(.A1(G168), .A2(G16), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(G16), .B2(G21), .ZN(new_n753));
  INV_X1    g328(.A(G1966), .ZN(new_n754));
  OR2_X1    g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n753), .A2(new_n754), .ZN(new_n756));
  OR2_X1    g331(.A1(new_n631), .A2(new_n745), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT30), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n745), .B1(new_n758), .B2(G28), .ZN(new_n759));
  OR2_X1    g334(.A1(new_n759), .A2(KEYINPUT100), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n758), .A2(G28), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n759), .A2(KEYINPUT100), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n760), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  NAND4_X1  g338(.A1(new_n755), .A2(new_n756), .A3(new_n757), .A4(new_n763), .ZN(new_n764));
  OR4_X1    g339(.A1(new_n728), .A2(new_n749), .A3(new_n751), .A4(new_n764), .ZN(new_n765));
  AND2_X1   g340(.A1(new_n688), .A2(G19), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(new_n613), .B2(G16), .ZN(new_n767));
  MUX2_X1   g342(.A(new_n766), .B(new_n767), .S(KEYINPUT95), .Z(new_n768));
  INV_X1    g343(.A(new_n768), .ZN(new_n769));
  XOR2_X1   g344(.A(KEYINPUT97), .B(KEYINPUT28), .Z(new_n770));
  NAND2_X1  g345(.A1(new_n745), .A2(G26), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  OR2_X1    g347(.A1(G104), .A2(G2105), .ZN(new_n773));
  OAI211_X1 g348(.A(new_n773), .B(G2104), .C1(G116), .C2(new_n486), .ZN(new_n774));
  INV_X1    g349(.A(G128), .ZN(new_n775));
  INV_X1    g350(.A(G140), .ZN(new_n776));
  OAI221_X1 g351(.A(new_n774), .B1(new_n492), .B2(new_n775), .C1(new_n776), .C2(new_n487), .ZN(new_n777));
  OR2_X1    g352(.A1(new_n777), .A2(KEYINPUT96), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n777), .A2(KEYINPUT96), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(new_n780), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n772), .B1(new_n781), .B2(new_n745), .ZN(new_n782));
  AOI22_X1  g357(.A1(new_n769), .A2(G1341), .B1(new_n782), .B2(G2067), .ZN(new_n783));
  INV_X1    g358(.A(G2090), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n745), .A2(G35), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(G162), .B2(new_n745), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(KEYINPUT29), .Z(new_n787));
  OAI221_X1 g362(.A(new_n783), .B1(G1341), .B2(new_n769), .C1(new_n784), .C2(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n627), .A2(G139), .ZN(new_n789));
  NAND3_X1  g364(.A1(new_n486), .A2(G103), .A3(G2104), .ZN(new_n790));
  XOR2_X1   g365(.A(new_n790), .B(KEYINPUT25), .Z(new_n791));
  NAND2_X1  g366(.A1(G115), .A2(G2104), .ZN(new_n792));
  INV_X1    g367(.A(G127), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n792), .B1(new_n480), .B2(new_n793), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT98), .Z(new_n795));
  OAI211_X1 g370(.A(new_n789), .B(new_n791), .C1(new_n795), .C2(new_n486), .ZN(new_n796));
  MUX2_X1   g371(.A(G33), .B(new_n796), .S(G29), .Z(new_n797));
  XOR2_X1   g372(.A(new_n797), .B(KEYINPUT99), .Z(new_n798));
  OR2_X1    g373(.A1(new_n798), .A2(G2072), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n787), .A2(new_n784), .ZN(new_n800));
  OR2_X1    g375(.A1(new_n782), .A2(G2067), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n798), .A2(G2072), .ZN(new_n802));
  NAND4_X1  g377(.A1(new_n799), .A2(new_n800), .A3(new_n801), .A4(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n688), .A2(G20), .ZN(new_n804));
  OAI211_X1 g379(.A(KEYINPUT23), .B(new_n804), .C1(new_n607), .C2(new_n688), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(KEYINPUT23), .B2(new_n804), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(G1956), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n688), .A2(G4), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(new_n601), .B2(new_n688), .ZN(new_n809));
  XOR2_X1   g384(.A(KEYINPUT94), .B(G1348), .Z(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n807), .A2(new_n811), .ZN(new_n812));
  NOR4_X1   g387(.A1(new_n765), .A2(new_n788), .A3(new_n803), .A4(new_n812), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n723), .A2(new_n724), .A3(new_n813), .ZN(G150));
  INV_X1    g389(.A(G150), .ZN(G311));
  INV_X1    g390(.A(G55), .ZN(new_n816));
  INV_X1    g391(.A(G93), .ZN(new_n817));
  OAI22_X1  g392(.A1(new_n540), .A2(new_n816), .B1(new_n551), .B2(new_n817), .ZN(new_n818));
  AOI22_X1  g393(.A1(new_n521), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n819), .A2(new_n523), .ZN(new_n820));
  OR2_X1    g395(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n821), .A2(G860), .ZN(new_n822));
  XOR2_X1   g397(.A(new_n822), .B(KEYINPUT37), .Z(new_n823));
  NAND2_X1  g398(.A1(new_n601), .A2(G559), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT38), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n821), .A2(new_n563), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n818), .A2(new_n820), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n613), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT39), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n825), .B(new_n830), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n823), .B1(new_n831), .B2(G860), .ZN(G145));
  XNOR2_X1  g407(.A(new_n780), .B(new_n621), .ZN(new_n833));
  INV_X1    g408(.A(new_n496), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n834), .B1(new_n473), .B2(G126), .ZN(new_n835));
  OAI211_X1 g410(.A(new_n503), .B(new_n507), .C1(new_n835), .C2(new_n486), .ZN(new_n836));
  XOR2_X1   g411(.A(new_n734), .B(new_n836), .Z(new_n837));
  XNOR2_X1  g412(.A(new_n833), .B(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n701), .B(new_n796), .ZN(new_n839));
  XOR2_X1   g414(.A(new_n838), .B(new_n839), .Z(new_n840));
  XNOR2_X1  g415(.A(new_n631), .B(G160), .ZN(new_n841));
  XOR2_X1   g416(.A(new_n841), .B(G162), .Z(new_n842));
  NAND3_X1  g417(.A1(new_n627), .A2(KEYINPUT102), .A3(G142), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n493), .A2(G130), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT102), .ZN(new_n845));
  INV_X1    g420(.A(G142), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n845), .B1(new_n487), .B2(new_n846), .ZN(new_n847));
  OR2_X1    g422(.A1(G106), .A2(G2105), .ZN(new_n848));
  OAI211_X1 g423(.A(new_n848), .B(G2104), .C1(G118), .C2(new_n486), .ZN(new_n849));
  NAND4_X1  g424(.A1(new_n843), .A2(new_n844), .A3(new_n847), .A4(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n842), .B(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n840), .A2(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(G37), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n838), .B(new_n839), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n855), .A2(new_n851), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n853), .A2(new_n854), .A3(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g433(.A(new_n607), .B(new_n600), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(KEYINPUT41), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n859), .B(KEYINPUT104), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  XOR2_X1   g437(.A(new_n829), .B(KEYINPUT103), .Z(new_n863));
  XNOR2_X1  g438(.A(new_n616), .B(new_n863), .ZN(new_n864));
  MUX2_X1   g439(.A(new_n860), .B(new_n862), .S(new_n864), .Z(new_n865));
  XNOR2_X1  g440(.A(G290), .B(new_n715), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(G303), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(new_n706), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(KEYINPUT42), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n865), .B(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n870), .A2(G868), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n871), .B1(G868), .B2(new_n827), .ZN(G295));
  OAI21_X1  g447(.A(new_n871), .B1(G868), .B2(new_n827), .ZN(G331));
  INV_X1    g448(.A(KEYINPUT44), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n829), .B(G301), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(G286), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n876), .A2(new_n860), .ZN(new_n877));
  OR2_X1    g452(.A1(new_n875), .A2(G168), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n875), .A2(G168), .ZN(new_n879));
  AND3_X1   g454(.A1(new_n878), .A2(new_n859), .A3(new_n879), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n877), .A2(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(G37), .B1(new_n881), .B2(new_n868), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT105), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT43), .ZN(new_n884));
  INV_X1    g459(.A(new_n868), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n885), .B1(new_n877), .B2(new_n880), .ZN(new_n886));
  NAND4_X1  g461(.A1(new_n882), .A2(new_n883), .A3(new_n884), .A4(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n876), .A2(new_n859), .ZN(new_n888));
  OAI211_X1 g463(.A(new_n888), .B(new_n868), .C1(new_n860), .C2(new_n876), .ZN(new_n889));
  NAND4_X1  g464(.A1(new_n886), .A2(new_n889), .A3(new_n884), .A4(new_n854), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n890), .A2(KEYINPUT105), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n874), .B1(new_n887), .B2(new_n891), .ZN(new_n892));
  AND2_X1   g467(.A1(new_n876), .A2(new_n861), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n885), .B1(new_n893), .B2(new_n877), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n882), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n895), .A2(KEYINPUT43), .ZN(new_n896));
  AND3_X1   g471(.A1(new_n892), .A2(KEYINPUT106), .A3(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(KEYINPUT106), .B1(new_n892), .B2(new_n896), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n889), .A2(new_n854), .ZN(new_n899));
  INV_X1    g474(.A(new_n886), .ZN(new_n900));
  OAI21_X1  g475(.A(KEYINPUT43), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n882), .A2(new_n884), .A3(new_n894), .ZN(new_n902));
  AND2_X1   g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  OAI22_X1  g478(.A1(new_n897), .A2(new_n898), .B1(KEYINPUT44), .B2(new_n903), .ZN(G397));
  INV_X1    g479(.A(G1384), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n905), .B1(new_n510), .B2(new_n511), .ZN(new_n906));
  XNOR2_X1  g481(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  AOI22_X1  g484(.A1(new_n473), .A2(G137), .B1(G101), .B2(new_n475), .ZN(new_n910));
  OAI211_X1 g485(.A(G40), .B(new_n483), .C1(new_n910), .C2(G2105), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(G2067), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n780), .B(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(G1996), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n734), .B(new_n916), .ZN(new_n917));
  AND2_X1   g492(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n701), .A2(new_n703), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n781), .A2(new_n914), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n913), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n912), .A2(new_n916), .ZN(new_n923));
  XOR2_X1   g498(.A(new_n923), .B(KEYINPUT46), .Z(new_n924));
  NAND2_X1  g499(.A1(new_n915), .A2(new_n735), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n924), .B1(new_n925), .B2(new_n912), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n926), .B(KEYINPUT47), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n701), .A2(new_n703), .ZN(new_n928));
  INV_X1    g503(.A(new_n919), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n918), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n930), .A2(new_n912), .ZN(new_n931));
  OR2_X1    g506(.A1(G290), .A2(G1986), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n913), .A2(new_n932), .ZN(new_n933));
  XOR2_X1   g508(.A(new_n933), .B(KEYINPUT48), .Z(new_n934));
  AOI211_X1 g509(.A(new_n922), .B(new_n927), .C1(new_n931), .C2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT125), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n531), .A2(G8), .A3(new_n533), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(KEYINPUT55), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT55), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n531), .A2(new_n939), .A3(G8), .A4(new_n533), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(new_n941), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n508), .A2(new_n905), .A3(new_n512), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(KEYINPUT50), .ZN(new_n944));
  INV_X1    g519(.A(new_n911), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT50), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n836), .A2(new_n946), .A3(new_n905), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n944), .A2(new_n945), .A3(new_n947), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n948), .A2(G2090), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n836), .A2(KEYINPUT45), .A3(new_n905), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(new_n945), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n951), .B1(new_n943), .B2(new_n908), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n952), .A2(G1971), .ZN(new_n953));
  OAI211_X1 g528(.A(new_n942), .B(G8), .C1(new_n949), .C2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(G8), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n943), .A2(new_n908), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n956), .A2(new_n945), .A3(new_n950), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(new_n712), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT114), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n946), .B1(new_n836), .B2(new_n905), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n959), .B1(new_n960), .B2(new_n911), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n508), .A2(new_n512), .A3(new_n946), .A4(new_n905), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n906), .A2(KEYINPUT50), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n963), .A2(KEYINPUT114), .A3(new_n945), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n961), .A2(new_n784), .A3(new_n962), .A4(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n955), .B1(new_n958), .B2(new_n965), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n954), .B1(new_n942), .B2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT110), .ZN(new_n968));
  NAND3_X1  g543(.A1(G305), .A2(new_n968), .A3(G1981), .ZN(new_n969));
  INV_X1    g544(.A(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n968), .B1(G305), .B2(G1981), .ZN(new_n971));
  XNOR2_X1  g546(.A(KEYINPUT109), .B(G1981), .ZN(new_n972));
  NOR2_X1   g547(.A1(G305), .A2(new_n972), .ZN(new_n973));
  NOR3_X1   g548(.A1(new_n970), .A2(new_n971), .A3(new_n973), .ZN(new_n974));
  OAI21_X1  g549(.A(KEYINPUT49), .B1(new_n974), .B2(KEYINPUT111), .ZN(new_n975));
  OR2_X1    g550(.A1(new_n906), .A2(new_n911), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(G8), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT108), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  OAI211_X1 g554(.A(KEYINPUT108), .B(G8), .C1(new_n906), .C2(new_n911), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(new_n971), .ZN(new_n982));
  INV_X1    g557(.A(new_n973), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n982), .A2(new_n983), .A3(new_n969), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT111), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT49), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n984), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n975), .A2(new_n981), .A3(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n706), .A2(G1976), .ZN(new_n989));
  INV_X1    g564(.A(G1976), .ZN(new_n990));
  AOI21_X1  g565(.A(KEYINPUT52), .B1(G288), .B2(new_n990), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n981), .A2(new_n989), .A3(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(KEYINPUT108), .B1(new_n976), .B2(G8), .ZN(new_n993));
  INV_X1    g568(.A(new_n980), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n989), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(KEYINPUT52), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n988), .A2(new_n992), .A3(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(KEYINPUT115), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT115), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n988), .A2(new_n992), .A3(new_n996), .A4(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n967), .B1(new_n998), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT53), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n1002), .B1(new_n957), .B2(G2078), .ZN(new_n1003));
  INV_X1    g578(.A(G1961), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n948), .A2(new_n1004), .ZN(new_n1005));
  AND2_X1   g580(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n508), .A2(new_n512), .A3(new_n905), .A4(new_n907), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT45), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n906), .A2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1007), .A2(new_n1009), .A3(new_n945), .ZN(new_n1010));
  OR3_X1    g585(.A1(new_n1010), .A2(new_n1002), .A3(G2078), .ZN(new_n1011));
  AOI21_X1  g586(.A(G301), .B1(new_n1006), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1010), .A2(new_n754), .ZN(new_n1013));
  INV_X1    g588(.A(G2084), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n944), .A2(new_n1014), .A3(new_n945), .A4(new_n947), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(G8), .ZN(new_n1017));
  NAND2_X1  g592(.A1(G286), .A2(G8), .ZN(new_n1018));
  AOI21_X1  g593(.A(KEYINPUT51), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n955), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT51), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1018), .ZN(new_n1022));
  NOR3_X1   g597(.A1(new_n1020), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1019), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT123), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1025), .B1(new_n1016), .B2(new_n1022), .ZN(new_n1026));
  AOI211_X1 g601(.A(KEYINPUT123), .B(new_n1018), .C1(new_n1013), .C2(new_n1015), .ZN(new_n1027));
  OR2_X1    g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(KEYINPUT62), .B1(new_n1024), .B2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1017), .A2(KEYINPUT51), .A3(new_n1018), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1021), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT62), .ZN(new_n1034));
  NOR3_X1   g609(.A1(new_n1032), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  OAI211_X1 g610(.A(new_n1001), .B(new_n1012), .C1(new_n1029), .C2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n988), .A2(new_n990), .A3(new_n706), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(new_n983), .ZN(new_n1038));
  XNOR2_X1  g613(.A(new_n981), .B(KEYINPUT112), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1038), .A2(new_n1040), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n997), .A2(new_n954), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1041), .A2(new_n1043), .A3(KEYINPUT113), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT113), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1039), .B1(new_n983), .B2(new_n1037), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1045), .B1(new_n1046), .B2(new_n1042), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1044), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1036), .A2(new_n1048), .ZN(new_n1049));
  AND2_X1   g624(.A1(new_n954), .A2(KEYINPUT63), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1017), .A2(G286), .ZN(new_n1051));
  INV_X1    g626(.A(new_n997), .ZN(new_n1052));
  OAI21_X1  g627(.A(G8), .B1(new_n953), .B2(new_n949), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(new_n941), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1050), .A2(new_n1051), .A3(new_n1052), .A4(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n998), .A2(new_n1000), .ZN(new_n1056));
  INV_X1    g631(.A(new_n967), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1056), .A2(new_n1057), .A3(new_n1051), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(KEYINPUT116), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT116), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1001), .A2(new_n1060), .A3(new_n1051), .ZN(new_n1061));
  XNOR2_X1  g636(.A(KEYINPUT117), .B(KEYINPUT63), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1059), .A2(new_n1061), .A3(new_n1062), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1049), .B1(new_n1055), .B2(new_n1063), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1002), .A2(G2078), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n950), .A2(new_n909), .A3(new_n945), .A4(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1003), .A2(new_n1005), .A3(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(KEYINPUT124), .B1(new_n1067), .B2(G171), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT54), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1006), .A2(new_n1011), .A3(G301), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1067), .A2(KEYINPUT124), .A3(G171), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1070), .A2(new_n1071), .A3(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1024), .A2(new_n1028), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1067), .A2(G171), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1069), .B1(new_n1012), .B2(new_n1075), .ZN(new_n1076));
  AND4_X1   g651(.A1(new_n1001), .A2(new_n1073), .A3(new_n1074), .A4(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n961), .A2(new_n962), .A3(new_n964), .ZN(new_n1078));
  INV_X1    g653(.A(G1956), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  XNOR2_X1  g655(.A(KEYINPUT118), .B(KEYINPUT57), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1081), .B1(new_n605), .B2(new_n606), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT119), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(G299), .A2(KEYINPUT119), .A3(new_n1081), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n607), .A2(KEYINPUT57), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1084), .A2(new_n1085), .A3(new_n1086), .ZN(new_n1087));
  XNOR2_X1  g662(.A(KEYINPUT56), .B(G2072), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n952), .A2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1080), .A2(new_n1087), .A3(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(KEYINPUT120), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1080), .A2(new_n1089), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1087), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT120), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1080), .A2(new_n1089), .A3(new_n1095), .A4(new_n1087), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1091), .A2(new_n1094), .A3(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT61), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT122), .ZN(new_n1100));
  AOI22_X1  g675(.A1(new_n1079), .A2(new_n1078), .B1(new_n952), .B2(new_n1088), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1098), .B1(new_n1101), .B2(new_n1087), .ZN(new_n1102));
  XOR2_X1   g677(.A(KEYINPUT58), .B(G1341), .Z(new_n1103));
  AND2_X1   g678(.A1(new_n976), .A2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1104), .B1(new_n952), .B2(new_n916), .ZN(new_n1105));
  OAI21_X1  g680(.A(KEYINPUT59), .B1(new_n1105), .B2(new_n613), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT59), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n957), .A2(G1996), .ZN(new_n1108));
  OAI211_X1 g683(.A(new_n1107), .B(new_n563), .C1(new_n1108), .C2(new_n1104), .ZN(new_n1109));
  AOI22_X1  g684(.A1(new_n1102), .A2(new_n1094), .B1(new_n1106), .B2(new_n1109), .ZN(new_n1110));
  AND3_X1   g685(.A1(new_n1099), .A2(new_n1100), .A3(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1100), .B1(new_n1099), .B2(new_n1110), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n976), .A2(G2067), .ZN(new_n1113));
  INV_X1    g688(.A(G1348), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1113), .B1(new_n948), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT121), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  AOI211_X1 g692(.A(KEYINPUT121), .B(new_n1113), .C1(new_n948), .C2(new_n1114), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT60), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n601), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  OAI211_X1 g696(.A(KEYINPUT60), .B(new_n600), .C1(new_n1117), .C2(new_n1118), .ZN(new_n1122));
  AOI22_X1  g697(.A1(new_n1121), .A2(new_n1122), .B1(new_n1120), .B2(new_n1119), .ZN(new_n1123));
  NOR3_X1   g698(.A1(new_n1111), .A2(new_n1112), .A3(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1091), .A2(new_n1096), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1119), .A2(new_n601), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1125), .B1(new_n1126), .B2(new_n1094), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1077), .B1(new_n1124), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1064), .A2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n930), .B1(G1986), .B2(G290), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n913), .B1(new_n1130), .B2(new_n932), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1131), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n936), .B1(new_n1129), .B2(new_n1132), .ZN(new_n1133));
  AOI211_X1 g708(.A(KEYINPUT125), .B(new_n1131), .C1(new_n1064), .C2(new_n1128), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n935), .B1(new_n1133), .B2(new_n1134), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g710(.A1(G401), .A2(G227), .ZN(new_n1137));
  AND2_X1   g711(.A1(new_n857), .A2(new_n1137), .ZN(new_n1138));
  NOR2_X1   g712(.A1(G229), .A2(new_n463), .ZN(new_n1139));
  INV_X1    g713(.A(new_n1139), .ZN(new_n1140));
  AOI21_X1  g714(.A(new_n1140), .B1(new_n901), .B2(new_n902), .ZN(new_n1141));
  NAND3_X1  g715(.A1(new_n1138), .A2(new_n1141), .A3(KEYINPUT126), .ZN(new_n1142));
  INV_X1    g716(.A(new_n1142), .ZN(new_n1143));
  AOI21_X1  g717(.A(KEYINPUT126), .B1(new_n1138), .B2(new_n1141), .ZN(new_n1144));
  NOR2_X1   g718(.A1(new_n1143), .A2(new_n1144), .ZN(G308));
  INV_X1    g719(.A(new_n1144), .ZN(new_n1146));
  NAND2_X1  g720(.A1(new_n1146), .A2(new_n1142), .ZN(G225));
endmodule


