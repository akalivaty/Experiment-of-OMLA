

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U553 ( .A1(G651), .A2(n636), .ZN(n641) );
  NOR2_X4 U554 ( .A1(n538), .A2(G2105), .ZN(n547) );
  XOR2_X1 U555 ( .A(KEYINPUT1), .B(n521), .Z(n645) );
  NOR2_X1 U556 ( .A1(n749), .A2(n748), .ZN(n751) );
  AND2_X1 U557 ( .A1(n762), .A2(n731), .ZN(n730) );
  NOR2_X2 U558 ( .A1(n636), .A2(n526), .ZN(n639) );
  XNOR2_X1 U559 ( .A(KEYINPUT23), .B(KEYINPUT65), .ZN(n548) );
  INV_X1 U560 ( .A(n981), .ZN(n758) );
  NOR2_X1 U561 ( .A1(n781), .A2(n780), .ZN(n782) );
  XOR2_X1 U562 ( .A(G543), .B(KEYINPUT0), .Z(n636) );
  XNOR2_X1 U563 ( .A(n549), .B(n548), .ZN(n550) );
  AND2_X1 U564 ( .A1(G137), .A2(n545), .ZN(n518) );
  NOR2_X1 U565 ( .A1(n820), .A2(n813), .ZN(n519) );
  NOR2_X1 U566 ( .A1(n759), .A2(n758), .ZN(n520) );
  INV_X1 U567 ( .A(n779), .ZN(n752) );
  OR2_X1 U568 ( .A1(n709), .A2(n708), .ZN(n710) );
  INV_X1 U569 ( .A(KEYINPUT94), .ZN(n712) );
  XNOR2_X1 U570 ( .A(n713), .B(n712), .ZN(n720) );
  INV_X1 U571 ( .A(KEYINPUT29), .ZN(n726) );
  INV_X1 U572 ( .A(KEYINPUT31), .ZN(n690) );
  XNOR2_X1 U573 ( .A(n691), .B(n690), .ZN(n762) );
  INV_X1 U574 ( .A(KEYINPUT96), .ZN(n750) );
  NOR2_X1 U575 ( .A1(n761), .A2(n766), .ZN(n769) );
  INV_X1 U576 ( .A(n824), .ZN(n813) );
  XNOR2_X1 U577 ( .A(n681), .B(KEYINPUT86), .ZN(n783) );
  XNOR2_X1 U578 ( .A(n527), .B(KEYINPUT74), .ZN(n528) );
  NOR2_X1 U579 ( .A1(G2105), .A2(G2104), .ZN(n535) );
  NOR2_X1 U580 ( .A1(G164), .A2(G1384), .ZN(n784) );
  INV_X1 U581 ( .A(G2104), .ZN(n538) );
  AND2_X1 U582 ( .A1(n814), .A2(n519), .ZN(n816) );
  BUF_X1 U583 ( .A(n545), .Z(n897) );
  XOR2_X1 U584 ( .A(KEYINPUT15), .B(n585), .Z(n991) );
  NOR2_X1 U585 ( .A1(n532), .A2(n531), .ZN(n533) );
  AND2_X1 U586 ( .A1(n551), .A2(n550), .ZN(n552) );
  XOR2_X1 U587 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U588 ( .A1(G51), .A2(n641), .ZN(n523) );
  INV_X1 U589 ( .A(G651), .ZN(n526) );
  NOR2_X1 U590 ( .A1(G543), .A2(n526), .ZN(n521) );
  NAND2_X1 U591 ( .A1(G63), .A2(n645), .ZN(n522) );
  NAND2_X1 U592 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U593 ( .A(KEYINPUT6), .B(n524), .ZN(n532) );
  NOR2_X1 U594 ( .A1(G651), .A2(G543), .ZN(n642) );
  NAND2_X1 U595 ( .A1(n642), .A2(G89), .ZN(n525) );
  XNOR2_X1 U596 ( .A(KEYINPUT4), .B(n525), .ZN(n529) );
  NAND2_X1 U597 ( .A1(n639), .A2(G76), .ZN(n527) );
  NAND2_X1 U598 ( .A1(n529), .A2(n528), .ZN(n530) );
  XOR2_X1 U599 ( .A(n530), .B(KEYINPUT5), .Z(n531) );
  XOR2_X1 U600 ( .A(KEYINPUT75), .B(n533), .Z(n534) );
  XOR2_X1 U601 ( .A(KEYINPUT7), .B(n534), .Z(G168) );
  XOR2_X1 U602 ( .A(KEYINPUT17), .B(n535), .Z(n545) );
  NAND2_X1 U603 ( .A1(G138), .A2(n897), .ZN(n537) );
  NAND2_X1 U604 ( .A1(G102), .A2(n547), .ZN(n536) );
  NAND2_X1 U605 ( .A1(n537), .A2(n536), .ZN(n542) );
  AND2_X2 U606 ( .A1(n538), .A2(G2105), .ZN(n892) );
  NAND2_X1 U607 ( .A1(G126), .A2(n892), .ZN(n540) );
  AND2_X1 U608 ( .A1(G2105), .A2(G2104), .ZN(n893) );
  NAND2_X1 U609 ( .A1(G114), .A2(n893), .ZN(n539) );
  NAND2_X1 U610 ( .A1(n540), .A2(n539), .ZN(n541) );
  NOR2_X1 U611 ( .A1(n542), .A2(n541), .ZN(G164) );
  NAND2_X1 U612 ( .A1(G125), .A2(n892), .ZN(n544) );
  NAND2_X1 U613 ( .A1(G113), .A2(n893), .ZN(n543) );
  NAND2_X1 U614 ( .A1(n544), .A2(n543), .ZN(n546) );
  NOR2_X1 U615 ( .A1(n546), .A2(n518), .ZN(n551) );
  NAND2_X1 U616 ( .A1(G101), .A2(n547), .ZN(n549) );
  XNOR2_X1 U617 ( .A(n552), .B(KEYINPUT64), .ZN(n680) );
  BUF_X1 U618 ( .A(n680), .Z(G160) );
  NAND2_X1 U619 ( .A1(G52), .A2(n641), .ZN(n554) );
  NAND2_X1 U620 ( .A1(G64), .A2(n645), .ZN(n553) );
  NAND2_X1 U621 ( .A1(n554), .A2(n553), .ZN(n560) );
  NAND2_X1 U622 ( .A1(G77), .A2(n639), .ZN(n556) );
  NAND2_X1 U623 ( .A1(G90), .A2(n642), .ZN(n555) );
  NAND2_X1 U624 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U625 ( .A(KEYINPUT69), .B(n557), .ZN(n558) );
  XNOR2_X1 U626 ( .A(KEYINPUT9), .B(n558), .ZN(n559) );
  NOR2_X1 U627 ( .A1(n560), .A2(n559), .ZN(G171) );
  INV_X1 U628 ( .A(G57), .ZN(G237) );
  NAND2_X1 U629 ( .A1(G75), .A2(n639), .ZN(n562) );
  NAND2_X1 U630 ( .A1(G88), .A2(n642), .ZN(n561) );
  NAND2_X1 U631 ( .A1(n562), .A2(n561), .ZN(n566) );
  NAND2_X1 U632 ( .A1(G50), .A2(n641), .ZN(n564) );
  NAND2_X1 U633 ( .A1(G62), .A2(n645), .ZN(n563) );
  NAND2_X1 U634 ( .A1(n564), .A2(n563), .ZN(n565) );
  NOR2_X1 U635 ( .A1(n566), .A2(n565), .ZN(G166) );
  NAND2_X1 U636 ( .A1(G94), .A2(G452), .ZN(n567) );
  XOR2_X1 U637 ( .A(KEYINPUT70), .B(n567), .Z(G173) );
  NAND2_X1 U638 ( .A1(G7), .A2(G661), .ZN(n568) );
  XNOR2_X1 U639 ( .A(n568), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U640 ( .A(G223), .ZN(n844) );
  NAND2_X1 U641 ( .A1(n844), .A2(G567), .ZN(n569) );
  XOR2_X1 U642 ( .A(KEYINPUT11), .B(n569), .Z(G234) );
  NAND2_X1 U643 ( .A1(G56), .A2(n645), .ZN(n570) );
  XOR2_X1 U644 ( .A(KEYINPUT14), .B(n570), .Z(n576) );
  NAND2_X1 U645 ( .A1(n642), .A2(G81), .ZN(n571) );
  XNOR2_X1 U646 ( .A(n571), .B(KEYINPUT12), .ZN(n573) );
  NAND2_X1 U647 ( .A1(G68), .A2(n639), .ZN(n572) );
  NAND2_X1 U648 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U649 ( .A(KEYINPUT13), .B(n574), .Z(n575) );
  NOR2_X1 U650 ( .A1(n576), .A2(n575), .ZN(n578) );
  NAND2_X1 U651 ( .A1(n641), .A2(G43), .ZN(n577) );
  NAND2_X1 U652 ( .A1(n578), .A2(n577), .ZN(n994) );
  INV_X1 U653 ( .A(G860), .ZN(n598) );
  OR2_X1 U654 ( .A1(n994), .A2(n598), .ZN(G153) );
  XNOR2_X1 U655 ( .A(G171), .B(KEYINPUT73), .ZN(G301) );
  NAND2_X1 U656 ( .A1(G868), .A2(G301), .ZN(n587) );
  NAND2_X1 U657 ( .A1(G66), .A2(n645), .ZN(n580) );
  NAND2_X1 U658 ( .A1(G92), .A2(n642), .ZN(n579) );
  NAND2_X1 U659 ( .A1(n580), .A2(n579), .ZN(n584) );
  NAND2_X1 U660 ( .A1(G79), .A2(n639), .ZN(n582) );
  NAND2_X1 U661 ( .A1(G54), .A2(n641), .ZN(n581) );
  NAND2_X1 U662 ( .A1(n582), .A2(n581), .ZN(n583) );
  NOR2_X1 U663 ( .A1(n584), .A2(n583), .ZN(n585) );
  INV_X1 U664 ( .A(n991), .ZN(n708) );
  INV_X1 U665 ( .A(G868), .ZN(n660) );
  NAND2_X1 U666 ( .A1(n708), .A2(n660), .ZN(n586) );
  NAND2_X1 U667 ( .A1(n587), .A2(n586), .ZN(G284) );
  NAND2_X1 U668 ( .A1(n645), .A2(G65), .ZN(n588) );
  XOR2_X1 U669 ( .A(KEYINPUT71), .B(n588), .Z(n590) );
  NAND2_X1 U670 ( .A1(n641), .A2(G53), .ZN(n589) );
  NAND2_X1 U671 ( .A1(n590), .A2(n589), .ZN(n591) );
  XOR2_X1 U672 ( .A(KEYINPUT72), .B(n591), .Z(n595) );
  NAND2_X1 U673 ( .A1(n639), .A2(G78), .ZN(n593) );
  NAND2_X1 U674 ( .A1(G91), .A2(n642), .ZN(n592) );
  AND2_X1 U675 ( .A1(n593), .A2(n592), .ZN(n594) );
  NAND2_X1 U676 ( .A1(n595), .A2(n594), .ZN(G299) );
  NOR2_X1 U677 ( .A1(G286), .A2(n660), .ZN(n597) );
  NOR2_X1 U678 ( .A1(G868), .A2(G299), .ZN(n596) );
  NOR2_X1 U679 ( .A1(n597), .A2(n596), .ZN(G297) );
  NAND2_X1 U680 ( .A1(n598), .A2(G559), .ZN(n599) );
  NAND2_X1 U681 ( .A1(n599), .A2(n991), .ZN(n600) );
  XNOR2_X1 U682 ( .A(n600), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U683 ( .A1(G868), .A2(n994), .ZN(n603) );
  NAND2_X1 U684 ( .A1(n991), .A2(G868), .ZN(n601) );
  NOR2_X1 U685 ( .A1(G559), .A2(n601), .ZN(n602) );
  NOR2_X1 U686 ( .A1(n603), .A2(n602), .ZN(G282) );
  NAND2_X1 U687 ( .A1(G123), .A2(n892), .ZN(n604) );
  XNOR2_X1 U688 ( .A(n604), .B(KEYINPUT76), .ZN(n605) );
  XNOR2_X1 U689 ( .A(n605), .B(KEYINPUT18), .ZN(n607) );
  NAND2_X1 U690 ( .A1(G111), .A2(n893), .ZN(n606) );
  NAND2_X1 U691 ( .A1(n607), .A2(n606), .ZN(n611) );
  NAND2_X1 U692 ( .A1(G135), .A2(n897), .ZN(n609) );
  NAND2_X1 U693 ( .A1(G99), .A2(n547), .ZN(n608) );
  NAND2_X1 U694 ( .A1(n609), .A2(n608), .ZN(n610) );
  NOR2_X1 U695 ( .A1(n611), .A2(n610), .ZN(n933) );
  XNOR2_X1 U696 ( .A(n933), .B(G2096), .ZN(n613) );
  INV_X1 U697 ( .A(G2100), .ZN(n612) );
  NAND2_X1 U698 ( .A1(n613), .A2(n612), .ZN(G156) );
  NAND2_X1 U699 ( .A1(G80), .A2(n639), .ZN(n615) );
  NAND2_X1 U700 ( .A1(G93), .A2(n642), .ZN(n614) );
  NAND2_X1 U701 ( .A1(n615), .A2(n614), .ZN(n616) );
  XNOR2_X1 U702 ( .A(KEYINPUT78), .B(n616), .ZN(n620) );
  NAND2_X1 U703 ( .A1(G55), .A2(n641), .ZN(n618) );
  NAND2_X1 U704 ( .A1(G67), .A2(n645), .ZN(n617) );
  NAND2_X1 U705 ( .A1(n618), .A2(n617), .ZN(n619) );
  OR2_X1 U706 ( .A1(n620), .A2(n619), .ZN(n659) );
  NAND2_X1 U707 ( .A1(G559), .A2(n991), .ZN(n621) );
  XNOR2_X1 U708 ( .A(n621), .B(n994), .ZN(n656) );
  XOR2_X1 U709 ( .A(KEYINPUT77), .B(n656), .Z(n622) );
  NOR2_X1 U710 ( .A1(G860), .A2(n622), .ZN(n623) );
  XOR2_X1 U711 ( .A(n659), .B(n623), .Z(G145) );
  NAND2_X1 U712 ( .A1(n642), .A2(G85), .ZN(n631) );
  NAND2_X1 U713 ( .A1(G72), .A2(n639), .ZN(n624) );
  XNOR2_X1 U714 ( .A(n624), .B(KEYINPUT66), .ZN(n626) );
  NAND2_X1 U715 ( .A1(n645), .A2(G60), .ZN(n625) );
  NAND2_X1 U716 ( .A1(n626), .A2(n625), .ZN(n629) );
  NAND2_X1 U717 ( .A1(G47), .A2(n641), .ZN(n627) );
  XNOR2_X1 U718 ( .A(KEYINPUT67), .B(n627), .ZN(n628) );
  NOR2_X1 U719 ( .A1(n629), .A2(n628), .ZN(n630) );
  NAND2_X1 U720 ( .A1(n631), .A2(n630), .ZN(n632) );
  XNOR2_X1 U721 ( .A(n632), .B(KEYINPUT68), .ZN(G290) );
  NAND2_X1 U722 ( .A1(G49), .A2(n641), .ZN(n634) );
  NAND2_X1 U723 ( .A1(G74), .A2(G651), .ZN(n633) );
  NAND2_X1 U724 ( .A1(n634), .A2(n633), .ZN(n635) );
  NOR2_X1 U725 ( .A1(n645), .A2(n635), .ZN(n638) );
  NAND2_X1 U726 ( .A1(n636), .A2(G87), .ZN(n637) );
  NAND2_X1 U727 ( .A1(n638), .A2(n637), .ZN(G288) );
  NAND2_X1 U728 ( .A1(G73), .A2(n639), .ZN(n640) );
  XNOR2_X1 U729 ( .A(n640), .B(KEYINPUT2), .ZN(n650) );
  NAND2_X1 U730 ( .A1(G48), .A2(n641), .ZN(n644) );
  NAND2_X1 U731 ( .A1(G86), .A2(n642), .ZN(n643) );
  NAND2_X1 U732 ( .A1(n644), .A2(n643), .ZN(n648) );
  NAND2_X1 U733 ( .A1(G61), .A2(n645), .ZN(n646) );
  XNOR2_X1 U734 ( .A(KEYINPUT79), .B(n646), .ZN(n647) );
  NOR2_X1 U735 ( .A1(n648), .A2(n647), .ZN(n649) );
  NAND2_X1 U736 ( .A1(n650), .A2(n649), .ZN(G305) );
  XNOR2_X1 U737 ( .A(KEYINPUT19), .B(n659), .ZN(n652) );
  INV_X1 U738 ( .A(G299), .ZN(n721) );
  XNOR2_X1 U739 ( .A(G166), .B(n721), .ZN(n651) );
  XNOR2_X1 U740 ( .A(n652), .B(n651), .ZN(n653) );
  XOR2_X1 U741 ( .A(n653), .B(G305), .Z(n654) );
  XNOR2_X1 U742 ( .A(G288), .B(n654), .ZN(n655) );
  XNOR2_X1 U743 ( .A(G290), .B(n655), .ZN(n919) );
  XNOR2_X1 U744 ( .A(KEYINPUT80), .B(n656), .ZN(n657) );
  XNOR2_X1 U745 ( .A(n919), .B(n657), .ZN(n658) );
  NAND2_X1 U746 ( .A1(n658), .A2(G868), .ZN(n662) );
  NAND2_X1 U747 ( .A1(n660), .A2(n659), .ZN(n661) );
  NAND2_X1 U748 ( .A1(n662), .A2(n661), .ZN(G295) );
  NAND2_X1 U749 ( .A1(G2084), .A2(G2078), .ZN(n663) );
  XNOR2_X1 U750 ( .A(n663), .B(KEYINPUT20), .ZN(n664) );
  XNOR2_X1 U751 ( .A(KEYINPUT81), .B(n664), .ZN(n665) );
  NAND2_X1 U752 ( .A1(n665), .A2(G2090), .ZN(n666) );
  XNOR2_X1 U753 ( .A(KEYINPUT21), .B(n666), .ZN(n667) );
  NAND2_X1 U754 ( .A1(n667), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U755 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U756 ( .A1(G483), .A2(G661), .ZN(n677) );
  NAND2_X1 U757 ( .A1(G69), .A2(G120), .ZN(n668) );
  NOR2_X1 U758 ( .A1(G237), .A2(n668), .ZN(n669) );
  NAND2_X1 U759 ( .A1(G108), .A2(n669), .ZN(n849) );
  NAND2_X1 U760 ( .A1(G567), .A2(n849), .ZN(n670) );
  XOR2_X1 U761 ( .A(KEYINPUT83), .B(n670), .Z(n676) );
  NAND2_X1 U762 ( .A1(G132), .A2(G82), .ZN(n671) );
  XNOR2_X1 U763 ( .A(n671), .B(KEYINPUT82), .ZN(n672) );
  XNOR2_X1 U764 ( .A(n672), .B(KEYINPUT22), .ZN(n673) );
  NOR2_X1 U765 ( .A1(G218), .A2(n673), .ZN(n674) );
  NAND2_X1 U766 ( .A1(G96), .A2(n674), .ZN(n850) );
  NAND2_X1 U767 ( .A1(G2106), .A2(n850), .ZN(n675) );
  NAND2_X1 U768 ( .A1(n676), .A2(n675), .ZN(n851) );
  NOR2_X1 U769 ( .A1(n677), .A2(n851), .ZN(n678) );
  XNOR2_X1 U770 ( .A(n678), .B(KEYINPUT84), .ZN(n847) );
  NAND2_X1 U771 ( .A1(n847), .A2(G36), .ZN(n679) );
  XOR2_X1 U772 ( .A(KEYINPUT85), .B(n679), .Z(G176) );
  INV_X1 U773 ( .A(G166), .ZN(G303) );
  NAND2_X1 U774 ( .A1(n680), .A2(G40), .ZN(n681) );
  INV_X1 U775 ( .A(n784), .ZN(n682) );
  NOR2_X2 U776 ( .A1(n783), .A2(n682), .ZN(n697) );
  INV_X2 U777 ( .A(n697), .ZN(n714) );
  NAND2_X2 U778 ( .A1(n714), .A2(G8), .ZN(n779) );
  NOR2_X1 U779 ( .A1(G1966), .A2(n779), .ZN(n740) );
  NOR2_X1 U780 ( .A1(G2084), .A2(n714), .ZN(n739) );
  NOR2_X1 U781 ( .A1(n740), .A2(n739), .ZN(n683) );
  NAND2_X1 U782 ( .A1(n683), .A2(G8), .ZN(n684) );
  XNOR2_X1 U783 ( .A(n684), .B(KEYINPUT30), .ZN(n685) );
  NOR2_X1 U784 ( .A1(G168), .A2(n685), .ZN(n689) );
  XNOR2_X1 U785 ( .A(G2078), .B(KEYINPUT25), .ZN(n956) );
  NOR2_X1 U786 ( .A1(n714), .A2(n956), .ZN(n687) );
  AND2_X1 U787 ( .A1(n714), .A2(G1961), .ZN(n686) );
  NOR2_X1 U788 ( .A1(n687), .A2(n686), .ZN(n696) );
  NOR2_X1 U789 ( .A1(G171), .A2(n696), .ZN(n688) );
  NOR2_X1 U790 ( .A1(n689), .A2(n688), .ZN(n691) );
  NOR2_X1 U791 ( .A1(G1971), .A2(n779), .ZN(n693) );
  NOR2_X1 U792 ( .A1(G2090), .A2(n714), .ZN(n692) );
  NOR2_X1 U793 ( .A1(n693), .A2(n692), .ZN(n694) );
  NAND2_X1 U794 ( .A1(n694), .A2(G303), .ZN(n695) );
  XOR2_X1 U795 ( .A(KEYINPUT95), .B(n695), .Z(n731) );
  NAND2_X1 U796 ( .A1(G171), .A2(n696), .ZN(n729) );
  AND2_X1 U797 ( .A1(n697), .A2(G1996), .ZN(n698) );
  XNOR2_X1 U798 ( .A(n698), .B(KEYINPUT26), .ZN(n702) );
  NAND2_X1 U799 ( .A1(n714), .A2(G1341), .ZN(n700) );
  INV_X1 U800 ( .A(n994), .ZN(n699) );
  NAND2_X1 U801 ( .A1(n700), .A2(n699), .ZN(n701) );
  NOR2_X1 U802 ( .A1(n702), .A2(n701), .ZN(n707) );
  INV_X1 U803 ( .A(G2067), .ZN(n703) );
  AND2_X1 U804 ( .A1(n703), .A2(n697), .ZN(n705) );
  NOR2_X1 U805 ( .A1(n697), .A2(G1348), .ZN(n704) );
  NOR2_X1 U806 ( .A1(n705), .A2(n704), .ZN(n709) );
  NAND2_X1 U807 ( .A1(n708), .A2(n709), .ZN(n706) );
  NAND2_X1 U808 ( .A1(n707), .A2(n706), .ZN(n711) );
  NAND2_X1 U809 ( .A1(n711), .A2(n710), .ZN(n713) );
  NAND2_X1 U810 ( .A1(G1956), .A2(n714), .ZN(n715) );
  XNOR2_X1 U811 ( .A(KEYINPUT93), .B(n715), .ZN(n718) );
  NAND2_X1 U812 ( .A1(n697), .A2(G2072), .ZN(n716) );
  XNOR2_X1 U813 ( .A(KEYINPUT27), .B(n716), .ZN(n717) );
  NOR2_X1 U814 ( .A1(n718), .A2(n717), .ZN(n722) );
  NAND2_X1 U815 ( .A1(n722), .A2(n721), .ZN(n719) );
  NAND2_X1 U816 ( .A1(n720), .A2(n719), .ZN(n725) );
  NOR2_X1 U817 ( .A1(n722), .A2(n721), .ZN(n723) );
  XOR2_X1 U818 ( .A(n723), .B(KEYINPUT28), .Z(n724) );
  NAND2_X1 U819 ( .A1(n725), .A2(n724), .ZN(n727) );
  XNOR2_X1 U820 ( .A(n727), .B(n726), .ZN(n728) );
  NAND2_X1 U821 ( .A1(n729), .A2(n728), .ZN(n763) );
  NAND2_X1 U822 ( .A1(n730), .A2(n763), .ZN(n735) );
  INV_X1 U823 ( .A(n731), .ZN(n732) );
  OR2_X1 U824 ( .A1(n732), .A2(G286), .ZN(n733) );
  AND2_X1 U825 ( .A1(n733), .A2(G8), .ZN(n734) );
  NAND2_X1 U826 ( .A1(n735), .A2(n734), .ZN(n737) );
  INV_X1 U827 ( .A(KEYINPUT32), .ZN(n736) );
  XNOR2_X1 U828 ( .A(n737), .B(n736), .ZN(n761) );
  NAND2_X1 U829 ( .A1(G1976), .A2(G288), .ZN(n984) );
  AND2_X1 U830 ( .A1(n762), .A2(n984), .ZN(n738) );
  AND2_X1 U831 ( .A1(n763), .A2(n738), .ZN(n744) );
  NAND2_X1 U832 ( .A1(G8), .A2(n739), .ZN(n742) );
  INV_X1 U833 ( .A(n740), .ZN(n741) );
  NAND2_X1 U834 ( .A1(n742), .A2(n741), .ZN(n764) );
  AND2_X1 U835 ( .A1(n984), .A2(n764), .ZN(n743) );
  NOR2_X1 U836 ( .A1(n744), .A2(n743), .ZN(n745) );
  NOR2_X1 U837 ( .A1(n761), .A2(n745), .ZN(n749) );
  INV_X1 U838 ( .A(n984), .ZN(n747) );
  NOR2_X1 U839 ( .A1(G1976), .A2(G288), .ZN(n756) );
  NOR2_X1 U840 ( .A1(G1971), .A2(G303), .ZN(n746) );
  NOR2_X1 U841 ( .A1(n756), .A2(n746), .ZN(n985) );
  NOR2_X1 U842 ( .A1(n747), .A2(n985), .ZN(n748) );
  XNOR2_X1 U843 ( .A(n751), .B(n750), .ZN(n753) );
  NAND2_X1 U844 ( .A1(n753), .A2(n752), .ZN(n755) );
  INV_X1 U845 ( .A(KEYINPUT33), .ZN(n754) );
  NAND2_X1 U846 ( .A1(n755), .A2(n754), .ZN(n760) );
  NAND2_X1 U847 ( .A1(n756), .A2(KEYINPUT33), .ZN(n757) );
  NOR2_X1 U848 ( .A1(n757), .A2(n779), .ZN(n759) );
  XOR2_X1 U849 ( .A(G1981), .B(G305), .Z(n981) );
  NAND2_X1 U850 ( .A1(n760), .A2(n520), .ZN(n773) );
  AND2_X1 U851 ( .A1(n763), .A2(n762), .ZN(n765) );
  NOR2_X1 U852 ( .A1(n765), .A2(n764), .ZN(n766) );
  NAND2_X1 U853 ( .A1(G166), .A2(G8), .ZN(n767) );
  NOR2_X1 U854 ( .A1(G2090), .A2(n767), .ZN(n768) );
  NOR2_X1 U855 ( .A1(n769), .A2(n768), .ZN(n770) );
  NOR2_X1 U856 ( .A1(n752), .A2(n770), .ZN(n771) );
  XNOR2_X1 U857 ( .A(n771), .B(KEYINPUT97), .ZN(n772) );
  NAND2_X1 U858 ( .A1(n773), .A2(n772), .ZN(n774) );
  XNOR2_X1 U859 ( .A(n774), .B(KEYINPUT98), .ZN(n781) );
  NOR2_X1 U860 ( .A1(G1981), .A2(G305), .ZN(n777) );
  XNOR2_X1 U861 ( .A(KEYINPUT24), .B(KEYINPUT92), .ZN(n775) );
  XNOR2_X1 U862 ( .A(n775), .B(KEYINPUT91), .ZN(n776) );
  XNOR2_X1 U863 ( .A(n777), .B(n776), .ZN(n778) );
  NOR2_X1 U864 ( .A1(n779), .A2(n778), .ZN(n780) );
  XNOR2_X1 U865 ( .A(n782), .B(KEYINPUT99), .ZN(n814) );
  NOR2_X1 U866 ( .A1(n783), .A2(n784), .ZN(n829) );
  INV_X1 U867 ( .A(n829), .ZN(n802) );
  XOR2_X1 U868 ( .A(KEYINPUT88), .B(KEYINPUT38), .Z(n786) );
  NAND2_X1 U869 ( .A1(G105), .A2(n547), .ZN(n785) );
  XNOR2_X1 U870 ( .A(n786), .B(n785), .ZN(n790) );
  NAND2_X1 U871 ( .A1(G141), .A2(n897), .ZN(n788) );
  NAND2_X1 U872 ( .A1(G129), .A2(n892), .ZN(n787) );
  NAND2_X1 U873 ( .A1(n788), .A2(n787), .ZN(n789) );
  NOR2_X1 U874 ( .A1(n790), .A2(n789), .ZN(n792) );
  NAND2_X1 U875 ( .A1(n893), .A2(G117), .ZN(n791) );
  NAND2_X1 U876 ( .A1(n792), .A2(n791), .ZN(n911) );
  NAND2_X1 U877 ( .A1(G1996), .A2(n911), .ZN(n793) );
  XNOR2_X1 U878 ( .A(n793), .B(KEYINPUT89), .ZN(n801) );
  XNOR2_X1 U879 ( .A(KEYINPUT87), .B(G1991), .ZN(n967) );
  NAND2_X1 U880 ( .A1(G131), .A2(n897), .ZN(n795) );
  NAND2_X1 U881 ( .A1(G95), .A2(n547), .ZN(n794) );
  NAND2_X1 U882 ( .A1(n795), .A2(n794), .ZN(n799) );
  NAND2_X1 U883 ( .A1(G119), .A2(n892), .ZN(n797) );
  NAND2_X1 U884 ( .A1(G107), .A2(n893), .ZN(n796) );
  NAND2_X1 U885 ( .A1(n797), .A2(n796), .ZN(n798) );
  NOR2_X1 U886 ( .A1(n799), .A2(n798), .ZN(n891) );
  NOR2_X1 U887 ( .A1(n967), .A2(n891), .ZN(n800) );
  NOR2_X1 U888 ( .A1(n801), .A2(n800), .ZN(n935) );
  NOR2_X1 U889 ( .A1(n802), .A2(n935), .ZN(n803) );
  XNOR2_X1 U890 ( .A(n803), .B(KEYINPUT90), .ZN(n820) );
  XNOR2_X1 U891 ( .A(G2067), .B(KEYINPUT37), .ZN(n817) );
  NAND2_X1 U892 ( .A1(G128), .A2(n892), .ZN(n805) );
  NAND2_X1 U893 ( .A1(G116), .A2(n893), .ZN(n804) );
  NAND2_X1 U894 ( .A1(n805), .A2(n804), .ZN(n806) );
  XNOR2_X1 U895 ( .A(n806), .B(KEYINPUT35), .ZN(n811) );
  NAND2_X1 U896 ( .A1(G140), .A2(n897), .ZN(n808) );
  NAND2_X1 U897 ( .A1(G104), .A2(n547), .ZN(n807) );
  NAND2_X1 U898 ( .A1(n808), .A2(n807), .ZN(n809) );
  XOR2_X1 U899 ( .A(KEYINPUT34), .B(n809), .Z(n810) );
  NAND2_X1 U900 ( .A1(n811), .A2(n810), .ZN(n812) );
  XOR2_X1 U901 ( .A(n812), .B(KEYINPUT36), .Z(n916) );
  NOR2_X1 U902 ( .A1(n817), .A2(n916), .ZN(n931) );
  NAND2_X1 U903 ( .A1(n829), .A2(n931), .ZN(n824) );
  XNOR2_X1 U904 ( .A(G1986), .B(G290), .ZN(n990) );
  NAND2_X1 U905 ( .A1(n990), .A2(n829), .ZN(n815) );
  NAND2_X1 U906 ( .A1(n816), .A2(n815), .ZN(n832) );
  AND2_X1 U907 ( .A1(n817), .A2(n916), .ZN(n930) );
  NOR2_X1 U908 ( .A1(G1996), .A2(n911), .ZN(n945) );
  AND2_X1 U909 ( .A1(n967), .A2(n891), .ZN(n937) );
  NOR2_X1 U910 ( .A1(G1986), .A2(G290), .ZN(n818) );
  XNOR2_X1 U911 ( .A(KEYINPUT100), .B(n818), .ZN(n819) );
  NOR2_X1 U912 ( .A1(n937), .A2(n819), .ZN(n821) );
  NOR2_X1 U913 ( .A1(n821), .A2(n820), .ZN(n822) );
  NOR2_X1 U914 ( .A1(n945), .A2(n822), .ZN(n823) );
  XNOR2_X1 U915 ( .A(n823), .B(KEYINPUT39), .ZN(n825) );
  NAND2_X1 U916 ( .A1(n825), .A2(n824), .ZN(n826) );
  XNOR2_X1 U917 ( .A(KEYINPUT101), .B(n826), .ZN(n827) );
  NOR2_X1 U918 ( .A1(n930), .A2(n827), .ZN(n828) );
  XOR2_X1 U919 ( .A(KEYINPUT102), .B(n828), .Z(n830) );
  NAND2_X1 U920 ( .A1(n830), .A2(n829), .ZN(n831) );
  NAND2_X1 U921 ( .A1(n832), .A2(n831), .ZN(n833) );
  XNOR2_X1 U922 ( .A(KEYINPUT40), .B(n833), .ZN(G329) );
  XOR2_X1 U923 ( .A(G2430), .B(G2451), .Z(n835) );
  XNOR2_X1 U924 ( .A(G2446), .B(G2427), .ZN(n834) );
  XNOR2_X1 U925 ( .A(n835), .B(n834), .ZN(n842) );
  XOR2_X1 U926 ( .A(G2438), .B(G2435), .Z(n837) );
  XNOR2_X1 U927 ( .A(G2443), .B(KEYINPUT103), .ZN(n836) );
  XNOR2_X1 U928 ( .A(n837), .B(n836), .ZN(n838) );
  XOR2_X1 U929 ( .A(n838), .B(G2454), .Z(n840) );
  XNOR2_X1 U930 ( .A(G1348), .B(G1341), .ZN(n839) );
  XNOR2_X1 U931 ( .A(n840), .B(n839), .ZN(n841) );
  XNOR2_X1 U932 ( .A(n842), .B(n841), .ZN(n843) );
  NAND2_X1 U933 ( .A1(n843), .A2(G14), .ZN(n924) );
  XOR2_X1 U934 ( .A(KEYINPUT104), .B(n924), .Z(G401) );
  NAND2_X1 U935 ( .A1(G2106), .A2(n844), .ZN(G217) );
  AND2_X1 U936 ( .A1(G15), .A2(G2), .ZN(n845) );
  NAND2_X1 U937 ( .A1(G661), .A2(n845), .ZN(G259) );
  NAND2_X1 U938 ( .A1(G3), .A2(G1), .ZN(n846) );
  XOR2_X1 U939 ( .A(KEYINPUT105), .B(n846), .Z(n848) );
  NAND2_X1 U940 ( .A1(n848), .A2(n847), .ZN(G188) );
  INV_X1 U942 ( .A(G132), .ZN(G219) );
  INV_X1 U943 ( .A(G120), .ZN(G236) );
  INV_X1 U944 ( .A(G82), .ZN(G220) );
  INV_X1 U945 ( .A(G69), .ZN(G235) );
  NOR2_X1 U946 ( .A1(n850), .A2(n849), .ZN(G325) );
  INV_X1 U947 ( .A(G325), .ZN(G261) );
  XOR2_X1 U948 ( .A(KEYINPUT106), .B(n851), .Z(G319) );
  XOR2_X1 U949 ( .A(KEYINPUT42), .B(G2090), .Z(n853) );
  XNOR2_X1 U950 ( .A(G2067), .B(G2084), .ZN(n852) );
  XNOR2_X1 U951 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U952 ( .A(n854), .B(G2100), .Z(n856) );
  XNOR2_X1 U953 ( .A(G2078), .B(G2072), .ZN(n855) );
  XNOR2_X1 U954 ( .A(n856), .B(n855), .ZN(n860) );
  XOR2_X1 U955 ( .A(G2096), .B(KEYINPUT43), .Z(n858) );
  XNOR2_X1 U956 ( .A(KEYINPUT107), .B(G2678), .ZN(n857) );
  XNOR2_X1 U957 ( .A(n858), .B(n857), .ZN(n859) );
  XOR2_X1 U958 ( .A(n860), .B(n859), .Z(G227) );
  XOR2_X1 U959 ( .A(G2474), .B(G1956), .Z(n862) );
  XNOR2_X1 U960 ( .A(G1981), .B(G1961), .ZN(n861) );
  XNOR2_X1 U961 ( .A(n862), .B(n861), .ZN(n863) );
  XOR2_X1 U962 ( .A(n863), .B(KEYINPUT108), .Z(n865) );
  XNOR2_X1 U963 ( .A(G1991), .B(G1996), .ZN(n864) );
  XNOR2_X1 U964 ( .A(n865), .B(n864), .ZN(n869) );
  XOR2_X1 U965 ( .A(G1966), .B(G1971), .Z(n867) );
  XNOR2_X1 U966 ( .A(G1986), .B(G1976), .ZN(n866) );
  XNOR2_X1 U967 ( .A(n867), .B(n866), .ZN(n868) );
  XOR2_X1 U968 ( .A(n869), .B(n868), .Z(n871) );
  XNOR2_X1 U969 ( .A(KEYINPUT41), .B(KEYINPUT109), .ZN(n870) );
  XNOR2_X1 U970 ( .A(n871), .B(n870), .ZN(G229) );
  NAND2_X1 U971 ( .A1(G124), .A2(n892), .ZN(n872) );
  XNOR2_X1 U972 ( .A(n872), .B(KEYINPUT110), .ZN(n873) );
  XNOR2_X1 U973 ( .A(n873), .B(KEYINPUT44), .ZN(n875) );
  NAND2_X1 U974 ( .A1(G112), .A2(n893), .ZN(n874) );
  NAND2_X1 U975 ( .A1(n875), .A2(n874), .ZN(n879) );
  NAND2_X1 U976 ( .A1(G136), .A2(n897), .ZN(n877) );
  NAND2_X1 U977 ( .A1(G100), .A2(n547), .ZN(n876) );
  NAND2_X1 U978 ( .A1(n877), .A2(n876), .ZN(n878) );
  NOR2_X1 U979 ( .A1(n879), .A2(n878), .ZN(G162) );
  NAND2_X1 U980 ( .A1(G127), .A2(n892), .ZN(n881) );
  NAND2_X1 U981 ( .A1(G115), .A2(n893), .ZN(n880) );
  NAND2_X1 U982 ( .A1(n881), .A2(n880), .ZN(n882) );
  XNOR2_X1 U983 ( .A(n882), .B(KEYINPUT47), .ZN(n884) );
  NAND2_X1 U984 ( .A1(G103), .A2(n547), .ZN(n883) );
  NAND2_X1 U985 ( .A1(n884), .A2(n883), .ZN(n887) );
  NAND2_X1 U986 ( .A1(G139), .A2(n897), .ZN(n885) );
  XNOR2_X1 U987 ( .A(KEYINPUT113), .B(n885), .ZN(n886) );
  NOR2_X1 U988 ( .A1(n887), .A2(n886), .ZN(n888) );
  XOR2_X1 U989 ( .A(KEYINPUT114), .B(n888), .Z(n940) );
  XOR2_X1 U990 ( .A(G164), .B(n940), .Z(n889) );
  XNOR2_X1 U991 ( .A(G160), .B(n889), .ZN(n890) );
  XNOR2_X1 U992 ( .A(n891), .B(n890), .ZN(n915) );
  NAND2_X1 U993 ( .A1(G130), .A2(n892), .ZN(n895) );
  NAND2_X1 U994 ( .A1(G118), .A2(n893), .ZN(n894) );
  NAND2_X1 U995 ( .A1(n895), .A2(n894), .ZN(n896) );
  XOR2_X1 U996 ( .A(KEYINPUT111), .B(n896), .Z(n903) );
  NAND2_X1 U997 ( .A1(n897), .A2(G142), .ZN(n898) );
  XNOR2_X1 U998 ( .A(n898), .B(KEYINPUT112), .ZN(n900) );
  NAND2_X1 U999 ( .A1(G106), .A2(n547), .ZN(n899) );
  NAND2_X1 U1000 ( .A1(n900), .A2(n899), .ZN(n901) );
  XOR2_X1 U1001 ( .A(KEYINPUT45), .B(n901), .Z(n902) );
  NOR2_X1 U1002 ( .A1(n903), .A2(n902), .ZN(n910) );
  XOR2_X1 U1003 ( .A(KEYINPUT115), .B(KEYINPUT117), .Z(n905) );
  XNOR2_X1 U1004 ( .A(KEYINPUT116), .B(KEYINPUT46), .ZN(n904) );
  XNOR2_X1 U1005 ( .A(n905), .B(n904), .ZN(n906) );
  XOR2_X1 U1006 ( .A(n906), .B(KEYINPUT48), .Z(n908) );
  XNOR2_X1 U1007 ( .A(n933), .B(KEYINPUT118), .ZN(n907) );
  XNOR2_X1 U1008 ( .A(n908), .B(n907), .ZN(n909) );
  XNOR2_X1 U1009 ( .A(n910), .B(n909), .ZN(n913) );
  XNOR2_X1 U1010 ( .A(n911), .B(G162), .ZN(n912) );
  XNOR2_X1 U1011 ( .A(n913), .B(n912), .ZN(n914) );
  XNOR2_X1 U1012 ( .A(n915), .B(n914), .ZN(n917) );
  XOR2_X1 U1013 ( .A(n917), .B(n916), .Z(n918) );
  NOR2_X1 U1014 ( .A1(G37), .A2(n918), .ZN(G395) );
  XOR2_X1 U1015 ( .A(n919), .B(G286), .Z(n921) );
  XNOR2_X1 U1016 ( .A(G171), .B(n991), .ZN(n920) );
  XNOR2_X1 U1017 ( .A(n921), .B(n920), .ZN(n922) );
  XNOR2_X1 U1018 ( .A(n922), .B(n994), .ZN(n923) );
  NOR2_X1 U1019 ( .A1(G37), .A2(n923), .ZN(G397) );
  NAND2_X1 U1020 ( .A1(G319), .A2(n924), .ZN(n927) );
  NOR2_X1 U1021 ( .A1(G227), .A2(G229), .ZN(n925) );
  XNOR2_X1 U1022 ( .A(KEYINPUT49), .B(n925), .ZN(n926) );
  NOR2_X1 U1023 ( .A1(n927), .A2(n926), .ZN(n929) );
  NOR2_X1 U1024 ( .A1(G395), .A2(G397), .ZN(n928) );
  NAND2_X1 U1025 ( .A1(n929), .A2(n928), .ZN(G225) );
  INV_X1 U1026 ( .A(G225), .ZN(G308) );
  INV_X1 U1027 ( .A(G96), .ZN(G221) );
  INV_X1 U1028 ( .A(G108), .ZN(G238) );
  NOR2_X1 U1029 ( .A1(n931), .A2(n930), .ZN(n939) );
  XOR2_X1 U1030 ( .A(G2084), .B(G160), .Z(n932) );
  NOR2_X1 U1031 ( .A1(n933), .A2(n932), .ZN(n934) );
  NAND2_X1 U1032 ( .A1(n935), .A2(n934), .ZN(n936) );
  NOR2_X1 U1033 ( .A1(n937), .A2(n936), .ZN(n938) );
  NAND2_X1 U1034 ( .A1(n939), .A2(n938), .ZN(n950) );
  XOR2_X1 U1035 ( .A(G164), .B(G2078), .Z(n942) );
  XNOR2_X1 U1036 ( .A(G2072), .B(n940), .ZN(n941) );
  NOR2_X1 U1037 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1038 ( .A(KEYINPUT50), .B(n943), .ZN(n948) );
  XOR2_X1 U1039 ( .A(G2090), .B(G162), .Z(n944) );
  NOR2_X1 U1040 ( .A1(n945), .A2(n944), .ZN(n946) );
  XOR2_X1 U1041 ( .A(KEYINPUT51), .B(n946), .Z(n947) );
  NAND2_X1 U1042 ( .A1(n948), .A2(n947), .ZN(n949) );
  NOR2_X1 U1043 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1044 ( .A(KEYINPUT52), .B(n951), .ZN(n952) );
  INV_X1 U1045 ( .A(KEYINPUT55), .ZN(n976) );
  NAND2_X1 U1046 ( .A1(n952), .A2(n976), .ZN(n953) );
  NAND2_X1 U1047 ( .A1(n953), .A2(G29), .ZN(n1035) );
  XNOR2_X1 U1048 ( .A(KEYINPUT54), .B(G34), .ZN(n954) );
  XNOR2_X1 U1049 ( .A(n954), .B(KEYINPUT121), .ZN(n955) );
  XNOR2_X1 U1050 ( .A(G2084), .B(n955), .ZN(n974) );
  XNOR2_X1 U1051 ( .A(G2090), .B(G35), .ZN(n972) );
  XNOR2_X1 U1052 ( .A(n956), .B(G27), .ZN(n959) );
  INV_X1 U1053 ( .A(G1996), .ZN(n957) );
  XNOR2_X1 U1054 ( .A(n957), .B(G32), .ZN(n958) );
  NAND2_X1 U1055 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1056 ( .A(KEYINPUT119), .B(n960), .ZN(n962) );
  XOR2_X1 U1057 ( .A(G2072), .B(G33), .Z(n961) );
  NAND2_X1 U1058 ( .A1(n962), .A2(n961), .ZN(n964) );
  XNOR2_X1 U1059 ( .A(G26), .B(G2067), .ZN(n963) );
  NOR2_X1 U1060 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1061 ( .A(KEYINPUT120), .B(n965), .ZN(n966) );
  NAND2_X1 U1062 ( .A1(n966), .A2(G28), .ZN(n969) );
  XOR2_X1 U1063 ( .A(G25), .B(n967), .Z(n968) );
  NOR2_X1 U1064 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1065 ( .A(KEYINPUT53), .B(n970), .ZN(n971) );
  NOR2_X1 U1066 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1067 ( .A1(n974), .A2(n973), .ZN(n975) );
  XNOR2_X1 U1068 ( .A(n976), .B(n975), .ZN(n978) );
  INV_X1 U1069 ( .A(G29), .ZN(n977) );
  NAND2_X1 U1070 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1071 ( .A1(G11), .A2(n979), .ZN(n1033) );
  INV_X1 U1072 ( .A(G16), .ZN(n1029) );
  XOR2_X1 U1073 ( .A(KEYINPUT56), .B(KEYINPUT122), .Z(n980) );
  XNOR2_X1 U1074 ( .A(n1029), .B(n980), .ZN(n1004) );
  XNOR2_X1 U1075 ( .A(G1966), .B(G168), .ZN(n982) );
  NAND2_X1 U1076 ( .A1(n982), .A2(n981), .ZN(n983) );
  XNOR2_X1 U1077 ( .A(n983), .B(KEYINPUT57), .ZN(n1002) );
  AND2_X1 U1078 ( .A1(G303), .A2(G1971), .ZN(n987) );
  NAND2_X1 U1079 ( .A1(n985), .A2(n984), .ZN(n986) );
  NOR2_X1 U1080 ( .A1(n987), .A2(n986), .ZN(n988) );
  XNOR2_X1 U1081 ( .A(KEYINPUT123), .B(n988), .ZN(n989) );
  NOR2_X1 U1082 ( .A1(n990), .A2(n989), .ZN(n998) );
  XNOR2_X1 U1083 ( .A(G1348), .B(n991), .ZN(n993) );
  XNOR2_X1 U1084 ( .A(G171), .B(G1961), .ZN(n992) );
  NAND2_X1 U1085 ( .A1(n993), .A2(n992), .ZN(n996) );
  XNOR2_X1 U1086 ( .A(G1341), .B(n994), .ZN(n995) );
  NOR2_X1 U1087 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1088 ( .A1(n998), .A2(n997), .ZN(n1000) );
  XNOR2_X1 U1089 ( .A(G1956), .B(G299), .ZN(n999) );
  NOR2_X1 U1090 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1091 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1092 ( .A1(n1004), .A2(n1003), .ZN(n1031) );
  XNOR2_X1 U1093 ( .A(G1348), .B(KEYINPUT59), .ZN(n1005) );
  XNOR2_X1 U1094 ( .A(n1005), .B(G4), .ZN(n1009) );
  XNOR2_X1 U1095 ( .A(G1981), .B(G6), .ZN(n1007) );
  XNOR2_X1 U1096 ( .A(G1341), .B(G19), .ZN(n1006) );
  NOR2_X1 U1097 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1098 ( .A1(n1009), .A2(n1008), .ZN(n1011) );
  XNOR2_X1 U1099 ( .A(G20), .B(G1956), .ZN(n1010) );
  NOR2_X1 U1100 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1101 ( .A(n1012), .B(KEYINPUT60), .ZN(n1015) );
  XOR2_X1 U1102 ( .A(G1966), .B(G21), .Z(n1013) );
  XNOR2_X1 U1103 ( .A(KEYINPUT124), .B(n1013), .ZN(n1014) );
  NAND2_X1 U1104 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1105 ( .A(n1016), .B(KEYINPUT125), .ZN(n1024) );
  XOR2_X1 U1106 ( .A(G1986), .B(KEYINPUT126), .Z(n1017) );
  XNOR2_X1 U1107 ( .A(G24), .B(n1017), .ZN(n1021) );
  XNOR2_X1 U1108 ( .A(G1976), .B(G23), .ZN(n1019) );
  XNOR2_X1 U1109 ( .A(G1971), .B(G22), .ZN(n1018) );
  NOR2_X1 U1110 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1111 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XOR2_X1 U1112 ( .A(KEYINPUT58), .B(n1022), .Z(n1023) );
  NAND2_X1 U1113 ( .A1(n1024), .A2(n1023), .ZN(n1026) );
  XNOR2_X1 U1114 ( .A(G5), .B(G1961), .ZN(n1025) );
  NOR2_X1 U1115 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XNOR2_X1 U1116 ( .A(KEYINPUT61), .B(n1027), .ZN(n1028) );
  NAND2_X1 U1117 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NAND2_X1 U1118 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  NOR2_X1 U1119 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  NAND2_X1 U1120 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  XOR2_X1 U1121 ( .A(KEYINPUT62), .B(n1036), .Z(G311) );
  INV_X1 U1122 ( .A(G311), .ZN(G150) );
endmodule

