

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580;

  XNOR2_X1 U320 ( .A(KEYINPUT113), .B(n438), .ZN(n533) );
  INV_X1 U321 ( .A(n554), .ZN(n524) );
  XOR2_X1 U322 ( .A(n390), .B(n389), .Z(n548) );
  XOR2_X1 U323 ( .A(n401), .B(KEYINPUT17), .Z(n288) );
  NOR2_X1 U324 ( .A1(n549), .A2(n464), .ZN(n465) );
  INV_X1 U325 ( .A(n397), .ZN(n326) );
  XNOR2_X1 U326 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U327 ( .A(G183GAT), .B(KEYINPUT18), .ZN(n400) );
  XNOR2_X1 U328 ( .A(n329), .B(n328), .ZN(n331) );
  NOR2_X1 U329 ( .A1(n548), .A2(n469), .ZN(n470) );
  XNOR2_X1 U330 ( .A(n572), .B(KEYINPUT41), .ZN(n557) );
  XNOR2_X1 U331 ( .A(n443), .B(G134GAT), .ZN(n444) );
  XNOR2_X1 U332 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U333 ( .A(n445), .B(n444), .ZN(G1343GAT) );
  XNOR2_X1 U334 ( .A(KEYINPUT111), .B(KEYINPUT48), .ZN(n370) );
  XOR2_X1 U335 ( .A(KEYINPUT72), .B(KEYINPUT11), .Z(n290) );
  NAND2_X1 U336 ( .A1(G232GAT), .A2(G233GAT), .ZN(n289) );
  XNOR2_X1 U337 ( .A(n290), .B(n289), .ZN(n291) );
  XOR2_X1 U338 ( .A(n291), .B(KEYINPUT10), .Z(n296) );
  XOR2_X1 U339 ( .A(G50GAT), .B(KEYINPUT71), .Z(n292) );
  XOR2_X1 U340 ( .A(G162GAT), .B(n292), .Z(n435) );
  XOR2_X1 U341 ( .A(G92GAT), .B(G218GAT), .Z(n294) );
  XNOR2_X1 U342 ( .A(G36GAT), .B(G190GAT), .ZN(n293) );
  XNOR2_X1 U343 ( .A(n294), .B(n293), .ZN(n391) );
  XNOR2_X1 U344 ( .A(n435), .B(n391), .ZN(n295) );
  XNOR2_X1 U345 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U346 ( .A(n297), .B(KEYINPUT9), .Z(n299) );
  XOR2_X1 U347 ( .A(G43GAT), .B(G134GAT), .Z(n417) );
  XNOR2_X1 U348 ( .A(n417), .B(KEYINPUT73), .ZN(n298) );
  XNOR2_X1 U349 ( .A(n299), .B(n298), .ZN(n305) );
  XOR2_X1 U350 ( .A(G29GAT), .B(KEYINPUT7), .Z(n301) );
  XNOR2_X1 U351 ( .A(KEYINPUT66), .B(KEYINPUT8), .ZN(n300) );
  XNOR2_X1 U352 ( .A(n301), .B(n300), .ZN(n316) );
  XOR2_X1 U353 ( .A(KEYINPUT68), .B(G85GAT), .Z(n303) );
  XNOR2_X1 U354 ( .A(G99GAT), .B(G106GAT), .ZN(n302) );
  XNOR2_X1 U355 ( .A(n303), .B(n302), .ZN(n334) );
  XOR2_X1 U356 ( .A(n316), .B(n334), .Z(n304) );
  XNOR2_X1 U357 ( .A(n305), .B(n304), .ZN(n546) );
  XOR2_X1 U358 ( .A(G43GAT), .B(G36GAT), .Z(n307) );
  NAND2_X1 U359 ( .A1(G229GAT), .A2(G233GAT), .ZN(n306) );
  XNOR2_X1 U360 ( .A(n307), .B(n306), .ZN(n320) );
  XOR2_X1 U361 ( .A(KEYINPUT65), .B(KEYINPUT29), .Z(n309) );
  XNOR2_X1 U362 ( .A(G113GAT), .B(KEYINPUT30), .ZN(n308) );
  XNOR2_X1 U363 ( .A(n309), .B(n308), .ZN(n313) );
  XOR2_X1 U364 ( .A(G141GAT), .B(G197GAT), .Z(n311) );
  XNOR2_X1 U365 ( .A(G169GAT), .B(G50GAT), .ZN(n310) );
  XNOR2_X1 U366 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U367 ( .A(n313), .B(n312), .Z(n318) );
  XOR2_X1 U368 ( .A(G1GAT), .B(G8GAT), .Z(n315) );
  XNOR2_X1 U369 ( .A(G22GAT), .B(G15GAT), .ZN(n314) );
  XNOR2_X1 U370 ( .A(n315), .B(n314), .ZN(n345) );
  XNOR2_X1 U371 ( .A(n316), .B(n345), .ZN(n317) );
  XNOR2_X1 U372 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U373 ( .A(n320), .B(n319), .Z(n505) );
  INV_X1 U374 ( .A(n505), .ZN(n568) );
  XOR2_X1 U375 ( .A(G57GAT), .B(KEYINPUT13), .Z(n342) );
  XOR2_X1 U376 ( .A(G148GAT), .B(G78GAT), .Z(n421) );
  XOR2_X1 U377 ( .A(n342), .B(n421), .Z(n322) );
  NAND2_X1 U378 ( .A1(G230GAT), .A2(G233GAT), .ZN(n321) );
  XNOR2_X1 U379 ( .A(n322), .B(n321), .ZN(n329) );
  XOR2_X1 U380 ( .A(G120GAT), .B(G71GAT), .Z(n414) );
  XOR2_X1 U381 ( .A(KEYINPUT32), .B(KEYINPUT67), .Z(n324) );
  XNOR2_X1 U382 ( .A(KEYINPUT70), .B(KEYINPUT69), .ZN(n323) );
  XNOR2_X1 U383 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U384 ( .A(n414), .B(n325), .ZN(n327) );
  XOR2_X1 U385 ( .A(G204GAT), .B(G64GAT), .Z(n397) );
  XNOR2_X1 U386 ( .A(G176GAT), .B(G92GAT), .ZN(n330) );
  XNOR2_X1 U387 ( .A(n331), .B(n330), .ZN(n333) );
  INV_X1 U388 ( .A(KEYINPUT33), .ZN(n332) );
  XNOR2_X1 U389 ( .A(n333), .B(n332), .ZN(n336) );
  XNOR2_X1 U390 ( .A(n334), .B(KEYINPUT31), .ZN(n335) );
  XNOR2_X1 U391 ( .A(n336), .B(n335), .ZN(n572) );
  NAND2_X1 U392 ( .A1(n568), .A2(n557), .ZN(n338) );
  INV_X1 U393 ( .A(KEYINPUT46), .ZN(n337) );
  XNOR2_X1 U394 ( .A(n338), .B(n337), .ZN(n358) );
  XOR2_X1 U395 ( .A(G155GAT), .B(G211GAT), .Z(n340) );
  XNOR2_X1 U396 ( .A(G127GAT), .B(G71GAT), .ZN(n339) );
  XNOR2_X1 U397 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U398 ( .A(n342), .B(n341), .Z(n344) );
  XNOR2_X1 U399 ( .A(G183GAT), .B(G78GAT), .ZN(n343) );
  XNOR2_X1 U400 ( .A(n344), .B(n343), .ZN(n349) );
  XOR2_X1 U401 ( .A(n345), .B(KEYINPUT12), .Z(n347) );
  NAND2_X1 U402 ( .A1(G231GAT), .A2(G233GAT), .ZN(n346) );
  XNOR2_X1 U403 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U404 ( .A(n349), .B(n348), .Z(n357) );
  XOR2_X1 U405 ( .A(KEYINPUT75), .B(KEYINPUT79), .Z(n351) );
  XNOR2_X1 U406 ( .A(KEYINPUT78), .B(KEYINPUT77), .ZN(n350) );
  XNOR2_X1 U407 ( .A(n351), .B(n350), .ZN(n355) );
  XOR2_X1 U408 ( .A(KEYINPUT76), .B(KEYINPUT15), .Z(n353) );
  XNOR2_X1 U409 ( .A(G64GAT), .B(KEYINPUT14), .ZN(n352) );
  XNOR2_X1 U410 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U411 ( .A(n355), .B(n354), .ZN(n356) );
  XNOR2_X1 U412 ( .A(n357), .B(n356), .ZN(n577) );
  NOR2_X1 U413 ( .A1(n358), .A2(n577), .ZN(n359) );
  XNOR2_X1 U414 ( .A(n359), .B(KEYINPUT109), .ZN(n360) );
  NOR2_X1 U415 ( .A1(n546), .A2(n360), .ZN(n361) );
  XNOR2_X1 U416 ( .A(n361), .B(KEYINPUT47), .ZN(n368) );
  XNOR2_X1 U417 ( .A(KEYINPUT74), .B(n546), .ZN(n564) );
  XNOR2_X1 U418 ( .A(KEYINPUT36), .B(n564), .ZN(n490) );
  NAND2_X1 U419 ( .A1(n490), .A2(n577), .ZN(n363) );
  XOR2_X1 U420 ( .A(KEYINPUT64), .B(KEYINPUT45), .Z(n362) );
  XNOR2_X1 U421 ( .A(n363), .B(n362), .ZN(n364) );
  NAND2_X1 U422 ( .A1(n364), .A2(n572), .ZN(n365) );
  XOR2_X1 U423 ( .A(KEYINPUT110), .B(n365), .Z(n366) );
  NAND2_X1 U424 ( .A1(n366), .A2(n505), .ZN(n367) );
  NAND2_X1 U425 ( .A1(n368), .A2(n367), .ZN(n369) );
  XNOR2_X1 U426 ( .A(n370), .B(n369), .ZN(n447) );
  XOR2_X1 U427 ( .A(G148GAT), .B(G162GAT), .Z(n372) );
  XNOR2_X1 U428 ( .A(G134GAT), .B(G120GAT), .ZN(n371) );
  XNOR2_X1 U429 ( .A(n372), .B(n371), .ZN(n374) );
  XOR2_X1 U430 ( .A(G29GAT), .B(G85GAT), .Z(n373) );
  XNOR2_X1 U431 ( .A(n374), .B(n373), .ZN(n388) );
  XOR2_X1 U432 ( .A(KEYINPUT5), .B(KEYINPUT4), .Z(n376) );
  XNOR2_X1 U433 ( .A(KEYINPUT6), .B(KEYINPUT90), .ZN(n375) );
  XNOR2_X1 U434 ( .A(n376), .B(n375), .ZN(n380) );
  XOR2_X1 U435 ( .A(KEYINPUT89), .B(KEYINPUT1), .Z(n378) );
  XNOR2_X1 U436 ( .A(G1GAT), .B(G57GAT), .ZN(n377) );
  XNOR2_X1 U437 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X1 U438 ( .A(n380), .B(n379), .Z(n386) );
  XOR2_X1 U439 ( .A(G127GAT), .B(KEYINPUT81), .Z(n382) );
  XNOR2_X1 U440 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n381) );
  XNOR2_X1 U441 ( .A(n382), .B(n381), .ZN(n416) );
  XOR2_X1 U442 ( .A(G155GAT), .B(KEYINPUT2), .Z(n384) );
  XNOR2_X1 U443 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n383) );
  XNOR2_X1 U444 ( .A(n384), .B(n383), .ZN(n420) );
  XNOR2_X1 U445 ( .A(n416), .B(n420), .ZN(n385) );
  XNOR2_X1 U446 ( .A(n386), .B(n385), .ZN(n387) );
  XNOR2_X1 U447 ( .A(n388), .B(n387), .ZN(n390) );
  NAND2_X1 U448 ( .A1(G225GAT), .A2(G233GAT), .ZN(n389) );
  XOR2_X1 U449 ( .A(KEYINPUT91), .B(n391), .Z(n395) );
  XOR2_X1 U450 ( .A(G211GAT), .B(KEYINPUT21), .Z(n393) );
  XNOR2_X1 U451 ( .A(G197GAT), .B(KEYINPUT88), .ZN(n392) );
  XNOR2_X1 U452 ( .A(n393), .B(n392), .ZN(n434) );
  XNOR2_X1 U453 ( .A(G8GAT), .B(n434), .ZN(n394) );
  XNOR2_X1 U454 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X1 U455 ( .A(n397), .B(n396), .Z(n399) );
  NAND2_X1 U456 ( .A1(G226GAT), .A2(G233GAT), .ZN(n398) );
  XNOR2_X1 U457 ( .A(n399), .B(n398), .ZN(n403) );
  XNOR2_X1 U458 ( .A(n400), .B(KEYINPUT19), .ZN(n401) );
  XNOR2_X1 U459 ( .A(G169GAT), .B(G176GAT), .ZN(n402) );
  XOR2_X1 U460 ( .A(n288), .B(n402), .Z(n411) );
  XNOR2_X1 U461 ( .A(n403), .B(n411), .ZN(n522) );
  XNOR2_X1 U462 ( .A(n522), .B(KEYINPUT27), .ZN(n461) );
  NAND2_X1 U463 ( .A1(n548), .A2(n461), .ZN(n472) );
  NOR2_X1 U464 ( .A1(n447), .A2(n472), .ZN(n404) );
  XOR2_X1 U465 ( .A(n404), .B(KEYINPUT112), .Z(n536) );
  XOR2_X1 U466 ( .A(KEYINPUT84), .B(KEYINPUT20), .Z(n406) );
  NAND2_X1 U467 ( .A1(G227GAT), .A2(G233GAT), .ZN(n405) );
  XNOR2_X1 U468 ( .A(n406), .B(n405), .ZN(n410) );
  XOR2_X1 U469 ( .A(KEYINPUT83), .B(KEYINPUT82), .Z(n408) );
  XNOR2_X1 U470 ( .A(G99GAT), .B(G190GAT), .ZN(n407) );
  XNOR2_X1 U471 ( .A(n408), .B(n407), .ZN(n409) );
  XOR2_X1 U472 ( .A(n410), .B(n409), .Z(n413) );
  XOR2_X1 U473 ( .A(G15GAT), .B(n411), .Z(n412) );
  XNOR2_X1 U474 ( .A(n413), .B(n412), .ZN(n415) );
  XNOR2_X1 U475 ( .A(n415), .B(n414), .ZN(n419) );
  XOR2_X1 U476 ( .A(n417), .B(n416), .Z(n418) );
  XNOR2_X1 U477 ( .A(n419), .B(n418), .ZN(n554) );
  XOR2_X1 U478 ( .A(n421), .B(n420), .Z(n423) );
  XNOR2_X1 U479 ( .A(G218GAT), .B(G106GAT), .ZN(n422) );
  XNOR2_X1 U480 ( .A(n423), .B(n422), .ZN(n427) );
  XOR2_X1 U481 ( .A(G204GAT), .B(KEYINPUT24), .Z(n425) );
  NAND2_X1 U482 ( .A1(G228GAT), .A2(G233GAT), .ZN(n424) );
  XNOR2_X1 U483 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U484 ( .A(n427), .B(n426), .Z(n432) );
  XOR2_X1 U485 ( .A(KEYINPUT22), .B(KEYINPUT86), .Z(n429) );
  XNOR2_X1 U486 ( .A(KEYINPUT87), .B(KEYINPUT23), .ZN(n428) );
  XNOR2_X1 U487 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U488 ( .A(G22GAT), .B(n430), .ZN(n431) );
  XNOR2_X1 U489 ( .A(n432), .B(n431), .ZN(n433) );
  XOR2_X1 U490 ( .A(n434), .B(n433), .Z(n436) );
  XNOR2_X1 U491 ( .A(n436), .B(n435), .ZN(n549) );
  XOR2_X1 U492 ( .A(KEYINPUT28), .B(n549), .Z(n471) );
  NAND2_X1 U493 ( .A1(n524), .A2(n471), .ZN(n437) );
  OR2_X1 U494 ( .A1(n536), .A2(n437), .ZN(n438) );
  NAND2_X1 U495 ( .A1(n533), .A2(n577), .ZN(n442) );
  XOR2_X1 U496 ( .A(KEYINPUT114), .B(KEYINPUT50), .Z(n440) );
  XNOR2_X1 U497 ( .A(G127GAT), .B(KEYINPUT115), .ZN(n439) );
  XNOR2_X1 U498 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U499 ( .A(n442), .B(n441), .ZN(G1342GAT) );
  NAND2_X1 U500 ( .A1(n533), .A2(n564), .ZN(n445) );
  XOR2_X1 U501 ( .A(KEYINPUT51), .B(KEYINPUT116), .Z(n443) );
  INV_X1 U502 ( .A(G218GAT), .ZN(n457) );
  XNOR2_X1 U503 ( .A(KEYINPUT62), .B(KEYINPUT126), .ZN(n455) );
  INV_X1 U504 ( .A(KEYINPUT123), .ZN(n453) );
  XNOR2_X1 U505 ( .A(n522), .B(KEYINPUT119), .ZN(n446) );
  NOR2_X1 U506 ( .A1(n447), .A2(n446), .ZN(n448) );
  XNOR2_X1 U507 ( .A(n448), .B(KEYINPUT54), .ZN(n551) );
  NAND2_X1 U508 ( .A1(n549), .A2(n554), .ZN(n450) );
  INV_X1 U509 ( .A(KEYINPUT26), .ZN(n449) );
  XNOR2_X1 U510 ( .A(n450), .B(n449), .ZN(n462) );
  INV_X1 U511 ( .A(n462), .ZN(n537) );
  NOR2_X1 U512 ( .A1(n537), .A2(n548), .ZN(n451) );
  AND2_X1 U513 ( .A1(n551), .A2(n451), .ZN(n452) );
  XNOR2_X1 U514 ( .A(n453), .B(n452), .ZN(n578) );
  AND2_X1 U515 ( .A1(n578), .A2(n490), .ZN(n454) );
  XNOR2_X1 U516 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U517 ( .A(n457), .B(n456), .ZN(G1355GAT) );
  XOR2_X1 U518 ( .A(KEYINPUT96), .B(KEYINPUT34), .Z(n480) );
  NAND2_X1 U519 ( .A1(n572), .A2(n568), .ZN(n493) );
  INV_X1 U520 ( .A(n577), .ZN(n458) );
  NOR2_X1 U521 ( .A1(n564), .A2(n458), .ZN(n460) );
  XNOR2_X1 U522 ( .A(KEYINPUT80), .B(KEYINPUT16), .ZN(n459) );
  XNOR2_X1 U523 ( .A(n460), .B(n459), .ZN(n478) );
  NAND2_X1 U524 ( .A1(n462), .A2(n461), .ZN(n463) );
  XNOR2_X1 U525 ( .A(KEYINPUT93), .B(n463), .ZN(n467) );
  AND2_X1 U526 ( .A1(n524), .A2(n522), .ZN(n464) );
  XOR2_X1 U527 ( .A(KEYINPUT25), .B(n465), .Z(n466) );
  NOR2_X1 U528 ( .A1(n467), .A2(n466), .ZN(n468) );
  XNOR2_X1 U529 ( .A(n468), .B(KEYINPUT94), .ZN(n469) );
  XNOR2_X1 U530 ( .A(n470), .B(KEYINPUT95), .ZN(n477) );
  XOR2_X1 U531 ( .A(n554), .B(KEYINPUT85), .Z(n475) );
  INV_X1 U532 ( .A(n471), .ZN(n526) );
  NOR2_X1 U533 ( .A1(n526), .A2(n472), .ZN(n473) );
  XNOR2_X1 U534 ( .A(n473), .B(KEYINPUT92), .ZN(n474) );
  NAND2_X1 U535 ( .A1(n475), .A2(n474), .ZN(n476) );
  NAND2_X1 U536 ( .A1(n477), .A2(n476), .ZN(n489) );
  NAND2_X1 U537 ( .A1(n478), .A2(n489), .ZN(n507) );
  NOR2_X1 U538 ( .A1(n493), .A2(n507), .ZN(n486) );
  NAND2_X1 U539 ( .A1(n486), .A2(n548), .ZN(n479) );
  XNOR2_X1 U540 ( .A(n480), .B(n479), .ZN(n481) );
  XOR2_X1 U541 ( .A(G1GAT), .B(n481), .Z(G1324GAT) );
  XOR2_X1 U542 ( .A(G8GAT), .B(KEYINPUT97), .Z(n483) );
  NAND2_X1 U543 ( .A1(n486), .A2(n522), .ZN(n482) );
  XNOR2_X1 U544 ( .A(n483), .B(n482), .ZN(G1325GAT) );
  XOR2_X1 U545 ( .A(G15GAT), .B(KEYINPUT35), .Z(n485) );
  NAND2_X1 U546 ( .A1(n486), .A2(n524), .ZN(n484) );
  XNOR2_X1 U547 ( .A(n485), .B(n484), .ZN(G1326GAT) );
  NAND2_X1 U548 ( .A1(n486), .A2(n526), .ZN(n487) );
  XNOR2_X1 U549 ( .A(n487), .B(KEYINPUT98), .ZN(n488) );
  XNOR2_X1 U550 ( .A(G22GAT), .B(n488), .ZN(G1327GAT) );
  XOR2_X1 U551 ( .A(G29GAT), .B(KEYINPUT39), .Z(n496) );
  NAND2_X1 U552 ( .A1(n490), .A2(n489), .ZN(n491) );
  NOR2_X1 U553 ( .A1(n577), .A2(n491), .ZN(n492) );
  XNOR2_X1 U554 ( .A(n492), .B(KEYINPUT37), .ZN(n519) );
  NOR2_X1 U555 ( .A1(n519), .A2(n493), .ZN(n494) );
  XNOR2_X1 U556 ( .A(n494), .B(KEYINPUT38), .ZN(n503) );
  NAND2_X1 U557 ( .A1(n503), .A2(n548), .ZN(n495) );
  XNOR2_X1 U558 ( .A(n496), .B(n495), .ZN(G1328GAT) );
  NAND2_X1 U559 ( .A1(n503), .A2(n522), .ZN(n498) );
  XOR2_X1 U560 ( .A(KEYINPUT99), .B(KEYINPUT100), .Z(n497) );
  XNOR2_X1 U561 ( .A(G36GAT), .B(n499), .ZN(G1329GAT) );
  XOR2_X1 U562 ( .A(KEYINPUT101), .B(KEYINPUT40), .Z(n501) );
  NAND2_X1 U563 ( .A1(n503), .A2(n524), .ZN(n500) );
  XNOR2_X1 U564 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U565 ( .A(G43GAT), .B(n502), .ZN(G1330GAT) );
  NAND2_X1 U566 ( .A1(n503), .A2(n526), .ZN(n504) );
  XNOR2_X1 U567 ( .A(n504), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U568 ( .A(KEYINPUT42), .B(KEYINPUT103), .Z(n509) );
  NAND2_X1 U569 ( .A1(n557), .A2(n505), .ZN(n506) );
  XNOR2_X1 U570 ( .A(n506), .B(KEYINPUT102), .ZN(n520) );
  NOR2_X1 U571 ( .A1(n520), .A2(n507), .ZN(n515) );
  NAND2_X1 U572 ( .A1(n515), .A2(n548), .ZN(n508) );
  XNOR2_X1 U573 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U574 ( .A(G57GAT), .B(n510), .ZN(G1332GAT) );
  NAND2_X1 U575 ( .A1(n515), .A2(n522), .ZN(n511) );
  XNOR2_X1 U576 ( .A(n511), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U577 ( .A(KEYINPUT104), .B(KEYINPUT105), .Z(n513) );
  NAND2_X1 U578 ( .A1(n515), .A2(n524), .ZN(n512) );
  XNOR2_X1 U579 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U580 ( .A(G71GAT), .B(n514), .ZN(G1334GAT) );
  XOR2_X1 U581 ( .A(KEYINPUT43), .B(KEYINPUT106), .Z(n517) );
  NAND2_X1 U582 ( .A1(n515), .A2(n526), .ZN(n516) );
  XNOR2_X1 U583 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U584 ( .A(G78GAT), .B(n518), .ZN(G1335GAT) );
  NOR2_X1 U585 ( .A1(n520), .A2(n519), .ZN(n527) );
  NAND2_X1 U586 ( .A1(n527), .A2(n548), .ZN(n521) );
  XNOR2_X1 U587 ( .A(G85GAT), .B(n521), .ZN(G1336GAT) );
  NAND2_X1 U588 ( .A1(n527), .A2(n522), .ZN(n523) );
  XNOR2_X1 U589 ( .A(n523), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U590 ( .A1(n524), .A2(n527), .ZN(n525) );
  XNOR2_X1 U591 ( .A(n525), .B(G99GAT), .ZN(G1338GAT) );
  XNOR2_X1 U592 ( .A(G106GAT), .B(KEYINPUT107), .ZN(n531) );
  XOR2_X1 U593 ( .A(KEYINPUT108), .B(KEYINPUT44), .Z(n529) );
  NAND2_X1 U594 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U595 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U596 ( .A(n531), .B(n530), .ZN(G1339GAT) );
  NAND2_X1 U597 ( .A1(n533), .A2(n568), .ZN(n532) );
  XNOR2_X1 U598 ( .A(G113GAT), .B(n532), .ZN(G1340GAT) );
  XOR2_X1 U599 ( .A(G120GAT), .B(KEYINPUT49), .Z(n535) );
  NAND2_X1 U600 ( .A1(n557), .A2(n533), .ZN(n534) );
  XNOR2_X1 U601 ( .A(n535), .B(n534), .ZN(G1341GAT) );
  NOR2_X1 U602 ( .A1(n537), .A2(n536), .ZN(n545) );
  NAND2_X1 U603 ( .A1(n545), .A2(n568), .ZN(n538) );
  XNOR2_X1 U604 ( .A(G141GAT), .B(n538), .ZN(G1344GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT52), .B(KEYINPUT117), .Z(n540) );
  NAND2_X1 U606 ( .A1(n545), .A2(n557), .ZN(n539) );
  XNOR2_X1 U607 ( .A(n540), .B(n539), .ZN(n542) );
  XOR2_X1 U608 ( .A(G148GAT), .B(KEYINPUT53), .Z(n541) );
  XNOR2_X1 U609 ( .A(n542), .B(n541), .ZN(G1345GAT) );
  NAND2_X1 U610 ( .A1(n545), .A2(n577), .ZN(n543) );
  XNOR2_X1 U611 ( .A(n543), .B(KEYINPUT118), .ZN(n544) );
  XNOR2_X1 U612 ( .A(G155GAT), .B(n544), .ZN(G1346GAT) );
  NAND2_X1 U613 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U614 ( .A(n547), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U615 ( .A1(n549), .A2(n548), .ZN(n550) );
  AND2_X1 U616 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U617 ( .A(n552), .B(KEYINPUT55), .ZN(n553) );
  NOR2_X1 U618 ( .A1(n554), .A2(n553), .ZN(n565) );
  NAND2_X1 U619 ( .A1(n568), .A2(n565), .ZN(n555) );
  XNOR2_X1 U620 ( .A(n555), .B(KEYINPUT120), .ZN(n556) );
  XNOR2_X1 U621 ( .A(G169GAT), .B(n556), .ZN(G1348GAT) );
  XOR2_X1 U622 ( .A(G176GAT), .B(KEYINPUT121), .Z(n559) );
  NAND2_X1 U623 ( .A1(n565), .A2(n557), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n559), .B(n558), .ZN(n561) );
  XOR2_X1 U625 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n560) );
  XNOR2_X1 U626 ( .A(n561), .B(n560), .ZN(G1349GAT) );
  NAND2_X1 U627 ( .A1(n565), .A2(n577), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n562), .B(KEYINPUT122), .ZN(n563) );
  XNOR2_X1 U629 ( .A(G183GAT), .B(n563), .ZN(G1350GAT) );
  NAND2_X1 U630 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U631 ( .A(n566), .B(KEYINPUT58), .ZN(n567) );
  XNOR2_X1 U632 ( .A(G190GAT), .B(n567), .ZN(G1351GAT) );
  XOR2_X1 U633 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n570) );
  NAND2_X1 U634 ( .A1(n578), .A2(n568), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U636 ( .A(G197GAT), .B(n571), .ZN(G1352GAT) );
  XOR2_X1 U637 ( .A(KEYINPUT124), .B(KEYINPUT61), .Z(n575) );
  INV_X1 U638 ( .A(n572), .ZN(n573) );
  NAND2_X1 U639 ( .A1(n578), .A2(n573), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U641 ( .A(G204GAT), .B(n576), .ZN(G1353GAT) );
  XOR2_X1 U642 ( .A(G211GAT), .B(KEYINPUT125), .Z(n580) );
  NAND2_X1 U643 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n580), .B(n579), .ZN(G1354GAT) );
endmodule

