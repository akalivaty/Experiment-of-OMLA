//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 1 0 1 0 0 0 0 1 0 1 1 0 0 0 1 0 0 1 1 1 1 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:00 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n687, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n726, new_n727, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n907, new_n908, new_n909, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004;
  INV_X1    g000(.A(KEYINPUT17), .ZN(new_n187));
  NOR2_X1   g001(.A1(G237), .A2(G953), .ZN(new_n188));
  AND3_X1   g002(.A1(new_n188), .A2(G143), .A3(G214), .ZN(new_n189));
  AOI21_X1  g003(.A(G143), .B1(new_n188), .B2(G214), .ZN(new_n190));
  OAI21_X1  g004(.A(G131), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT84), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G237), .ZN(new_n194));
  INV_X1    g008(.A(G953), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n194), .A2(new_n195), .A3(G214), .ZN(new_n196));
  INV_X1    g010(.A(G143), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n188), .A2(G143), .A3(G214), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n200), .A2(KEYINPUT84), .A3(G131), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n187), .B1(new_n193), .B2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT16), .ZN(new_n203));
  INV_X1    g017(.A(G140), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n203), .A2(new_n204), .A3(G125), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(G125), .ZN(new_n206));
  INV_X1    g020(.A(G125), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G140), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n205), .B1(new_n209), .B2(new_n203), .ZN(new_n210));
  INV_X1    g024(.A(G146), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  OAI211_X1 g026(.A(G146), .B(new_n205), .C1(new_n209), .C2(new_n203), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  OAI21_X1  g028(.A(KEYINPUT85), .B1(new_n202), .B2(new_n214), .ZN(new_n215));
  AOI21_X1  g029(.A(KEYINPUT84), .B1(new_n200), .B2(G131), .ZN(new_n216));
  INV_X1    g030(.A(G131), .ZN(new_n217));
  AOI211_X1 g031(.A(new_n192), .B(new_n217), .C1(new_n198), .C2(new_n199), .ZN(new_n218));
  OAI21_X1  g032(.A(KEYINPUT17), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT85), .ZN(new_n220));
  AND2_X1   g034(.A1(new_n212), .A2(new_n213), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n219), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n216), .A2(new_n218), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT86), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n198), .A2(new_n217), .A3(new_n199), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n223), .A2(new_n224), .A3(new_n187), .A4(new_n225), .ZN(new_n226));
  NAND4_X1  g040(.A1(new_n193), .A2(new_n201), .A3(new_n187), .A4(new_n225), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(KEYINPUT86), .ZN(new_n228));
  NAND4_X1  g042(.A1(new_n215), .A2(new_n222), .A3(new_n226), .A4(new_n228), .ZN(new_n229));
  XNOR2_X1  g043(.A(G113), .B(G122), .ZN(new_n230));
  INV_X1    g044(.A(G104), .ZN(new_n231));
  XNOR2_X1  g045(.A(new_n230), .B(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(new_n209), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(new_n211), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n209), .A2(G146), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT18), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n237), .A2(new_n217), .ZN(new_n238));
  OAI221_X1 g052(.A(new_n236), .B1(new_n200), .B2(new_n238), .C1(new_n191), .C2(new_n237), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n229), .A2(new_n232), .A3(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT87), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n229), .A2(KEYINPUT87), .A3(new_n232), .A4(new_n239), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n223), .A2(new_n225), .ZN(new_n245));
  XOR2_X1   g059(.A(new_n209), .B(KEYINPUT19), .Z(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(new_n211), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n245), .A2(new_n213), .A3(new_n247), .ZN(new_n248));
  AND2_X1   g062(.A1(new_n248), .A2(new_n239), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n249), .A2(new_n232), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n244), .A2(new_n251), .ZN(new_n252));
  NOR2_X1   g066(.A1(G475), .A2(G902), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n252), .A2(KEYINPUT20), .A3(new_n253), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n232), .B1(new_n229), .B2(new_n239), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n255), .B1(new_n242), .B2(new_n243), .ZN(new_n256));
  OAI21_X1  g070(.A(G475), .B1(new_n256), .B2(G902), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT20), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n250), .B1(new_n242), .B2(new_n243), .ZN(new_n259));
  INV_X1    g073(.A(new_n253), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n258), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  AND3_X1   g075(.A1(new_n254), .A2(new_n257), .A3(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT90), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n195), .A2(G952), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n264), .B1(G234), .B2(G237), .ZN(new_n265));
  XOR2_X1   g079(.A(KEYINPUT21), .B(G898), .Z(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(G234), .A2(G237), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n268), .A2(G902), .A3(G953), .ZN(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n265), .B1(new_n267), .B2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(G902), .ZN(new_n273));
  XNOR2_X1  g087(.A(G116), .B(G122), .ZN(new_n274));
  INV_X1    g088(.A(G107), .ZN(new_n275));
  XNOR2_X1  g089(.A(new_n274), .B(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n197), .A2(G128), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT13), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(G128), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(G143), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n277), .A2(new_n278), .ZN(new_n283));
  OAI21_X1  g097(.A(G134), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(G134), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n277), .A2(new_n281), .A3(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n276), .A2(new_n284), .A3(new_n286), .ZN(new_n287));
  XNOR2_X1  g101(.A(new_n287), .B(KEYINPUT88), .ZN(new_n288));
  INV_X1    g102(.A(new_n274), .ZN(new_n289));
  INV_X1    g103(.A(G116), .ZN(new_n290));
  OAI21_X1  g104(.A(KEYINPUT14), .B1(new_n290), .B2(G122), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n289), .A2(G107), .A3(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n274), .B1(KEYINPUT14), .B2(new_n275), .ZN(new_n293));
  INV_X1    g107(.A(new_n286), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n285), .B1(new_n277), .B2(new_n281), .ZN(new_n295));
  OAI211_X1 g109(.A(new_n292), .B(new_n293), .C1(new_n294), .C2(new_n295), .ZN(new_n296));
  XOR2_X1   g110(.A(KEYINPUT9), .B(G234), .Z(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  XNOR2_X1  g112(.A(KEYINPUT70), .B(G217), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  NOR3_X1   g114(.A1(new_n298), .A2(G953), .A3(new_n300), .ZN(new_n301));
  AND3_X1   g115(.A1(new_n288), .A2(new_n296), .A3(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n301), .B1(new_n288), .B2(new_n296), .ZN(new_n303));
  OAI211_X1 g117(.A(KEYINPUT89), .B(new_n273), .C1(new_n302), .C2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(G478), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n305), .A2(KEYINPUT15), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  XNOR2_X1  g121(.A(new_n304), .B(new_n307), .ZN(new_n308));
  NAND4_X1  g122(.A1(new_n262), .A2(new_n263), .A3(new_n272), .A4(new_n308), .ZN(new_n309));
  NAND4_X1  g123(.A1(new_n254), .A2(new_n257), .A3(new_n261), .A4(new_n308), .ZN(new_n310));
  OAI21_X1  g124(.A(KEYINPUT90), .B1(new_n310), .B2(new_n271), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(G469), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n231), .A2(G107), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n231), .A2(G107), .ZN(new_n316));
  OAI21_X1  g130(.A(G101), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  OAI21_X1  g131(.A(KEYINPUT3), .B1(new_n231), .B2(G107), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT3), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n319), .A2(new_n275), .A3(G104), .ZN(new_n320));
  INV_X1    g134(.A(G101), .ZN(new_n321));
  NAND4_X1  g135(.A1(new_n318), .A2(new_n320), .A3(new_n321), .A4(new_n314), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n317), .A2(new_n322), .ZN(new_n323));
  OAI21_X1  g137(.A(KEYINPUT64), .B1(new_n211), .B2(G143), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n211), .A2(G143), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n211), .A2(KEYINPUT64), .A3(G143), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n197), .A2(G146), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT1), .ZN(new_n330));
  OAI21_X1  g144(.A(G128), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n328), .A2(new_n331), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n326), .A2(new_n330), .A3(G128), .A4(new_n327), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n323), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  OR2_X1    g148(.A1(new_n334), .A2(KEYINPUT10), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT11), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n336), .B1(new_n285), .B2(G137), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n285), .A2(G137), .ZN(new_n338));
  INV_X1    g152(.A(G137), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n339), .A2(KEYINPUT11), .A3(G134), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n337), .A2(new_n338), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(G131), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n337), .A2(new_n340), .A3(new_n217), .A4(new_n338), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT64), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n346), .B1(new_n197), .B2(G146), .ZN(new_n347));
  OAI211_X1 g161(.A(G128), .B(new_n327), .C1(new_n347), .C2(new_n329), .ZN(new_n348));
  XNOR2_X1  g162(.A(KEYINPUT0), .B(G128), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n197), .A2(G146), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n325), .A2(new_n351), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n352), .A2(new_n349), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n350), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n318), .A2(new_n320), .A3(new_n314), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(G101), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n357), .A2(KEYINPUT4), .A3(new_n322), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT4), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n356), .A2(new_n359), .A3(G101), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n355), .A2(new_n358), .A3(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n323), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n331), .A2(new_n352), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n333), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n362), .A2(new_n364), .A3(KEYINPUT10), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n335), .A2(new_n345), .A3(new_n361), .A4(new_n365), .ZN(new_n366));
  XNOR2_X1  g180(.A(G110), .B(G140), .ZN(new_n367));
  AND2_X1   g181(.A1(new_n195), .A2(G227), .ZN(new_n368));
  XOR2_X1   g182(.A(new_n367), .B(new_n368), .Z(new_n369));
  NOR2_X1   g183(.A1(new_n362), .A2(new_n364), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n344), .B1(new_n370), .B2(new_n334), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(KEYINPUT12), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT12), .ZN(new_n373));
  OAI211_X1 g187(.A(new_n373), .B(new_n344), .C1(new_n370), .C2(new_n334), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n366), .A2(new_n369), .A3(new_n372), .A4(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n361), .A2(new_n365), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n334), .A2(KEYINPUT10), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n344), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(new_n366), .ZN(new_n379));
  INV_X1    g193(.A(new_n369), .ZN(new_n380));
  AOI22_X1  g194(.A1(new_n375), .A2(KEYINPUT78), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  AND3_X1   g195(.A1(new_n379), .A2(KEYINPUT78), .A3(new_n380), .ZN(new_n382));
  OAI211_X1 g196(.A(new_n313), .B(new_n273), .C1(new_n381), .C2(new_n382), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n366), .A2(new_n372), .A3(new_n374), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(KEYINPUT77), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT77), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n366), .A2(new_n386), .A3(new_n372), .A4(new_n374), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n385), .A2(new_n380), .A3(new_n387), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n378), .A2(new_n366), .A3(new_n369), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n388), .A2(G469), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(G469), .A2(G902), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n383), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  OAI21_X1  g206(.A(G221), .B1(new_n298), .B2(G902), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  AOI21_X1  g208(.A(G125), .B1(new_n333), .B2(new_n363), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n395), .B1(G125), .B2(new_n355), .ZN(new_n396));
  INV_X1    g210(.A(G224), .ZN(new_n397));
  OAI21_X1  g211(.A(KEYINPUT7), .B1(new_n397), .B2(G953), .ZN(new_n398));
  AOI21_X1  g212(.A(KEYINPUT82), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n353), .B1(new_n348), .B2(new_n349), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n400), .A2(new_n207), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT82), .ZN(new_n402));
  INV_X1    g216(.A(new_n398), .ZN(new_n403));
  NOR4_X1   g217(.A1(new_n401), .A2(new_n395), .A3(new_n402), .A4(new_n403), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n399), .A2(new_n404), .ZN(new_n405));
  XOR2_X1   g219(.A(G110), .B(G122), .Z(new_n406));
  XOR2_X1   g220(.A(new_n406), .B(KEYINPUT8), .Z(new_n407));
  INV_X1    g221(.A(KEYINPUT5), .ZN(new_n408));
  INV_X1    g222(.A(G119), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n408), .A2(new_n409), .A3(G116), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT79), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n408), .A2(new_n409), .A3(KEYINPUT79), .A4(G116), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  XNOR2_X1  g228(.A(G116), .B(G119), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(KEYINPUT5), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n414), .A2(G113), .A3(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT80), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(new_n415), .ZN(new_n420));
  XNOR2_X1  g234(.A(KEYINPUT2), .B(G113), .ZN(new_n421));
  OR2_X1    g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND4_X1  g236(.A1(new_n414), .A2(KEYINPUT80), .A3(G113), .A4(new_n416), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n419), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  AND2_X1   g238(.A1(new_n424), .A2(new_n323), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n362), .A2(new_n422), .A3(new_n417), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT81), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND4_X1  g242(.A1(new_n362), .A2(KEYINPUT81), .A3(new_n417), .A4(new_n422), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n407), .B1(new_n425), .B2(new_n430), .ZN(new_n431));
  NAND4_X1  g245(.A1(new_n419), .A2(new_n422), .A3(new_n362), .A4(new_n423), .ZN(new_n432));
  XNOR2_X1  g246(.A(new_n415), .B(new_n421), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n434), .A2(new_n358), .A3(new_n360), .ZN(new_n435));
  INV_X1    g249(.A(new_n406), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n432), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n403), .B1(new_n401), .B2(new_n395), .ZN(new_n438));
  NAND4_X1  g252(.A1(new_n405), .A2(new_n431), .A3(new_n437), .A4(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n432), .A2(new_n435), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(new_n406), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n441), .A2(KEYINPUT6), .A3(new_n437), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT6), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n440), .A2(new_n443), .A3(new_n406), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n397), .A2(G953), .ZN(new_n445));
  XNOR2_X1  g259(.A(new_n396), .B(new_n445), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n442), .A2(new_n444), .A3(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n439), .A2(new_n447), .A3(new_n273), .ZN(new_n448));
  OAI21_X1  g262(.A(G210), .B1(G237), .B2(G902), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT83), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n439), .A2(new_n447), .A3(new_n273), .A4(new_n449), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n451), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n448), .A2(KEYINPUT83), .A3(new_n450), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  OAI21_X1  g270(.A(G214), .B1(G237), .B2(G902), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  NOR3_X1   g272(.A1(new_n394), .A2(new_n456), .A3(new_n458), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n300), .B1(G234), .B2(new_n273), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT75), .ZN(new_n461));
  OAI21_X1  g275(.A(KEYINPUT72), .B1(new_n409), .B2(G128), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(KEYINPUT23), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n409), .A2(G128), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT23), .ZN(new_n465));
  OAI211_X1 g279(.A(KEYINPUT72), .B(new_n465), .C1(new_n409), .C2(G128), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n463), .A2(new_n464), .A3(new_n466), .ZN(new_n467));
  OR2_X1    g281(.A1(new_n467), .A2(G110), .ZN(new_n468));
  OAI21_X1  g282(.A(KEYINPUT71), .B1(new_n280), .B2(G119), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT71), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n470), .A2(new_n409), .A3(G128), .ZN(new_n471));
  OAI211_X1 g285(.A(new_n469), .B(new_n471), .C1(new_n409), .C2(G128), .ZN(new_n472));
  XNOR2_X1  g286(.A(KEYINPUT24), .B(G110), .ZN(new_n473));
  AOI21_X1  g287(.A(KEYINPUT73), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n472), .A2(KEYINPUT73), .A3(new_n473), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n468), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n234), .A2(new_n213), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n472), .A2(new_n473), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n480), .B1(new_n212), .B2(new_n213), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n467), .A2(G110), .ZN(new_n482));
  AOI22_X1  g296(.A1(new_n477), .A2(new_n479), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT74), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n195), .A2(G221), .A3(G234), .ZN(new_n485));
  OR2_X1    g299(.A1(new_n485), .A2(KEYINPUT22), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(KEYINPUT22), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n486), .A2(G137), .A3(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(G137), .B1(new_n486), .B2(new_n487), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n484), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(new_n490), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n492), .A2(KEYINPUT74), .A3(new_n488), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n461), .B1(new_n483), .B2(new_n494), .ZN(new_n495));
  AND2_X1   g309(.A1(new_n491), .A2(new_n493), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n481), .A2(new_n482), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(new_n476), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n499), .A2(new_n474), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n478), .B1(new_n500), .B2(new_n468), .ZN(new_n501));
  OAI211_X1 g315(.A(KEYINPUT75), .B(new_n496), .C1(new_n498), .C2(new_n501), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n483), .A2(new_n488), .A3(new_n492), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n495), .A2(new_n502), .A3(new_n273), .A4(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT25), .ZN(new_n505));
  AND2_X1   g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n504), .A2(new_n505), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n460), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  AND2_X1   g322(.A1(new_n495), .A2(new_n502), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n509), .A2(KEYINPUT76), .A3(new_n503), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n460), .A2(G902), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n495), .A2(new_n502), .A3(new_n503), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT76), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n510), .A2(new_n511), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n508), .A2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT32), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n339), .A2(G134), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n285), .A2(G137), .ZN(new_n519));
  OAI21_X1  g333(.A(G131), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n343), .A2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n364), .A2(new_n522), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n523), .B(new_n433), .C1(new_n345), .C2(new_n400), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT28), .ZN(new_n525));
  AND3_X1   g339(.A1(new_n524), .A2(KEYINPUT66), .A3(new_n525), .ZN(new_n526));
  AOI21_X1  g340(.A(KEYINPUT66), .B1(new_n524), .B2(new_n525), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  AOI22_X1  g342(.A1(new_n350), .A2(new_n354), .B1(new_n342), .B2(new_n343), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n521), .B1(new_n363), .B2(new_n333), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n434), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n524), .A2(new_n531), .ZN(new_n532));
  AOI21_X1  g346(.A(KEYINPUT65), .B1(new_n532), .B2(KEYINPUT28), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT65), .ZN(new_n534));
  AOI211_X1 g348(.A(new_n534), .B(new_n525), .C1(new_n524), .C2(new_n531), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n528), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n188), .A2(G210), .ZN(new_n537));
  XNOR2_X1  g351(.A(new_n537), .B(KEYINPUT27), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(KEYINPUT26), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT27), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n537), .B(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT26), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AND3_X1   g357(.A1(new_n539), .A2(new_n543), .A3(G101), .ZN(new_n544));
  AOI21_X1  g358(.A(G101), .B1(new_n539), .B2(new_n543), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n355), .A2(new_n344), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n548), .A2(KEYINPUT30), .A3(new_n523), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT30), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n550), .B1(new_n529), .B2(new_n530), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n549), .A2(new_n551), .A3(new_n434), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n552), .A2(new_n546), .A3(new_n524), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT31), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND4_X1  g369(.A1(new_n552), .A2(KEYINPUT31), .A3(new_n546), .A4(new_n524), .ZN(new_n556));
  AOI22_X1  g370(.A1(new_n536), .A2(new_n547), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NOR2_X1   g371(.A1(G472), .A2(G902), .ZN(new_n558));
  XOR2_X1   g372(.A(new_n558), .B(KEYINPUT67), .Z(new_n559));
  OAI21_X1  g373(.A(new_n517), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT68), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n555), .A2(new_n556), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT66), .ZN(new_n563));
  NOR3_X1   g377(.A1(new_n529), .A2(new_n530), .A3(new_n434), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n563), .B1(new_n564), .B2(KEYINPUT28), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n524), .A2(KEYINPUT66), .A3(new_n525), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n433), .B1(new_n548), .B2(new_n523), .ZN(new_n568));
  OAI21_X1  g382(.A(KEYINPUT28), .B1(new_n568), .B2(new_n564), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(new_n534), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n532), .A2(KEYINPUT65), .A3(KEYINPUT28), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n567), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n562), .B1(new_n572), .B2(new_n546), .ZN(new_n573));
  INV_X1    g387(.A(new_n559), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n573), .A2(KEYINPUT32), .A3(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n560), .A2(new_n561), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n573), .A2(new_n574), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n577), .A2(KEYINPUT68), .A3(new_n517), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  OAI211_X1 g393(.A(new_n528), .B(new_n546), .C1(new_n533), .C2(new_n535), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT29), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n552), .A2(new_n524), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(new_n547), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n580), .A2(new_n581), .A3(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT69), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n528), .A2(KEYINPUT29), .A3(new_n546), .A4(new_n569), .ZN(new_n587));
  AND2_X1   g401(.A1(new_n587), .A2(new_n273), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n580), .A2(KEYINPUT69), .A3(new_n581), .A4(new_n583), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n586), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(G472), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n516), .B1(new_n579), .B2(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n312), .A2(new_n459), .A3(new_n592), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n593), .B(G101), .ZN(G3));
  INV_X1    g408(.A(KEYINPUT91), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n595), .B1(new_n557), .B2(G902), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n573), .A2(KEYINPUT91), .A3(new_n273), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n596), .A2(G472), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(new_n577), .ZN(new_n599));
  NOR3_X1   g413(.A1(new_n599), .A2(new_n516), .A3(new_n394), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n254), .A2(new_n257), .A3(new_n261), .ZN(new_n601));
  NAND2_X1  g415(.A1(KEYINPUT92), .A2(G478), .ZN(new_n602));
  OR2_X1    g416(.A1(KEYINPUT92), .A2(G478), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n302), .A2(new_n303), .ZN(new_n604));
  OAI211_X1 g418(.A(new_n602), .B(new_n603), .C1(new_n604), .C2(G902), .ZN(new_n605));
  OR2_X1    g419(.A1(new_n604), .A2(KEYINPUT33), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n604), .A2(KEYINPUT33), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n273), .A2(G478), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n605), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n601), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n451), .A2(new_n453), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(new_n457), .ZN(new_n613));
  NOR3_X1   g427(.A1(new_n611), .A2(new_n271), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n600), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(KEYINPUT93), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n616), .B(KEYINPUT34), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n617), .B(new_n231), .ZN(G6));
  XNOR2_X1  g432(.A(new_n304), .B(new_n306), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n254), .A2(new_n257), .A3(new_n261), .A4(new_n619), .ZN(new_n620));
  NOR3_X1   g434(.A1(new_n620), .A2(new_n613), .A3(new_n271), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n600), .A2(new_n621), .ZN(new_n622));
  XOR2_X1   g436(.A(KEYINPUT35), .B(G107), .Z(new_n623));
  XNOR2_X1  g437(.A(new_n622), .B(new_n623), .ZN(G9));
  INV_X1    g438(.A(new_n599), .ZN(new_n625));
  INV_X1    g439(.A(new_n460), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n509), .A2(KEYINPUT25), .A3(new_n273), .A4(new_n503), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n504), .A2(new_n505), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n626), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT36), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n494), .A2(new_n630), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n631), .B1(new_n501), .B2(new_n498), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n483), .A2(new_n630), .A3(new_n494), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n632), .A2(new_n633), .A3(new_n511), .ZN(new_n634));
  XOR2_X1   g448(.A(new_n634), .B(KEYINPUT94), .Z(new_n635));
  OAI21_X1  g449(.A(KEYINPUT95), .B1(new_n629), .B2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT95), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n634), .B(KEYINPUT94), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n508), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n636), .A2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n312), .A2(new_n459), .A3(new_n625), .A4(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(KEYINPUT37), .ZN(new_n643));
  XOR2_X1   g457(.A(new_n643), .B(G110), .Z(G12));
  AOI21_X1  g458(.A(new_n640), .B1(new_n579), .B2(new_n591), .ZN(new_n645));
  INV_X1    g459(.A(new_n394), .ZN(new_n646));
  XNOR2_X1  g460(.A(KEYINPUT96), .B(G900), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n265), .B1(new_n270), .B2(new_n647), .ZN(new_n648));
  NOR3_X1   g462(.A1(new_n620), .A2(new_n613), .A3(new_n648), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n645), .A2(new_n646), .A3(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(G128), .ZN(G30));
  NAND2_X1  g465(.A1(new_n456), .A2(KEYINPUT97), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT97), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n454), .A2(new_n653), .A3(new_n455), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT38), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n648), .B(KEYINPUT39), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n646), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(KEYINPUT40), .ZN(new_n661));
  OR3_X1    g475(.A1(new_n394), .A2(KEYINPUT40), .A3(new_n658), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n652), .A2(KEYINPUT38), .A3(new_n654), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n657), .A2(new_n661), .A3(new_n662), .A4(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n582), .A2(new_n546), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n273), .B1(new_n532), .B2(new_n546), .ZN(new_n667));
  OAI21_X1  g481(.A(G472), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n579), .A2(new_n668), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n262), .A2(new_n308), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n669), .A2(new_n457), .A3(new_n640), .A4(new_n670), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n664), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(new_n197), .ZN(G45));
  AOI21_X1  g487(.A(new_n458), .B1(new_n451), .B2(new_n453), .ZN(new_n674));
  INV_X1    g488(.A(new_n648), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n601), .A2(new_n610), .A3(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n645), .A2(new_n646), .A3(new_n674), .A4(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G146), .ZN(G48));
  OAI21_X1  g493(.A(new_n273), .B1(new_n381), .B2(new_n382), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(G469), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n681), .A2(new_n393), .A3(new_n383), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n614), .A2(new_n592), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(KEYINPUT41), .B(G113), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(G15));
  NAND3_X1  g500(.A1(new_n592), .A2(new_n621), .A3(new_n683), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G116), .ZN(G18));
  AND2_X1   g502(.A1(new_n681), .A2(new_n383), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n689), .A2(KEYINPUT98), .A3(new_n393), .A4(new_n674), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT98), .ZN(new_n691));
  OAI21_X1  g505(.A(new_n691), .B1(new_n682), .B2(new_n613), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n312), .A2(new_n645), .A3(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G119), .ZN(G21));
  OAI21_X1  g509(.A(G472), .B1(new_n557), .B2(G902), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n559), .B(KEYINPUT99), .ZN(new_n697));
  INV_X1    g511(.A(new_n562), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n546), .B1(new_n528), .B2(new_n569), .ZN(new_n699));
  OAI21_X1  g513(.A(new_n697), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n696), .A2(new_n700), .ZN(new_n701));
  NOR3_X1   g515(.A1(new_n682), .A2(new_n701), .A3(new_n516), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n702), .A2(new_n670), .A3(new_n272), .A4(new_n674), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G122), .ZN(G24));
  NAND4_X1  g518(.A1(new_n636), .A2(new_n639), .A3(new_n696), .A4(new_n700), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n705), .A2(new_n676), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n693), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G125), .ZN(G27));
  NAND2_X1  g522(.A1(new_n456), .A2(new_n457), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n389), .B(KEYINPUT100), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(new_n388), .ZN(new_n711));
  OAI211_X1 g525(.A(new_n383), .B(new_n391), .C1(new_n711), .C2(new_n313), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(new_n393), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n709), .A2(new_n713), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n676), .A2(KEYINPUT42), .ZN(new_n715));
  AND3_X1   g529(.A1(new_n592), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT101), .ZN(new_n717));
  AND2_X1   g531(.A1(new_n560), .A2(new_n575), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n591), .A2(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(new_n516), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n717), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  AOI211_X1 g535(.A(KEYINPUT101), .B(new_n516), .C1(new_n591), .C2(new_n718), .ZN(new_n722));
  OAI211_X1 g536(.A(new_n677), .B(new_n714), .C1(new_n721), .C2(new_n722), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n716), .B1(new_n723), .B2(KEYINPUT42), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G131), .ZN(G33));
  INV_X1    g539(.A(new_n620), .ZN(new_n726));
  AND4_X1   g540(.A1(new_n592), .A2(new_n726), .A3(new_n675), .A4(new_n714), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(new_n285), .ZN(G36));
  INV_X1    g542(.A(KEYINPUT102), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT45), .ZN(new_n730));
  OAI21_X1  g544(.A(G469), .B1(new_n711), .B2(new_n730), .ZN(new_n731));
  AOI21_X1  g545(.A(KEYINPUT45), .B1(new_n388), .B2(new_n389), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n391), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT46), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  OAI211_X1 g549(.A(KEYINPUT46), .B(new_n391), .C1(new_n731), .C2(new_n732), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n735), .A2(new_n383), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(new_n393), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n729), .B1(new_n738), .B2(new_n658), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n737), .A2(KEYINPUT102), .A3(new_n393), .A4(new_n659), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n709), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n262), .A2(new_n610), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT103), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT43), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n742), .A2(new_n743), .A3(KEYINPUT43), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n746), .A2(KEYINPUT104), .A3(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT104), .ZN(new_n749));
  AOI21_X1  g563(.A(KEYINPUT43), .B1(new_n742), .B2(new_n743), .ZN(new_n750));
  AOI211_X1 g564(.A(KEYINPUT103), .B(new_n745), .C1(new_n262), .C2(new_n610), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n749), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n625), .A2(new_n640), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n748), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT44), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n748), .A2(new_n752), .A3(KEYINPUT44), .A4(new_n753), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n741), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G137), .ZN(G39));
  NAND2_X1  g573(.A1(new_n579), .A2(new_n591), .ZN(new_n760));
  NOR4_X1   g574(.A1(new_n760), .A2(new_n720), .A3(new_n676), .A4(new_n709), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT105), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n761), .B(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT47), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n737), .A2(new_n764), .A3(new_n393), .ZN(new_n765));
  INV_X1    g579(.A(new_n765), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n764), .B1(new_n737), .B2(new_n393), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n763), .A2(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G140), .ZN(G42));
  INV_X1    g584(.A(new_n669), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(new_n265), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n709), .A2(new_n682), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(new_n720), .ZN(new_n774));
  OR3_X1    g588(.A1(new_n772), .A2(new_n774), .A3(new_n611), .ZN(new_n775));
  NOR2_X1   g589(.A1(KEYINPUT114), .A2(KEYINPUT48), .ZN(new_n776));
  AND2_X1   g590(.A1(KEYINPUT114), .A2(KEYINPUT48), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n746), .A2(new_n773), .A3(new_n265), .A4(new_n747), .ZN(new_n778));
  OR2_X1    g592(.A1(new_n778), .A2(KEYINPUT112), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(KEYINPUT112), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n721), .A2(new_n722), .ZN(new_n782));
  INV_X1    g596(.A(new_n782), .ZN(new_n783));
  AOI211_X1 g597(.A(new_n776), .B(new_n777), .C1(new_n781), .C2(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(new_n780), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n778), .A2(KEYINPUT112), .ZN(new_n786));
  OAI211_X1 g600(.A(new_n783), .B(new_n777), .C1(new_n785), .C2(new_n786), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n701), .A2(new_n516), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n746), .A2(new_n265), .A3(new_n788), .A4(new_n747), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n789), .B1(new_n692), .B2(new_n690), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n790), .A2(new_n264), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n787), .A2(new_n791), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n784), .A2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT51), .ZN(new_n794));
  INV_X1    g608(.A(new_n767), .ZN(new_n795));
  INV_X1    g609(.A(new_n393), .ZN(new_n796));
  AOI22_X1  g610(.A1(new_n795), .A2(new_n765), .B1(new_n796), .B2(new_n689), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n789), .A2(new_n709), .ZN(new_n798));
  INV_X1    g612(.A(new_n798), .ZN(new_n799));
  OAI21_X1  g613(.A(KEYINPUT111), .B1(new_n797), .B2(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(new_n689), .ZN(new_n801));
  OAI22_X1  g615(.A1(new_n766), .A2(new_n767), .B1(new_n393), .B2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT111), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n802), .A2(new_n803), .A3(new_n798), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n800), .A2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(new_n705), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n806), .B1(new_n785), .B2(new_n786), .ZN(new_n807));
  AND3_X1   g621(.A1(new_n746), .A2(new_n265), .A3(new_n747), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n457), .B1(new_n657), .B2(new_n663), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n808), .A2(KEYINPUT50), .A3(new_n702), .A4(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT50), .ZN(new_n811));
  INV_X1    g625(.A(new_n809), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n746), .A2(new_n265), .A3(new_n702), .A4(new_n747), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n811), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n810), .A2(new_n814), .ZN(new_n815));
  NOR4_X1   g629(.A1(new_n772), .A2(new_n774), .A3(new_n601), .A4(new_n610), .ZN(new_n816));
  INV_X1    g630(.A(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n807), .A2(new_n815), .A3(new_n817), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n794), .B1(new_n805), .B2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT113), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n797), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n802), .A2(KEYINPUT113), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n821), .A2(new_n798), .A3(new_n822), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n816), .B1(new_n781), .B2(new_n806), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n823), .A2(new_n824), .A3(KEYINPUT51), .A4(new_n815), .ZN(new_n825));
  AND4_X1   g639(.A1(new_n775), .A2(new_n793), .A3(new_n819), .A4(new_n825), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n714), .A2(new_n601), .A3(new_n806), .A4(new_n610), .ZN(new_n827));
  INV_X1    g641(.A(new_n310), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n645), .A2(new_n828), .A3(new_n646), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n827), .B1(new_n829), .B2(new_n709), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n830), .A2(new_n675), .ZN(new_n831));
  INV_X1    g645(.A(new_n727), .ZN(new_n832));
  AND3_X1   g646(.A1(new_n724), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n694), .A2(new_n684), .A3(new_n687), .A4(new_n703), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n456), .A2(new_n458), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n611), .A2(new_n620), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n600), .A2(new_n272), .A3(new_n835), .A4(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n642), .A2(new_n837), .A3(new_n593), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n838), .A2(KEYINPUT108), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT108), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n642), .A2(new_n837), .A3(new_n593), .A4(new_n840), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n834), .B1(new_n839), .B2(new_n841), .ZN(new_n842));
  AND2_X1   g656(.A1(new_n833), .A2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT110), .ZN(new_n844));
  XNOR2_X1  g658(.A(new_n648), .B(KEYINPUT109), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n713), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n629), .A2(new_n635), .ZN(new_n847));
  AND3_X1   g661(.A1(new_n601), .A2(new_n619), .A3(new_n674), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n669), .A2(new_n846), .A3(new_n847), .A4(new_n848), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n678), .A2(new_n650), .A3(new_n707), .A4(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT52), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n844), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n850), .A2(new_n851), .ZN(new_n853));
  XNOR2_X1  g667(.A(new_n852), .B(new_n853), .ZN(new_n854));
  AOI21_X1  g668(.A(KEYINPUT53), .B1(new_n843), .B2(new_n854), .ZN(new_n855));
  XNOR2_X1  g669(.A(new_n850), .B(new_n851), .ZN(new_n856));
  AND4_X1   g670(.A1(KEYINPUT53), .A2(new_n833), .A3(new_n842), .A4(new_n856), .ZN(new_n857));
  OAI21_X1  g671(.A(KEYINPUT54), .B1(new_n855), .B2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT54), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT53), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n860), .B1(new_n843), .B2(new_n854), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n833), .A2(new_n842), .A3(new_n856), .A4(new_n860), .ZN(new_n862));
  INV_X1    g676(.A(new_n862), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n859), .B1(new_n861), .B2(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n826), .A2(new_n858), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n865), .A2(KEYINPUT115), .ZN(new_n866));
  OR2_X1    g680(.A1(G952), .A2(G953), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT115), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n826), .A2(new_n858), .A3(new_n864), .A4(new_n868), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n866), .A2(new_n867), .A3(new_n869), .ZN(new_n870));
  NOR4_X1   g684(.A1(new_n742), .A2(new_n516), .A3(new_n796), .A4(new_n458), .ZN(new_n871));
  XOR2_X1   g685(.A(new_n871), .B(KEYINPUT106), .Z(new_n872));
  NOR2_X1   g686(.A1(new_n801), .A2(KEYINPUT49), .ZN(new_n873));
  XNOR2_X1  g687(.A(new_n873), .B(KEYINPUT107), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n874), .B1(KEYINPUT49), .B2(new_n801), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n657), .A2(new_n663), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n872), .A2(new_n875), .A3(new_n771), .A4(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n870), .A2(new_n877), .ZN(G75));
  NOR3_X1   g692(.A1(new_n861), .A2(new_n273), .A3(new_n863), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(G210), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT56), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n442), .A2(new_n444), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n882), .B(new_n446), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n883), .B(KEYINPUT55), .ZN(new_n884));
  INV_X1    g698(.A(new_n884), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n885), .B1(KEYINPUT116), .B2(new_n881), .ZN(new_n886));
  AND3_X1   g700(.A1(new_n880), .A2(new_n881), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n886), .B1(new_n880), .B2(new_n881), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n195), .A2(G952), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n887), .A2(new_n888), .A3(new_n889), .ZN(G51));
  XOR2_X1   g704(.A(new_n391), .B(KEYINPUT57), .Z(new_n891));
  NOR2_X1   g705(.A1(new_n852), .A2(new_n853), .ZN(new_n892));
  NOR3_X1   g706(.A1(new_n850), .A2(new_n844), .A3(new_n851), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n839), .A2(new_n841), .ZN(new_n895));
  AOI211_X1 g709(.A(new_n716), .B(new_n727), .C1(new_n723), .C2(KEYINPUT42), .ZN(new_n896));
  INV_X1    g710(.A(new_n834), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n895), .A2(new_n896), .A3(new_n831), .A4(new_n897), .ZN(new_n898));
  OAI21_X1  g712(.A(KEYINPUT53), .B1(new_n894), .B2(new_n898), .ZN(new_n899));
  AND3_X1   g713(.A1(new_n899), .A2(KEYINPUT54), .A3(new_n862), .ZN(new_n900));
  AOI21_X1  g714(.A(KEYINPUT54), .B1(new_n899), .B2(new_n862), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n891), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n902), .B1(new_n381), .B2(new_n382), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n731), .A2(new_n732), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n879), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n889), .B1(new_n903), .B2(new_n905), .ZN(G54));
  NAND3_X1  g720(.A1(new_n879), .A2(KEYINPUT58), .A3(G475), .ZN(new_n907));
  AND2_X1   g721(.A1(new_n907), .A2(new_n259), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n907), .A2(new_n259), .ZN(new_n909));
  NOR3_X1   g723(.A1(new_n908), .A2(new_n909), .A3(new_n889), .ZN(G60));
  INV_X1    g724(.A(KEYINPUT117), .ZN(new_n911));
  INV_X1    g725(.A(new_n608), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n858), .A2(new_n864), .ZN(new_n913));
  NAND2_X1  g727(.A1(G478), .A2(G902), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n914), .B(KEYINPUT59), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n912), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  AND2_X1   g730(.A1(new_n912), .A2(new_n915), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n917), .B1(new_n900), .B2(new_n901), .ZN(new_n918));
  INV_X1    g732(.A(new_n889), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n911), .B1(new_n916), .B2(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(new_n857), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n860), .B1(new_n894), .B2(new_n898), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n859), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n915), .B1(new_n924), .B2(new_n901), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n925), .A2(new_n608), .ZN(new_n926));
  NAND4_X1  g740(.A1(new_n926), .A2(KEYINPUT117), .A3(new_n919), .A4(new_n918), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n921), .A2(new_n927), .ZN(G63));
  NOR2_X1   g742(.A1(new_n861), .A2(new_n863), .ZN(new_n929));
  NAND2_X1  g743(.A1(G217), .A2(G902), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n930), .B(KEYINPUT60), .Z(new_n931));
  INV_X1    g745(.A(KEYINPUT118), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n632), .A2(new_n633), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n932), .B1(new_n933), .B2(KEYINPUT119), .ZN(new_n934));
  OR2_X1    g748(.A1(new_n933), .A2(KEYINPUT119), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n929), .A2(new_n931), .A3(new_n934), .A4(new_n935), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n899), .A2(new_n862), .A3(new_n931), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n510), .A2(new_n514), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n889), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n936), .B1(new_n939), .B2(new_n932), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT61), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n940), .B(new_n941), .ZN(G66));
  OAI21_X1  g756(.A(G953), .B1(new_n267), .B2(new_n397), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n842), .B(KEYINPUT120), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n943), .B1(new_n944), .B2(G953), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n882), .B1(G898), .B2(new_n195), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n946), .B(KEYINPUT121), .Z(new_n947));
  XNOR2_X1  g761(.A(new_n945), .B(new_n947), .ZN(G69));
  INV_X1    g762(.A(new_n672), .ZN(new_n949));
  AND2_X1   g763(.A1(new_n650), .A2(new_n707), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n949), .A2(KEYINPUT62), .A3(new_n678), .A4(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT62), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n950), .A2(new_n678), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n952), .B1(new_n953), .B2(new_n672), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n951), .A2(new_n954), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n660), .A2(new_n709), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n956), .A2(new_n592), .A3(new_n836), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n957), .B(KEYINPUT122), .ZN(new_n958));
  INV_X1    g772(.A(new_n958), .ZN(new_n959));
  NAND4_X1  g773(.A1(new_n955), .A2(new_n769), .A3(new_n758), .A4(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n960), .A2(new_n195), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n549), .A2(new_n551), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n962), .B(new_n246), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n963), .B1(G900), .B2(G953), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n953), .B1(new_n763), .B2(new_n768), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n739), .A2(new_n740), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n967), .A2(new_n783), .A3(new_n848), .ZN(new_n968));
  NAND4_X1  g782(.A1(new_n758), .A2(new_n966), .A3(new_n896), .A4(new_n968), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n965), .B1(new_n969), .B2(G953), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n970), .A2(KEYINPUT124), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT124), .ZN(new_n972));
  OAI211_X1 g786(.A(new_n972), .B(new_n965), .C1(new_n969), .C2(G953), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n964), .A2(new_n971), .A3(new_n973), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n195), .B1(G227), .B2(G900), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  AND2_X1   g790(.A1(new_n758), .A2(new_n769), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n958), .B1(new_n951), .B2(new_n954), .ZN(new_n978));
  AOI21_X1  g792(.A(G953), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(new_n963), .ZN(new_n980));
  OAI21_X1  g794(.A(KEYINPUT123), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(KEYINPUT123), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n961), .A2(new_n982), .A3(new_n963), .ZN(new_n983));
  INV_X1    g797(.A(new_n975), .ZN(new_n984));
  NAND4_X1  g798(.A1(new_n981), .A2(new_n983), .A3(new_n984), .A4(new_n970), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n976), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n986), .A2(KEYINPUT125), .ZN(new_n987));
  INV_X1    g801(.A(KEYINPUT125), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n976), .A2(new_n988), .A3(new_n985), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n987), .A2(new_n989), .ZN(G72));
  NAND2_X1  g804(.A1(G472), .A2(G902), .ZN(new_n991));
  XOR2_X1   g805(.A(new_n991), .B(KEYINPUT63), .Z(new_n992));
  INV_X1    g806(.A(new_n992), .ZN(new_n993));
  INV_X1    g807(.A(new_n960), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n993), .B1(new_n994), .B2(new_n944), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n919), .B1(new_n995), .B2(new_n665), .ZN(new_n996));
  AND3_X1   g810(.A1(new_n758), .A2(new_n966), .A3(new_n896), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n944), .A2(new_n968), .A3(new_n997), .ZN(new_n998));
  AOI211_X1 g812(.A(new_n546), .B(new_n582), .C1(new_n998), .C2(new_n992), .ZN(new_n999));
  XNOR2_X1  g813(.A(new_n583), .B(KEYINPUT126), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n1000), .A2(new_n553), .ZN(new_n1001));
  OAI211_X1 g815(.A(new_n992), .B(new_n1001), .C1(new_n855), .C2(new_n857), .ZN(new_n1002));
  OR2_X1    g816(.A1(new_n1002), .A2(KEYINPUT127), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1002), .A2(KEYINPUT127), .ZN(new_n1004));
  AOI211_X1 g818(.A(new_n996), .B(new_n999), .C1(new_n1003), .C2(new_n1004), .ZN(G57));
endmodule


