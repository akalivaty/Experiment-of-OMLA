//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 1 0 0 0 1 0 0 0 0 1 0 0 1 0 1 0 0 0 1 1 1 1 1 1 0 1 0 0 1 1 0 1 1 0 1 0 1 1 0 1 1 1 0 0 0 0 1 0 0 1 0 0 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:41 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n705, new_n706, new_n707, new_n708, new_n709, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n754, new_n755, new_n756, new_n757,
    new_n759, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n779, new_n780, new_n781, new_n783,
    new_n784, new_n785, new_n786, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n827,
    new_n829, new_n831, new_n832, new_n833, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n862, new_n863, new_n864, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n927, new_n928, new_n929, new_n930,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n939,
    new_n940, new_n941, new_n942;
  INV_X1    g000(.A(KEYINPUT1), .ZN(new_n202));
  INV_X1    g001(.A(G113gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n203), .A2(G120gat), .ZN(new_n204));
  INV_X1    g003(.A(G120gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n205), .A2(G113gat), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n202), .B1(new_n204), .B2(new_n206), .ZN(new_n207));
  NOR2_X1   g006(.A1(KEYINPUT68), .A2(KEYINPUT1), .ZN(new_n208));
  OR2_X1    g007(.A1(G127gat), .A2(G134gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(G127gat), .A2(G134gat), .ZN(new_n210));
  AOI21_X1  g009(.A(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n207), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n205), .A2(G113gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n203), .A2(G120gat), .ZN(new_n214));
  AOI21_X1  g013(.A(KEYINPUT1), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  AND2_X1   g014(.A1(G127gat), .A2(G134gat), .ZN(new_n216));
  NOR2_X1   g015(.A1(G127gat), .A2(G134gat), .ZN(new_n217));
  OAI22_X1  g016(.A1(new_n216), .A2(new_n217), .B1(KEYINPUT68), .B2(KEYINPUT1), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n212), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g019(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(KEYINPUT66), .ZN(new_n222));
  NAND2_X1  g021(.A1(G169gat), .A2(G176gat), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT66), .ZN(new_n224));
  OAI211_X1 g023(.A(new_n224), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n222), .A2(new_n223), .A3(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(KEYINPUT67), .ZN(new_n227));
  OR3_X1    g026(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT67), .ZN(new_n229));
  NAND4_X1  g028(.A1(new_n222), .A2(new_n229), .A3(new_n225), .A4(new_n223), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n227), .A2(new_n228), .A3(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(G183gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(KEYINPUT27), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT27), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(G183gat), .ZN(new_n235));
  INV_X1    g034(.A(G190gat), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n233), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT28), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  XNOR2_X1  g038(.A(KEYINPUT27), .B(G183gat), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n240), .A2(KEYINPUT28), .A3(new_n236), .ZN(new_n241));
  AOI22_X1  g040(.A1(new_n239), .A2(new_n241), .B1(G183gat), .B2(G190gat), .ZN(new_n242));
  AND2_X1   g041(.A1(new_n231), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(G169gat), .ZN(new_n244));
  INV_X1    g043(.A(G176gat), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n244), .A2(new_n245), .A3(KEYINPUT23), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT23), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n247), .B1(G169gat), .B2(G176gat), .ZN(new_n248));
  NAND4_X1  g047(.A1(new_n246), .A2(new_n248), .A3(KEYINPUT25), .A4(new_n223), .ZN(new_n249));
  NOR2_X1   g048(.A1(G183gat), .A2(G190gat), .ZN(new_n250));
  AND2_X1   g049(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n250), .B1(new_n251), .B2(G190gat), .ZN(new_n252));
  NAND2_X1  g051(.A1(G183gat), .A2(G190gat), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT64), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT24), .ZN(new_n255));
  AND3_X1   g054(.A1(new_n253), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n254), .B1(new_n253), .B2(new_n255), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n252), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT65), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n249), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  OAI211_X1 g059(.A(new_n252), .B(KEYINPUT65), .C1(new_n256), .C2(new_n257), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT25), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n253), .A2(new_n255), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n252), .A2(new_n263), .ZN(new_n264));
  AND3_X1   g063(.A1(new_n246), .A2(new_n248), .A3(new_n223), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  AOI22_X1  g065(.A1(new_n260), .A2(new_n261), .B1(new_n262), .B2(new_n266), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n220), .B1(new_n243), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n266), .A2(new_n262), .ZN(new_n269));
  INV_X1    g068(.A(new_n249), .ZN(new_n270));
  NAND3_X1  g069(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n271), .B1(G183gat), .B2(G190gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n263), .A2(KEYINPUT64), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n253), .A2(new_n254), .A3(new_n255), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n272), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n270), .B1(new_n275), .B2(KEYINPUT65), .ZN(new_n276));
  INV_X1    g075(.A(new_n261), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n269), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n231), .A2(new_n242), .ZN(new_n279));
  INV_X1    g078(.A(new_n220), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n278), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n268), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(G227gat), .ZN(new_n283));
  INV_X1    g082(.A(G233gat), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n282), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(KEYINPUT34), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT34), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n282), .A2(new_n289), .A3(new_n286), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT32), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n268), .A2(new_n285), .A3(new_n281), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(KEYINPUT69), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT69), .ZN(new_n295));
  NAND4_X1  g094(.A1(new_n268), .A2(new_n295), .A3(new_n285), .A4(new_n281), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n292), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(G15gat), .B(G43gat), .ZN(new_n298));
  XNOR2_X1  g097(.A(G71gat), .B(G99gat), .ZN(new_n299));
  XNOR2_X1  g098(.A(new_n298), .B(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  AND2_X1   g100(.A1(new_n301), .A2(KEYINPUT70), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n301), .A2(KEYINPUT70), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT33), .ZN(new_n304));
  NOR3_X1   g103(.A1(new_n302), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n294), .A2(new_n296), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n300), .B1(new_n307), .B2(KEYINPUT32), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n304), .ZN(new_n309));
  AOI221_X4 g108(.A(new_n291), .B1(new_n297), .B2(new_n306), .C1(new_n308), .C2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(new_n291), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n308), .A2(new_n309), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n297), .A2(new_n306), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n311), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n310), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(G225gat), .A2(G233gat), .ZN(new_n316));
  XNOR2_X1  g115(.A(new_n316), .B(KEYINPUT77), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT75), .ZN(new_n319));
  NAND2_X1  g118(.A1(G155gat), .A2(G162gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(KEYINPUT2), .ZN(new_n321));
  INV_X1    g120(.A(G141gat), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n322), .A2(G148gat), .ZN(new_n323));
  INV_X1    g122(.A(G148gat), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n324), .A2(G141gat), .ZN(new_n325));
  OAI211_X1 g124(.A(new_n319), .B(new_n321), .C1(new_n323), .C2(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(G155gat), .B(G162gat), .ZN(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n324), .A2(G141gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n322), .A2(G148gat), .ZN(new_n331));
  AOI21_X1  g130(.A(KEYINPUT75), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n327), .B1(new_n332), .B2(new_n321), .ZN(new_n333));
  OAI211_X1 g132(.A(new_n219), .B(new_n212), .C1(new_n329), .C2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n326), .A2(new_n328), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n332), .A2(new_n327), .A3(new_n321), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n207), .A2(new_n211), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n215), .A2(new_n218), .ZN(new_n338));
  OAI211_X1 g137(.A(new_n335), .B(new_n336), .C1(new_n337), .C2(new_n338), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n318), .B1(new_n334), .B2(new_n339), .ZN(new_n340));
  OR2_X1    g139(.A1(new_n340), .A2(KEYINPUT78), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT5), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n342), .B1(new_n340), .B2(KEYINPUT78), .ZN(new_n343));
  OAI21_X1  g142(.A(KEYINPUT3), .B1(new_n329), .B2(new_n333), .ZN(new_n344));
  XNOR2_X1  g143(.A(KEYINPUT76), .B(KEYINPUT3), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n335), .A2(new_n336), .A3(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n344), .A2(new_n280), .A3(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT4), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n339), .A2(new_n348), .ZN(new_n349));
  NAND4_X1  g148(.A1(new_n220), .A2(KEYINPUT4), .A3(new_n335), .A4(new_n336), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n347), .A2(new_n349), .A3(new_n318), .A4(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n341), .A2(new_n343), .A3(new_n351), .ZN(new_n352));
  OR2_X1    g151(.A1(new_n351), .A2(KEYINPUT5), .ZN(new_n353));
  XOR2_X1   g152(.A(G1gat), .B(G29gat), .Z(new_n354));
  XNOR2_X1  g153(.A(new_n354), .B(KEYINPUT0), .ZN(new_n355));
  XNOR2_X1  g154(.A(G57gat), .B(G85gat), .ZN(new_n356));
  XNOR2_X1  g155(.A(new_n355), .B(new_n356), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n352), .A2(new_n353), .A3(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT6), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n357), .B1(new_n352), .B2(new_n353), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  AOI211_X1 g161(.A(new_n359), .B(new_n357), .C1(new_n352), .C2(new_n353), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT73), .ZN(new_n365));
  AOI21_X1  g164(.A(KEYINPUT29), .B1(new_n278), .B2(new_n279), .ZN(new_n366));
  NAND2_X1  g165(.A1(G226gat), .A2(G233gat), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n365), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  AND2_X1   g168(.A1(G211gat), .A2(G218gat), .ZN(new_n370));
  NOR2_X1   g169(.A1(G211gat), .A2(G218gat), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  AND2_X1   g171(.A1(G197gat), .A2(G204gat), .ZN(new_n373));
  NOR2_X1   g172(.A1(G197gat), .A2(G204gat), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  AOI21_X1  g174(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n372), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  XNOR2_X1  g176(.A(G211gat), .B(G218gat), .ZN(new_n378));
  XNOR2_X1  g177(.A(G197gat), .B(G204gat), .ZN(new_n379));
  INV_X1    g178(.A(new_n376), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n378), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n377), .A2(new_n381), .ZN(new_n382));
  XNOR2_X1  g181(.A(new_n367), .B(KEYINPUT72), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n383), .B1(new_n243), .B2(new_n267), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n258), .A2(new_n259), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n385), .A2(new_n261), .A3(new_n270), .ZN(new_n386));
  AOI22_X1  g185(.A1(new_n386), .A2(new_n269), .B1(new_n231), .B2(new_n242), .ZN(new_n387));
  OAI211_X1 g186(.A(KEYINPUT73), .B(new_n367), .C1(new_n387), .C2(KEYINPUT29), .ZN(new_n388));
  NAND4_X1  g187(.A1(new_n369), .A2(new_n382), .A3(new_n384), .A4(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(new_n382), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n366), .A2(new_n383), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n387), .A2(new_n367), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n390), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  XNOR2_X1  g192(.A(G8gat), .B(G36gat), .ZN(new_n394));
  XNOR2_X1  g193(.A(G64gat), .B(G92gat), .ZN(new_n395));
  XOR2_X1   g194(.A(new_n394), .B(new_n395), .Z(new_n396));
  NAND3_X1  g195(.A1(new_n389), .A2(new_n393), .A3(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT30), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND4_X1  g198(.A1(new_n389), .A2(new_n393), .A3(KEYINPUT30), .A4(new_n396), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n389), .A2(new_n393), .ZN(new_n401));
  XNOR2_X1  g200(.A(new_n396), .B(KEYINPUT74), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n399), .A2(new_n400), .A3(new_n403), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n364), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n335), .A2(new_n336), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT3), .ZN(new_n407));
  AOI21_X1  g206(.A(KEYINPUT29), .B1(new_n377), .B2(new_n381), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n407), .B1(new_n408), .B2(KEYINPUT81), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT81), .ZN(new_n410));
  AOI211_X1 g209(.A(new_n410), .B(KEYINPUT29), .C1(new_n377), .C2(new_n381), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n406), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(KEYINPUT82), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT82), .ZN(new_n414));
  OAI211_X1 g213(.A(new_n414), .B(new_n406), .C1(new_n409), .C2(new_n411), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT29), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n382), .B1(new_n346), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(G228gat), .A2(G233gat), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n413), .A2(new_n415), .A3(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(G22gat), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n382), .A2(new_n416), .ZN(new_n422));
  AOI22_X1  g221(.A1(new_n422), .A2(new_n345), .B1(new_n335), .B2(new_n336), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n418), .B1(new_n423), .B2(new_n417), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(KEYINPUT80), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT80), .ZN(new_n426));
  OAI211_X1 g225(.A(new_n426), .B(new_n418), .C1(new_n423), .C2(new_n417), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n420), .A2(new_n421), .A3(new_n425), .A4(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT83), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n346), .A2(new_n416), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(new_n390), .ZN(new_n432));
  INV_X1    g231(.A(new_n345), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n406), .B1(new_n408), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n426), .B1(new_n435), .B2(new_n418), .ZN(new_n436));
  INV_X1    g235(.A(new_n427), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n438), .A2(KEYINPUT83), .A3(new_n421), .A4(new_n420), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n420), .A2(new_n425), .A3(new_n427), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(G22gat), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n430), .A2(new_n439), .A3(new_n441), .ZN(new_n442));
  XNOR2_X1  g241(.A(G78gat), .B(G106gat), .ZN(new_n443));
  XNOR2_X1  g242(.A(KEYINPUT31), .B(G50gat), .ZN(new_n444));
  XOR2_X1   g243(.A(new_n443), .B(new_n444), .Z(new_n445));
  XOR2_X1   g244(.A(new_n445), .B(KEYINPUT79), .Z(new_n446));
  NAND2_X1  g245(.A1(new_n442), .A2(new_n446), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n445), .B1(new_n440), .B2(G22gat), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(new_n428), .ZN(new_n449));
  AOI21_X1  g248(.A(KEYINPUT84), .B1(new_n447), .B2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT84), .ZN(new_n451));
  AOI221_X4 g250(.A(new_n451), .B1(new_n448), .B2(new_n428), .C1(new_n442), .C2(new_n446), .ZN(new_n452));
  OAI211_X1 g251(.A(new_n315), .B(new_n405), .C1(new_n450), .C2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT87), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n454), .A2(KEYINPUT35), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n447), .A2(new_n449), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(new_n451), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n447), .A2(KEYINPUT84), .A3(new_n449), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  XNOR2_X1  g259(.A(KEYINPUT87), .B(KEYINPUT35), .ZN(new_n461));
  NAND4_X1  g260(.A1(new_n460), .A2(new_n405), .A3(new_n315), .A4(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT37), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n389), .A2(new_n393), .A3(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(new_n396), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n463), .B1(new_n389), .B2(new_n393), .ZN(new_n467));
  OAI21_X1  g266(.A(KEYINPUT38), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n369), .A2(new_n390), .A3(new_n384), .A4(new_n388), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n382), .B1(new_n391), .B2(new_n392), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n469), .A2(KEYINPUT37), .A3(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT38), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n464), .A2(new_n471), .A3(new_n472), .A4(new_n402), .ZN(new_n473));
  NAND4_X1  g272(.A1(new_n364), .A2(new_n468), .A3(new_n397), .A4(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT40), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n347), .A2(new_n350), .A3(new_n349), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(new_n317), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n334), .A2(new_n318), .A3(new_n339), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT85), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n334), .A2(new_n339), .A3(KEYINPUT85), .A4(new_n318), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  AND3_X1   g281(.A1(new_n477), .A2(new_n482), .A3(KEYINPUT39), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT39), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n476), .A2(new_n484), .A3(new_n317), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(new_n357), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n475), .B1(new_n483), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n352), .A2(new_n353), .ZN(new_n488));
  INV_X1    g287(.A(new_n357), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n477), .A2(new_n482), .A3(KEYINPUT39), .ZN(new_n491));
  NAND4_X1  g290(.A1(new_n491), .A2(KEYINPUT40), .A3(new_n357), .A4(new_n485), .ZN(new_n492));
  AND3_X1   g291(.A1(new_n487), .A2(new_n490), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n404), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(KEYINPUT86), .ZN(new_n495));
  OAI211_X1 g294(.A(new_n474), .B(new_n495), .C1(new_n452), .C2(new_n450), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n494), .A2(KEYINPUT86), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AND2_X1   g297(.A1(new_n399), .A2(new_n403), .ZN(new_n499));
  OAI211_X1 g298(.A(new_n499), .B(new_n400), .C1(new_n363), .C2(new_n362), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n458), .A2(new_n459), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n312), .A2(new_n313), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(new_n291), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT71), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n312), .A2(new_n311), .A3(new_n313), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT36), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n503), .A2(new_n504), .A3(new_n505), .A4(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n504), .A2(new_n506), .ZN(new_n508));
  NAND2_X1  g307(.A1(KEYINPUT71), .A2(KEYINPUT36), .ZN(new_n509));
  OAI211_X1 g308(.A(new_n508), .B(new_n509), .C1(new_n310), .C2(new_n314), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n501), .A2(new_n507), .A3(new_n510), .ZN(new_n511));
  OAI211_X1 g310(.A(new_n456), .B(new_n462), .C1(new_n498), .C2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  XNOR2_X1  g312(.A(KEYINPUT95), .B(KEYINPUT13), .ZN(new_n514));
  NAND2_X1  g313(.A1(G229gat), .A2(G233gat), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n514), .B(new_n515), .ZN(new_n516));
  OAI21_X1  g315(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT14), .ZN(new_n518));
  INV_X1    g317(.A(G29gat), .ZN(new_n519));
  INV_X1    g318(.A(G36gat), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n518), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n521), .A2(KEYINPUT89), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT89), .ZN(new_n523));
  NOR2_X1   g322(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n523), .B1(new_n524), .B2(new_n520), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n517), .B1(new_n522), .B2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT90), .ZN(new_n527));
  AOI22_X1  g326(.A1(new_n526), .A2(new_n527), .B1(G29gat), .B2(G36gat), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n528), .B1(new_n527), .B2(new_n526), .ZN(new_n529));
  INV_X1    g328(.A(G50gat), .ZN(new_n530));
  OAI21_X1  g329(.A(KEYINPUT15), .B1(new_n530), .B2(G43gat), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n531), .B1(G43gat), .B2(new_n530), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n529), .A2(new_n532), .ZN(new_n533));
  AND2_X1   g332(.A1(new_n521), .A2(KEYINPUT92), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n521), .A2(KEYINPUT92), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n517), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n532), .B1(G29gat), .B2(G36gat), .ZN(new_n537));
  INV_X1    g336(.A(G43gat), .ZN(new_n538));
  AOI21_X1  g337(.A(KEYINPUT91), .B1(new_n538), .B2(G50gat), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT91), .ZN(new_n540));
  NOR3_X1   g339(.A1(new_n540), .A2(new_n530), .A3(G43gat), .ZN(new_n541));
  AOI211_X1 g340(.A(new_n539), .B(new_n541), .C1(G43gat), .C2(new_n530), .ZN(new_n542));
  OAI211_X1 g341(.A(new_n536), .B(new_n537), .C1(new_n542), .C2(KEYINPUT15), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n533), .A2(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(G15gat), .B(G22gat), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT16), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n545), .B1(new_n546), .B2(G1gat), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n547), .B1(G1gat), .B2(new_n545), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(G8gat), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n544), .A2(new_n549), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n550), .B(KEYINPUT93), .ZN(new_n551));
  INV_X1    g350(.A(new_n544), .ZN(new_n552));
  INV_X1    g351(.A(new_n549), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n516), .B1(new_n551), .B2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT96), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  OAI211_X1 g357(.A(KEYINPUT96), .B(new_n516), .C1(new_n551), .C2(new_n555), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT93), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n550), .B(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT17), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n544), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n533), .A2(KEYINPUT17), .A3(new_n543), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n564), .A2(new_n553), .A3(new_n565), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n562), .A2(new_n515), .A3(new_n566), .ZN(new_n567));
  AND3_X1   g366(.A1(new_n567), .A2(KEYINPUT94), .A3(KEYINPUT18), .ZN(new_n568));
  AOI21_X1  g367(.A(KEYINPUT18), .B1(new_n567), .B2(KEYINPUT94), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n560), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  XOR2_X1   g369(.A(G113gat), .B(G141gat), .Z(new_n571));
  XNOR2_X1  g370(.A(KEYINPUT88), .B(KEYINPUT11), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(G169gat), .B(G197gat), .ZN(new_n574));
  XOR2_X1   g373(.A(new_n573), .B(new_n574), .Z(new_n575));
  XOR2_X1   g374(.A(new_n575), .B(KEYINPUT12), .Z(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n570), .A2(new_n577), .ZN(new_n578));
  OAI211_X1 g377(.A(new_n560), .B(new_n576), .C1(new_n568), .C2(new_n569), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  XOR2_X1   g380(.A(G57gat), .B(G64gat), .Z(new_n582));
  INV_X1    g381(.A(G71gat), .ZN(new_n583));
  INV_X1    g382(.A(G78gat), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n582), .B1(KEYINPUT9), .B2(new_n585), .ZN(new_n586));
  XOR2_X1   g385(.A(G71gat), .B(G78gat), .Z(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(KEYINPUT100), .B(KEYINPUT7), .ZN(new_n589));
  INV_X1    g388(.A(G85gat), .ZN(new_n590));
  INV_X1    g389(.A(G92gat), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  OR2_X1    g391(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n589), .A2(new_n592), .ZN(new_n594));
  NAND2_X1  g393(.A1(G99gat), .A2(G106gat), .ZN(new_n595));
  AOI22_X1  g394(.A1(KEYINPUT8), .A2(new_n595), .B1(new_n590), .B2(new_n591), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n593), .A2(new_n594), .A3(new_n596), .ZN(new_n597));
  XOR2_X1   g396(.A(G99gat), .B(G106gat), .Z(new_n598));
  XNOR2_X1  g397(.A(new_n597), .B(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT102), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n588), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n599), .A2(new_n600), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n603), .A2(KEYINPUT10), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n599), .B(KEYINPUT101), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT10), .ZN(new_n606));
  NOR3_X1   g405(.A1(new_n605), .A2(new_n606), .A3(new_n588), .ZN(new_n607));
  INV_X1    g406(.A(G230gat), .ZN(new_n608));
  OAI22_X1  g407(.A1(new_n604), .A2(new_n607), .B1(new_n608), .B2(new_n284), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n608), .A2(new_n284), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n603), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(G120gat), .B(G148gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(G176gat), .B(G204gat), .ZN(new_n614));
  XOR2_X1   g413(.A(new_n613), .B(new_n614), .Z(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n612), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n609), .A2(new_n611), .A3(new_n615), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT103), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n617), .A2(KEYINPUT103), .A3(new_n618), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT21), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n588), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(G231gat), .A2(G233gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XOR2_X1   g426(.A(new_n627), .B(KEYINPUT20), .Z(new_n628));
  XNOR2_X1  g427(.A(G183gat), .B(G211gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n553), .B1(new_n624), .B2(new_n588), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n631), .B(KEYINPUT99), .ZN(new_n632));
  XOR2_X1   g431(.A(KEYINPUT97), .B(KEYINPUT19), .Z(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(KEYINPUT98), .ZN(new_n634));
  XOR2_X1   g433(.A(G127gat), .B(G155gat), .Z(new_n635));
  XNOR2_X1  g434(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n632), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n630), .B(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n605), .A2(new_n564), .A3(new_n565), .ZN(new_n640));
  AND2_X1   g439(.A1(G232gat), .A2(G233gat), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n641), .A2(KEYINPUT41), .ZN(new_n642));
  OAI211_X1 g441(.A(new_n640), .B(new_n642), .C1(new_n552), .C2(new_n605), .ZN(new_n643));
  XNOR2_X1  g442(.A(G190gat), .B(G218gat), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n643), .B(new_n644), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n641), .A2(KEYINPUT41), .ZN(new_n646));
  XNOR2_X1  g445(.A(G134gat), .B(G162gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(new_n648));
  OR2_X1    g447(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n645), .A2(new_n648), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n623), .A2(new_n639), .A3(new_n651), .ZN(new_n652));
  NOR3_X1   g451(.A1(new_n513), .A2(new_n581), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n653), .A2(new_n364), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g454(.A(KEYINPUT16), .B(G8gat), .Z(new_n656));
  NAND3_X1  g455(.A1(new_n653), .A2(new_n404), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n653), .A2(new_n404), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n658), .A2(G8gat), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(new_n657), .ZN(new_n660));
  MUX2_X1   g459(.A(new_n657), .B(new_n660), .S(KEYINPUT42), .Z(G1325gat));
  INV_X1    g460(.A(G15gat), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n653), .A2(new_n662), .A3(new_n315), .ZN(new_n663));
  AND2_X1   g462(.A1(new_n510), .A2(new_n507), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  AND2_X1   g464(.A1(new_n653), .A2(new_n665), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n663), .B1(new_n666), .B2(new_n662), .ZN(G1326gat));
  INV_X1    g466(.A(new_n460), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n653), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g468(.A(KEYINPUT43), .B(G22gat), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n669), .B(new_n670), .ZN(G1327gat));
  INV_X1    g470(.A(new_n651), .ZN(new_n672));
  AND2_X1   g471(.A1(new_n512), .A2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n623), .ZN(new_n674));
  NOR3_X1   g473(.A1(new_n581), .A2(new_n674), .A3(new_n639), .ZN(new_n675));
  AND2_X1   g474(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n676), .A2(new_n519), .A3(new_n364), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(KEYINPUT45), .ZN(new_n678));
  XOR2_X1   g477(.A(KEYINPUT105), .B(KEYINPUT44), .Z(new_n679));
  NAND2_X1  g478(.A1(new_n672), .A2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT104), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n681), .B1(new_n498), .B2(new_n511), .ZN(new_n682));
  INV_X1    g481(.A(new_n497), .ZN(new_n683));
  NAND4_X1  g482(.A1(new_n460), .A2(new_n683), .A3(new_n495), .A4(new_n474), .ZN(new_n684));
  NAND4_X1  g483(.A1(new_n684), .A2(new_n664), .A3(KEYINPUT104), .A4(new_n501), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n456), .A2(new_n462), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n680), .B1(new_n686), .B2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT44), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n690), .B1(new_n512), .B2(new_n672), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n675), .B1(new_n689), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(KEYINPUT106), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n687), .B1(new_n682), .B2(new_n685), .ZN(new_n694));
  OAI22_X1  g493(.A1(new_n673), .A2(new_n690), .B1(new_n694), .B2(new_n680), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT106), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n695), .A2(new_n696), .A3(new_n675), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n693), .A2(new_n364), .A3(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(G29gat), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n678), .A2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT107), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n678), .A2(new_n699), .A3(KEYINPUT107), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(G1328gat));
  NAND3_X1  g503(.A1(new_n676), .A2(new_n520), .A3(new_n404), .ZN(new_n705));
  AND2_X1   g504(.A1(KEYINPUT108), .A2(KEYINPUT46), .ZN(new_n706));
  NOR2_X1   g505(.A1(KEYINPUT108), .A2(KEYINPUT46), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n705), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  AND3_X1   g507(.A1(new_n693), .A2(new_n404), .A3(new_n697), .ZN(new_n709));
  OAI221_X1 g508(.A(new_n708), .B1(new_n706), .B2(new_n705), .C1(new_n709), .C2(new_n520), .ZN(G1329gat));
  NAND3_X1  g509(.A1(new_n693), .A2(new_n665), .A3(new_n697), .ZN(new_n711));
  INV_X1    g510(.A(new_n315), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n712), .A2(G43gat), .ZN(new_n713));
  AOI22_X1  g512(.A1(new_n711), .A2(G43gat), .B1(new_n676), .B2(new_n713), .ZN(new_n714));
  XNOR2_X1  g513(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n715));
  INV_X1    g514(.A(new_n692), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n538), .B1(new_n716), .B2(new_n665), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n676), .A2(new_n713), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(KEYINPUT47), .ZN(new_n719));
  OAI22_X1  g518(.A1(new_n714), .A2(new_n715), .B1(new_n717), .B2(new_n719), .ZN(G1330gat));
  OAI211_X1 g519(.A(new_n668), .B(new_n675), .C1(new_n689), .C2(new_n691), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT110), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND4_X1  g522(.A1(new_n695), .A2(KEYINPUT110), .A3(new_n668), .A4(new_n675), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n723), .A2(G50gat), .A3(new_n724), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n460), .A2(G50gat), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n676), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(KEYINPUT48), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT111), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n693), .A2(new_n668), .A3(new_n697), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(G50gat), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT48), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n727), .A2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n729), .A2(new_n730), .A3(new_n736), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n733), .B1(new_n725), .B2(new_n727), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n734), .B1(new_n731), .B2(G50gat), .ZN(new_n739));
  OAI21_X1  g538(.A(KEYINPUT111), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n737), .A2(new_n740), .ZN(G1331gat));
  NAND2_X1  g540(.A1(new_n686), .A2(new_n688), .ZN(new_n742));
  NOR4_X1   g541(.A1(new_n580), .A2(new_n623), .A3(new_n672), .A4(new_n638), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(new_n364), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(G57gat), .ZN(G1332gat));
  INV_X1    g546(.A(new_n404), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n744), .A2(new_n748), .ZN(new_n749));
  NOR2_X1   g548(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n750));
  AND2_X1   g549(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n749), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n752), .B1(new_n749), .B2(new_n750), .ZN(G1333gat));
  NOR3_X1   g552(.A1(new_n744), .A2(G71gat), .A3(new_n712), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n745), .A2(new_n665), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n754), .B1(G71gat), .B2(new_n755), .ZN(new_n756));
  XOR2_X1   g555(.A(KEYINPUT112), .B(KEYINPUT50), .Z(new_n757));
  XNOR2_X1  g556(.A(new_n756), .B(new_n757), .ZN(G1334gat));
  NOR2_X1   g557(.A1(new_n744), .A2(new_n460), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n759), .B(new_n584), .ZN(G1335gat));
  NOR3_X1   g559(.A1(new_n580), .A2(new_n623), .A3(new_n639), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n695), .A2(new_n364), .A3(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(G85gat), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n581), .A2(new_n638), .A3(new_n672), .ZN(new_n764));
  INV_X1    g563(.A(new_n764), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n742), .A2(KEYINPUT51), .A3(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(new_n766), .ZN(new_n767));
  AOI21_X1  g566(.A(KEYINPUT51), .B1(new_n742), .B2(new_n765), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n674), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n364), .A2(new_n590), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n763), .B1(new_n769), .B2(new_n770), .ZN(G1336gat));
  NOR2_X1   g570(.A1(new_n767), .A2(new_n768), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n772), .A2(new_n623), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n748), .A2(G92gat), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n695), .A2(new_n404), .A3(new_n761), .ZN(new_n775));
  AOI22_X1  g574(.A1(new_n773), .A2(new_n774), .B1(G92gat), .B2(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT52), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n776), .B(new_n777), .ZN(G1337gat));
  NOR2_X1   g577(.A1(new_n712), .A2(G99gat), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n695), .A2(new_n665), .A3(new_n761), .ZN(new_n780));
  AOI22_X1  g579(.A1(new_n773), .A2(new_n779), .B1(G99gat), .B2(new_n780), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n781), .B(KEYINPUT113), .ZN(G1338gat));
  NOR2_X1   g581(.A1(new_n460), .A2(G106gat), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n695), .A2(new_n668), .A3(new_n761), .ZN(new_n784));
  AOI22_X1  g583(.A1(new_n773), .A2(new_n783), .B1(G106gat), .B2(new_n784), .ZN(new_n785));
  XNOR2_X1  g584(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n785), .B(new_n786), .ZN(G1339gat));
  NOR2_X1   g586(.A1(new_n652), .A2(new_n580), .ZN(new_n788));
  INV_X1    g587(.A(new_n575), .ZN(new_n789));
  NOR3_X1   g588(.A1(new_n551), .A2(new_n555), .A3(new_n516), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n515), .B1(new_n562), .B2(new_n566), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n789), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT115), .ZN(new_n793));
  OR2_X1    g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n792), .A2(new_n793), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n579), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n651), .B1(new_n623), .B2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(new_n603), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n607), .B1(new_n799), .B2(new_n606), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n800), .A2(new_n610), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT54), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n615), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n800), .A2(new_n610), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n804), .A2(KEYINPUT54), .A3(new_n609), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT55), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n803), .A2(KEYINPUT55), .A3(new_n805), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n808), .A2(new_n618), .A3(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(new_n580), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n639), .B1(new_n798), .B2(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(new_n796), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(KEYINPUT116), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT116), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n796), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n815), .A2(new_n811), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(new_n672), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n788), .B1(new_n813), .B2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(new_n364), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n668), .A2(new_n712), .ZN(new_n822));
  INV_X1    g621(.A(new_n822), .ZN(new_n823));
  NOR4_X1   g622(.A1(new_n820), .A2(new_n821), .A3(new_n404), .A4(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(new_n580), .ZN(new_n825));
  XNOR2_X1  g624(.A(new_n825), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g625(.A1(new_n824), .A2(new_n674), .ZN(new_n827));
  XNOR2_X1  g626(.A(new_n827), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g627(.A1(new_n824), .A2(new_n639), .ZN(new_n829));
  XNOR2_X1  g628(.A(new_n829), .B(G127gat), .ZN(G1342gat));
  AOI21_X1  g629(.A(new_n651), .B1(KEYINPUT56), .B2(G134gat), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n824), .A2(new_n831), .ZN(new_n832));
  NOR2_X1   g631(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n833));
  XOR2_X1   g632(.A(new_n832), .B(new_n833), .Z(G1343gat));
  OAI21_X1  g633(.A(KEYINPUT57), .B1(new_n820), .B2(new_n460), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n810), .B1(new_n816), .B2(new_n796), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n651), .B1(new_n836), .B2(new_n815), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n581), .A2(new_n810), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n638), .B1(new_n838), .B2(new_n797), .ZN(new_n839));
  OAI22_X1  g638(.A1(new_n837), .A2(new_n839), .B1(new_n580), .B2(new_n652), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT57), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n840), .A2(new_n841), .A3(new_n668), .ZN(new_n842));
  NOR3_X1   g641(.A1(new_n665), .A2(new_n821), .A3(new_n404), .ZN(new_n843));
  XOR2_X1   g642(.A(new_n843), .B(KEYINPUT117), .Z(new_n844));
  NAND4_X1  g643(.A1(new_n835), .A2(new_n842), .A3(new_n580), .A4(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(G141gat), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n820), .A2(new_n460), .ZN(new_n847));
  NAND4_X1  g646(.A1(new_n847), .A2(new_n322), .A3(new_n580), .A4(new_n843), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(KEYINPUT58), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT58), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n846), .A2(new_n848), .A3(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n850), .A2(new_n852), .ZN(G1344gat));
  NAND2_X1  g652(.A1(new_n847), .A2(new_n843), .ZN(new_n854));
  INV_X1    g653(.A(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n855), .A2(new_n324), .A3(new_n674), .ZN(new_n856));
  NAND4_X1  g655(.A1(new_n835), .A2(new_n842), .A3(new_n674), .A4(new_n844), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT59), .ZN(new_n858));
  AND3_X1   g657(.A1(new_n857), .A2(new_n858), .A3(G148gat), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n858), .B1(new_n857), .B2(G148gat), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n856), .B1(new_n859), .B2(new_n860), .ZN(G1345gat));
  NAND4_X1  g660(.A1(new_n835), .A2(new_n842), .A3(new_n639), .A4(new_n844), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(G155gat), .ZN(new_n863));
  OR2_X1    g662(.A1(new_n638), .A2(G155gat), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n863), .B1(new_n854), .B2(new_n864), .ZN(G1346gat));
  INV_X1    g664(.A(G162gat), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n835), .A2(new_n842), .A3(new_n672), .A4(new_n844), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT118), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n866), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n869), .B1(new_n868), .B2(new_n867), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n855), .A2(new_n866), .A3(new_n672), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(G1347gat));
  NOR2_X1   g671(.A1(new_n748), .A2(new_n364), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n840), .A2(new_n822), .A3(new_n873), .ZN(new_n874));
  OAI21_X1  g673(.A(G169gat), .B1(new_n874), .B2(new_n581), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT120), .ZN(new_n876));
  AND2_X1   g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n875), .A2(new_n876), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n820), .A2(new_n823), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n879), .A2(KEYINPUT119), .A3(new_n873), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT119), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n874), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n580), .A2(new_n244), .ZN(new_n884));
  OAI22_X1  g683(.A1(new_n877), .A2(new_n878), .B1(new_n883), .B2(new_n884), .ZN(G1348gat));
  NAND4_X1  g684(.A1(new_n880), .A2(new_n882), .A3(new_n245), .A4(new_n674), .ZN(new_n886));
  OAI21_X1  g685(.A(G176gat), .B1(new_n874), .B2(new_n623), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT121), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n886), .A2(KEYINPUT121), .A3(new_n887), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n890), .A2(new_n891), .ZN(G1349gat));
  OAI21_X1  g691(.A(new_n232), .B1(new_n874), .B2(new_n638), .ZN(new_n893));
  INV_X1    g692(.A(new_n240), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n879), .A2(new_n894), .A3(new_n639), .A4(new_n873), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n893), .A2(new_n895), .A3(KEYINPUT122), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT123), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n897), .B1(new_n893), .B2(new_n895), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n896), .B1(new_n898), .B2(KEYINPUT60), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT122), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(KEYINPUT60), .ZN(new_n901));
  AOI211_X1 g700(.A(new_n897), .B(new_n901), .C1(new_n893), .C2(new_n895), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n899), .A2(new_n902), .ZN(G1350gat));
  OAI21_X1  g702(.A(G190gat), .B1(new_n874), .B2(new_n651), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT124), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  OAI211_X1 g705(.A(KEYINPUT124), .B(G190gat), .C1(new_n874), .C2(new_n651), .ZN(new_n907));
  OR2_X1    g706(.A1(KEYINPUT125), .A2(KEYINPUT61), .ZN(new_n908));
  NAND2_X1  g707(.A1(KEYINPUT125), .A2(KEYINPUT61), .ZN(new_n909));
  NAND4_X1  g708(.A1(new_n906), .A2(new_n907), .A3(new_n908), .A4(new_n909), .ZN(new_n910));
  NAND4_X1  g709(.A1(new_n880), .A2(new_n882), .A3(new_n236), .A4(new_n672), .ZN(new_n911));
  AND2_X1   g710(.A1(new_n906), .A2(new_n907), .ZN(new_n912));
  OAI211_X1 g711(.A(new_n910), .B(new_n911), .C1(new_n912), .C2(new_n908), .ZN(G1351gat));
  NOR3_X1   g712(.A1(new_n820), .A2(KEYINPUT57), .A3(new_n460), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n841), .B1(new_n840), .B2(new_n668), .ZN(new_n915));
  OAI21_X1  g714(.A(KEYINPUT126), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT126), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n835), .A2(new_n842), .A3(new_n917), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n664), .A2(new_n873), .ZN(new_n919));
  INV_X1    g718(.A(G197gat), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n581), .A2(new_n920), .ZN(new_n921));
  NAND4_X1  g720(.A1(new_n916), .A2(new_n918), .A3(new_n919), .A4(new_n921), .ZN(new_n922));
  AND3_X1   g721(.A1(new_n664), .A2(new_n668), .A3(new_n873), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n840), .A2(new_n923), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n920), .B1(new_n924), .B2(new_n581), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n922), .A2(new_n925), .ZN(G1352gat));
  NAND3_X1  g725(.A1(new_n916), .A2(new_n918), .A3(new_n919), .ZN(new_n927));
  OAI21_X1  g726(.A(G204gat), .B1(new_n927), .B2(new_n623), .ZN(new_n928));
  NOR3_X1   g727(.A1(new_n924), .A2(G204gat), .A3(new_n623), .ZN(new_n929));
  XNOR2_X1  g728(.A(new_n929), .B(KEYINPUT62), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n928), .A2(new_n930), .ZN(G1353gat));
  AND4_X1   g730(.A1(new_n639), .A2(new_n835), .A3(new_n842), .A4(new_n919), .ZN(new_n932));
  INV_X1    g731(.A(G211gat), .ZN(new_n933));
  OR3_X1    g732(.A1(new_n932), .A2(KEYINPUT63), .A3(new_n933), .ZN(new_n934));
  NAND4_X1  g733(.A1(new_n840), .A2(new_n933), .A3(new_n639), .A4(new_n923), .ZN(new_n935));
  XNOR2_X1  g734(.A(new_n935), .B(KEYINPUT127), .ZN(new_n936));
  OAI21_X1  g735(.A(KEYINPUT63), .B1(new_n932), .B2(new_n933), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n934), .A2(new_n936), .A3(new_n937), .ZN(G1354gat));
  INV_X1    g737(.A(G218gat), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n651), .A2(new_n939), .ZN(new_n940));
  NAND4_X1  g739(.A1(new_n916), .A2(new_n918), .A3(new_n919), .A4(new_n940), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n939), .B1(new_n924), .B2(new_n651), .ZN(new_n942));
  AND2_X1   g741(.A1(new_n941), .A2(new_n942), .ZN(G1355gat));
endmodule


