

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791;

  AND2_X1 U372 ( .A1(n643), .A2(n642), .ZN(n389) );
  AND2_X1 U373 ( .A1(n424), .A2(n423), .ZN(n420) );
  AND2_X1 U374 ( .A1(n409), .A2(n413), .ZN(n572) );
  XNOR2_X1 U375 ( .A(n615), .B(KEYINPUT107), .ZN(n622) );
  NOR2_X1 U376 ( .A1(n568), .A2(n711), .ZN(n569) );
  AND2_X1 U377 ( .A1(n614), .A2(n613), .ZN(n615) );
  XNOR2_X1 U378 ( .A(n633), .B(n351), .ZN(n598) );
  INV_X1 U379 ( .A(KEYINPUT87), .ZN(n351) );
  INV_X1 U380 ( .A(n601), .ZN(n496) );
  OR2_X1 U381 ( .A1(n392), .A2(n390), .ZN(n612) );
  XNOR2_X1 U382 ( .A(n495), .B(n494), .ZN(n601) );
  AND2_X1 U383 ( .A1(n439), .A2(n516), .ZN(n376) );
  XNOR2_X1 U384 ( .A(n446), .B(n445), .ZN(n749) );
  XNOR2_X1 U385 ( .A(n395), .B(n447), .ZN(n446) );
  XNOR2_X1 U386 ( .A(n411), .B(n489), .ZN(n499) );
  XNOR2_X1 U387 ( .A(n488), .B(n487), .ZN(n411) );
  NOR2_X2 U388 ( .A1(n649), .A2(n707), .ZN(n650) );
  XNOR2_X2 U389 ( .A(n584), .B(n583), .ZN(n763) );
  AND2_X2 U390 ( .A1(n409), .A2(n566), .ZN(n570) );
  INV_X2 U391 ( .A(KEYINPUT67), .ZN(n478) );
  XNOR2_X1 U392 ( .A(n482), .B(G104), .ZN(n498) );
  XNOR2_X1 U393 ( .A(n500), .B(n499), .ZN(n760) );
  NOR2_X1 U394 ( .A1(n718), .A2(n552), .ZN(n553) );
  XNOR2_X2 U395 ( .A(n396), .B(n522), .ZN(n563) );
  NAND2_X2 U396 ( .A1(n378), .A2(n377), .ZN(n396) );
  AND2_X2 U397 ( .A1(n375), .A2(n397), .ZN(n378) );
  INV_X1 U398 ( .A(n709), .ZN(n633) );
  XNOR2_X2 U399 ( .A(n387), .B(n647), .ZN(n386) );
  XNOR2_X1 U400 ( .A(G146), .B(G125), .ZN(n503) );
  NOR2_X1 U401 ( .A1(n661), .A2(n758), .ZN(n663) );
  NOR2_X1 U402 ( .A1(n655), .A2(n758), .ZN(n657) );
  INV_X1 U403 ( .A(n386), .ZN(n352) );
  NOR2_X1 U404 ( .A1(n380), .A2(n379), .ZN(n437) );
  XNOR2_X1 U405 ( .A(n619), .B(n618), .ZN(n787) );
  AND2_X1 U406 ( .A1(n607), .A2(n455), .ZN(n423) );
  XNOR2_X1 U407 ( .A(n567), .B(KEYINPUT99), .ZN(n379) );
  AND2_X1 U408 ( .A1(n405), .A2(n404), .ZN(n403) );
  OR2_X1 U409 ( .A1(n602), .A2(n429), .ZN(n617) );
  NOR2_X1 U410 ( .A1(n596), .A2(n595), .ZN(n597) );
  XNOR2_X1 U411 ( .A(n374), .B(n457), .ZN(n430) );
  NOR2_X2 U412 ( .A1(n556), .A2(n559), .ZN(n693) );
  XNOR2_X1 U413 ( .A(n483), .B(n775), .ZN(n445) );
  INV_X1 U414 ( .A(n589), .ZN(n573) );
  XNOR2_X1 U415 ( .A(n426), .B(n475), .ZN(n658) );
  XNOR2_X1 U416 ( .A(n431), .B(G137), .ZN(n449) );
  NAND2_X2 U417 ( .A1(n442), .A2(n439), .ZN(n604) );
  AND2_X1 U418 ( .A1(n438), .A2(n443), .ZN(n442) );
  INV_X1 U419 ( .A(G237), .ZN(n513) );
  XNOR2_X1 U420 ( .A(KEYINPUT3), .B(G119), .ZN(n489) );
  NAND2_X1 U421 ( .A1(n514), .A2(n644), .ZN(n443) );
  XNOR2_X1 U422 ( .A(G902), .B(KEYINPUT15), .ZN(n512) );
  AND2_X1 U423 ( .A1(n630), .A2(n629), .ZN(n424) );
  INV_X1 U424 ( .A(KEYINPUT34), .ZN(n406) );
  OR2_X1 U425 ( .A1(n651), .A2(G902), .ZN(n495) );
  INV_X1 U426 ( .A(KEYINPUT45), .ZN(n583) );
  XOR2_X1 U427 ( .A(KEYINPUT23), .B(G140), .Z(n471) );
  XNOR2_X1 U428 ( .A(n365), .B(n364), .ZN(n525) );
  NAND2_X1 U429 ( .A1(n464), .A2(n463), .ZN(n364) );
  XNOR2_X1 U430 ( .A(n366), .B(n465), .ZN(n365) );
  INV_X1 U431 ( .A(KEYINPUT69), .ZN(n466) );
  XNOR2_X1 U432 ( .A(n501), .B(G134), .ZN(n528) );
  XOR2_X1 U433 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n508) );
  XNOR2_X1 U434 ( .A(n591), .B(n410), .ZN(n608) );
  INV_X1 U435 ( .A(KEYINPUT70), .ZN(n410) );
  NAND2_X1 U436 ( .A1(n441), .A2(n512), .ZN(n440) );
  XNOR2_X1 U437 ( .A(n609), .B(KEYINPUT106), .ZN(n610) );
  NAND2_X1 U438 ( .A1(n394), .A2(n393), .ZN(n392) );
  NAND2_X1 U439 ( .A1(n355), .A2(G902), .ZN(n393) );
  INV_X1 U440 ( .A(KEYINPUT48), .ZN(n421) );
  XNOR2_X1 U441 ( .A(KEYINPUT16), .B(G122), .ZN(n497) );
  AND2_X1 U442 ( .A1(n525), .A2(G217), .ZN(n526) );
  XNOR2_X1 U443 ( .A(G116), .B(G107), .ZN(n523) );
  NAND2_X1 U444 ( .A1(n430), .A2(n603), .ZN(n429) );
  AND2_X1 U445 ( .A1(n373), .A2(n371), .ZN(n370) );
  XNOR2_X1 U446 ( .A(n533), .B(n412), .ZN(n556) );
  XNOR2_X1 U447 ( .A(G478), .B(KEYINPUT97), .ZN(n412) );
  INV_X1 U448 ( .A(KEYINPUT84), .ZN(n433) );
  NAND2_X1 U449 ( .A1(n779), .A2(G234), .ZN(n366) );
  INV_X1 U450 ( .A(KEYINPUT8), .ZN(n462) );
  OR2_X1 U451 ( .A1(n355), .A2(G902), .ZN(n391) );
  NAND2_X1 U452 ( .A1(n749), .A2(n355), .ZN(n394) );
  AND2_X1 U453 ( .A1(n358), .A2(n398), .ZN(n397) );
  NAND2_X1 U454 ( .A1(n399), .A2(n516), .ZN(n398) );
  INV_X1 U455 ( .A(n723), .ZN(n399) );
  XNOR2_X1 U456 ( .A(G131), .B(KEYINPUT73), .ZN(n484) );
  NOR2_X1 U457 ( .A1(n787), .A2(n790), .ZN(n422) );
  NOR2_X1 U458 ( .A1(G953), .A2(G237), .ZN(n541) );
  XNOR2_X1 U459 ( .A(G143), .B(G113), .ZN(n536) );
  XNOR2_X1 U460 ( .A(G104), .B(G122), .ZN(n537) );
  XOR2_X1 U461 ( .A(G131), .B(G140), .Z(n534) );
  NAND2_X1 U462 ( .A1(G234), .A2(G237), .ZN(n517) );
  NAND2_X1 U463 ( .A1(n372), .A2(KEYINPUT102), .ZN(n371) );
  XNOR2_X1 U464 ( .A(KEYINPUT103), .B(KEYINPUT30), .ZN(n457) );
  NAND2_X1 U465 ( .A1(n601), .A2(n723), .ZN(n374) );
  NAND2_X1 U466 ( .A1(n369), .A2(n360), .ZN(n367) );
  INV_X1 U467 ( .A(KEYINPUT102), .ZN(n368) );
  INV_X1 U468 ( .A(G902), .ZN(n545) );
  NAND2_X1 U469 ( .A1(n573), .A2(n712), .ZN(n417) );
  XNOR2_X1 U470 ( .A(n468), .B(n774), .ZN(n426) );
  XNOR2_X1 U471 ( .A(n534), .B(n481), .ZN(n775) );
  INV_X1 U472 ( .A(KEYINPUT90), .ZN(n481) );
  XNOR2_X1 U473 ( .A(n448), .B(n356), .ZN(n447) );
  XNOR2_X1 U474 ( .A(n480), .B(n479), .ZN(n448) );
  INV_X1 U475 ( .A(G146), .ZN(n479) );
  XNOR2_X1 U476 ( .A(n511), .B(n760), .ZN(n667) );
  NAND2_X1 U477 ( .A1(n452), .A2(n450), .ZN(n631) );
  NAND2_X1 U478 ( .A1(n451), .A2(n354), .ZN(n450) );
  AND2_X1 U479 ( .A1(n454), .A2(n453), .ZN(n452) );
  XNOR2_X1 U480 ( .A(n407), .B(KEYINPUT35), .ZN(n577) );
  NAND2_X1 U481 ( .A1(n402), .A2(n555), .ZN(n401) );
  XNOR2_X1 U482 ( .A(n611), .B(n610), .ZN(n614) );
  INV_X1 U483 ( .A(n612), .ZN(n416) );
  INV_X1 U484 ( .A(n417), .ZN(n369) );
  INV_X2 U485 ( .A(n496), .ZN(n715) );
  INV_X1 U486 ( .A(KEYINPUT83), .ZN(n415) );
  BUF_X1 U487 ( .A(n709), .Z(n413) );
  NAND2_X1 U488 ( .A1(n352), .A2(n382), .ZN(n653) );
  INV_X1 U489 ( .A(G472), .ZN(n383) );
  XNOR2_X1 U490 ( .A(n651), .B(KEYINPUT62), .ZN(n652) );
  INV_X2 U491 ( .A(G953), .ZN(n779) );
  NAND2_X1 U492 ( .A1(n352), .A2(n384), .ZN(n660) );
  INV_X1 U493 ( .A(G217), .ZN(n385) );
  XNOR2_X1 U494 ( .A(n658), .B(KEYINPUT120), .ZN(n659) );
  XNOR2_X1 U495 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U496 ( .A(n571), .B(KEYINPUT32), .ZN(n791) );
  NAND2_X1 U497 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U498 ( .A(n428), .B(n427), .ZN(n789) );
  INV_X1 U499 ( .A(KEYINPUT104), .ZN(n427) );
  NOR2_X1 U500 ( .A1(n617), .A2(n606), .ZN(n428) );
  XNOR2_X1 U501 ( .A(n751), .B(n750), .ZN(n752) );
  XNOR2_X1 U502 ( .A(n379), .B(n363), .ZN(G3) );
  AND2_X1 U503 ( .A1(G217), .A2(n476), .ZN(n353) );
  NOR2_X1 U504 ( .A1(n620), .A2(KEYINPUT39), .ZN(n354) );
  XNOR2_X1 U505 ( .A(KEYINPUT71), .B(G469), .ZN(n355) );
  XOR2_X1 U506 ( .A(KEYINPUT74), .B(KEYINPUT91), .Z(n356) );
  XOR2_X1 U507 ( .A(n595), .B(KEYINPUT19), .Z(n357) );
  NAND2_X1 U508 ( .A1(n588), .A2(n521), .ZN(n358) );
  AND2_X1 U509 ( .A1(n723), .A2(KEYINPUT19), .ZN(n359) );
  AND2_X1 U510 ( .A1(n416), .A2(n368), .ZN(n360) );
  AND2_X1 U511 ( .A1(n413), .A2(n711), .ZN(n361) );
  XOR2_X1 U512 ( .A(KEYINPUT86), .B(KEYINPUT33), .Z(n362) );
  XOR2_X1 U513 ( .A(G101), .B(KEYINPUT110), .Z(n363) );
  NAND2_X1 U514 ( .A1(n525), .A2(G221), .ZN(n468) );
  NAND2_X1 U515 ( .A1(n369), .A2(n416), .ZN(n600) );
  NAND2_X1 U516 ( .A1(n370), .A2(n367), .ZN(n602) );
  INV_X1 U517 ( .A(n416), .ZN(n372) );
  NAND2_X1 U518 ( .A1(n417), .A2(KEYINPUT102), .ZN(n373) );
  NAND2_X1 U519 ( .A1(n376), .A2(n442), .ZN(n375) );
  NAND2_X1 U520 ( .A1(n604), .A2(n359), .ZN(n377) );
  NAND2_X1 U521 ( .A1(n381), .A2(n558), .ZN(n380) );
  NAND2_X1 U522 ( .A1(n577), .A2(KEYINPUT44), .ZN(n381) );
  NOR2_X2 U523 ( .A1(n386), .A2(n650), .ZN(n753) );
  NOR2_X1 U524 ( .A1(n650), .A2(n383), .ZN(n382) );
  NOR2_X1 U525 ( .A1(n650), .A2(n385), .ZN(n384) );
  NAND2_X1 U526 ( .A1(n753), .A2(G210), .ZN(n669) );
  NAND2_X1 U527 ( .A1(n753), .A2(G475), .ZN(n677) );
  NAND2_X1 U528 ( .A1(n389), .A2(n388), .ZN(n387) );
  NAND2_X1 U529 ( .A1(n646), .A2(n645), .ZN(n388) );
  XNOR2_X2 U530 ( .A(n612), .B(KEYINPUT1), .ZN(n709) );
  NOR2_X1 U531 ( .A1(n749), .A2(n391), .ZN(n390) );
  XNOR2_X1 U532 ( .A(n395), .B(G146), .ZN(n492) );
  XNOR2_X1 U533 ( .A(n395), .B(n775), .ZN(n776) );
  XNOR2_X2 U534 ( .A(n449), .B(n528), .ZN(n395) );
  NAND2_X1 U535 ( .A1(n604), .A2(n723), .ZN(n595) );
  BUF_X1 U536 ( .A(n648), .Z(n706) );
  NOR2_X1 U537 ( .A1(n722), .A2(n406), .ZN(n402) );
  NAND2_X1 U538 ( .A1(n550), .A2(n592), .ZN(n444) );
  NAND2_X1 U539 ( .A1(n420), .A2(n419), .ZN(n418) );
  BUF_X1 U540 ( .A(n563), .Z(n555) );
  NAND2_X1 U541 ( .A1(n408), .A2(n605), .ZN(n407) );
  NAND2_X1 U542 ( .A1(n403), .A2(n401), .ZN(n408) );
  XNOR2_X1 U543 ( .A(n570), .B(n415), .ZN(n414) );
  BUF_X1 U544 ( .A(n791), .Z(n400) );
  NAND2_X1 U545 ( .A1(n563), .A2(n562), .ZN(n565) );
  NAND2_X1 U546 ( .A1(n722), .A2(n406), .ZN(n404) );
  NAND2_X1 U547 ( .A1(n552), .A2(n406), .ZN(n405) );
  XNOR2_X2 U548 ( .A(n565), .B(n564), .ZN(n409) );
  NAND2_X1 U549 ( .A1(n608), .A2(n715), .ZN(n611) );
  NOR2_X2 U550 ( .A1(n622), .A2(n357), .ZN(n694) );
  NAND2_X1 U551 ( .A1(n437), .A2(n435), .ZN(n434) );
  XNOR2_X1 U552 ( .A(n434), .B(n433), .ZN(n432) );
  NAND2_X1 U553 ( .A1(n414), .A2(n361), .ZN(n567) );
  XNOR2_X1 U554 ( .A(n431), .B(n501), .ZN(n505) );
  XNOR2_X1 U555 ( .A(n532), .B(n531), .ZN(n754) );
  NOR2_X2 U556 ( .A1(n709), .A2(n417), .ZN(n550) );
  NAND2_X1 U557 ( .A1(n413), .A2(n417), .ZN(n710) );
  XNOR2_X1 U558 ( .A(n418), .B(n421), .ZN(n640) );
  XNOR2_X1 U559 ( .A(n422), .B(KEYINPUT46), .ZN(n419) );
  XNOR2_X2 U560 ( .A(n425), .B(n477), .ZN(n589) );
  NOR2_X2 U561 ( .A1(n658), .A2(G902), .ZN(n425) );
  XNOR2_X2 U562 ( .A(n478), .B(KEYINPUT4), .ZN(n431) );
  NAND2_X1 U563 ( .A1(n432), .A2(n582), .ZN(n584) );
  XNOR2_X1 U564 ( .A(n576), .B(n436), .ZN(n435) );
  INV_X1 U565 ( .A(KEYINPUT65), .ZN(n436) );
  NAND2_X1 U566 ( .A1(n667), .A2(n514), .ZN(n438) );
  OR2_X1 U567 ( .A1(n667), .A2(n440), .ZN(n439) );
  INV_X1 U568 ( .A(n514), .ZN(n441) );
  XNOR2_X2 U569 ( .A(n444), .B(n362), .ZN(n722) );
  XNOR2_X2 U570 ( .A(n496), .B(KEYINPUT6), .ZN(n592) );
  INV_X1 U571 ( .A(n617), .ZN(n451) );
  NAND2_X1 U572 ( .A1(n620), .A2(KEYINPUT39), .ZN(n453) );
  NAND2_X1 U573 ( .A1(n617), .A2(KEYINPUT39), .ZN(n454) );
  NOR2_X1 U574 ( .A1(n616), .A2(n456), .ZN(n455) );
  INV_X1 U575 ( .A(n789), .ZN(n456) );
  XNOR2_X2 U576 ( .A(G110), .B(G107), .ZN(n482) );
  NOR2_X2 U577 ( .A1(n763), .A2(n773), .ZN(n648) );
  AND2_X1 U578 ( .A1(n608), .A2(n693), .ZN(n593) );
  INV_X1 U579 ( .A(KEYINPUT109), .ZN(n594) );
  XNOR2_X1 U580 ( .A(n749), .B(n748), .ZN(n750) );
  INV_X1 U581 ( .A(KEYINPUT63), .ZN(n656) );
  INV_X1 U582 ( .A(KEYINPUT121), .ZN(n662) );
  NAND2_X1 U583 ( .A1(n512), .A2(G234), .ZN(n458) );
  XNOR2_X1 U584 ( .A(n458), .B(KEYINPUT20), .ZN(n459) );
  XNOR2_X1 U585 ( .A(KEYINPUT92), .B(n459), .ZN(n476) );
  AND2_X1 U586 ( .A1(n476), .A2(G221), .ZN(n460) );
  XNOR2_X1 U587 ( .A(n460), .B(KEYINPUT21), .ZN(n712) );
  INV_X1 U588 ( .A(KEYINPUT68), .ZN(n461) );
  NAND2_X1 U589 ( .A1(KEYINPUT8), .A2(n461), .ZN(n464) );
  NAND2_X1 U590 ( .A1(n462), .A2(KEYINPUT68), .ZN(n463) );
  INV_X1 U591 ( .A(KEYINPUT79), .ZN(n465) );
  XNOR2_X1 U592 ( .A(n466), .B(KEYINPUT10), .ZN(n467) );
  XNOR2_X1 U593 ( .A(n503), .B(n467), .ZN(n774) );
  XNOR2_X1 U594 ( .A(G137), .B(G110), .ZN(n470) );
  INV_X1 U595 ( .A(KEYINPUT24), .ZN(n469) );
  XNOR2_X1 U596 ( .A(n470), .B(n469), .ZN(n472) );
  XNOR2_X1 U597 ( .A(n472), .B(n471), .ZN(n474) );
  XNOR2_X1 U598 ( .A(G128), .B(G119), .ZN(n473) );
  XNOR2_X1 U599 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X1 U600 ( .A(KEYINPUT25), .B(n353), .ZN(n477) );
  XNOR2_X2 U601 ( .A(G143), .B(G128), .ZN(n501) );
  NAND2_X1 U602 ( .A1(G227), .A2(n779), .ZN(n480) );
  XNOR2_X1 U603 ( .A(n498), .B(G101), .ZN(n483) );
  XNOR2_X1 U604 ( .A(n484), .B(KEYINPUT5), .ZN(n486) );
  AND2_X1 U605 ( .A1(n541), .A2(G210), .ZN(n485) );
  XNOR2_X1 U606 ( .A(n486), .B(n485), .ZN(n490) );
  XNOR2_X2 U607 ( .A(G116), .B(G113), .ZN(n488) );
  XNOR2_X2 U608 ( .A(G101), .B(KEYINPUT72), .ZN(n487) );
  XNOR2_X1 U609 ( .A(n499), .B(n490), .ZN(n491) );
  XNOR2_X1 U610 ( .A(n492), .B(n491), .ZN(n651) );
  INV_X1 U611 ( .A(KEYINPUT93), .ZN(n493) );
  XNOR2_X1 U612 ( .A(n493), .B(G472), .ZN(n494) );
  XNOR2_X1 U613 ( .A(n498), .B(n497), .ZN(n500) );
  XNOR2_X1 U614 ( .A(KEYINPUT75), .B(KEYINPUT76), .ZN(n502) );
  XNOR2_X1 U615 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U616 ( .A(n505), .B(n504), .ZN(n510) );
  NAND2_X1 U617 ( .A1(G224), .A2(n779), .ZN(n506) );
  XNOR2_X1 U618 ( .A(n506), .B(KEYINPUT88), .ZN(n507) );
  XNOR2_X1 U619 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U620 ( .A(n510), .B(n509), .ZN(n511) );
  INV_X1 U621 ( .A(n512), .ZN(n644) );
  NAND2_X1 U622 ( .A1(n545), .A2(n513), .ZN(n515) );
  AND2_X1 U623 ( .A1(n515), .A2(G210), .ZN(n514) );
  NAND2_X1 U624 ( .A1(n515), .A2(G214), .ZN(n723) );
  INV_X1 U625 ( .A(KEYINPUT19), .ZN(n516) );
  XNOR2_X1 U626 ( .A(n517), .B(KEYINPUT14), .ZN(n519) );
  NAND2_X1 U627 ( .A1(n519), .A2(G952), .ZN(n518) );
  XNOR2_X1 U628 ( .A(n518), .B(KEYINPUT89), .ZN(n735) );
  NAND2_X1 U629 ( .A1(n735), .A2(n779), .ZN(n588) );
  NAND2_X1 U630 ( .A1(G902), .A2(n519), .ZN(n585) );
  INV_X1 U631 ( .A(n585), .ZN(n520) );
  NOR2_X1 U632 ( .A1(G898), .A2(n779), .ZN(n761) );
  NAND2_X1 U633 ( .A1(n520), .A2(n761), .ZN(n521) );
  INV_X1 U634 ( .A(KEYINPUT0), .ZN(n522) );
  INV_X1 U635 ( .A(n555), .ZN(n552) );
  XOR2_X1 U636 ( .A(KEYINPUT96), .B(G122), .Z(n524) );
  XNOR2_X1 U637 ( .A(n524), .B(n523), .ZN(n527) );
  XNOR2_X1 U638 ( .A(n527), .B(n526), .ZN(n532) );
  BUF_X1 U639 ( .A(n528), .Z(n530) );
  XNOR2_X1 U640 ( .A(KEYINPUT9), .B(KEYINPUT7), .ZN(n529) );
  NOR2_X1 U641 ( .A1(n754), .A2(G902), .ZN(n533) );
  INV_X1 U642 ( .A(n556), .ZN(n560) );
  INV_X1 U643 ( .A(n534), .ZN(n535) );
  XOR2_X1 U644 ( .A(n536), .B(n535), .Z(n540) );
  XOR2_X1 U645 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n538) );
  XNOR2_X1 U646 ( .A(n538), .B(n537), .ZN(n539) );
  XOR2_X1 U647 ( .A(n540), .B(n539), .Z(n544) );
  AND2_X1 U648 ( .A1(G214), .A2(n541), .ZN(n542) );
  XNOR2_X1 U649 ( .A(n774), .B(n542), .ZN(n543) );
  XNOR2_X1 U650 ( .A(n544), .B(n543), .ZN(n675) );
  NAND2_X1 U651 ( .A1(n675), .A2(n545), .ZN(n549) );
  XOR2_X1 U652 ( .A(KEYINPUT95), .B(KEYINPUT13), .Z(n547) );
  XNOR2_X1 U653 ( .A(KEYINPUT94), .B(G475), .ZN(n546) );
  XNOR2_X1 U654 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U655 ( .A(n549), .B(n548), .ZN(n559) );
  NOR2_X1 U656 ( .A1(n560), .A2(n559), .ZN(n605) );
  BUF_X1 U657 ( .A(n550), .Z(n551) );
  NAND2_X1 U658 ( .A1(n551), .A2(n715), .ZN(n718) );
  XNOR2_X1 U659 ( .A(n553), .B(KEYINPUT31), .ZN(n698) );
  NOR2_X1 U660 ( .A1(n600), .A2(n715), .ZN(n554) );
  NAND2_X1 U661 ( .A1(n555), .A2(n554), .ZN(n686) );
  NAND2_X1 U662 ( .A1(n698), .A2(n686), .ZN(n557) );
  AND2_X1 U663 ( .A1(n556), .A2(n559), .ZN(n689) );
  NOR2_X1 U664 ( .A1(n689), .A2(n693), .ZN(n728) );
  INV_X1 U665 ( .A(n728), .ZN(n626) );
  NAND2_X1 U666 ( .A1(n557), .A2(n626), .ZN(n558) );
  NAND2_X1 U667 ( .A1(n560), .A2(n559), .ZN(n726) );
  INV_X1 U668 ( .A(n712), .ZN(n561) );
  NOR2_X1 U669 ( .A1(n726), .A2(n561), .ZN(n562) );
  INV_X1 U670 ( .A(KEYINPUT22), .ZN(n564) );
  INV_X1 U671 ( .A(n592), .ZN(n566) );
  XOR2_X1 U672 ( .A(KEYINPUT98), .B(n589), .Z(n711) );
  INV_X1 U673 ( .A(n598), .ZN(n568) );
  XNOR2_X1 U674 ( .A(n572), .B(KEYINPUT100), .ZN(n575) );
  NOR2_X1 U675 ( .A1(n715), .A2(n573), .ZN(n574) );
  NAND2_X1 U676 ( .A1(n575), .A2(n574), .ZN(n673) );
  NAND2_X1 U677 ( .A1(n791), .A2(n673), .ZN(n578) );
  NAND2_X1 U678 ( .A1(n578), .A2(KEYINPUT44), .ZN(n576) );
  BUF_X1 U679 ( .A(n577), .Z(n788) );
  NOR2_X1 U680 ( .A1(n788), .A2(KEYINPUT44), .ZN(n581) );
  BUF_X1 U681 ( .A(n578), .Z(n579) );
  INV_X1 U682 ( .A(n579), .ZN(n580) );
  NAND2_X1 U683 ( .A1(n581), .A2(n580), .ZN(n582) );
  NOR2_X1 U684 ( .A1(G900), .A2(n585), .ZN(n586) );
  NAND2_X1 U685 ( .A1(G953), .A2(n586), .ZN(n587) );
  NAND2_X1 U686 ( .A1(n588), .A2(n587), .ZN(n603) );
  AND2_X1 U687 ( .A1(n712), .A2(n603), .ZN(n590) );
  NAND2_X1 U688 ( .A1(n590), .A2(n589), .ZN(n591) );
  NAND2_X1 U689 ( .A1(n593), .A2(n592), .ZN(n632) );
  XNOR2_X1 U690 ( .A(n632), .B(n594), .ZN(n596) );
  XNOR2_X1 U691 ( .A(n597), .B(KEYINPUT36), .ZN(n599) );
  NAND2_X1 U692 ( .A1(n599), .A2(n598), .ZN(n704) );
  XNOR2_X1 U693 ( .A(n704), .B(KEYINPUT82), .ZN(n607) );
  NAND2_X1 U694 ( .A1(n605), .A2(n604), .ZN(n606) );
  INV_X1 U695 ( .A(KEYINPUT28), .ZN(n609) );
  XNOR2_X1 U696 ( .A(n372), .B(KEYINPUT105), .ZN(n613) );
  INV_X1 U697 ( .A(KEYINPUT78), .ZN(n627) );
  AND2_X1 U698 ( .A1(n694), .A2(n627), .ZN(n616) );
  XOR2_X1 U699 ( .A(KEYINPUT108), .B(KEYINPUT40), .Z(n619) );
  XNOR2_X1 U700 ( .A(n604), .B(KEYINPUT38), .ZN(n620) );
  NAND2_X1 U701 ( .A1(n631), .A2(n693), .ZN(n618) );
  INV_X1 U702 ( .A(n620), .ZN(n724) );
  NAND2_X1 U703 ( .A1(n724), .A2(n723), .ZN(n727) );
  NOR2_X1 U704 ( .A1(n727), .A2(n726), .ZN(n621) );
  XNOR2_X1 U705 ( .A(n621), .B(KEYINPUT41), .ZN(n737) );
  NOR2_X1 U706 ( .A1(n737), .A2(n622), .ZN(n623) );
  XNOR2_X1 U707 ( .A(n623), .B(KEYINPUT42), .ZN(n790) );
  NAND2_X1 U708 ( .A1(n694), .A2(n626), .ZN(n624) );
  XNOR2_X1 U709 ( .A(n624), .B(KEYINPUT47), .ZN(n625) );
  NAND2_X1 U710 ( .A1(n625), .A2(KEYINPUT78), .ZN(n630) );
  NAND2_X1 U711 ( .A1(n626), .A2(KEYINPUT47), .ZN(n628) );
  NAND2_X1 U712 ( .A1(n628), .A2(n627), .ZN(n629) );
  NAND2_X1 U713 ( .A1(n631), .A2(n689), .ZN(n705) );
  XOR2_X1 U714 ( .A(KEYINPUT43), .B(KEYINPUT101), .Z(n636) );
  NOR2_X1 U715 ( .A1(n633), .A2(n632), .ZN(n634) );
  NAND2_X1 U716 ( .A1(n634), .A2(n723), .ZN(n635) );
  XNOR2_X1 U717 ( .A(n636), .B(n635), .ZN(n638) );
  INV_X1 U718 ( .A(n604), .ZN(n637) );
  NAND2_X1 U719 ( .A1(n638), .A2(n637), .ZN(n664) );
  AND2_X1 U720 ( .A1(n705), .A2(n664), .ZN(n639) );
  NAND2_X1 U721 ( .A1(n640), .A2(n639), .ZN(n773) );
  AND2_X1 U722 ( .A1(KEYINPUT80), .A2(n644), .ZN(n641) );
  NAND2_X1 U723 ( .A1(n648), .A2(n641), .ZN(n643) );
  INV_X1 U724 ( .A(KEYINPUT2), .ZN(n707) );
  OR2_X1 U725 ( .A1(n512), .A2(n707), .ZN(n642) );
  NAND2_X1 U726 ( .A1(n648), .A2(n644), .ZN(n646) );
  INV_X1 U727 ( .A(KEYINPUT80), .ZN(n645) );
  INV_X1 U728 ( .A(KEYINPUT64), .ZN(n647) );
  INV_X1 U729 ( .A(n706), .ZN(n649) );
  XNOR2_X1 U730 ( .A(n653), .B(n652), .ZN(n655) );
  INV_X1 U731 ( .A(G952), .ZN(n654) );
  AND2_X1 U732 ( .A1(n654), .A2(G953), .ZN(n758) );
  XNOR2_X1 U733 ( .A(n657), .B(n656), .ZN(G57) );
  XNOR2_X1 U734 ( .A(n660), .B(n659), .ZN(n661) );
  XNOR2_X1 U735 ( .A(n663), .B(n662), .ZN(G66) );
  XNOR2_X1 U736 ( .A(n664), .B(G140), .ZN(G42) );
  XOR2_X1 U737 ( .A(KEYINPUT85), .B(KEYINPUT54), .Z(n665) );
  XNOR2_X1 U738 ( .A(n665), .B(KEYINPUT55), .ZN(n666) );
  XNOR2_X1 U739 ( .A(n667), .B(n666), .ZN(n668) );
  XNOR2_X1 U740 ( .A(n669), .B(n668), .ZN(n670) );
  INV_X1 U741 ( .A(n758), .ZN(n678) );
  NAND2_X1 U742 ( .A1(n670), .A2(n678), .ZN(n672) );
  XNOR2_X1 U743 ( .A(KEYINPUT81), .B(KEYINPUT56), .ZN(n671) );
  XNOR2_X1 U744 ( .A(n672), .B(n671), .ZN(G51) );
  XNOR2_X1 U745 ( .A(n673), .B(G110), .ZN(G12) );
  XOR2_X1 U746 ( .A(KEYINPUT66), .B(KEYINPUT59), .Z(n674) );
  XNOR2_X1 U747 ( .A(n675), .B(n674), .ZN(n676) );
  XNOR2_X1 U748 ( .A(n677), .B(n676), .ZN(n679) );
  NAND2_X1 U749 ( .A1(n679), .A2(n678), .ZN(n681) );
  INV_X1 U750 ( .A(KEYINPUT60), .ZN(n680) );
  XNOR2_X1 U751 ( .A(n681), .B(n680), .ZN(G60) );
  INV_X1 U752 ( .A(n693), .ZN(n696) );
  NOR2_X1 U753 ( .A1(n696), .A2(n686), .ZN(n683) );
  XNOR2_X1 U754 ( .A(G104), .B(KEYINPUT111), .ZN(n682) );
  XNOR2_X1 U755 ( .A(n683), .B(n682), .ZN(G6) );
  XOR2_X1 U756 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n685) );
  XNOR2_X1 U757 ( .A(G107), .B(KEYINPUT112), .ZN(n684) );
  XNOR2_X1 U758 ( .A(n685), .B(n684), .ZN(n688) );
  INV_X1 U759 ( .A(n689), .ZN(n699) );
  NOR2_X1 U760 ( .A1(n686), .A2(n699), .ZN(n687) );
  XOR2_X1 U761 ( .A(n688), .B(n687), .Z(G9) );
  XOR2_X1 U762 ( .A(KEYINPUT113), .B(KEYINPUT29), .Z(n691) );
  NAND2_X1 U763 ( .A1(n694), .A2(n689), .ZN(n690) );
  XNOR2_X1 U764 ( .A(n691), .B(n690), .ZN(n692) );
  XOR2_X1 U765 ( .A(G128), .B(n692), .Z(G30) );
  NAND2_X1 U766 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U767 ( .A(n695), .B(G146), .ZN(G48) );
  NOR2_X1 U768 ( .A1(n696), .A2(n698), .ZN(n697) );
  XOR2_X1 U769 ( .A(G113), .B(n697), .Z(G15) );
  NOR2_X1 U770 ( .A1(n699), .A2(n698), .ZN(n701) );
  XNOR2_X1 U771 ( .A(KEYINPUT114), .B(KEYINPUT115), .ZN(n700) );
  XNOR2_X1 U772 ( .A(n701), .B(n700), .ZN(n702) );
  XNOR2_X1 U773 ( .A(G116), .B(n702), .ZN(G18) );
  XOR2_X1 U774 ( .A(G125), .B(KEYINPUT37), .Z(n703) );
  XNOR2_X1 U775 ( .A(n704), .B(n703), .ZN(G27) );
  XNOR2_X1 U776 ( .A(G134), .B(n705), .ZN(G36) );
  NOR2_X1 U777 ( .A1(n706), .A2(KEYINPUT77), .ZN(n708) );
  XNOR2_X1 U778 ( .A(n708), .B(n707), .ZN(n744) );
  XNOR2_X1 U779 ( .A(n710), .B(KEYINPUT50), .ZN(n717) );
  NOR2_X1 U780 ( .A1(n712), .A2(n711), .ZN(n713) );
  XOR2_X1 U781 ( .A(KEYINPUT49), .B(n713), .Z(n714) );
  NOR2_X1 U782 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U783 ( .A1(n717), .A2(n716), .ZN(n719) );
  NAND2_X1 U784 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U785 ( .A(KEYINPUT51), .B(n720), .ZN(n721) );
  NOR2_X1 U786 ( .A1(n737), .A2(n721), .ZN(n733) );
  BUF_X1 U787 ( .A(n722), .Z(n738) );
  NOR2_X1 U788 ( .A1(n724), .A2(n723), .ZN(n725) );
  NOR2_X1 U789 ( .A1(n726), .A2(n725), .ZN(n730) );
  NOR2_X1 U790 ( .A1(n728), .A2(n727), .ZN(n729) );
  NOR2_X1 U791 ( .A1(n730), .A2(n729), .ZN(n731) );
  NOR2_X1 U792 ( .A1(n738), .A2(n731), .ZN(n732) );
  NOR2_X1 U793 ( .A1(n733), .A2(n732), .ZN(n734) );
  XOR2_X1 U794 ( .A(KEYINPUT52), .B(n734), .Z(n736) );
  NAND2_X1 U795 ( .A1(n736), .A2(n735), .ZN(n741) );
  NOR2_X1 U796 ( .A1(n738), .A2(n737), .ZN(n739) );
  XOR2_X1 U797 ( .A(KEYINPUT116), .B(n739), .Z(n740) );
  NAND2_X1 U798 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U799 ( .A(n742), .B(KEYINPUT117), .ZN(n743) );
  NAND2_X1 U800 ( .A1(n744), .A2(n743), .ZN(n745) );
  NOR2_X1 U801 ( .A1(G953), .A2(n745), .ZN(n747) );
  XNOR2_X1 U802 ( .A(KEYINPUT53), .B(KEYINPUT118), .ZN(n746) );
  XNOR2_X1 U803 ( .A(n747), .B(n746), .ZN(G75) );
  NAND2_X1 U804 ( .A1(n753), .A2(G469), .ZN(n751) );
  XOR2_X1 U805 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n748) );
  NOR2_X1 U806 ( .A1(n758), .A2(n752), .ZN(G54) );
  NAND2_X1 U807 ( .A1(n753), .A2(G478), .ZN(n756) );
  XOR2_X1 U808 ( .A(n754), .B(KEYINPUT119), .Z(n755) );
  XNOR2_X1 U809 ( .A(n756), .B(n755), .ZN(n757) );
  NOR2_X1 U810 ( .A1(n758), .A2(n757), .ZN(G63) );
  XNOR2_X1 U811 ( .A(KEYINPUT125), .B(KEYINPUT122), .ZN(n772) );
  XOR2_X1 U812 ( .A(KEYINPUT123), .B(KEYINPUT124), .Z(n759) );
  XNOR2_X1 U813 ( .A(n760), .B(n759), .ZN(n762) );
  NOR2_X1 U814 ( .A1(n762), .A2(n761), .ZN(n770) );
  BUF_X1 U815 ( .A(n763), .Z(n764) );
  NOR2_X1 U816 ( .A1(n764), .A2(G953), .ZN(n768) );
  NAND2_X1 U817 ( .A1(G953), .A2(G224), .ZN(n765) );
  XNOR2_X1 U818 ( .A(KEYINPUT61), .B(n765), .ZN(n766) );
  AND2_X1 U819 ( .A1(n766), .A2(G898), .ZN(n767) );
  NOR2_X1 U820 ( .A1(n768), .A2(n767), .ZN(n769) );
  XNOR2_X1 U821 ( .A(n770), .B(n769), .ZN(n771) );
  XNOR2_X1 U822 ( .A(n772), .B(n771), .ZN(G69) );
  BUF_X1 U823 ( .A(n773), .Z(n778) );
  XOR2_X1 U824 ( .A(KEYINPUT126), .B(n774), .Z(n777) );
  XNOR2_X1 U825 ( .A(n777), .B(n776), .ZN(n781) );
  XNOR2_X1 U826 ( .A(n778), .B(n781), .ZN(n780) );
  NAND2_X1 U827 ( .A1(n780), .A2(n779), .ZN(n786) );
  XNOR2_X1 U828 ( .A(G227), .B(n781), .ZN(n782) );
  NAND2_X1 U829 ( .A1(n782), .A2(G900), .ZN(n783) );
  XOR2_X1 U830 ( .A(KEYINPUT127), .B(n783), .Z(n784) );
  NAND2_X1 U831 ( .A1(G953), .A2(n784), .ZN(n785) );
  NAND2_X1 U832 ( .A1(n786), .A2(n785), .ZN(G72) );
  XOR2_X1 U833 ( .A(n787), .B(G131), .Z(G33) );
  XOR2_X1 U834 ( .A(G122), .B(n788), .Z(G24) );
  XNOR2_X1 U835 ( .A(G143), .B(n789), .ZN(G45) );
  XOR2_X1 U836 ( .A(G137), .B(n790), .Z(G39) );
  XNOR2_X1 U837 ( .A(n400), .B(G119), .ZN(G21) );
endmodule

