

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583;

  XNOR2_X1 U322 ( .A(n381), .B(n380), .ZN(n523) );
  XNOR2_X1 U323 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U324 ( .A(n449), .B(n448), .Z(n290) );
  XOR2_X1 U325 ( .A(n419), .B(n361), .Z(n291) );
  XNOR2_X1 U326 ( .A(n379), .B(KEYINPUT48), .ZN(n380) );
  XNOR2_X1 U327 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U328 ( .A(KEYINPUT55), .B(KEYINPUT116), .ZN(n425) );
  NOR2_X1 U329 ( .A1(n407), .A2(n482), .ZN(n562) );
  XNOR2_X1 U330 ( .A(n426), .B(n425), .ZN(n445) );
  XOR2_X1 U331 ( .A(KEYINPUT77), .B(n550), .Z(n537) );
  XOR2_X1 U332 ( .A(G211GAT), .B(G71GAT), .Z(n293) );
  XNOR2_X1 U333 ( .A(G127GAT), .B(G183GAT), .ZN(n292) );
  XNOR2_X1 U334 ( .A(n293), .B(n292), .ZN(n306) );
  XOR2_X1 U335 ( .A(KEYINPUT13), .B(G57GAT), .Z(n340) );
  XOR2_X1 U336 ( .A(G8GAT), .B(KEYINPUT78), .Z(n315) );
  XOR2_X1 U337 ( .A(n340), .B(n315), .Z(n295) );
  NAND2_X1 U338 ( .A1(G231GAT), .A2(G233GAT), .ZN(n294) );
  XNOR2_X1 U339 ( .A(n295), .B(n294), .ZN(n299) );
  XOR2_X1 U340 ( .A(G64GAT), .B(KEYINPUT15), .Z(n297) );
  XNOR2_X1 U341 ( .A(KEYINPUT12), .B(KEYINPUT79), .ZN(n296) );
  XNOR2_X1 U342 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U343 ( .A(n299), .B(n298), .Z(n304) );
  XOR2_X1 U344 ( .A(G15GAT), .B(G1GAT), .Z(n323) );
  XOR2_X1 U345 ( .A(KEYINPUT14), .B(G78GAT), .Z(n301) );
  XNOR2_X1 U346 ( .A(G22GAT), .B(G155GAT), .ZN(n300) );
  XNOR2_X1 U347 ( .A(n301), .B(n300), .ZN(n302) );
  XNOR2_X1 U348 ( .A(n323), .B(n302), .ZN(n303) );
  XNOR2_X1 U349 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U350 ( .A(n306), .B(n305), .ZN(n576) );
  INV_X1 U351 ( .A(n576), .ZN(n547) );
  XNOR2_X1 U352 ( .A(KEYINPUT54), .B(KEYINPUT115), .ZN(n383) );
  XNOR2_X1 U353 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n307) );
  XNOR2_X1 U354 ( .A(n307), .B(G211GAT), .ZN(n412) );
  XNOR2_X1 U355 ( .A(G36GAT), .B(G190GAT), .ZN(n308) );
  XNOR2_X1 U356 ( .A(n308), .B(G218GAT), .ZN(n357) );
  XNOR2_X1 U357 ( .A(n412), .B(n357), .ZN(n319) );
  XOR2_X1 U358 ( .A(G176GAT), .B(G64GAT), .Z(n341) );
  XOR2_X1 U359 ( .A(n341), .B(G92GAT), .Z(n313) );
  XOR2_X1 U360 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n310) );
  XNOR2_X1 U361 ( .A(KEYINPUT19), .B(G183GAT), .ZN(n309) );
  XNOR2_X1 U362 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U363 ( .A(G169GAT), .B(n311), .Z(n440) );
  XNOR2_X1 U364 ( .A(n440), .B(G204GAT), .ZN(n312) );
  XNOR2_X1 U365 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U366 ( .A(n315), .B(n314), .Z(n317) );
  NAND2_X1 U367 ( .A1(G226GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U368 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U369 ( .A(n319), .B(n318), .ZN(n487) );
  XOR2_X1 U370 ( .A(KEYINPUT107), .B(KEYINPUT108), .Z(n371) );
  XOR2_X1 U371 ( .A(KEYINPUT46), .B(KEYINPUT106), .Z(n355) );
  XOR2_X1 U372 ( .A(G8GAT), .B(G197GAT), .Z(n321) );
  XNOR2_X1 U373 ( .A(G50GAT), .B(G36GAT), .ZN(n320) );
  XNOR2_X1 U374 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U375 ( .A(n322), .B(G113GAT), .Z(n325) );
  XNOR2_X1 U376 ( .A(G169GAT), .B(n323), .ZN(n324) );
  XNOR2_X1 U377 ( .A(n325), .B(n324), .ZN(n331) );
  XOR2_X1 U378 ( .A(G29GAT), .B(G43GAT), .Z(n327) );
  XNOR2_X1 U379 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n326) );
  XNOR2_X1 U380 ( .A(n327), .B(n326), .ZN(n358) );
  XOR2_X1 U381 ( .A(G141GAT), .B(G22GAT), .Z(n420) );
  XOR2_X1 U382 ( .A(n358), .B(n420), .Z(n329) );
  NAND2_X1 U383 ( .A1(G229GAT), .A2(G233GAT), .ZN(n328) );
  XNOR2_X1 U384 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U385 ( .A(n331), .B(n330), .Z(n339) );
  XOR2_X1 U386 ( .A(KEYINPUT69), .B(KEYINPUT74), .Z(n333) );
  XNOR2_X1 U387 ( .A(KEYINPUT73), .B(KEYINPUT72), .ZN(n332) );
  XNOR2_X1 U388 ( .A(n333), .B(n332), .ZN(n337) );
  XOR2_X1 U389 ( .A(KEYINPUT71), .B(KEYINPUT29), .Z(n335) );
  XNOR2_X1 U390 ( .A(KEYINPUT30), .B(KEYINPUT70), .ZN(n334) );
  XNOR2_X1 U391 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U392 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U393 ( .A(n339), .B(n338), .ZN(n563) );
  XOR2_X1 U394 ( .A(n341), .B(n340), .Z(n346) );
  XNOR2_X1 U395 ( .A(G78GAT), .B(G204GAT), .ZN(n342) );
  XNOR2_X1 U396 ( .A(n342), .B(G148GAT), .ZN(n411) );
  XOR2_X1 U397 ( .A(G85GAT), .B(G92GAT), .Z(n344) );
  XNOR2_X1 U398 ( .A(G99GAT), .B(G106GAT), .ZN(n343) );
  XNOR2_X1 U399 ( .A(n344), .B(n343), .ZN(n364) );
  XNOR2_X1 U400 ( .A(n411), .B(n364), .ZN(n345) );
  XNOR2_X1 U401 ( .A(n346), .B(n345), .ZN(n353) );
  XOR2_X1 U402 ( .A(G120GAT), .B(G71GAT), .Z(n436) );
  XOR2_X1 U403 ( .A(KEYINPUT33), .B(KEYINPUT75), .Z(n348) );
  XNOR2_X1 U404 ( .A(KEYINPUT31), .B(KEYINPUT32), .ZN(n347) );
  XNOR2_X1 U405 ( .A(n348), .B(n347), .ZN(n349) );
  XOR2_X1 U406 ( .A(n436), .B(n349), .Z(n351) );
  NAND2_X1 U407 ( .A1(G230GAT), .A2(G233GAT), .ZN(n350) );
  XNOR2_X1 U408 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U409 ( .A(n353), .B(n352), .ZN(n571) );
  XNOR2_X1 U410 ( .A(KEYINPUT41), .B(n571), .ZN(n558) );
  NOR2_X1 U411 ( .A1(n563), .A2(n558), .ZN(n354) );
  XOR2_X1 U412 ( .A(n355), .B(n354), .Z(n356) );
  NOR2_X1 U413 ( .A1(n576), .A2(n356), .ZN(n369) );
  XNOR2_X1 U414 ( .A(n358), .B(n357), .ZN(n368) );
  XOR2_X1 U415 ( .A(G50GAT), .B(G162GAT), .Z(n419) );
  XOR2_X1 U416 ( .A(KEYINPUT76), .B(KEYINPUT9), .Z(n360) );
  XNOR2_X1 U417 ( .A(KEYINPUT67), .B(KEYINPUT10), .ZN(n359) );
  XNOR2_X1 U418 ( .A(n360), .B(n359), .ZN(n361) );
  NAND2_X1 U419 ( .A1(G232GAT), .A2(G233GAT), .ZN(n362) );
  XNOR2_X1 U420 ( .A(n291), .B(n362), .ZN(n366) );
  XOR2_X1 U421 ( .A(G134GAT), .B(KEYINPUT11), .Z(n363) );
  XNOR2_X1 U422 ( .A(n368), .B(n367), .ZN(n550) );
  NAND2_X1 U423 ( .A1(n369), .A2(n550), .ZN(n370) );
  XNOR2_X1 U424 ( .A(n371), .B(n370), .ZN(n372) );
  XNOR2_X1 U425 ( .A(n372), .B(KEYINPUT47), .ZN(n378) );
  XNOR2_X1 U426 ( .A(KEYINPUT36), .B(n537), .ZN(n581) );
  NOR2_X1 U427 ( .A1(n547), .A2(n581), .ZN(n374) );
  XNOR2_X1 U428 ( .A(KEYINPUT66), .B(KEYINPUT45), .ZN(n373) );
  XNOR2_X1 U429 ( .A(n374), .B(n373), .ZN(n375) );
  NAND2_X1 U430 ( .A1(n375), .A2(n563), .ZN(n376) );
  NOR2_X1 U431 ( .A1(n571), .A2(n376), .ZN(n377) );
  NOR2_X1 U432 ( .A1(n378), .A2(n377), .ZN(n381) );
  INV_X1 U433 ( .A(KEYINPUT64), .ZN(n379) );
  AND2_X1 U434 ( .A1(n487), .A2(n523), .ZN(n382) );
  XNOR2_X1 U435 ( .A(n383), .B(n382), .ZN(n407) );
  XOR2_X1 U436 ( .A(KEYINPUT81), .B(G134GAT), .Z(n385) );
  XNOR2_X1 U437 ( .A(KEYINPUT0), .B(G127GAT), .ZN(n384) );
  XNOR2_X1 U438 ( .A(n385), .B(n384), .ZN(n386) );
  XNOR2_X1 U439 ( .A(G113GAT), .B(n386), .ZN(n443) );
  INV_X1 U440 ( .A(n443), .ZN(n406) );
  XOR2_X1 U441 ( .A(G57GAT), .B(G148GAT), .Z(n388) );
  XNOR2_X1 U442 ( .A(G141GAT), .B(G1GAT), .ZN(n387) );
  XNOR2_X1 U443 ( .A(n388), .B(n387), .ZN(n392) );
  XOR2_X1 U444 ( .A(KEYINPUT4), .B(KEYINPUT91), .Z(n390) );
  XNOR2_X1 U445 ( .A(KEYINPUT6), .B(KEYINPUT1), .ZN(n389) );
  XNOR2_X1 U446 ( .A(n390), .B(n389), .ZN(n391) );
  XOR2_X1 U447 ( .A(n392), .B(n391), .Z(n404) );
  XOR2_X1 U448 ( .A(KEYINPUT90), .B(KEYINPUT89), .Z(n394) );
  XNOR2_X1 U449 ( .A(KEYINPUT3), .B(G155GAT), .ZN(n393) );
  XNOR2_X1 U450 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U451 ( .A(KEYINPUT2), .B(n395), .ZN(n423) );
  INV_X1 U452 ( .A(n423), .ZN(n402) );
  XOR2_X1 U453 ( .A(G85GAT), .B(G162GAT), .Z(n397) );
  XNOR2_X1 U454 ( .A(G29GAT), .B(G120GAT), .ZN(n396) );
  XNOR2_X1 U455 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U456 ( .A(KEYINPUT5), .B(n398), .Z(n400) );
  NAND2_X1 U457 ( .A1(G225GAT), .A2(G233GAT), .ZN(n399) );
  XNOR2_X1 U458 ( .A(n400), .B(n399), .ZN(n401) );
  XNOR2_X1 U459 ( .A(n402), .B(n401), .ZN(n403) );
  XNOR2_X1 U460 ( .A(n404), .B(n403), .ZN(n405) );
  XOR2_X1 U461 ( .A(n406), .B(n405), .Z(n507) );
  INV_X1 U462 ( .A(n507), .ZN(n482) );
  XOR2_X1 U463 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n409) );
  NAND2_X1 U464 ( .A1(G228GAT), .A2(G233GAT), .ZN(n408) );
  XNOR2_X1 U465 ( .A(n409), .B(n408), .ZN(n410) );
  XOR2_X1 U466 ( .A(n410), .B(KEYINPUT88), .Z(n414) );
  XNOR2_X1 U467 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U468 ( .A(n414), .B(n413), .ZN(n418) );
  XOR2_X1 U469 ( .A(KEYINPUT87), .B(KEYINPUT22), .Z(n416) );
  XNOR2_X1 U470 ( .A(G218GAT), .B(G106GAT), .ZN(n415) );
  XNOR2_X1 U471 ( .A(n416), .B(n415), .ZN(n417) );
  XOR2_X1 U472 ( .A(n418), .B(n417), .Z(n422) );
  XNOR2_X1 U473 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U474 ( .A(n422), .B(n421), .ZN(n424) );
  XNOR2_X1 U475 ( .A(n424), .B(n423), .ZN(n461) );
  NAND2_X1 U476 ( .A1(n562), .A2(n461), .ZN(n426) );
  XOR2_X1 U477 ( .A(KEYINPUT83), .B(KEYINPUT20), .Z(n428) );
  XNOR2_X1 U478 ( .A(G15GAT), .B(KEYINPUT84), .ZN(n427) );
  XNOR2_X1 U479 ( .A(n428), .B(n427), .ZN(n432) );
  XOR2_X1 U480 ( .A(KEYINPUT86), .B(KEYINPUT65), .Z(n430) );
  XNOR2_X1 U481 ( .A(KEYINPUT82), .B(KEYINPUT85), .ZN(n429) );
  XNOR2_X1 U482 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U483 ( .A(n432), .B(n431), .Z(n442) );
  XOR2_X1 U484 ( .A(G176GAT), .B(G190GAT), .Z(n434) );
  XNOR2_X1 U485 ( .A(G43GAT), .B(G99GAT), .ZN(n433) );
  XNOR2_X1 U486 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U487 ( .A(n436), .B(n435), .Z(n438) );
  NAND2_X1 U488 ( .A1(G227GAT), .A2(G233GAT), .ZN(n437) );
  XNOR2_X1 U489 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U490 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U491 ( .A(n442), .B(n441), .ZN(n444) );
  XOR2_X1 U492 ( .A(n444), .B(n443), .Z(n514) );
  INV_X1 U493 ( .A(n514), .ZN(n526) );
  NAND2_X1 U494 ( .A1(n445), .A2(n526), .ZN(n557) );
  NOR2_X1 U495 ( .A1(n547), .A2(n557), .ZN(n447) );
  INV_X1 U496 ( .A(G183GAT), .ZN(n446) );
  XNOR2_X1 U497 ( .A(n447), .B(n446), .ZN(G1350GAT) );
  NOR2_X1 U498 ( .A1(n537), .A2(n557), .ZN(n450) );
  XOR2_X1 U499 ( .A(KEYINPUT119), .B(KEYINPUT58), .Z(n449) );
  XNOR2_X1 U500 ( .A(G190GAT), .B(KEYINPUT120), .ZN(n448) );
  XNOR2_X1 U501 ( .A(n450), .B(n290), .ZN(G1351GAT) );
  NOR2_X1 U502 ( .A1(n563), .A2(n571), .ZN(n480) );
  XOR2_X1 U503 ( .A(KEYINPUT80), .B(KEYINPUT16), .Z(n452) );
  NAND2_X1 U504 ( .A1(n537), .A2(n576), .ZN(n451) );
  XNOR2_X1 U505 ( .A(n452), .B(n451), .ZN(n468) );
  XNOR2_X1 U506 ( .A(n487), .B(KEYINPUT27), .ZN(n463) );
  NOR2_X1 U507 ( .A1(n526), .A2(n461), .ZN(n453) );
  XOR2_X1 U508 ( .A(KEYINPUT93), .B(n453), .Z(n454) );
  XNOR2_X1 U509 ( .A(KEYINPUT26), .B(n454), .ZN(n561) );
  NAND2_X1 U510 ( .A1(n463), .A2(n561), .ZN(n459) );
  NAND2_X1 U511 ( .A1(n487), .A2(n526), .ZN(n455) );
  NAND2_X1 U512 ( .A1(n455), .A2(n461), .ZN(n456) );
  XNOR2_X1 U513 ( .A(n456), .B(KEYINPUT25), .ZN(n457) );
  XOR2_X1 U514 ( .A(KEYINPUT94), .B(n457), .Z(n458) );
  NAND2_X1 U515 ( .A1(n459), .A2(n458), .ZN(n460) );
  NAND2_X1 U516 ( .A1(n460), .A2(n507), .ZN(n467) );
  XNOR2_X1 U517 ( .A(n461), .B(KEYINPUT68), .ZN(n462) );
  XNOR2_X1 U518 ( .A(n462), .B(KEYINPUT28), .ZN(n519) );
  NAND2_X1 U519 ( .A1(n463), .A2(n482), .ZN(n464) );
  XOR2_X1 U520 ( .A(n464), .B(KEYINPUT92), .Z(n522) );
  AND2_X1 U521 ( .A1(n522), .A2(n514), .ZN(n465) );
  NAND2_X1 U522 ( .A1(n519), .A2(n465), .ZN(n466) );
  NAND2_X1 U523 ( .A1(n467), .A2(n466), .ZN(n477) );
  AND2_X1 U524 ( .A1(n468), .A2(n477), .ZN(n495) );
  NAND2_X1 U525 ( .A1(n480), .A2(n495), .ZN(n475) );
  NOR2_X1 U526 ( .A1(n507), .A2(n475), .ZN(n470) );
  XNOR2_X1 U527 ( .A(KEYINPUT95), .B(KEYINPUT34), .ZN(n469) );
  XNOR2_X1 U528 ( .A(n470), .B(n469), .ZN(n471) );
  XNOR2_X1 U529 ( .A(G1GAT), .B(n471), .ZN(G1324GAT) );
  INV_X1 U530 ( .A(n487), .ZN(n510) );
  NOR2_X1 U531 ( .A1(n510), .A2(n475), .ZN(n472) );
  XOR2_X1 U532 ( .A(G8GAT), .B(n472), .Z(G1325GAT) );
  NOR2_X1 U533 ( .A1(n514), .A2(n475), .ZN(n474) );
  XNOR2_X1 U534 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n473) );
  XNOR2_X1 U535 ( .A(n474), .B(n473), .ZN(G1326GAT) );
  NOR2_X1 U536 ( .A1(n519), .A2(n475), .ZN(n476) );
  XOR2_X1 U537 ( .A(G22GAT), .B(n476), .Z(G1327GAT) );
  XOR2_X1 U538 ( .A(G29GAT), .B(KEYINPUT96), .Z(n484) );
  NAND2_X1 U539 ( .A1(n547), .A2(n477), .ZN(n478) );
  NOR2_X1 U540 ( .A1(n581), .A2(n478), .ZN(n479) );
  XOR2_X1 U541 ( .A(KEYINPUT37), .B(n479), .Z(n506) );
  NAND2_X1 U542 ( .A1(n480), .A2(n506), .ZN(n481) );
  XOR2_X1 U543 ( .A(KEYINPUT38), .B(n481), .Z(n491) );
  NAND2_X1 U544 ( .A1(n491), .A2(n482), .ZN(n483) );
  XNOR2_X1 U545 ( .A(n484), .B(n483), .ZN(n486) );
  XOR2_X1 U546 ( .A(KEYINPUT39), .B(KEYINPUT97), .Z(n485) );
  XNOR2_X1 U547 ( .A(n486), .B(n485), .ZN(G1328GAT) );
  NAND2_X1 U548 ( .A1(n491), .A2(n487), .ZN(n488) );
  XNOR2_X1 U549 ( .A(n488), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U550 ( .A1(n491), .A2(n526), .ZN(n489) );
  XNOR2_X1 U551 ( .A(n489), .B(KEYINPUT40), .ZN(n490) );
  XNOR2_X1 U552 ( .A(G43GAT), .B(n490), .ZN(G1330GAT) );
  INV_X1 U553 ( .A(n519), .ZN(n524) );
  NAND2_X1 U554 ( .A1(n524), .A2(n491), .ZN(n492) );
  XNOR2_X1 U555 ( .A(G50GAT), .B(n492), .ZN(G1331GAT) );
  INV_X1 U556 ( .A(n563), .ZN(n493) );
  NOR2_X1 U557 ( .A1(n493), .A2(n558), .ZN(n494) );
  XNOR2_X1 U558 ( .A(n494), .B(KEYINPUT98), .ZN(n505) );
  NAND2_X1 U559 ( .A1(n495), .A2(n505), .ZN(n502) );
  NOR2_X1 U560 ( .A1(n507), .A2(n502), .ZN(n496) );
  XOR2_X1 U561 ( .A(G57GAT), .B(n496), .Z(n497) );
  XNOR2_X1 U562 ( .A(KEYINPUT42), .B(n497), .ZN(G1332GAT) );
  NOR2_X1 U563 ( .A1(n510), .A2(n502), .ZN(n499) );
  XNOR2_X1 U564 ( .A(G64GAT), .B(KEYINPUT99), .ZN(n498) );
  XNOR2_X1 U565 ( .A(n499), .B(n498), .ZN(G1333GAT) );
  NOR2_X1 U566 ( .A1(n514), .A2(n502), .ZN(n500) );
  XOR2_X1 U567 ( .A(KEYINPUT100), .B(n500), .Z(n501) );
  XNOR2_X1 U568 ( .A(G71GAT), .B(n501), .ZN(G1334GAT) );
  NOR2_X1 U569 ( .A1(n519), .A2(n502), .ZN(n504) );
  XNOR2_X1 U570 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n503) );
  XNOR2_X1 U571 ( .A(n504), .B(n503), .ZN(G1335GAT) );
  NAND2_X1 U572 ( .A1(n506), .A2(n505), .ZN(n518) );
  NOR2_X1 U573 ( .A1(n507), .A2(n518), .ZN(n509) );
  XNOR2_X1 U574 ( .A(G85GAT), .B(KEYINPUT101), .ZN(n508) );
  XNOR2_X1 U575 ( .A(n509), .B(n508), .ZN(G1336GAT) );
  NOR2_X1 U576 ( .A1(n510), .A2(n518), .ZN(n512) );
  XNOR2_X1 U577 ( .A(KEYINPUT102), .B(KEYINPUT103), .ZN(n511) );
  XNOR2_X1 U578 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U579 ( .A(G92GAT), .B(n513), .ZN(G1337GAT) );
  NOR2_X1 U580 ( .A1(n514), .A2(n518), .ZN(n516) );
  XNOR2_X1 U581 ( .A(KEYINPUT104), .B(KEYINPUT105), .ZN(n515) );
  XNOR2_X1 U582 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X1 U583 ( .A(G99GAT), .B(n517), .ZN(G1338GAT) );
  NOR2_X1 U584 ( .A1(n519), .A2(n518), .ZN(n520) );
  XOR2_X1 U585 ( .A(KEYINPUT44), .B(n520), .Z(n521) );
  XNOR2_X1 U586 ( .A(G106GAT), .B(n521), .ZN(G1339GAT) );
  NAND2_X1 U587 ( .A1(n523), .A2(n522), .ZN(n540) );
  NOR2_X1 U588 ( .A1(n524), .A2(n540), .ZN(n525) );
  NAND2_X1 U589 ( .A1(n526), .A2(n525), .ZN(n536) );
  NOR2_X1 U590 ( .A1(n563), .A2(n536), .ZN(n528) );
  XNOR2_X1 U591 ( .A(G113GAT), .B(KEYINPUT109), .ZN(n527) );
  XNOR2_X1 U592 ( .A(n528), .B(n527), .ZN(G1340GAT) );
  NOR2_X1 U593 ( .A1(n536), .A2(n558), .ZN(n532) );
  XOR2_X1 U594 ( .A(KEYINPUT110), .B(KEYINPUT111), .Z(n530) );
  XNOR2_X1 U595 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n529) );
  XNOR2_X1 U596 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U597 ( .A(n532), .B(n531), .ZN(G1341GAT) );
  NOR2_X1 U598 ( .A1(n547), .A2(n536), .ZN(n534) );
  XNOR2_X1 U599 ( .A(KEYINPUT112), .B(KEYINPUT50), .ZN(n533) );
  XNOR2_X1 U600 ( .A(n534), .B(n533), .ZN(n535) );
  XOR2_X1 U601 ( .A(G127GAT), .B(n535), .Z(G1342GAT) );
  NOR2_X1 U602 ( .A1(n537), .A2(n536), .ZN(n539) );
  XNOR2_X1 U603 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n538) );
  XNOR2_X1 U604 ( .A(n539), .B(n538), .ZN(G1343GAT) );
  INV_X1 U605 ( .A(n540), .ZN(n541) );
  NAND2_X1 U606 ( .A1(n541), .A2(n561), .ZN(n549) );
  NOR2_X1 U607 ( .A1(n563), .A2(n549), .ZN(n542) );
  XOR2_X1 U608 ( .A(G141GAT), .B(n542), .Z(G1344GAT) );
  NOR2_X1 U609 ( .A1(n549), .A2(n558), .ZN(n546) );
  XOR2_X1 U610 ( .A(KEYINPUT113), .B(KEYINPUT53), .Z(n544) );
  XNOR2_X1 U611 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n543) );
  XNOR2_X1 U612 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U613 ( .A(n546), .B(n545), .ZN(G1345GAT) );
  NOR2_X1 U614 ( .A1(n547), .A2(n549), .ZN(n548) );
  XOR2_X1 U615 ( .A(G155GAT), .B(n548), .Z(G1346GAT) );
  NOR2_X1 U616 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U617 ( .A(KEYINPUT114), .B(n551), .Z(n552) );
  XNOR2_X1 U618 ( .A(G162GAT), .B(n552), .ZN(G1347GAT) );
  NOR2_X1 U619 ( .A1(n563), .A2(n557), .ZN(n554) );
  XNOR2_X1 U620 ( .A(G169GAT), .B(KEYINPUT117), .ZN(n553) );
  XNOR2_X1 U621 ( .A(n554), .B(n553), .ZN(G1348GAT) );
  XOR2_X1 U622 ( .A(KEYINPUT56), .B(KEYINPUT118), .Z(n556) );
  XNOR2_X1 U623 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n555) );
  XNOR2_X1 U624 ( .A(n556), .B(n555), .ZN(n560) );
  NOR2_X1 U625 ( .A1(n558), .A2(n557), .ZN(n559) );
  XOR2_X1 U626 ( .A(n560), .B(n559), .Z(G1349GAT) );
  NAND2_X1 U627 ( .A1(n562), .A2(n561), .ZN(n580) );
  NOR2_X1 U628 ( .A1(n563), .A2(n580), .ZN(n568) );
  XOR2_X1 U629 ( .A(KEYINPUT60), .B(KEYINPUT122), .Z(n565) );
  XNOR2_X1 U630 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n565), .B(n564), .ZN(n566) );
  XNOR2_X1 U632 ( .A(KEYINPUT121), .B(n566), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n568), .B(n567), .ZN(G1352GAT) );
  XOR2_X1 U634 ( .A(KEYINPUT61), .B(KEYINPUT125), .Z(n570) );
  XNOR2_X1 U635 ( .A(G204GAT), .B(KEYINPUT124), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(n574) );
  INV_X1 U637 ( .A(n580), .ZN(n575) );
  NAND2_X1 U638 ( .A1(n571), .A2(n575), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n572), .B(KEYINPUT123), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(G1353GAT) );
  NAND2_X1 U641 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U642 ( .A(n577), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U643 ( .A(KEYINPUT126), .B(KEYINPUT127), .Z(n579) );
  XNOR2_X1 U644 ( .A(G218GAT), .B(KEYINPUT62), .ZN(n578) );
  XNOR2_X1 U645 ( .A(n579), .B(n578), .ZN(n583) );
  NOR2_X1 U646 ( .A1(n581), .A2(n580), .ZN(n582) );
  XOR2_X1 U647 ( .A(n583), .B(n582), .Z(G1355GAT) );
endmodule

