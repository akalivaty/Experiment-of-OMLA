//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 1 0 1 0 0 1 1 0 0 1 0 1 0 1 1 1 0 0 0 0 0 1 1 1 0 1 0 0 1 1 0 0 0 1 1 1 0 0 1 1 1 0 0 1 0 0 1 0 0 0 0 0 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:22 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1269, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n201), .A2(G77), .A3(new_n203), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n206), .B(KEYINPUT65), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XOR2_X1   g0009(.A(new_n209), .B(KEYINPUT0), .Z(new_n210));
  INV_X1    g0010(.A(G68), .ZN(new_n211));
  INV_X1    g0011(.A(G238), .ZN(new_n212));
  INV_X1    g0012(.A(G97), .ZN(new_n213));
  INV_X1    g0013(.A(G257), .ZN(new_n214));
  OAI22_X1  g0014(.A1(new_n211), .A2(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(G50), .ZN(new_n216));
  INV_X1    g0016(.A(G226), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g0018(.A(G58), .ZN(new_n219));
  INV_X1    g0019(.A(G232), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  AND2_X1   g0021(.A1(G116), .A2(G270), .ZN(new_n222));
  NOR4_X1   g0022(.A1(new_n215), .A2(new_n218), .A3(new_n221), .A4(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(G77), .ZN(new_n224));
  INV_X1    g0024(.A(G244), .ZN(new_n225));
  INV_X1    g0025(.A(G87), .ZN(new_n226));
  INV_X1    g0026(.A(G250), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n223), .B1(new_n224), .B2(new_n225), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  INV_X1    g0028(.A(G107), .ZN(new_n229));
  INV_X1    g0029(.A(G264), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n207), .B1(new_n228), .B2(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT1), .ZN(new_n233));
  NAND2_X1  g0033(.A1(G1), .A2(G13), .ZN(new_n234));
  INV_X1    g0034(.A(G20), .ZN(new_n235));
  NOR2_X1   g0035(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g0036(.A1(new_n203), .A2(G50), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT66), .ZN(new_n238));
  AOI211_X1 g0038(.A(new_n210), .B(new_n233), .C1(new_n236), .C2(new_n238), .ZN(G361));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G232), .ZN(new_n241));
  XNOR2_X1  g0041(.A(KEYINPUT2), .B(G226), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G250), .B(G257), .Z(new_n244));
  XNOR2_X1  g0044(.A(G264), .B(G270), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G358));
  XNOR2_X1  g0047(.A(G87), .B(G97), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G107), .B(G116), .ZN(new_n249));
  XOR2_X1   g0049(.A(new_n248), .B(new_n249), .Z(new_n250));
  XNOR2_X1  g0050(.A(G68), .B(G77), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G50), .B(G58), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XOR2_X1   g0053(.A(new_n250), .B(new_n253), .Z(G351));
  AND2_X1   g0054(.A1(KEYINPUT3), .A2(G33), .ZN(new_n255));
  NOR2_X1   g0055(.A1(KEYINPUT3), .A2(G33), .ZN(new_n256));
  OAI21_X1  g0056(.A(KEYINPUT67), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT3), .ZN(new_n258));
  INV_X1    g0058(.A(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT67), .ZN(new_n261));
  NAND2_X1  g0061(.A1(KEYINPUT3), .A2(G33), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n260), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  AOI22_X1  g0063(.A1(new_n257), .A2(new_n263), .B1(new_n220), .B2(G1698), .ZN(new_n264));
  INV_X1    g0064(.A(G1698), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n217), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(G33), .A2(G97), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G41), .ZN(new_n270));
  OAI211_X1 g0070(.A(G1), .B(G13), .C1(new_n259), .C2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n269), .A2(KEYINPUT71), .A3(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT71), .ZN(new_n274));
  AOI22_X1  g0074(.A1(new_n264), .A2(new_n266), .B1(G33), .B2(G97), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n274), .B1(new_n275), .B2(new_n271), .ZN(new_n276));
  INV_X1    g0076(.A(G1), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n277), .B1(G41), .B2(G45), .ZN(new_n278));
  INV_X1    g0078(.A(G274), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  AND2_X1   g0080(.A1(new_n271), .A2(new_n278), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n280), .B1(new_n281), .B2(G238), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n273), .A2(new_n276), .A3(new_n282), .ZN(new_n283));
  OR2_X1    g0083(.A1(new_n283), .A2(KEYINPUT13), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(KEYINPUT13), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G190), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NOR2_X1   g0088(.A1(G20), .A2(G33), .ZN(new_n289));
  AOI22_X1  g0089(.A1(new_n289), .A2(G50), .B1(G20), .B2(new_n211), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n259), .A2(G20), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n290), .B1(new_n292), .B2(new_n224), .ZN(new_n293));
  NAND3_X1  g0093(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(new_n234), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  XOR2_X1   g0096(.A(new_n296), .B(KEYINPUT11), .Z(new_n297));
  INV_X1    g0097(.A(new_n295), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n298), .B1(G1), .B2(new_n235), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT12), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n277), .A2(G13), .A3(G20), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n300), .B1(new_n302), .B2(new_n211), .ZN(new_n303));
  NOR3_X1   g0103(.A1(new_n301), .A2(KEYINPUT12), .A3(G68), .ZN(new_n304));
  OAI22_X1  g0104(.A1(new_n299), .A2(new_n211), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n297), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G200), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n308), .B1(new_n284), .B2(new_n285), .ZN(new_n309));
  NOR3_X1   g0109(.A1(new_n288), .A2(new_n307), .A3(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n286), .A2(G169), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(KEYINPUT14), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n284), .A2(G179), .A3(new_n285), .ZN(new_n313));
  INV_X1    g0113(.A(G169), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n314), .B1(new_n284), .B2(new_n285), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT14), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n312), .A2(new_n313), .A3(new_n317), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n310), .B1(new_n318), .B2(new_n307), .ZN(new_n319));
  OAI21_X1  g0119(.A(G20), .B1(new_n201), .B2(new_n203), .ZN(new_n320));
  INV_X1    g0120(.A(G150), .ZN(new_n321));
  INV_X1    g0121(.A(new_n289), .ZN(new_n322));
  XOR2_X1   g0122(.A(KEYINPUT8), .B(G58), .Z(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  OAI221_X1 g0124(.A(new_n320), .B1(new_n321), .B2(new_n322), .C1(new_n324), .C2(new_n292), .ZN(new_n325));
  AOI22_X1  g0125(.A1(new_n325), .A2(new_n295), .B1(new_n216), .B2(new_n302), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n326), .B1(new_n216), .B2(new_n299), .ZN(new_n327));
  XNOR2_X1  g0127(.A(new_n327), .B(KEYINPUT9), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT70), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n281), .A2(G226), .ZN(new_n330));
  INV_X1    g0130(.A(new_n280), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n257), .A2(new_n263), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  MUX2_X1   g0133(.A(G222), .B(G223), .S(G1698), .Z(new_n334));
  OAI21_X1  g0134(.A(new_n272), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n332), .A2(G77), .ZN(new_n336));
  OAI211_X1 g0136(.A(new_n330), .B(new_n331), .C1(new_n335), .C2(new_n336), .ZN(new_n337));
  OR2_X1    g0137(.A1(new_n337), .A2(new_n287), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(G200), .ZN(new_n339));
  NAND4_X1  g0139(.A1(new_n328), .A2(new_n329), .A3(new_n338), .A4(new_n339), .ZN(new_n340));
  XNOR2_X1  g0140(.A(new_n340), .B(KEYINPUT10), .ZN(new_n341));
  OR2_X1    g0141(.A1(new_n322), .A2(KEYINPUT69), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n322), .A2(KEYINPUT69), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n342), .A2(new_n323), .A3(new_n343), .ZN(new_n344));
  XNOR2_X1  g0144(.A(KEYINPUT15), .B(G87), .ZN(new_n345));
  OAI221_X1 g0145(.A(new_n344), .B1(new_n235), .B2(new_n224), .C1(new_n292), .C2(new_n345), .ZN(new_n346));
  AOI22_X1  g0146(.A1(new_n346), .A2(new_n295), .B1(new_n224), .B2(new_n302), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n347), .B1(new_n224), .B2(new_n299), .ZN(new_n348));
  AOI21_X1  g0148(.A(G1698), .B1(new_n257), .B2(new_n263), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(G232), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n332), .A2(G1698), .ZN(new_n351));
  OAI221_X1 g0151(.A(new_n350), .B1(new_n229), .B2(new_n332), .C1(new_n351), .C2(new_n212), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(new_n272), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n281), .A2(G244), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n353), .A2(new_n331), .A3(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n348), .B1(new_n355), .B2(G200), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n356), .B1(new_n287), .B2(new_n355), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n319), .A2(new_n341), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n337), .A2(new_n314), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n327), .B(new_n359), .C1(G179), .C2(new_n337), .ZN(new_n360));
  XOR2_X1   g0160(.A(new_n360), .B(KEYINPUT68), .Z(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n355), .ZN(new_n363));
  INV_X1    g0163(.A(G179), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  OAI211_X1 g0165(.A(new_n365), .B(new_n348), .C1(G169), .C2(new_n363), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT72), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n323), .A2(new_n302), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n369), .B1(new_n299), .B2(new_n323), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n217), .A2(G1698), .ZN(new_n371));
  OAI221_X1 g0171(.A(new_n371), .B1(G223), .B2(G1698), .C1(new_n255), .C2(new_n256), .ZN(new_n372));
  NAND2_X1  g0172(.A1(G33), .A2(G87), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n280), .B1(new_n374), .B2(new_n272), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n281), .A2(G232), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n308), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n219), .A2(new_n211), .ZN(new_n378));
  OAI21_X1  g0178(.A(G20), .B1(new_n378), .B2(new_n202), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n289), .A2(G159), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT7), .ZN(new_n383));
  NOR4_X1   g0183(.A1(new_n255), .A2(new_n256), .A3(new_n383), .A4(G20), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n257), .A2(new_n263), .A3(new_n235), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n384), .B1(new_n385), .B2(new_n383), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n382), .B1(new_n386), .B2(new_n211), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT16), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n260), .A2(new_n262), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n383), .B1(new_n390), .B2(G20), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n255), .A2(new_n256), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n392), .A2(KEYINPUT7), .A3(new_n235), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n381), .B1(new_n394), .B2(G68), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n298), .B1(new_n395), .B2(KEYINPUT16), .ZN(new_n396));
  AOI211_X1 g0196(.A(new_n370), .B(new_n377), .C1(new_n389), .C2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n375), .A2(new_n376), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(G190), .ZN(new_n400));
  AOI21_X1  g0200(.A(KEYINPUT17), .B1(new_n397), .B2(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n370), .B1(new_n389), .B2(new_n396), .ZN(new_n402));
  INV_X1    g0202(.A(new_n377), .ZN(new_n403));
  AND4_X1   g0203(.A1(KEYINPUT17), .A2(new_n402), .A3(new_n400), .A4(new_n403), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n368), .B1(new_n401), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n389), .A2(new_n396), .ZN(new_n406));
  INV_X1    g0206(.A(new_n370), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n314), .B1(new_n375), .B2(new_n376), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n409), .B1(new_n399), .B2(G179), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT18), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n408), .A2(new_n411), .A3(KEYINPUT18), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n402), .A2(new_n400), .A3(new_n403), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT17), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n397), .A2(KEYINPUT17), .A3(new_n400), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n419), .A2(new_n420), .A3(KEYINPUT72), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n405), .A2(new_n416), .A3(new_n421), .ZN(new_n422));
  NOR4_X1   g0222(.A1(new_n358), .A2(new_n362), .A3(new_n367), .A4(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT75), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT74), .ZN(new_n425));
  AND2_X1   g0225(.A1(KEYINPUT5), .A2(G41), .ZN(new_n426));
  NOR2_X1   g0226(.A1(KEYINPUT5), .A2(G41), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n277), .A2(G45), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n271), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  OR2_X1    g0230(.A1(new_n430), .A2(new_n214), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT73), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n277), .A2(G45), .A3(G274), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n432), .B1(new_n428), .B2(new_n433), .ZN(new_n434));
  XNOR2_X1  g0234(.A(KEYINPUT5), .B(G41), .ZN(new_n435));
  AND3_X1   g0235(.A1(new_n277), .A2(G45), .A3(G274), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n435), .A2(KEYINPUT73), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n434), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n431), .A2(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n265), .B1(new_n257), .B2(new_n263), .ZN(new_n440));
  AOI22_X1  g0240(.A1(new_n440), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT4), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n442), .B1(new_n349), .B2(G244), .ZN(new_n443));
  NOR4_X1   g0243(.A1(new_n392), .A2(KEYINPUT4), .A3(new_n225), .A4(G1698), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n441), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n439), .B1(new_n445), .B2(new_n272), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n425), .B1(new_n446), .B2(G190), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n332), .A2(G244), .A3(new_n265), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n444), .B1(new_n448), .B2(KEYINPUT4), .ZN(new_n449));
  NAND2_X1  g0249(.A1(G33), .A2(G283), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n450), .B1(new_n351), .B2(new_n227), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n272), .B1(new_n449), .B2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n439), .ZN(new_n453));
  AND4_X1   g0253(.A1(new_n425), .A2(new_n452), .A3(G190), .A4(new_n453), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n447), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n302), .A2(new_n213), .ZN(new_n456));
  OAI211_X1 g0256(.A(new_n298), .B(new_n301), .C1(G1), .C2(new_n259), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n457), .A2(new_n213), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT6), .ZN(new_n460));
  NOR3_X1   g0260(.A1(new_n460), .A2(new_n213), .A3(G107), .ZN(new_n461));
  XNOR2_X1  g0261(.A(G97), .B(G107), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n461), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  OAI22_X1  g0263(.A1(new_n463), .A2(new_n235), .B1(new_n224), .B2(new_n322), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n385), .A2(new_n383), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(new_n393), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n464), .B1(new_n466), .B2(G107), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n456), .B(new_n459), .C1(new_n467), .C2(new_n298), .ZN(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n469), .B1(new_n308), .B2(new_n446), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n424), .B1(new_n455), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n452), .A2(new_n364), .A3(new_n453), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n468), .B(new_n472), .C1(G169), .C2(new_n446), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT76), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n452), .A2(new_n453), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(new_n314), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n477), .A2(KEYINPUT76), .A3(new_n468), .A4(new_n472), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n475), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n468), .B1(G200), .B2(new_n476), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n480), .B(KEYINPUT75), .C1(new_n447), .C2(new_n454), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n471), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n390), .A2(new_n235), .A3(G87), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(KEYINPUT22), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT84), .ZN(new_n485));
  NOR2_X1   g0285(.A1(KEYINPUT22), .A2(G20), .ZN(new_n486));
  AND4_X1   g0286(.A1(new_n485), .A2(new_n332), .A3(G87), .A4(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n226), .B1(new_n257), .B2(new_n263), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n485), .B1(new_n488), .B2(new_n486), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n484), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  NOR3_X1   g0290(.A1(new_n235), .A2(KEYINPUT23), .A3(G107), .ZN(new_n491));
  XNOR2_X1  g0291(.A(new_n491), .B(KEYINPUT85), .ZN(new_n492));
  NAND2_X1  g0292(.A1(G33), .A2(G116), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  OR2_X1    g0294(.A1(new_n494), .A2(KEYINPUT23), .ZN(new_n495));
  AOI22_X1  g0295(.A1(new_n495), .A2(new_n235), .B1(KEYINPUT23), .B2(G107), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n490), .A2(new_n492), .A3(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT24), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n490), .A2(KEYINPUT24), .A3(new_n492), .A4(new_n496), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n499), .A2(new_n295), .A3(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(new_n457), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(G107), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n301), .A2(G107), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT86), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n504), .B1(new_n505), .B2(KEYINPUT25), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(KEYINPUT25), .ZN(new_n507));
  MUX2_X1   g0307(.A(new_n504), .B(new_n506), .S(new_n507), .Z(new_n508));
  NAND3_X1  g0308(.A1(new_n501), .A2(new_n503), .A3(new_n508), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n430), .A2(new_n230), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n390), .A2(G257), .A3(G1698), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(KEYINPUT87), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n390), .A2(G250), .A3(new_n265), .ZN(new_n513));
  NAND2_X1  g0313(.A1(G33), .A2(G294), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT87), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n390), .A2(new_n515), .A3(G257), .A4(G1698), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n512), .A2(new_n513), .A3(new_n514), .A4(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n510), .B1(new_n517), .B2(new_n272), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(new_n438), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n519), .A2(new_n287), .ZN(new_n520));
  INV_X1    g0320(.A(new_n519), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n521), .A2(new_n308), .ZN(new_n522));
  NOR3_X1   g0322(.A1(new_n509), .A2(new_n520), .A3(new_n522), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n482), .A2(new_n523), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n450), .B(new_n235), .C1(G33), .C2(new_n213), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT81), .ZN(new_n526));
  INV_X1    g0326(.A(G116), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(G20), .ZN(new_n528));
  AND3_X1   g0328(.A1(new_n295), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n526), .B1(new_n295), .B2(new_n528), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n525), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT82), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT20), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n502), .A2(G116), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n302), .A2(new_n527), .ZN(new_n536));
  AND3_X1   g0336(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  OR2_X1    g0337(.A1(new_n531), .A2(new_n533), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n531), .A2(new_n533), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n538), .A2(KEYINPUT82), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n537), .A2(new_n540), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n271), .B(G270), .C1(new_n428), .C2(new_n429), .ZN(new_n542));
  NOR3_X1   g0342(.A1(new_n428), .A2(new_n432), .A3(new_n433), .ZN(new_n543));
  AOI21_X1  g0343(.A(KEYINPUT73), .B1(new_n435), .B2(new_n436), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n542), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(KEYINPUT79), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT79), .ZN(new_n547));
  OAI211_X1 g0347(.A(new_n542), .B(new_n547), .C1(new_n543), .C2(new_n544), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n257), .A2(new_n263), .A3(G303), .ZN(new_n550));
  OAI211_X1 g0350(.A(G257), .B(new_n265), .C1(new_n255), .C2(new_n256), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT80), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n390), .A2(KEYINPUT80), .A3(G257), .A4(new_n265), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n390), .A2(G264), .A3(G1698), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n550), .A2(new_n553), .A3(new_n554), .A4(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(new_n272), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n314), .B1(new_n549), .B2(new_n557), .ZN(new_n558));
  AOI21_X1  g0358(.A(KEYINPUT21), .B1(new_n541), .B2(new_n558), .ZN(new_n559));
  AOI22_X1  g0359(.A1(new_n546), .A2(new_n548), .B1(new_n272), .B2(new_n556), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n558), .A2(KEYINPUT21), .B1(G179), .B2(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(new_n541), .ZN(new_n562));
  OAI21_X1  g0362(.A(KEYINPUT83), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(new_n548), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n547), .B1(new_n438), .B2(new_n542), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n557), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n566), .A2(KEYINPUT21), .A3(G169), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n560), .A2(G179), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT83), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n569), .A2(new_n570), .A3(new_n541), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n559), .B1(new_n563), .B2(new_n571), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n519), .A2(G179), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n573), .B1(new_n314), .B2(new_n519), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n509), .A2(new_n574), .ZN(new_n575));
  AND2_X1   g0375(.A1(G33), .A2(G41), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n429), .B(G250), .C1(new_n576), .C2(new_n234), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n433), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT77), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n212), .A2(new_n265), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n225), .A2(G1698), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n581), .B(new_n582), .C1(new_n255), .C2(new_n256), .ZN(new_n583));
  AND2_X1   g0383(.A1(new_n583), .A2(new_n493), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n579), .B(new_n580), .C1(new_n584), .C2(new_n271), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n271), .B1(new_n583), .B2(new_n493), .ZN(new_n586));
  OAI21_X1  g0386(.A(KEYINPUT77), .B1(new_n586), .B2(new_n578), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n585), .A2(G200), .A3(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT78), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n457), .A2(new_n226), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT19), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n235), .B1(new_n268), .B2(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n226), .A2(new_n213), .A3(new_n229), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n235), .A2(G33), .A3(G97), .ZN(new_n594));
  AOI22_X1  g0394(.A1(new_n592), .A2(new_n593), .B1(new_n591), .B2(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n390), .A2(new_n235), .A3(G68), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n298), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n345), .A2(new_n302), .ZN(new_n598));
  INV_X1    g0398(.A(new_n598), .ZN(new_n599));
  NOR3_X1   g0399(.A1(new_n590), .A2(new_n597), .A3(new_n599), .ZN(new_n600));
  AND3_X1   g0400(.A1(new_n588), .A2(new_n589), .A3(new_n600), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n589), .B1(new_n588), .B2(new_n600), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n585), .A2(new_n587), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(G190), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n585), .A2(new_n314), .A3(new_n587), .ZN(new_n606));
  AOI21_X1  g0406(.A(G179), .B1(new_n585), .B2(new_n587), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n457), .A2(new_n345), .ZN(new_n608));
  NOR3_X1   g0408(.A1(new_n608), .A2(new_n597), .A3(new_n599), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  AOI22_X1  g0410(.A1(new_n603), .A2(new_n605), .B1(new_n606), .B2(new_n610), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n541), .B1(G200), .B2(new_n566), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n612), .B1(new_n287), .B2(new_n566), .ZN(new_n613));
  AND4_X1   g0413(.A1(new_n572), .A2(new_n575), .A3(new_n611), .A4(new_n613), .ZN(new_n614));
  AND3_X1   g0414(.A1(new_n423), .A2(new_n524), .A3(new_n614), .ZN(G372));
  INV_X1    g0415(.A(new_n310), .ZN(new_n616));
  AND2_X1   g0416(.A1(new_n318), .A2(new_n307), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n616), .B1(new_n617), .B2(new_n367), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n405), .A2(new_n421), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n416), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n362), .B1(new_n620), .B2(new_n341), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n287), .B1(new_n585), .B2(new_n587), .ZN(new_n622));
  OR3_X1    g0422(.A1(new_n590), .A2(new_n597), .A3(new_n599), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n578), .A2(KEYINPUT88), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT88), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n577), .A2(new_n625), .A3(new_n433), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n586), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n308), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NOR3_X1   g0429(.A1(new_n622), .A2(new_n623), .A3(new_n629), .ZN(new_n630));
  AOI21_X1  g0430(.A(G169), .B1(new_n627), .B2(new_n628), .ZN(new_n631));
  NOR3_X1   g0431(.A1(new_n607), .A2(new_n631), .A3(new_n609), .ZN(new_n632));
  OAI21_X1  g0432(.A(KEYINPUT89), .B1(new_n630), .B2(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(new_n607), .ZN(new_n634));
  INV_X1    g0434(.A(new_n609), .ZN(new_n635));
  INV_X1    g0435(.A(new_n631), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n634), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n629), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n605), .A2(new_n638), .A3(new_n600), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT89), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n637), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n633), .A2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n642), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n559), .B1(new_n541), .B2(new_n569), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n643), .B1(new_n575), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n524), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n611), .A2(new_n475), .A3(new_n478), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(KEYINPUT26), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n473), .B1(new_n633), .B2(new_n641), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT26), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  AND3_X1   g0451(.A1(new_n648), .A2(new_n637), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n646), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n423), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n621), .A2(new_n654), .ZN(G369));
  INV_X1    g0455(.A(G13), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n656), .A2(G20), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  OR3_X1    g0458(.A1(new_n658), .A2(KEYINPUT27), .A3(G1), .ZN(new_n659));
  OAI21_X1  g0459(.A(KEYINPUT27), .B1(new_n658), .B2(G1), .ZN(new_n660));
  AND3_X1   g0460(.A1(new_n659), .A2(G213), .A3(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(G343), .ZN(new_n662));
  XOR2_X1   g0462(.A(new_n662), .B(KEYINPUT90), .Z(new_n663));
  NOR2_X1   g0463(.A1(new_n575), .A2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n501), .A2(new_n503), .ZN(new_n666));
  INV_X1    g0466(.A(new_n520), .ZN(new_n667));
  INV_X1    g0467(.A(new_n522), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n666), .A2(new_n667), .A3(new_n508), .A4(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n509), .A2(new_n663), .ZN(new_n670));
  AND2_X1   g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  AND2_X1   g0471(.A1(new_n509), .A2(new_n574), .ZN(new_n672));
  OAI211_X1 g0472(.A(KEYINPUT91), .B(new_n665), .C1(new_n671), .C2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT91), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n672), .B1(new_n669), .B2(new_n670), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n674), .B1(new_n675), .B2(new_n664), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n663), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n679), .A2(new_n562), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n572), .A2(new_n613), .A3(new_n681), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n682), .B1(new_n644), .B2(new_n681), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(G330), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n678), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n559), .ZN(new_n687));
  AOI221_X4 g0487(.A(KEYINPUT83), .B1(new_n540), .B2(new_n537), .C1(new_n567), .C2(new_n568), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n570), .B1(new_n569), .B2(new_n541), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n687), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(new_n679), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n691), .B1(new_n673), .B2(new_n676), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n692), .A2(new_n664), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n686), .A2(new_n693), .ZN(G399));
  INV_X1    g0494(.A(new_n208), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n695), .A2(G41), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n593), .A2(G116), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n697), .A2(G1), .A3(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n238), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n699), .B1(new_n700), .B2(new_n697), .ZN(new_n701));
  XNOR2_X1  g0501(.A(new_n701), .B(KEYINPUT28), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n614), .A2(new_n524), .A3(new_n679), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n566), .A2(new_n364), .ZN(new_n704));
  AND2_X1   g0504(.A1(new_n518), .A2(new_n604), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n704), .A2(new_n705), .A3(KEYINPUT30), .A4(new_n446), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(KEYINPUT92), .ZN(new_n707));
  AND4_X1   g0507(.A1(new_n452), .A2(new_n453), .A3(new_n518), .A4(new_n604), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT92), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n708), .A2(new_n709), .A3(KEYINPUT30), .A4(new_n704), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n707), .A2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT30), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n705), .A2(new_n446), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n712), .B1(new_n713), .B2(new_n568), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(KEYINPUT93), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n521), .A2(new_n560), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n627), .A2(new_n628), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n716), .A2(new_n364), .A3(new_n476), .A4(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT93), .ZN(new_n719));
  OAI211_X1 g0519(.A(new_n719), .B(new_n712), .C1(new_n713), .C2(new_n568), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n711), .A2(new_n715), .A3(new_n718), .A4(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(new_n663), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT31), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n711), .A2(new_n714), .A3(new_n718), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n725), .A2(KEYINPUT31), .A3(new_n663), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n703), .A2(new_n724), .A3(new_n726), .ZN(new_n727));
  AND2_X1   g0527(.A1(new_n727), .A2(G330), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT94), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n643), .B1(new_n572), .B2(new_n575), .ZN(new_n730));
  AND3_X1   g0530(.A1(new_n471), .A2(new_n481), .A3(new_n479), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n730), .A2(new_n731), .A3(new_n669), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n611), .A2(new_n650), .A3(new_n475), .A4(new_n478), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n637), .B1(new_n649), .B2(new_n650), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  AOI211_X1 g0536(.A(new_n729), .B(new_n663), .C1(new_n732), .C2(new_n736), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n669), .A2(new_n481), .A3(new_n471), .A4(new_n479), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n642), .B1(new_n672), .B2(new_n690), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n736), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  AOI21_X1  g0540(.A(KEYINPUT94), .B1(new_n740), .B2(new_n679), .ZN(new_n741));
  OAI21_X1  g0541(.A(KEYINPUT29), .B1(new_n737), .B2(new_n741), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n663), .B1(new_n646), .B2(new_n652), .ZN(new_n743));
  OR2_X1    g0543(.A1(new_n743), .A2(KEYINPUT29), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n728), .B1(new_n742), .B2(new_n744), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n702), .B1(new_n745), .B2(G1), .ZN(G364));
  NOR2_X1   g0546(.A1(G13), .A2(G33), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n748), .A2(G20), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n683), .A2(new_n750), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n234), .B1(G20), .B2(new_n314), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n749), .A2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n208), .A2(new_n332), .ZN(new_n755));
  INV_X1    g0555(.A(G355), .ZN(new_n756));
  OAI22_X1  g0556(.A1(new_n755), .A2(new_n756), .B1(G116), .B2(new_n208), .ZN(new_n757));
  XNOR2_X1  g0557(.A(new_n757), .B(KEYINPUT95), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n695), .A2(new_n390), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n253), .A2(G45), .ZN(new_n760));
  OAI211_X1 g0560(.A(new_n759), .B(new_n760), .C1(G45), .C2(new_n700), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n754), .B1(new_n758), .B2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n287), .A2(new_n308), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n235), .A2(G179), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(G87), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n308), .A2(G190), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n764), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(G107), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n767), .A2(new_n771), .A3(new_n332), .ZN(new_n772));
  XNOR2_X1  g0572(.A(new_n772), .B(KEYINPUT96), .ZN(new_n773));
  NOR2_X1   g0573(.A1(G190), .A2(G200), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n764), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(G159), .ZN(new_n777));
  XNOR2_X1  g0577(.A(new_n777), .B(KEYINPUT32), .ZN(new_n778));
  NOR3_X1   g0578(.A1(new_n287), .A2(G179), .A3(G200), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(new_n235), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(G97), .ZN(new_n782));
  NAND2_X1  g0582(.A1(G20), .A2(G179), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(new_n774), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n782), .B1(new_n224), .B2(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n778), .A2(new_n786), .ZN(new_n787));
  NOR3_X1   g0587(.A1(new_n783), .A2(new_n308), .A3(G190), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(G68), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n763), .A2(new_n784), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NOR3_X1   g0591(.A1(new_n783), .A2(new_n287), .A3(G200), .ZN(new_n792));
  AOI22_X1  g0592(.A1(new_n791), .A2(G50), .B1(G58), .B2(new_n792), .ZN(new_n793));
  NAND4_X1  g0593(.A1(new_n773), .A2(new_n787), .A3(new_n789), .A4(new_n793), .ZN(new_n794));
  AOI22_X1  g0594(.A1(G326), .A2(new_n791), .B1(new_n776), .B2(G329), .ZN(new_n795));
  INV_X1    g0595(.A(G283), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n795), .B1(new_n796), .B2(new_n769), .ZN(new_n797));
  AOI211_X1 g0597(.A(new_n332), .B(new_n797), .C1(G303), .C2(new_n766), .ZN(new_n798));
  INV_X1    g0598(.A(new_n785), .ZN(new_n799));
  XNOR2_X1  g0599(.A(KEYINPUT33), .B(G317), .ZN(new_n800));
  AOI22_X1  g0600(.A1(new_n799), .A2(G311), .B1(new_n788), .B2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(G294), .ZN(new_n802));
  OAI211_X1 g0602(.A(new_n798), .B(new_n801), .C1(new_n802), .C2(new_n780), .ZN(new_n803));
  INV_X1    g0603(.A(new_n792), .ZN(new_n804));
  INV_X1    g0604(.A(G322), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n794), .B1(new_n803), .B2(new_n806), .ZN(new_n807));
  AND2_X1   g0607(.A1(new_n807), .A2(new_n752), .ZN(new_n808));
  OR3_X1    g0608(.A1(new_n751), .A2(new_n762), .A3(new_n808), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n277), .B1(new_n657), .B2(G45), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n696), .A2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n683), .A2(G330), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n684), .A2(new_n813), .ZN(new_n815));
  OAI22_X1  g0615(.A1(new_n809), .A2(new_n813), .B1(new_n814), .B2(new_n815), .ZN(G396));
  NAND2_X1  g0616(.A1(new_n663), .A2(new_n348), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n357), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n818), .A2(new_n366), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n366), .A2(new_n663), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  OR2_X1    g0622(.A1(new_n743), .A2(new_n822), .ZN(new_n823));
  AND3_X1   g0623(.A1(new_n731), .A2(new_n645), .A3(new_n669), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n648), .A2(new_n637), .A3(new_n651), .ZN(new_n825));
  OAI211_X1 g0625(.A(new_n822), .B(new_n679), .C1(new_n824), .C2(new_n825), .ZN(new_n826));
  AND2_X1   g0626(.A1(new_n823), .A2(new_n826), .ZN(new_n827));
  XOR2_X1   g0627(.A(new_n827), .B(new_n728), .Z(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(new_n813), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n822), .A2(new_n748), .ZN(new_n830));
  INV_X1    g0630(.A(new_n752), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n390), .B1(new_n765), .B2(new_n216), .ZN(new_n832));
  XNOR2_X1  g0632(.A(KEYINPUT98), .B(G143), .ZN(new_n833));
  AOI22_X1  g0633(.A1(new_n792), .A2(new_n833), .B1(new_n788), .B2(G150), .ZN(new_n834));
  INV_X1    g0634(.A(G137), .ZN(new_n835));
  INV_X1    g0635(.A(G159), .ZN(new_n836));
  OAI221_X1 g0636(.A(new_n834), .B1(new_n835), .B2(new_n790), .C1(new_n836), .C2(new_n785), .ZN(new_n837));
  XOR2_X1   g0637(.A(new_n837), .B(KEYINPUT34), .Z(new_n838));
  AOI211_X1 g0638(.A(new_n832), .B(new_n838), .C1(G68), .C2(new_n770), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n776), .A2(G132), .ZN(new_n840));
  OAI211_X1 g0640(.A(new_n839), .B(new_n840), .C1(new_n219), .C2(new_n780), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n782), .B1(new_n229), .B2(new_n765), .ZN(new_n842));
  XNOR2_X1  g0642(.A(KEYINPUT97), .B(G283), .ZN(new_n843));
  AOI211_X1 g0643(.A(new_n332), .B(new_n842), .C1(new_n788), .C2(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n792), .A2(G294), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n791), .A2(G303), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n770), .A2(G87), .ZN(new_n847));
  INV_X1    g0647(.A(G311), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n847), .B1(new_n848), .B2(new_n775), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n849), .B1(G116), .B2(new_n799), .ZN(new_n850));
  NAND4_X1  g0650(.A1(new_n844), .A2(new_n845), .A3(new_n846), .A4(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n831), .B1(new_n841), .B2(new_n851), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n752), .A2(new_n747), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n854), .A2(G77), .ZN(new_n855));
  OR4_X1    g0655(.A1(new_n813), .A2(new_n830), .A3(new_n852), .A4(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n829), .A2(new_n856), .ZN(G384));
  INV_X1    g0657(.A(KEYINPUT101), .ZN(new_n858));
  XNOR2_X1  g0658(.A(new_n821), .B(KEYINPUT99), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n860), .B1(new_n743), .B2(new_n822), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n663), .A2(new_n307), .ZN(new_n862));
  XOR2_X1   g0662(.A(new_n862), .B(KEYINPUT100), .Z(new_n863));
  INV_X1    g0663(.A(new_n862), .ZN(new_n864));
  AOI22_X1  g0664(.A1(new_n319), .A2(new_n863), .B1(new_n318), .B2(new_n864), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n858), .B1(new_n861), .B2(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n396), .B1(KEYINPUT16), .B2(new_n395), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n407), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n422), .A2(new_n661), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n408), .A2(new_n661), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT37), .ZN(new_n871));
  NAND4_X1  g0671(.A1(new_n412), .A2(new_n870), .A3(new_n871), .A4(new_n417), .ZN(new_n872));
  AND3_X1   g0672(.A1(new_n402), .A2(new_n400), .A3(new_n403), .ZN(new_n873));
  INV_X1    g0673(.A(new_n661), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n410), .A2(new_n874), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n873), .B1(new_n868), .B2(new_n875), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n872), .B1(new_n876), .B2(new_n871), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n869), .A2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT38), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n869), .A2(KEYINPUT38), .A3(new_n877), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n826), .A2(new_n859), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n319), .A2(new_n863), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n318), .A2(new_n864), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n883), .A2(KEYINPUT101), .A3(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n866), .A2(new_n882), .A3(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n414), .A2(new_n415), .A3(new_n874), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(KEYINPUT102), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n402), .B1(new_n410), .B2(new_n874), .ZN(new_n892));
  OAI21_X1  g0692(.A(KEYINPUT37), .B1(new_n873), .B2(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n893), .A2(KEYINPUT103), .A3(new_n872), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT103), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n895), .B(KEYINPUT37), .C1(new_n873), .C2(new_n892), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n401), .A2(new_n404), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n870), .B1(new_n898), .B2(new_n416), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n879), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n881), .A2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT104), .ZN(new_n902));
  OR2_X1    g0702(.A1(new_n902), .A2(KEYINPUT39), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n900), .A2(new_n902), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n880), .A2(new_n881), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n904), .B1(KEYINPUT39), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n617), .A2(new_n679), .ZN(new_n908));
  OR2_X1    g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT102), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n888), .A2(new_n910), .A3(new_n889), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n891), .A2(new_n909), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n724), .A2(KEYINPUT105), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n721), .A2(KEYINPUT31), .A3(new_n663), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT105), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n722), .A2(new_n915), .A3(new_n723), .ZN(new_n916));
  NAND4_X1  g0716(.A1(new_n913), .A2(new_n703), .A3(new_n914), .A4(new_n916), .ZN(new_n917));
  NAND4_X1  g0717(.A1(new_n917), .A2(new_n822), .A3(new_n886), .A4(new_n901), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(KEYINPUT40), .ZN(new_n919));
  AOI21_X1  g0719(.A(KEYINPUT40), .B1(new_n880), .B2(new_n881), .ZN(new_n920));
  NAND4_X1  g0720(.A1(new_n920), .A2(new_n822), .A3(new_n917), .A4(new_n886), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  AND2_X1   g0722(.A1(new_n423), .A2(new_n917), .ZN(new_n923));
  OAI21_X1  g0723(.A(G330), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n924), .B1(new_n922), .B2(new_n923), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n912), .B(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n742), .A2(new_n423), .A3(new_n744), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(new_n621), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n926), .B(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n929), .B1(new_n277), .B2(new_n657), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT35), .ZN(new_n931));
  AOI211_X1 g0731(.A(new_n235), .B(new_n234), .C1(new_n463), .C2(new_n931), .ZN(new_n932));
  OAI211_X1 g0732(.A(new_n932), .B(G116), .C1(new_n931), .C2(new_n463), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n933), .B(KEYINPUT36), .ZN(new_n934));
  NOR3_X1   g0734(.A1(new_n700), .A2(new_n224), .A3(new_n378), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n201), .A2(new_n211), .ZN(new_n936));
  OAI211_X1 g0736(.A(G1), .B(new_n656), .C1(new_n935), .C2(new_n936), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n930), .A2(new_n934), .A3(new_n937), .ZN(G367));
  INV_X1    g0738(.A(new_n759), .ZN(new_n939));
  OAI221_X1 g0739(.A(new_n753), .B1(new_n208), .B2(new_n345), .C1(new_n939), .C2(new_n246), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n390), .B1(new_n776), .B2(G317), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n941), .B1(new_n213), .B2(new_n769), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n942), .B(KEYINPUT109), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n766), .A2(G116), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n944), .B(KEYINPUT46), .ZN(new_n945));
  INV_X1    g0745(.A(new_n788), .ZN(new_n946));
  OAI221_X1 g0746(.A(new_n945), .B1(new_n229), .B2(new_n780), .C1(new_n802), .C2(new_n946), .ZN(new_n947));
  AOI211_X1 g0747(.A(new_n943), .B(new_n947), .C1(G311), .C2(new_n791), .ZN(new_n948));
  INV_X1    g0748(.A(G303), .ZN(new_n949));
  INV_X1    g0749(.A(new_n843), .ZN(new_n950));
  OAI221_X1 g0750(.A(new_n948), .B1(new_n949), .B2(new_n804), .C1(new_n785), .C2(new_n950), .ZN(new_n951));
  XOR2_X1   g0751(.A(new_n951), .B(KEYINPUT110), .Z(new_n952));
  NOR2_X1   g0752(.A1(new_n780), .A2(new_n211), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n953), .B1(G150), .B2(new_n792), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n954), .B(KEYINPUT111), .ZN(new_n955));
  INV_X1    g0755(.A(new_n201), .ZN(new_n956));
  OAI22_X1  g0756(.A1(new_n956), .A2(new_n785), .B1(new_n765), .B2(new_n219), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n332), .B1(new_n835), .B2(new_n775), .ZN(new_n958));
  NOR3_X1   g0758(.A1(new_n955), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n791), .A2(new_n833), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n770), .A2(G77), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n788), .A2(G159), .ZN(new_n962));
  NAND4_X1  g0762(.A1(new_n959), .A2(new_n960), .A3(new_n961), .A4(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n952), .A2(new_n963), .ZN(new_n964));
  XOR2_X1   g0764(.A(new_n964), .B(KEYINPUT47), .Z(new_n965));
  OAI211_X1 g0765(.A(new_n812), .B(new_n940), .C1(new_n965), .C2(new_n831), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n663), .A2(new_n623), .ZN(new_n967));
  MUX2_X1   g0767(.A(new_n632), .B(new_n642), .S(new_n967), .Z(new_n968));
  NOR2_X1   g0768(.A1(new_n968), .A2(new_n750), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n966), .A2(new_n969), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n696), .B(KEYINPUT41), .ZN(new_n971));
  INV_X1    g0771(.A(new_n692), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n972), .A2(new_n684), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT107), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n678), .A2(new_n974), .A3(new_n691), .ZN(new_n975));
  INV_X1    g0775(.A(new_n975), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n974), .B1(new_n678), .B2(new_n691), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n973), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n977), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n979), .A2(new_n684), .A3(new_n975), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n978), .A2(new_n980), .A3(new_n745), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n731), .B1(new_n469), .B2(new_n679), .ZN(new_n982));
  OR2_X1    g0782(.A1(new_n679), .A2(new_n473), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n972), .A2(new_n665), .A3(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT45), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n693), .A2(KEYINPUT45), .A3(new_n984), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT44), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n990), .B1(new_n693), .B2(new_n984), .ZN(new_n991));
  INV_X1    g0791(.A(new_n984), .ZN(new_n992));
  OAI211_X1 g0792(.A(KEYINPUT44), .B(new_n992), .C1(new_n692), .C2(new_n664), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n991), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n989), .A2(new_n994), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n995), .A2(KEYINPUT108), .A3(new_n686), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n686), .A2(KEYINPUT108), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT108), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n685), .A2(new_n998), .ZN(new_n999));
  NAND4_X1  g0799(.A1(new_n989), .A2(new_n994), .A3(new_n997), .A4(new_n999), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n981), .B1(new_n996), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n745), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n971), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1003), .A2(new_n810), .ZN(new_n1004));
  OAI21_X1  g0804(.A(KEYINPUT42), .B1(new_n972), .B2(new_n482), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n479), .B1(new_n992), .B2(new_n575), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1006), .A2(new_n679), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT42), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n692), .A2(new_n1008), .A3(new_n731), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1005), .A2(new_n1007), .A3(new_n1009), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1010), .A2(KEYINPUT43), .A3(new_n968), .ZN(new_n1011));
  OR2_X1    g0811(.A1(new_n968), .A2(KEYINPUT43), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT106), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1010), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n686), .A2(new_n992), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n968), .A2(KEYINPUT43), .ZN(new_n1018));
  NAND4_X1  g0818(.A1(new_n1010), .A2(new_n1014), .A3(new_n1018), .A4(new_n1012), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1016), .A2(new_n1017), .A3(new_n1019), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n1017), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n1011), .A2(new_n1012), .B1(new_n1014), .B2(new_n1010), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n1019), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1021), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1020), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n1025), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n970), .B1(new_n1004), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n1027), .ZN(G387));
  NAND2_X1  g0828(.A1(new_n978), .A2(new_n980), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1029), .A2(new_n1002), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1030), .A2(new_n696), .A3(new_n981), .ZN(new_n1031));
  INV_X1    g0831(.A(G45), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n759), .B1(new_n243), .B2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n698), .B2(new_n755), .ZN(new_n1034));
  OR3_X1    g0834(.A1(new_n324), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1035));
  OAI21_X1  g0835(.A(KEYINPUT50), .B1(new_n324), .B2(G50), .ZN(new_n1036));
  AOI21_X1  g0836(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1035), .A2(new_n1036), .A3(new_n698), .A4(new_n1037), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n1034), .A2(new_n1038), .B1(new_n229), .B2(new_n695), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n780), .A2(new_n345), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n804), .A2(new_n216), .B1(new_n769), .B2(new_n213), .ZN(new_n1041));
  AOI211_X1 g0841(.A(new_n1040), .B(new_n1041), .C1(new_n323), .C2(new_n788), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n790), .A2(new_n836), .B1(new_n785), .B2(new_n211), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n765), .A2(new_n224), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n776), .A2(G150), .ZN(new_n1046));
  NAND4_X1  g0846(.A1(new_n1042), .A2(new_n390), .A3(new_n1045), .A4(new_n1046), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(G311), .A2(new_n788), .B1(new_n792), .B2(G317), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n1048), .B1(new_n949), .B2(new_n785), .C1(new_n805), .C2(new_n790), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT48), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n1050), .B1(new_n802), .B2(new_n765), .C1(new_n780), .C2(new_n950), .ZN(new_n1051));
  XOR2_X1   g0851(.A(new_n1051), .B(KEYINPUT49), .Z(new_n1052));
  AOI21_X1  g0852(.A(new_n390), .B1(new_n776), .B2(G326), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(new_n527), .B2(new_n769), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1047), .B1(new_n1052), .B2(new_n1054), .ZN(new_n1055));
  XOR2_X1   g0855(.A(new_n1055), .B(KEYINPUT112), .Z(new_n1056));
  OAI221_X1 g0856(.A(new_n812), .B1(new_n754), .B2(new_n1039), .C1(new_n1056), .C2(new_n831), .ZN(new_n1057));
  INV_X1    g0857(.A(KEYINPUT113), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n1057), .A2(new_n1058), .B1(new_n678), .B2(new_n749), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1059), .B1(new_n1058), .B2(new_n1057), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n1031), .B(new_n1060), .C1(new_n810), .C2(new_n1029), .ZN(G393));
  NAND3_X1  g0861(.A1(new_n996), .A2(new_n981), .A3(new_n1000), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n697), .B1(new_n1062), .B2(KEYINPUT118), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n981), .ZN(new_n1064));
  AOI211_X1 g0864(.A(new_n998), .B(new_n685), .C1(new_n989), .C2(new_n994), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n1000), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1064), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT118), .ZN(new_n1068));
  NAND4_X1  g0868(.A1(new_n996), .A2(new_n981), .A3(new_n1068), .A4(new_n1000), .ZN(new_n1069));
  AND2_X1   g0869(.A1(new_n1067), .A2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n810), .B1(new_n996), .B2(new_n1000), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n992), .A2(new_n749), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n766), .A2(G68), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n776), .A2(new_n833), .ZN(new_n1074));
  NAND4_X1  g0874(.A1(new_n1073), .A2(new_n847), .A3(new_n1074), .A4(new_n390), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n1075), .A2(KEYINPUT115), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT51), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n804), .A2(new_n836), .B1(new_n790), .B2(new_n321), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1076), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1079), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n781), .A2(G77), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n324), .A2(new_n785), .B1(new_n946), .B2(new_n956), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(new_n1083), .B(KEYINPUT116), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1075), .A2(KEYINPUT115), .ZN(new_n1085));
  NAND4_X1  g0885(.A1(new_n1081), .A2(new_n1082), .A3(new_n1084), .A4(new_n1085), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n949), .A2(new_n946), .B1(new_n950), .B2(new_n765), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n791), .A2(G317), .B1(G311), .B2(new_n792), .ZN(new_n1088));
  XNOR2_X1  g0888(.A(new_n1088), .B(KEYINPUT52), .ZN(new_n1089));
  AOI211_X1 g0889(.A(new_n1087), .B(new_n1089), .C1(G322), .C2(new_n776), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n332), .B1(G294), .B2(new_n799), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n781), .A2(G116), .ZN(new_n1092));
  NAND4_X1  g0892(.A1(new_n1090), .A2(new_n771), .A3(new_n1091), .A4(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n831), .B1(new_n1086), .B2(new_n1093), .ZN(new_n1094));
  OAI221_X1 g0894(.A(new_n753), .B1(new_n213), .B2(new_n208), .C1(new_n939), .C2(new_n250), .ZN(new_n1095));
  AND2_X1   g0895(.A1(new_n1095), .A2(KEYINPUT114), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n1095), .A2(KEYINPUT114), .ZN(new_n1097));
  NOR4_X1   g0897(.A1(new_n1094), .A2(new_n813), .A3(new_n1096), .A4(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1072), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  OAI21_X1  g0900(.A(KEYINPUT117), .B1(new_n1071), .B2(new_n1100), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n811), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1102));
  INV_X1    g0902(.A(KEYINPUT117), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1102), .A2(new_n1103), .A3(new_n1099), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n1063), .A2(new_n1070), .B1(new_n1101), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1105), .ZN(G390));
  NAND2_X1  g0906(.A1(new_n906), .A2(KEYINPUT39), .ZN(new_n1107));
  OR2_X1    g0907(.A1(new_n901), .A2(new_n903), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n865), .B1(new_n826), .B2(new_n859), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n908), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n1107), .B(new_n1108), .C1(new_n1109), .C2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n727), .A2(G330), .A3(new_n822), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n1112), .A2(new_n865), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n819), .B1(new_n737), .B2(new_n741), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n821), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n865), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n901), .A2(new_n908), .ZN(new_n1117));
  OAI211_X1 g0917(.A(new_n1111), .B(new_n1113), .C1(new_n1116), .C2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  NAND4_X1  g0919(.A1(new_n917), .A2(G330), .A3(new_n886), .A4(new_n822), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n733), .B(new_n637), .C1(new_n650), .C2(new_n649), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1122), .B1(new_n524), .B2(new_n730), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n729), .B1(new_n1123), .B2(new_n663), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n740), .A2(KEYINPUT94), .A3(new_n679), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n820), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n886), .B1(new_n1126), .B2(new_n821), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1117), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1121), .B1(new_n1129), .B2(new_n1111), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n1119), .A2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1112), .A2(new_n865), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(new_n1120), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1133), .A2(new_n883), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n821), .B1(new_n1135), .B2(new_n819), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n728), .A2(new_n822), .A3(new_n886), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n917), .A2(G330), .A3(new_n822), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1138), .A2(new_n865), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1136), .A2(new_n1137), .A3(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1134), .A2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n423), .A2(G330), .A3(new_n917), .ZN(new_n1142));
  AND3_X1   g0942(.A1(new_n927), .A2(new_n621), .A3(new_n1142), .ZN(new_n1143));
  AND3_X1   g0943(.A1(new_n1141), .A2(KEYINPUT120), .A3(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(KEYINPUT120), .B1(new_n1141), .B2(new_n1143), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1131), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n908), .B1(new_n861), .B2(new_n865), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(new_n1127), .A2(new_n1128), .B1(new_n907), .B2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1118), .B1(new_n1148), .B2(new_n1121), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n927), .A2(new_n621), .A3(new_n1142), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1150), .B1(new_n1134), .B2(new_n1140), .ZN(new_n1151));
  AND3_X1   g0951(.A1(new_n1149), .A2(KEYINPUT119), .A3(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(KEYINPUT119), .B1(new_n1149), .B2(new_n1151), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n1146), .B(new_n696), .C1(new_n1152), .C2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n907), .A2(new_n747), .ZN(new_n1155));
  XOR2_X1   g0955(.A(KEYINPUT54), .B(G143), .Z(new_n1156));
  AOI22_X1  g0956(.A1(G125), .A2(new_n776), .B1(new_n799), .B2(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(G128), .ZN(new_n1158));
  OAI211_X1 g0958(.A(new_n1157), .B(new_n332), .C1(new_n1158), .C2(new_n790), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n765), .A2(new_n321), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(new_n1160), .B(KEYINPUT53), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(new_n781), .A2(G159), .B1(new_n770), .B2(new_n201), .ZN(new_n1162));
  OAI211_X1 g0962(.A(new_n1161), .B(new_n1162), .C1(new_n835), .C2(new_n946), .ZN(new_n1163));
  AOI211_X1 g0963(.A(new_n1159), .B(new_n1163), .C1(G132), .C2(new_n792), .ZN(new_n1164));
  OAI221_X1 g0964(.A(new_n1082), .B1(new_n211), .B2(new_n769), .C1(new_n229), .C2(new_n946), .ZN(new_n1165));
  OAI221_X1 g0965(.A(new_n767), .B1(new_n527), .B2(new_n804), .C1(new_n796), .C2(new_n790), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n333), .B1(new_n802), .B2(new_n775), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n785), .A2(new_n213), .ZN(new_n1168));
  NOR4_X1   g0968(.A1(new_n1165), .A2(new_n1166), .A3(new_n1167), .A4(new_n1168), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n752), .B1(new_n1164), .B2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n853), .A2(new_n324), .ZN(new_n1171));
  AND4_X1   g0971(.A1(new_n812), .A2(new_n1155), .A3(new_n1170), .A4(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1172), .B1(new_n1149), .B2(new_n811), .ZN(new_n1173));
  AND3_X1   g0973(.A1(new_n1154), .A2(KEYINPUT121), .A3(new_n1173), .ZN(new_n1174));
  AOI21_X1  g0974(.A(KEYINPUT121), .B1(new_n1154), .B2(new_n1173), .ZN(new_n1175));
  OR2_X1    g0975(.A1(new_n1174), .A2(new_n1175), .ZN(G378));
  INV_X1    g0976(.A(KEYINPUT57), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1149), .A2(new_n1151), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT119), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1149), .A2(KEYINPUT119), .A3(new_n1151), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1150), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n327), .A2(new_n661), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n341), .A2(new_n360), .A3(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1183), .B1(new_n341), .B2(new_n360), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  XOR2_X1   g0987(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1188));
  XNOR2_X1  g0988(.A(new_n1187), .B(new_n1188), .ZN(new_n1189));
  AND3_X1   g0989(.A1(new_n917), .A2(new_n822), .A3(new_n886), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n1190), .A2(new_n920), .B1(new_n918), .B2(KEYINPUT40), .ZN(new_n1191));
  INV_X1    g0991(.A(G330), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1189), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1189), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n922), .A2(new_n1194), .A3(G330), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1193), .A2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n912), .B1(new_n1197), .B2(KEYINPUT122), .ZN(new_n1198));
  AOI21_X1  g0998(.A(KEYINPUT122), .B1(new_n1193), .B2(new_n1195), .ZN(new_n1199));
  NAND4_X1  g0999(.A1(new_n1199), .A2(new_n909), .A3(new_n891), .A4(new_n911), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1198), .A2(new_n1200), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1177), .B1(new_n1182), .B2(new_n1201), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1143), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT123), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n912), .A2(new_n1204), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n891), .A2(KEYINPUT123), .A3(new_n909), .A4(new_n911), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1205), .A2(new_n1196), .A3(new_n1206), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n912), .A2(new_n1197), .A3(new_n1204), .ZN(new_n1208));
  NAND4_X1  g1008(.A1(new_n1203), .A2(KEYINPUT57), .A3(new_n1207), .A4(new_n1208), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1202), .A2(new_n1209), .A3(new_n696), .ZN(new_n1210));
  XNOR2_X1  g1010(.A(new_n912), .B(new_n1199), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1211), .A2(new_n811), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n813), .B1(new_n1189), .B2(new_n747), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n270), .B1(new_n790), .B2(new_n527), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n804), .A2(new_n229), .B1(new_n785), .B2(new_n345), .ZN(new_n1215));
  AOI211_X1 g1015(.A(new_n1214), .B(new_n1215), .C1(G283), .C2(new_n776), .ZN(new_n1216));
  AOI211_X1 g1016(.A(new_n1044), .B(new_n953), .C1(G97), .C2(new_n788), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n770), .A2(G58), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1216), .A2(new_n1217), .A3(new_n392), .A4(new_n1218), .ZN(new_n1219));
  XNOR2_X1  g1019(.A(new_n1219), .B(KEYINPUT58), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n216), .B1(new_n255), .B2(G41), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n781), .A2(G150), .B1(new_n791), .B2(G125), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n799), .A2(G137), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n788), .A2(G132), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n766), .A2(new_n1156), .B1(G128), .B2(new_n792), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(new_n1222), .A2(new_n1223), .A3(new_n1224), .A4(new_n1225), .ZN(new_n1226));
  XOR2_X1   g1026(.A(new_n1226), .B(KEYINPUT59), .Z(new_n1227));
  OAI21_X1  g1027(.A(new_n270), .B1(new_n769), .B2(new_n836), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1228), .B1(G124), .B2(new_n776), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1227), .A2(new_n259), .A3(new_n1229), .ZN(new_n1230));
  AND3_X1   g1030(.A1(new_n1220), .A2(new_n1221), .A3(new_n1230), .ZN(new_n1231));
  OAI221_X1 g1031(.A(new_n1213), .B1(new_n201), .B2(new_n854), .C1(new_n831), .C2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1212), .A2(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1210), .A2(new_n1234), .ZN(G375));
  OAI221_X1 g1035(.A(new_n971), .B1(new_n1143), .B2(new_n1141), .C1(new_n1144), .C2(new_n1145), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1040), .B1(G97), .B2(new_n766), .ZN(new_n1237));
  OAI221_X1 g1037(.A(new_n1237), .B1(new_n229), .B2(new_n785), .C1(new_n949), .C2(new_n775), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n946), .A2(new_n527), .ZN(new_n1239));
  OAI221_X1 g1039(.A(new_n961), .B1(new_n796), .B2(new_n804), .C1(new_n802), .C2(new_n790), .ZN(new_n1240));
  NOR4_X1   g1040(.A1(new_n1238), .A2(new_n332), .A3(new_n1239), .A4(new_n1240), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n765), .A2(new_n836), .B1(new_n775), .B2(new_n1158), .ZN(new_n1242));
  XNOR2_X1  g1042(.A(new_n1242), .B(KEYINPUT124), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(new_n791), .A2(G132), .B1(new_n799), .B2(G150), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1244), .B1(new_n835), .B2(new_n804), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1156), .A2(new_n788), .ZN(new_n1246));
  OAI211_X1 g1046(.A(new_n1218), .B(new_n1246), .C1(new_n216), .C2(new_n780), .ZN(new_n1247));
  NOR4_X1   g1047(.A1(new_n1243), .A2(new_n1245), .A3(new_n392), .A4(new_n1247), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n752), .B1(new_n1241), .B2(new_n1248), .ZN(new_n1249));
  OAI211_X1 g1049(.A(new_n1249), .B(new_n812), .C1(G68), .C2(new_n854), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1250), .B1(new_n865), .B2(new_n747), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1251), .B1(new_n1141), .B2(new_n811), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1236), .A2(new_n1252), .ZN(G381));
  NAND2_X1  g1053(.A1(new_n1203), .A2(new_n1211), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n697), .B1(new_n1254), .B2(new_n1177), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1233), .B1(new_n1255), .B2(new_n1209), .ZN(new_n1256));
  AND2_X1   g1056(.A1(new_n1154), .A2(new_n1173), .ZN(new_n1257));
  AND2_X1   g1057(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(G381), .A2(G384), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n971), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1260), .B1(new_n1067), .B2(new_n745), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1026), .B1(new_n1261), .B2(new_n811), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n970), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1101), .A2(new_n1104), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1070), .A2(new_n1063), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1262), .A2(new_n1263), .A3(new_n1264), .A4(new_n1265), .ZN(new_n1266));
  NOR3_X1   g1066(.A1(new_n1266), .A2(G396), .A3(G393), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1258), .A2(new_n1259), .A3(new_n1267), .ZN(G407));
  INV_X1    g1068(.A(new_n1258), .ZN(new_n1269));
  OAI211_X1 g1069(.A(G407), .B(G213), .C1(G343), .C2(new_n1269), .ZN(G409));
  NAND3_X1  g1070(.A1(new_n1207), .A2(new_n811), .A3(new_n1208), .ZN(new_n1271));
  OAI211_X1 g1071(.A(new_n1232), .B(new_n1271), .C1(new_n1254), .C2(new_n1260), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1272), .A2(new_n1257), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1273), .B1(G375), .B2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(G213), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1276), .A2(G343), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1277), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1279), .A2(KEYINPUT60), .ZN(new_n1280));
  OAI21_X1  g1080(.A(KEYINPUT125), .B1(new_n1280), .B2(new_n1151), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n697), .B1(new_n1279), .B2(KEYINPUT60), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1151), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT125), .ZN(new_n1284));
  OAI211_X1 g1084(.A(new_n1283), .B(new_n1284), .C1(KEYINPUT60), .C2(new_n1279), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1281), .A2(new_n1282), .A3(new_n1285), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1286), .A2(G384), .A3(new_n1252), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(G384), .B1(new_n1286), .B2(new_n1252), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1275), .A2(new_n1278), .A3(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1291), .A2(KEYINPUT62), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT61), .ZN(new_n1293));
  OAI211_X1 g1093(.A(G2897), .B(new_n1277), .C1(new_n1288), .C2(new_n1289), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1289), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1277), .A2(G2897), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1295), .A2(new_n1287), .A3(new_n1296), .ZN(new_n1297));
  AND2_X1   g1097(.A1(new_n1294), .A2(new_n1297), .ZN(new_n1298));
  AOI22_X1  g1098(.A1(new_n1256), .A2(G378), .B1(new_n1257), .B2(new_n1272), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1298), .B1(new_n1299), .B2(new_n1277), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT62), .ZN(new_n1301));
  NAND4_X1  g1101(.A1(new_n1275), .A2(new_n1301), .A3(new_n1278), .A4(new_n1290), .ZN(new_n1302));
  NAND4_X1  g1102(.A1(new_n1292), .A2(new_n1293), .A3(new_n1300), .A4(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1264), .ZN(new_n1304));
  AND3_X1   g1104(.A1(new_n1063), .A2(new_n1067), .A3(new_n1069), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1025), .B1(new_n1003), .B2(new_n810), .ZN(new_n1306));
  OAI22_X1  g1106(.A1(new_n1304), .A2(new_n1305), .B1(new_n1306), .B2(new_n970), .ZN(new_n1307));
  XNOR2_X1  g1107(.A(G393), .B(G396), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1308), .ZN(new_n1309));
  AND4_X1   g1109(.A1(KEYINPUT126), .A2(new_n1307), .A3(new_n1266), .A4(new_n1309), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1308), .B1(new_n1027), .B2(new_n1105), .ZN(new_n1311));
  AOI21_X1  g1111(.A(KEYINPUT126), .B1(new_n1311), .B2(new_n1307), .ZN(new_n1312));
  NOR2_X1   g1112(.A1(new_n1310), .A2(new_n1312), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(G387), .A2(KEYINPUT127), .A3(new_n1105), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT127), .ZN(new_n1315));
  OAI21_X1  g1115(.A(G390), .B1(new_n1027), .B2(new_n1315), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1314), .A2(new_n1316), .A3(new_n1308), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1313), .A2(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1303), .A2(new_n1319), .ZN(new_n1320));
  AOI21_X1  g1120(.A(KEYINPUT61), .B1(new_n1313), .B2(new_n1317), .ZN(new_n1321));
  AND3_X1   g1121(.A1(new_n1275), .A2(new_n1278), .A3(new_n1290), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1322), .A2(KEYINPUT63), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT63), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1275), .A2(new_n1278), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1324), .B1(new_n1325), .B2(new_n1298), .ZN(new_n1326));
  OAI211_X1 g1126(.A(new_n1321), .B(new_n1323), .C1(new_n1326), .C2(new_n1322), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1320), .A2(new_n1327), .ZN(G405));
  NAND2_X1  g1128(.A1(new_n1256), .A2(G378), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(G375), .A2(new_n1257), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1329), .A2(new_n1330), .ZN(new_n1331));
  XNOR2_X1  g1131(.A(new_n1331), .B(new_n1290), .ZN(new_n1332));
  NOR2_X1   g1132(.A1(new_n1332), .A2(new_n1318), .ZN(new_n1333));
  OR2_X1    g1133(.A1(new_n1331), .A2(new_n1290), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1331), .A2(new_n1290), .ZN(new_n1335));
  AOI22_X1  g1135(.A1(new_n1334), .A2(new_n1335), .B1(new_n1313), .B2(new_n1317), .ZN(new_n1336));
  NOR2_X1   g1136(.A1(new_n1333), .A2(new_n1336), .ZN(G402));
endmodule


