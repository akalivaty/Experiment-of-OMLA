//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 0 0 0 1 0 1 1 1 1 1 1 0 0 1 0 1 0 0 1 1 1 1 0 1 1 1 0 1 1 0 1 0 1 0 1 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:48 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1271, new_n1272, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(KEYINPUT64), .ZN(new_n202));
  XNOR2_X1  g0002(.A(new_n201), .B(new_n202), .ZN(new_n203));
  INV_X1    g0003(.A(G77), .ZN(new_n204));
  AND2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n209), .B(KEYINPUT0), .ZN(new_n210));
  XNOR2_X1  g0010(.A(KEYINPUT65), .B(G20), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(G58), .ZN(new_n214));
  INV_X1    g0014(.A(G68), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(G50), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n213), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n220));
  INV_X1    g0020(.A(G244), .ZN(new_n221));
  INV_X1    g0021(.A(G107), .ZN(new_n222));
  INV_X1    g0022(.A(G264), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n220), .B1(new_n204), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n207), .B1(new_n224), .B2(new_n227), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n210), .B(new_n219), .C1(KEYINPUT1), .C2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT2), .B(G226), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G264), .B(G270), .Z(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XOR2_X1   g0039(.A(G107), .B(G116), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G50), .B(G68), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G58), .B(G77), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G351));
  NOR2_X1   g0045(.A1(G20), .A2(G33), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(G150), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n211), .A2(G33), .ZN(new_n248));
  XNOR2_X1  g0048(.A(KEYINPUT8), .B(G58), .ZN(new_n249));
  INV_X1    g0049(.A(G20), .ZN(new_n250));
  OAI221_X1 g0050(.A(new_n247), .B1(new_n248), .B2(new_n249), .C1(new_n203), .C2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT69), .ZN(new_n252));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n252), .B1(new_n207), .B2(new_n253), .ZN(new_n254));
  NAND4_X1  g0054(.A1(KEYINPUT69), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n254), .A2(new_n212), .A3(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G50), .ZN(new_n257));
  INV_X1    g0057(.A(G1), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n258), .A2(G13), .A3(G20), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  AOI22_X1  g0060(.A1(new_n251), .A2(new_n256), .B1(new_n257), .B2(new_n260), .ZN(new_n261));
  NAND4_X1  g0061(.A1(new_n254), .A2(new_n212), .A3(new_n255), .A4(new_n259), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(KEYINPUT70), .ZN(new_n263));
  AND2_X1   g0063(.A1(new_n255), .A2(new_n212), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT70), .ZN(new_n265));
  NAND4_X1  g0065(.A1(new_n264), .A2(new_n265), .A3(new_n254), .A4(new_n259), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n263), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n258), .A2(G20), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n267), .A2(G50), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n261), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(KEYINPUT9), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT9), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n261), .A2(new_n272), .A3(new_n269), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G274), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT67), .ZN(new_n276));
  NAND2_X1  g0076(.A1(G33), .A2(G41), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n212), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(KEYINPUT67), .A2(G33), .A3(G41), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n275), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT66), .ZN(new_n281));
  NOR2_X1   g0081(.A1(G41), .A2(G45), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n281), .B1(new_n282), .B2(G1), .ZN(new_n283));
  OAI211_X1 g0083(.A(new_n258), .B(KEYINPUT66), .C1(G41), .C2(G45), .ZN(new_n284));
  AND2_X1   g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n282), .A2(G1), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n286), .B1(new_n278), .B2(new_n279), .ZN(new_n287));
  AOI22_X1  g0087(.A1(new_n280), .A2(new_n285), .B1(new_n287), .B2(G226), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT3), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(new_n253), .ZN(new_n290));
  NAND2_X1  g0090(.A1(KEYINPUT3), .A2(G33), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n292), .A2(G223), .A3(G1698), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n293), .B1(new_n204), .B2(new_n292), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT68), .ZN(new_n295));
  AND2_X1   g0095(.A1(KEYINPUT3), .A2(G33), .ZN(new_n296));
  NOR2_X1   g0096(.A1(KEYINPUT3), .A2(G33), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G1698), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(G222), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n295), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  NAND4_X1  g0101(.A1(new_n292), .A2(KEYINPUT68), .A3(G222), .A4(new_n299), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n294), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(new_n212), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(new_n277), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n288), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(G200), .ZN(new_n307));
  OAI211_X1 g0107(.A(G190), .B(new_n288), .C1(new_n303), .C2(new_n305), .ZN(new_n308));
  AND2_X1   g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n274), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n307), .A2(KEYINPUT74), .A3(new_n308), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT10), .ZN(new_n312));
  AND2_X1   g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n310), .A2(new_n313), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n274), .B(new_n309), .C1(KEYINPUT74), .C2(KEYINPUT10), .ZN(new_n315));
  AND2_X1   g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n249), .B1(new_n258), .B2(G20), .ZN(new_n317));
  AOI22_X1  g0117(.A1(new_n267), .A2(new_n317), .B1(new_n260), .B2(new_n249), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT7), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n298), .A2(new_n211), .A3(new_n319), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n290), .A2(new_n250), .A3(new_n291), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(KEYINPUT7), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n320), .A2(new_n322), .A3(G68), .ZN(new_n323));
  NAND2_X1  g0123(.A1(G58), .A2(G68), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT77), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g0126(.A1(KEYINPUT77), .A2(G58), .A3(G68), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n326), .A2(new_n216), .A3(new_n327), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n250), .A2(new_n253), .A3(G159), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(KEYINPUT78), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT78), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n246), .A2(new_n331), .A3(G159), .ZN(new_n332));
  AOI22_X1  g0132(.A1(G20), .A2(new_n328), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n323), .A2(KEYINPUT16), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(new_n256), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n250), .A2(KEYINPUT65), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT65), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(G20), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  OAI21_X1  g0139(.A(KEYINPUT7), .B1(new_n339), .B2(new_n292), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n298), .A2(new_n319), .A3(new_n250), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n340), .A2(G68), .A3(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(KEYINPUT16), .B1(new_n342), .B2(new_n333), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n318), .B1(new_n335), .B2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT18), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n277), .A2(new_n276), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n346), .A2(new_n304), .A3(new_n279), .ZN(new_n347));
  NAND4_X1  g0147(.A1(new_n347), .A2(G274), .A3(new_n283), .A4(new_n284), .ZN(new_n348));
  INV_X1    g0148(.A(new_n286), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n349), .A2(new_n347), .A3(G232), .ZN(new_n350));
  MUX2_X1   g0150(.A(G223), .B(G226), .S(G1698), .Z(new_n351));
  AOI22_X1  g0151(.A1(new_n351), .A2(new_n292), .B1(G33), .B2(G87), .ZN(new_n352));
  OAI211_X1 g0152(.A(new_n348), .B(new_n350), .C1(new_n352), .C2(new_n305), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(G169), .ZN(new_n354));
  INV_X1    g0154(.A(G179), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n354), .B1(new_n355), .B2(new_n353), .ZN(new_n356));
  AND3_X1   g0156(.A1(new_n344), .A2(new_n345), .A3(new_n356), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n345), .B1(new_n344), .B2(new_n356), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  XNOR2_X1  g0159(.A(KEYINPUT15), .B(G87), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n248), .A2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(new_n246), .ZN(new_n362));
  OAI22_X1  g0162(.A1(new_n204), .A2(new_n211), .B1(new_n249), .B2(new_n362), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n256), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  XNOR2_X1  g0164(.A(new_n364), .B(KEYINPUT72), .ZN(new_n365));
  INV_X1    g0165(.A(new_n262), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n204), .B1(new_n258), .B2(G20), .ZN(new_n367));
  AOI22_X1  g0167(.A1(new_n366), .A2(new_n367), .B1(new_n204), .B2(new_n260), .ZN(new_n368));
  NOR2_X1   g0168(.A1(G232), .A2(G1698), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n299), .A2(G238), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n292), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(new_n305), .ZN(new_n372));
  OAI211_X1 g0172(.A(new_n371), .B(new_n372), .C1(G107), .C2(new_n292), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n287), .A2(G244), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n373), .A2(new_n348), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(G200), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n365), .A2(new_n368), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(KEYINPUT73), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT73), .ZN(new_n379));
  NAND4_X1  g0179(.A1(new_n365), .A2(new_n379), .A3(new_n368), .A4(new_n376), .ZN(new_n380));
  INV_X1    g0180(.A(G190), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n375), .A2(new_n381), .ZN(new_n382));
  XNOR2_X1  g0182(.A(new_n382), .B(KEYINPUT71), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n378), .A2(new_n380), .A3(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT17), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n351), .A2(new_n292), .ZN(new_n386));
  NAND2_X1  g0186(.A1(G33), .A2(G87), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(new_n372), .ZN(new_n389));
  NAND4_X1  g0189(.A1(new_n389), .A2(G190), .A3(new_n348), .A4(new_n350), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n353), .A2(G200), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n385), .B1(new_n344), .B2(new_n392), .ZN(new_n393));
  AND2_X1   g0193(.A1(new_n390), .A2(new_n391), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n342), .A2(new_n333), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT16), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n397), .A2(new_n256), .A3(new_n334), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n394), .A2(new_n398), .A3(KEYINPUT17), .A4(new_n318), .ZN(new_n399));
  AND2_X1   g0199(.A1(new_n393), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n365), .A2(new_n368), .ZN(new_n401));
  INV_X1    g0201(.A(G169), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n375), .A2(new_n402), .ZN(new_n403));
  OAI211_X1 g0203(.A(new_n401), .B(new_n403), .C1(G179), .C2(new_n375), .ZN(new_n404));
  AND4_X1   g0204(.A1(new_n359), .A2(new_n384), .A3(new_n400), .A4(new_n404), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n349), .A2(new_n347), .A3(G238), .ZN(new_n406));
  NOR2_X1   g0206(.A1(G226), .A2(G1698), .ZN(new_n407));
  INV_X1    g0207(.A(G232), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n407), .B1(new_n408), .B2(G1698), .ZN(new_n409));
  AOI22_X1  g0209(.A1(new_n409), .A2(new_n292), .B1(G33), .B2(G97), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n406), .B1(new_n410), .B2(new_n305), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n348), .A2(KEYINPUT75), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT75), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n285), .A2(new_n280), .A3(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n411), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT13), .ZN(new_n416));
  NOR3_X1   g0216(.A1(new_n415), .A2(KEYINPUT76), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n412), .A2(new_n414), .ZN(new_n418));
  NAND2_X1  g0218(.A1(G33), .A2(G97), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n408), .A2(G1698), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n420), .B1(G226), .B2(G1698), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n419), .B1(new_n421), .B2(new_n298), .ZN(new_n422));
  AOI22_X1  g0222(.A1(new_n422), .A2(new_n372), .B1(new_n287), .B2(G238), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n416), .B1(new_n418), .B2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT76), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n418), .A2(new_n423), .ZN(new_n427));
  OAI21_X1  g0227(.A(G190), .B1(new_n427), .B2(KEYINPUT13), .ZN(new_n428));
  NOR3_X1   g0228(.A1(new_n417), .A2(new_n426), .A3(new_n428), .ZN(new_n429));
  AND3_X1   g0229(.A1(new_n418), .A2(new_n416), .A3(new_n423), .ZN(new_n430));
  OAI21_X1  g0230(.A(G200), .B1(new_n430), .B2(new_n424), .ZN(new_n431));
  AOI22_X1  g0231(.A1(new_n246), .A2(G50), .B1(G20), .B2(new_n215), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n432), .B1(new_n248), .B2(new_n204), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(new_n256), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT11), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n260), .A2(new_n215), .ZN(new_n437));
  XNOR2_X1  g0237(.A(new_n437), .B(KEYINPUT12), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n366), .A2(G68), .A3(new_n268), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n440), .B1(new_n434), .B2(new_n435), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n431), .A2(new_n442), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n429), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n442), .ZN(new_n445));
  OAI21_X1  g0245(.A(G169), .B1(new_n430), .B2(new_n424), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(KEYINPUT14), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT14), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n448), .B(G169), .C1(new_n430), .C2(new_n424), .ZN(new_n449));
  OAI21_X1  g0249(.A(KEYINPUT76), .B1(new_n415), .B2(new_n416), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n355), .B1(new_n415), .B2(new_n416), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n424), .A2(new_n425), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n450), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n447), .A2(new_n449), .A3(new_n453), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n444), .B1(new_n445), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n306), .A2(new_n402), .ZN(new_n456));
  OAI211_X1 g0256(.A(new_n456), .B(new_n270), .C1(G179), .C2(new_n306), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n316), .A2(new_n405), .A3(new_n455), .A4(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT5), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(G41), .ZN(new_n461));
  INV_X1    g0261(.A(G41), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(KEYINPUT5), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n461), .A2(new_n463), .A3(new_n258), .A4(G45), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(new_n347), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n465), .A2(new_n223), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT87), .ZN(new_n467));
  INV_X1    g0267(.A(G257), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(G1698), .ZN(new_n469));
  OAI221_X1 g0269(.A(new_n469), .B1(G250), .B2(G1698), .C1(new_n296), .C2(new_n297), .ZN(new_n470));
  NAND2_X1  g0270(.A1(G33), .A2(G294), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n305), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n466), .B1(new_n467), .B2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT80), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n474), .B1(new_n460), .B2(G41), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n462), .A2(KEYINPUT80), .A3(KEYINPUT5), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n462), .A2(KEYINPUT5), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n258), .A2(G45), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n347), .A2(new_n477), .A3(new_n480), .A4(G274), .ZN(new_n481));
  NOR2_X1   g0281(.A1(G250), .A2(G1698), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n482), .B1(new_n468), .B2(G1698), .ZN(new_n483));
  AOI22_X1  g0283(.A1(new_n483), .A2(new_n292), .B1(G33), .B2(G294), .ZN(new_n484));
  OAI21_X1  g0284(.A(KEYINPUT87), .B1(new_n484), .B2(new_n305), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n473), .A2(new_n481), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(G169), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n466), .A2(new_n472), .ZN(new_n488));
  AND2_X1   g0288(.A1(new_n488), .A2(new_n481), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(G179), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n487), .A2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(new_n256), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n292), .A2(new_n211), .A3(G87), .ZN(new_n493));
  XNOR2_X1  g0293(.A(KEYINPUT84), .B(KEYINPUT22), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(KEYINPUT23), .A2(G107), .ZN(new_n497));
  AOI21_X1  g0297(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n497), .B1(new_n498), .B2(G20), .ZN(new_n499));
  NOR2_X1   g0299(.A1(KEYINPUT23), .A2(G107), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n499), .B1(new_n339), .B2(new_n500), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n211), .A2(new_n292), .A3(new_n494), .A4(G87), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n496), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(KEYINPUT24), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT24), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n496), .A2(new_n501), .A3(new_n505), .A4(new_n502), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n492), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(KEYINPUT85), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n260), .A2(new_n222), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT86), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n510), .A2(new_n511), .A3(KEYINPUT25), .ZN(new_n512));
  XOR2_X1   g0312(.A(KEYINPUT86), .B(KEYINPUT25), .Z(new_n513));
  OAI21_X1  g0313(.A(new_n512), .B1(new_n510), .B2(new_n513), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n253), .A2(G1), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n262), .A2(new_n515), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n514), .B1(G107), .B2(new_n516), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n517), .B1(new_n507), .B2(KEYINPUT85), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n491), .B1(new_n509), .B2(new_n518), .ZN(new_n519));
  OR2_X1    g0319(.A1(new_n507), .A2(KEYINPUT85), .ZN(new_n520));
  OAI22_X1  g0320(.A1(new_n486), .A2(G190), .B1(new_n489), .B2(G200), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n520), .A2(new_n521), .A3(new_n508), .A4(new_n517), .ZN(new_n522));
  AND2_X1   g0322(.A1(new_n519), .A2(new_n522), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n221), .A2(G1698), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n524), .B(KEYINPUT4), .C1(new_n297), .C2(new_n296), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(KEYINPUT79), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT79), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n292), .A2(new_n527), .A3(KEYINPUT4), .A4(new_n524), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  OAI211_X1 g0329(.A(G250), .B(G1698), .C1(new_n296), .C2(new_n297), .ZN(new_n530));
  NAND2_X1  g0330(.A1(G33), .A2(G283), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n299), .A2(G244), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n532), .B1(new_n290), .B2(new_n291), .ZN(new_n533));
  OAI211_X1 g0333(.A(new_n530), .B(new_n531), .C1(new_n533), .C2(KEYINPUT4), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n372), .B1(new_n529), .B2(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n464), .A2(new_n347), .A3(G257), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n481), .A2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n535), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(G200), .ZN(new_n540));
  AND2_X1   g0340(.A1(new_n530), .A2(new_n531), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT4), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n542), .B1(new_n298), .B2(new_n532), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n541), .A2(new_n543), .A3(new_n526), .A4(new_n528), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n537), .B1(new_n544), .B2(new_n372), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(G190), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n259), .A2(G97), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n362), .A2(new_n204), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT6), .ZN(new_n549));
  INV_X1    g0349(.A(G97), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n550), .A2(new_n222), .ZN(new_n551));
  NOR2_X1   g0351(.A1(G97), .A2(G107), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n549), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NOR3_X1   g0353(.A1(new_n549), .A2(new_n550), .A3(G107), .ZN(new_n554));
  INV_X1    g0354(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n548), .B1(new_n556), .B2(new_n339), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n340), .A2(G107), .A3(new_n341), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n547), .B1(new_n559), .B2(new_n256), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n516), .A2(G97), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n540), .A2(new_n546), .A3(new_n560), .A4(new_n561), .ZN(new_n562));
  AND3_X1   g0362(.A1(new_n340), .A2(G107), .A3(new_n341), .ZN(new_n563));
  XNOR2_X1  g0363(.A(G97), .B(G107), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n554), .B1(new_n549), .B2(new_n564), .ZN(new_n565));
  OAI22_X1  g0365(.A1(new_n565), .A2(new_n211), .B1(new_n204), .B2(new_n362), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n256), .B1(new_n563), .B2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(new_n547), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n567), .A2(new_n561), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n539), .A2(new_n402), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n545), .A2(new_n355), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n562), .A2(new_n572), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n336), .A2(new_n338), .A3(G33), .A4(G97), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT19), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(G87), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n552), .A2(new_n577), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n419), .A2(new_n575), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n578), .B1(new_n339), .B2(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n292), .A2(new_n211), .A3(G68), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n576), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n256), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n360), .A2(new_n260), .ZN(new_n584));
  INV_X1    g0384(.A(new_n360), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n516), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n583), .A2(new_n584), .A3(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(G250), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n479), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n258), .A2(new_n275), .A3(G45), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n347), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  NOR2_X1   g0391(.A1(G238), .A2(G1698), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n592), .B1(new_n221), .B2(G1698), .ZN(new_n593));
  AOI22_X1  g0393(.A1(new_n593), .A2(new_n292), .B1(G33), .B2(G116), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n591), .B1(new_n594), .B2(new_n305), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(new_n402), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n221), .A2(G1698), .ZN(new_n597));
  OAI221_X1 g0397(.A(new_n597), .B1(G238), .B2(G1698), .C1(new_n296), .C2(new_n297), .ZN(new_n598));
  NAND2_X1  g0398(.A1(G33), .A2(G116), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AND2_X1   g0400(.A1(new_n589), .A2(new_n590), .ZN(new_n601));
  AOI22_X1  g0401(.A1(new_n600), .A2(new_n372), .B1(new_n347), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(new_n355), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n587), .A2(new_n596), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n602), .A2(G190), .ZN(new_n605));
  AOI22_X1  g0405(.A1(new_n582), .A2(new_n256), .B1(new_n260), .B2(new_n360), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n595), .A2(G200), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n516), .A2(G87), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n605), .A2(new_n606), .A3(new_n607), .A4(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n604), .A2(new_n609), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n573), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n253), .A2(G97), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n211), .A2(new_n531), .A3(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(G116), .ZN(new_n614));
  AOI22_X1  g0414(.A1(new_n613), .A2(KEYINPUT82), .B1(G20), .B2(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT82), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n211), .A2(new_n616), .A3(new_n531), .A4(new_n612), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n615), .A2(KEYINPUT20), .A3(new_n256), .A4(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n612), .A2(new_n531), .ZN(new_n619));
  OAI21_X1  g0419(.A(KEYINPUT82), .B1(new_n339), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n614), .A2(G20), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n620), .A2(new_n617), .A3(new_n256), .A4(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT20), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  AOI22_X1  g0424(.A1(new_n618), .A2(new_n624), .B1(new_n614), .B2(new_n260), .ZN(new_n625));
  NOR3_X1   g0425(.A1(new_n262), .A2(new_n614), .A3(new_n515), .ZN(new_n626));
  XNOR2_X1  g0426(.A(new_n626), .B(KEYINPUT81), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  NOR2_X1   g0428(.A1(G257), .A2(G1698), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n299), .A2(G264), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n292), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(G303), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n298), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n631), .A2(new_n372), .A3(new_n633), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n464), .A2(new_n347), .A3(G270), .ZN(new_n635));
  AND4_X1   g0435(.A1(G179), .A2(new_n634), .A3(new_n481), .A4(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n628), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(KEYINPUT83), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT83), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n628), .A2(new_n639), .A3(new_n636), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n634), .A2(new_n481), .A3(new_n635), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(G169), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  AOI21_X1  g0444(.A(KEYINPUT21), .B1(new_n628), .B2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT21), .ZN(new_n646));
  AOI211_X1 g0446(.A(new_n646), .B(new_n643), .C1(new_n625), .C2(new_n627), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n628), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n642), .A2(G200), .ZN(new_n650));
  OAI211_X1 g0450(.A(new_n649), .B(new_n650), .C1(new_n381), .C2(new_n642), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n641), .A2(new_n648), .A3(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n459), .A2(new_n523), .A3(new_n611), .A4(new_n653), .ZN(new_n654));
  XNOR2_X1  g0454(.A(new_n654), .B(KEYINPUT88), .ZN(G372));
  INV_X1    g0455(.A(new_n573), .ZN(new_n656));
  AND3_X1   g0456(.A1(new_n605), .A2(new_n606), .A3(new_n608), .ZN(new_n657));
  NOR3_X1   g0457(.A1(new_n594), .A2(KEYINPUT89), .A3(new_n305), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT89), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n659), .B1(new_n600), .B2(new_n372), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n591), .B1(new_n658), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(G200), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n657), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n661), .A2(new_n402), .ZN(new_n664));
  AOI22_X1  g0464(.A1(new_n606), .A2(new_n586), .B1(new_n355), .B2(new_n602), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n509), .A2(new_n518), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n667), .B1(new_n668), .B2(new_n521), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n628), .A2(new_n644), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(new_n646), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n628), .A2(KEYINPUT21), .A3(new_n644), .ZN(new_n672));
  AND3_X1   g0472(.A1(new_n628), .A2(new_n639), .A3(new_n636), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n639), .B1(new_n628), .B2(new_n636), .ZN(new_n674));
  OAI211_X1 g0474(.A(new_n671), .B(new_n672), .C1(new_n673), .C2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n519), .ZN(new_n676));
  OAI211_X1 g0476(.A(new_n656), .B(new_n669), .C1(new_n675), .C2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT90), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n572), .A2(new_n678), .ZN(new_n679));
  AOI22_X1  g0479(.A1(new_n657), .A2(new_n662), .B1(new_n664), .B2(new_n665), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT26), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n569), .A2(new_n570), .A3(new_n571), .A4(KEYINPUT90), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n679), .A2(new_n680), .A3(new_n681), .A4(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(KEYINPUT26), .B1(new_n572), .B2(new_n610), .ZN(new_n684));
  AND3_X1   g0484(.A1(new_n683), .A2(new_n666), .A3(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n677), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n459), .A2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n400), .ZN(new_n688));
  INV_X1    g0488(.A(new_n404), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n450), .A2(new_n452), .ZN(new_n690));
  OAI211_X1 g0490(.A(new_n431), .B(new_n442), .C1(new_n690), .C2(new_n428), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n454), .A2(new_n445), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n688), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n359), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n316), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(new_n457), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n687), .A2(new_n698), .ZN(G369));
  INV_X1    g0499(.A(KEYINPUT91), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n211), .A2(new_n258), .A3(G13), .ZN(new_n701));
  OR2_X1    g0501(.A1(new_n701), .A2(KEYINPUT27), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(KEYINPUT27), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n702), .A2(G213), .A3(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(G343), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n649), .A2(new_n707), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n700), .B1(new_n675), .B2(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n709), .B1(new_n652), .B2(new_n708), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n675), .A2(new_n700), .A3(new_n708), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n710), .A2(G330), .A3(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n519), .A2(new_n522), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n668), .A2(new_n707), .ZN(new_n715));
  OAI22_X1  g0515(.A1(new_n714), .A2(new_n715), .B1(new_n519), .B2(new_n707), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n713), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n706), .B1(new_n641), .B2(new_n648), .ZN(new_n718));
  AOI22_X1  g0518(.A1(new_n718), .A2(new_n523), .B1(new_n676), .B2(new_n707), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n717), .A2(new_n719), .ZN(G399));
  INV_X1    g0520(.A(new_n208), .ZN(new_n721));
  OR3_X1    g0521(.A1(new_n721), .A2(KEYINPUT92), .A3(G41), .ZN(new_n722));
  OAI21_X1  g0522(.A(KEYINPUT92), .B1(new_n721), .B2(G41), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n552), .A2(new_n577), .A3(new_n614), .ZN(new_n726));
  NOR3_X1   g0526(.A1(new_n725), .A2(new_n258), .A3(new_n726), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n727), .B1(new_n218), .B2(new_n725), .ZN(new_n728));
  XOR2_X1   g0528(.A(new_n728), .B(KEYINPUT28), .Z(new_n729));
  NAND3_X1  g0529(.A1(new_n641), .A2(new_n648), .A3(new_n519), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT95), .ZN(new_n731));
  AND3_X1   g0531(.A1(new_n562), .A2(new_n572), .A3(new_n731), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n731), .B1(new_n562), .B2(new_n572), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n730), .A2(new_n669), .A3(new_n734), .ZN(new_n735));
  AND3_X1   g0535(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n736));
  INV_X1    g0536(.A(new_n610), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n736), .A2(new_n737), .A3(new_n681), .ZN(new_n738));
  AND3_X1   g0538(.A1(new_n664), .A2(new_n665), .A3(KEYINPUT94), .ZN(new_n739));
  AOI21_X1  g0539(.A(KEYINPUT94), .B1(new_n664), .B2(new_n665), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n738), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n679), .A2(new_n680), .A3(new_n682), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n742), .B1(KEYINPUT26), .B2(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n706), .B1(new_n735), .B2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT29), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT93), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n748), .B1(new_n686), .B2(new_n707), .ZN(new_n749));
  AOI211_X1 g0549(.A(KEYINPUT93), .B(new_n706), .C1(new_n677), .C2(new_n685), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n747), .B1(new_n751), .B2(new_n746), .ZN(new_n752));
  OAI22_X1  g0552(.A1(new_n484), .A2(new_n305), .B1(new_n465), .B2(new_n223), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n753), .A2(new_n595), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n545), .A2(new_n636), .A3(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT30), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND4_X1  g0557(.A1(new_n545), .A2(new_n754), .A3(new_n636), .A4(KEYINPUT30), .ZN(new_n758));
  AOI21_X1  g0558(.A(G179), .B1(new_n488), .B2(new_n481), .ZN(new_n759));
  NAND4_X1  g0559(.A1(new_n759), .A2(new_n661), .A3(new_n539), .A4(new_n642), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n757), .A2(new_n758), .A3(new_n760), .ZN(new_n761));
  AND3_X1   g0561(.A1(new_n761), .A2(KEYINPUT31), .A3(new_n706), .ZN(new_n762));
  AOI21_X1  g0562(.A(KEYINPUT31), .B1(new_n761), .B2(new_n706), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND4_X1  g0564(.A1(new_n611), .A2(new_n519), .A3(new_n522), .A4(new_n707), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n764), .B1(new_n765), .B2(new_n652), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(G330), .ZN(new_n767));
  AND2_X1   g0567(.A1(new_n752), .A2(new_n767), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n729), .B1(new_n768), .B2(G1), .ZN(G364));
  AND2_X1   g0569(.A1(new_n211), .A2(G13), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(G45), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(G1), .ZN(new_n772));
  OR3_X1    g0572(.A1(new_n725), .A2(KEYINPUT96), .A3(new_n772), .ZN(new_n773));
  OAI21_X1  g0573(.A(KEYINPUT96), .B1(new_n725), .B2(new_n772), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(G13), .A2(G33), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(G20), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n212), .B1(G20), .B2(new_n402), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g0581(.A(new_n781), .B(KEYINPUT98), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n721), .A2(new_n298), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(G355), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n784), .B1(G116), .B2(new_n208), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n721), .A2(new_n292), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(G45), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n787), .B1(new_n788), .B2(new_n218), .ZN(new_n789));
  OR2_X1    g0589(.A1(new_n789), .A2(KEYINPUT97), .ZN(new_n790));
  AOI22_X1  g0590(.A1(new_n789), .A2(KEYINPUT97), .B1(G45), .B2(new_n244), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n785), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n211), .A2(G190), .ZN(new_n793));
  INV_X1    g0593(.A(G200), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(G179), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  XNOR2_X1  g0596(.A(new_n796), .B(KEYINPUT100), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(new_n222), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n355), .A2(G200), .ZN(new_n800));
  AND3_X1   g0600(.A1(new_n793), .A2(KEYINPUT99), .A3(new_n800), .ZN(new_n801));
  AOI21_X1  g0601(.A(KEYINPUT99), .B1(new_n793), .B2(new_n800), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n803), .A2(new_n204), .ZN(new_n804));
  NOR2_X1   g0604(.A1(G179), .A2(G200), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n339), .B1(new_n381), .B2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n808), .A2(new_n550), .ZN(new_n809));
  AND3_X1   g0609(.A1(new_n339), .A2(G190), .A3(new_n800), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n355), .A2(new_n794), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n339), .A2(G190), .A3(new_n812), .ZN(new_n813));
  OAI22_X1  g0613(.A1(new_n811), .A2(new_n214), .B1(new_n257), .B2(new_n813), .ZN(new_n814));
  NOR4_X1   g0614(.A1(new_n799), .A2(new_n804), .A3(new_n809), .A4(new_n814), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n795), .A2(G20), .A3(G190), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n816), .A2(new_n577), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n793), .A2(new_n812), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  AOI211_X1 g0619(.A(new_n298), .B(new_n817), .C1(new_n819), .C2(G68), .ZN(new_n820));
  INV_X1    g0620(.A(new_n793), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n821), .A2(new_n806), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n822), .A2(G159), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n820), .B1(KEYINPUT32), .B2(new_n823), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n824), .B1(KEYINPUT32), .B2(new_n823), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n298), .B1(new_n816), .B2(new_n632), .ZN(new_n826));
  AOI22_X1  g0626(.A1(new_n822), .A2(G329), .B1(G294), .B2(new_n807), .ZN(new_n827));
  XNOR2_X1  g0627(.A(KEYINPUT33), .B(G317), .ZN(new_n828));
  INV_X1    g0628(.A(new_n813), .ZN(new_n829));
  AOI22_X1  g0629(.A1(new_n819), .A2(new_n828), .B1(G326), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n827), .A2(new_n830), .ZN(new_n831));
  AOI211_X1 g0631(.A(new_n826), .B(new_n831), .C1(G322), .C2(new_n810), .ZN(new_n832));
  INV_X1    g0632(.A(new_n803), .ZN(new_n833));
  AOI22_X1  g0633(.A1(new_n833), .A2(G311), .B1(new_n797), .B2(G283), .ZN(new_n834));
  AOI22_X1  g0634(.A1(new_n815), .A2(new_n825), .B1(new_n832), .B2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n780), .ZN(new_n836));
  OAI221_X1 g0636(.A(new_n776), .B1(new_n782), .B2(new_n792), .C1(new_n835), .C2(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n710), .A2(new_n711), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n837), .B1(new_n838), .B2(new_n779), .ZN(new_n839));
  XNOR2_X1  g0639(.A(new_n839), .B(KEYINPUT101), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n712), .B1(new_n725), .B2(new_n772), .ZN(new_n841));
  INV_X1    g0641(.A(G330), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n841), .B1(new_n842), .B2(new_n838), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n840), .A2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(G396));
  NOR2_X1   g0645(.A1(new_n725), .A2(new_n772), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n401), .A2(new_n706), .ZN(new_n847));
  NAND4_X1  g0647(.A1(new_n384), .A2(new_n404), .A3(new_n707), .A4(new_n847), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n848), .B1(new_n677), .B2(new_n685), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n404), .A2(new_n706), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n384), .A2(new_n847), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n851), .B1(new_n852), .B2(new_n404), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n850), .B1(new_n751), .B2(new_n853), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n846), .B1(new_n854), .B2(new_n767), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n855), .B1(new_n767), .B2(new_n854), .ZN(new_n856));
  INV_X1    g0656(.A(new_n816), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n298), .B1(new_n857), .B2(G50), .ZN(new_n858));
  INV_X1    g0658(.A(new_n822), .ZN(new_n859));
  INV_X1    g0659(.A(G132), .ZN(new_n860));
  OAI221_X1 g0660(.A(new_n858), .B1(new_n808), .B2(new_n214), .C1(new_n859), .C2(new_n860), .ZN(new_n861));
  AOI22_X1  g0661(.A1(G137), .A2(new_n829), .B1(new_n810), .B2(G143), .ZN(new_n862));
  INV_X1    g0662(.A(G150), .ZN(new_n863));
  INV_X1    g0663(.A(G159), .ZN(new_n864));
  OAI221_X1 g0664(.A(new_n862), .B1(new_n863), .B2(new_n818), .C1(new_n803), .C2(new_n864), .ZN(new_n865));
  XOR2_X1   g0665(.A(new_n865), .B(KEYINPUT34), .Z(new_n866));
  AOI211_X1 g0666(.A(new_n861), .B(new_n866), .C1(G68), .C2(new_n797), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n798), .A2(new_n577), .ZN(new_n868));
  AOI211_X1 g0668(.A(new_n292), .B(new_n809), .C1(G107), .C2(new_n857), .ZN(new_n869));
  AOI22_X1  g0669(.A1(new_n822), .A2(G311), .B1(G294), .B2(new_n810), .ZN(new_n870));
  AOI22_X1  g0670(.A1(new_n819), .A2(G283), .B1(G303), .B2(new_n829), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n869), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  AOI211_X1 g0672(.A(new_n868), .B(new_n872), .C1(G116), .C2(new_n833), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n780), .B1(new_n867), .B2(new_n873), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n780), .A2(new_n777), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n775), .B1(new_n204), .B2(new_n875), .ZN(new_n876));
  OAI211_X1 g0676(.A(new_n874), .B(new_n876), .C1(new_n778), .C2(new_n853), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n856), .A2(new_n877), .ZN(G384));
  OR2_X1    g0678(.A1(new_n556), .A2(KEYINPUT35), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n556), .A2(KEYINPUT35), .ZN(new_n880));
  NAND4_X1  g0680(.A1(new_n879), .A2(G116), .A3(new_n213), .A4(new_n880), .ZN(new_n881));
  XOR2_X1   g0681(.A(new_n881), .B(KEYINPUT36), .Z(new_n882));
  NAND4_X1  g0682(.A1(new_n218), .A2(G77), .A3(new_n326), .A4(new_n327), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n215), .A2(G50), .ZN(new_n884));
  XNOR2_X1  g0684(.A(new_n884), .B(KEYINPUT102), .ZN(new_n885));
  AOI211_X1 g0685(.A(new_n258), .B(G13), .C1(new_n883), .C2(new_n885), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n882), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n686), .A2(new_n707), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(KEYINPUT93), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n686), .A2(new_n748), .A3(new_n707), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n889), .A2(new_n746), .A3(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n747), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n697), .B1(new_n893), .B2(new_n459), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT39), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n394), .A2(new_n398), .A3(new_n318), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n344), .A2(new_n356), .ZN(new_n897));
  INV_X1    g0697(.A(new_n704), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n344), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n896), .A2(new_n897), .A3(new_n899), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n900), .A2(KEYINPUT37), .ZN(new_n901));
  AOI21_X1  g0701(.A(KEYINPUT16), .B1(new_n323), .B2(new_n333), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n318), .B1(new_n335), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(KEYINPUT103), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT103), .ZN(new_n905));
  OAI211_X1 g0705(.A(new_n905), .B(new_n318), .C1(new_n335), .C2(new_n902), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n904), .A2(new_n898), .A3(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n904), .A2(new_n356), .A3(new_n906), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n907), .A2(new_n908), .A3(new_n896), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n901), .B1(KEYINPUT37), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n897), .A2(KEYINPUT18), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n344), .A2(new_n345), .A3(new_n356), .ZN(new_n912));
  NAND4_X1  g0712(.A1(new_n911), .A2(new_n912), .A3(new_n393), .A4(new_n399), .ZN(new_n913));
  INV_X1    g0713(.A(new_n907), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(KEYINPUT38), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n910), .A2(new_n916), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n900), .B(KEYINPUT37), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n913), .A2(new_n344), .A3(new_n898), .ZN(new_n919));
  AOI21_X1  g0719(.A(KEYINPUT38), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n895), .B1(new_n917), .B2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT38), .ZN(new_n922));
  INV_X1    g0722(.A(new_n915), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n922), .B1(new_n910), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n909), .A2(KEYINPUT37), .ZN(new_n925));
  INV_X1    g0725(.A(new_n901), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n922), .B1(new_n913), .B2(new_n914), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n924), .A2(KEYINPUT39), .A3(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n454), .A2(new_n445), .A3(new_n707), .ZN(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n921), .A2(new_n930), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n924), .A2(new_n929), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n445), .A2(new_n706), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n693), .A2(new_n691), .A3(new_n935), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n445), .B(new_n706), .C1(new_n444), .C2(new_n454), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  OAI211_X1 g0738(.A(new_n934), .B(new_n938), .C1(new_n851), .C2(new_n849), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n695), .A2(new_n704), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n933), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n894), .B(new_n942), .ZN(new_n943));
  AND3_X1   g0743(.A1(new_n766), .A2(new_n938), .A3(new_n853), .ZN(new_n944));
  AOI21_X1  g0744(.A(KEYINPUT40), .B1(new_n944), .B2(new_n934), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT40), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT37), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n900), .B(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n899), .B1(new_n400), .B2(new_n359), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n922), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n946), .B1(new_n929), .B2(new_n950), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n945), .B1(new_n944), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n459), .A2(new_n766), .ZN(new_n953));
  INV_X1    g0753(.A(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n842), .B1(new_n952), .B2(new_n954), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(new_n952), .B2(new_n954), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n943), .A2(new_n956), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(new_n258), .B2(new_n770), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n943), .A2(new_n956), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n887), .B1(new_n958), .B2(new_n959), .ZN(G367));
  NAND2_X1  g0760(.A1(new_n606), .A2(new_n608), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(new_n706), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n680), .A2(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n963), .B1(new_n666), .B2(new_n962), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n964), .A2(KEYINPUT43), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n965), .B(KEYINPUT104), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n569), .A2(new_n706), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n734), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n736), .A2(new_n706), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n970), .A2(new_n523), .A3(new_n718), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(KEYINPUT42), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n572), .B1(new_n968), .B2(new_n519), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(new_n707), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n971), .A2(KEYINPUT42), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n966), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  OR2_X1    g0777(.A1(new_n964), .A2(KEYINPUT43), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n977), .B(new_n978), .ZN(new_n979));
  AND2_X1   g0779(.A1(new_n713), .A2(new_n716), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(new_n970), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n979), .B(new_n981), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n724), .B(KEYINPUT41), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n718), .A2(new_n523), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n984), .B1(new_n716), .B2(new_n718), .ZN(new_n985));
  INV_X1    g0785(.A(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n712), .A2(new_n986), .ZN(new_n987));
  NAND4_X1  g0787(.A1(new_n985), .A2(G330), .A3(new_n710), .A4(new_n711), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND4_X1  g0789(.A1(new_n989), .A2(new_n891), .A3(new_n767), .A4(new_n892), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(KEYINPUT107), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT107), .ZN(new_n992));
  NAND4_X1  g0792(.A1(new_n752), .A2(new_n992), .A3(new_n767), .A4(new_n989), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n719), .A2(new_n970), .ZN(new_n994));
  XNOR2_X1  g0794(.A(KEYINPUT105), .B(KEYINPUT45), .ZN(new_n995));
  INV_X1    g0795(.A(new_n995), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n994), .B(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT106), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT44), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  OAI211_X1 g0800(.A(new_n968), .B(new_n969), .C1(KEYINPUT106), .C2(KEYINPUT44), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1000), .B1(new_n1001), .B2(new_n719), .ZN(new_n1002));
  OR3_X1    g0802(.A1(new_n1001), .A2(new_n719), .A3(new_n1000), .ZN(new_n1003));
  NAND4_X1  g0803(.A1(new_n997), .A2(new_n717), .A3(new_n1002), .A4(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(new_n1002), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n994), .B(new_n995), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n980), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  NAND4_X1  g0807(.A1(new_n991), .A2(new_n993), .A3(new_n1004), .A4(new_n1007), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n983), .B1(new_n1008), .B2(new_n768), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n982), .B1(new_n1009), .B2(new_n772), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n782), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n1011), .B1(new_n208), .B2(new_n360), .C1(new_n237), .C2(new_n787), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n775), .B1(KEYINPUT108), .B2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(KEYINPUT108), .B2(new_n1012), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(G143), .A2(new_n829), .B1(new_n810), .B2(G150), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1015), .B1(new_n215), .B2(new_n808), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(G137), .A2(new_n822), .B1(new_n819), .B2(G159), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n298), .B1(new_n857), .B2(G58), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n1017), .B(new_n1018), .C1(new_n204), .C2(new_n796), .ZN(new_n1019));
  AOI211_X1 g0819(.A(new_n1016), .B(new_n1019), .C1(G50), .C2(new_n833), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n857), .A2(G116), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT46), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(G311), .A2(new_n829), .B1(new_n810), .B2(G303), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1022), .A2(new_n298), .A3(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n822), .A2(G317), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1025), .B1(new_n550), .B2(new_n796), .ZN(new_n1026));
  INV_X1    g0826(.A(G294), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n818), .A2(new_n1027), .B1(new_n808), .B2(new_n222), .ZN(new_n1028));
  NOR3_X1   g0828(.A1(new_n1024), .A2(new_n1026), .A3(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n833), .A2(G283), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1020), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  XOR2_X1   g0831(.A(new_n1031), .B(KEYINPUT47), .Z(new_n1032));
  AOI21_X1  g0832(.A(new_n1014), .B1(new_n1032), .B2(new_n780), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n779), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1033), .B1(new_n1034), .B2(new_n964), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1010), .A2(new_n1035), .ZN(G387));
  AOI22_X1  g0836(.A1(new_n783), .A2(new_n726), .B1(new_n222), .B2(new_n721), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n249), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1038), .A2(new_n257), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1039), .B(KEYINPUT50), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n788), .B1(new_n215), .B2(new_n204), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1041), .B1(new_n726), .B2(KEYINPUT109), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(KEYINPUT109), .B2(new_n726), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n786), .B1(new_n1040), .B2(new_n1043), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n1044), .A2(KEYINPUT110), .B1(new_n234), .B2(new_n788), .ZN(new_n1045));
  AND2_X1   g0845(.A1(new_n1044), .A2(KEYINPUT110), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1037), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n775), .B1(new_n1047), .B2(new_n1011), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1048), .B1(new_n716), .B2(new_n1034), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n807), .A2(new_n585), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n1050), .B1(new_n864), .B2(new_n813), .C1(new_n818), .C2(new_n249), .ZN(new_n1051));
  AOI211_X1 g0851(.A(new_n298), .B(new_n1051), .C1(G50), .C2(new_n810), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n822), .A2(G150), .B1(G77), .B2(new_n857), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(KEYINPUT111), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n797), .A2(G97), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n833), .A2(G68), .ZN(new_n1056));
  NAND4_X1  g0856(.A1(new_n1052), .A2(new_n1054), .A3(new_n1055), .A4(new_n1056), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n807), .A2(G283), .B1(new_n857), .B2(G294), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n819), .A2(G311), .B1(G317), .B2(new_n810), .ZN(new_n1059));
  INV_X1    g0859(.A(G322), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1059), .B1(new_n1060), .B2(new_n813), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1061), .B1(G303), .B2(new_n833), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n1062), .ZN(new_n1063));
  INV_X1    g0863(.A(KEYINPUT48), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1058), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  AND2_X1   g0865(.A1(new_n1065), .A2(KEYINPUT112), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n1065), .A2(KEYINPUT112), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n1066), .A2(new_n1067), .B1(KEYINPUT48), .B2(new_n1062), .ZN(new_n1068));
  OR2_X1    g0868(.A1(new_n1068), .A2(KEYINPUT113), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1068), .A2(KEYINPUT113), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1069), .A2(KEYINPUT49), .A3(new_n1070), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n292), .B1(new_n822), .B2(G326), .ZN(new_n1072));
  OAI211_X1 g0872(.A(new_n1071), .B(new_n1072), .C1(new_n614), .C2(new_n796), .ZN(new_n1073));
  AOI21_X1  g0873(.A(KEYINPUT49), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1057), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1049), .B1(new_n1075), .B2(new_n780), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1076), .B1(new_n772), .B2(new_n989), .ZN(new_n1077));
  AND2_X1   g0877(.A1(new_n990), .A2(new_n725), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1078), .B1(new_n768), .B2(new_n989), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1077), .A2(new_n1079), .ZN(G393));
  NAND3_X1  g0880(.A1(new_n1007), .A2(new_n1004), .A3(new_n772), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT114), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n241), .A2(new_n786), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n1011), .B(new_n1083), .C1(new_n550), .C2(new_n208), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n775), .B1(new_n1082), .B2(new_n1084), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1085), .B1(new_n1082), .B2(new_n1084), .ZN(new_n1086));
  INV_X1    g0886(.A(G283), .ZN(new_n1087));
  OAI221_X1 g0887(.A(new_n298), .B1(new_n1087), .B2(new_n816), .C1(new_n818), .C2(new_n632), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n859), .A2(new_n1060), .B1(new_n808), .B2(new_n614), .ZN(new_n1089));
  NOR3_X1   g0889(.A1(new_n799), .A2(new_n1088), .A3(new_n1089), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1090), .B1(new_n1027), .B2(new_n803), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(G317), .A2(new_n829), .B1(new_n810), .B2(G311), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(new_n1092), .B(KEYINPUT52), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n868), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n833), .A2(new_n1038), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n808), .A2(new_n204), .ZN(new_n1096));
  AOI211_X1 g0896(.A(new_n298), .B(new_n1096), .C1(G68), .C2(new_n857), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(G143), .A2(new_n822), .B1(new_n819), .B2(G50), .ZN(new_n1098));
  NAND4_X1  g0898(.A1(new_n1094), .A2(new_n1095), .A3(new_n1097), .A4(new_n1098), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(G150), .A2(new_n829), .B1(new_n810), .B2(G159), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(new_n1100), .B(KEYINPUT51), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n1091), .A2(new_n1093), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1086), .B1(new_n1102), .B2(new_n780), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1103), .B1(new_n970), .B2(new_n1034), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1081), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1007), .A2(new_n1004), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1106), .A2(new_n990), .ZN(new_n1107));
  INV_X1    g0907(.A(KEYINPUT115), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(new_n1107), .B(new_n1108), .ZN(new_n1109));
  AND2_X1   g0909(.A1(new_n1008), .A2(new_n725), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1105), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1111), .ZN(G390));
  AOI21_X1  g0912(.A(new_n775), .B1(new_n249), .B2(new_n875), .ZN(new_n1113));
  INV_X1    g0913(.A(G137), .ZN(new_n1114));
  OAI22_X1  g0914(.A1(new_n818), .A2(new_n1114), .B1(new_n808), .B2(new_n864), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n816), .A2(new_n863), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(new_n1116), .B(KEYINPUT53), .ZN(new_n1117));
  INV_X1    g0917(.A(G128), .ZN(new_n1118));
  OAI221_X1 g0918(.A(new_n1117), .B1(new_n1118), .B2(new_n813), .C1(new_n860), .C2(new_n811), .ZN(new_n1119));
  XOR2_X1   g0919(.A(KEYINPUT54), .B(G143), .Z(new_n1120));
  AOI211_X1 g0920(.A(new_n1115), .B(new_n1119), .C1(new_n833), .C2(new_n1120), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n292), .B1(new_n796), .B2(new_n257), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1122), .B1(G125), .B2(new_n822), .ZN(new_n1123));
  XOR2_X1   g0923(.A(new_n1123), .B(KEYINPUT117), .Z(new_n1124));
  AOI22_X1  g0924(.A1(new_n819), .A2(G107), .B1(G283), .B2(new_n829), .ZN(new_n1125));
  OAI221_X1 g0925(.A(new_n1125), .B1(new_n614), .B2(new_n811), .C1(new_n1027), .C2(new_n859), .ZN(new_n1126));
  NOR4_X1   g0926(.A1(new_n1126), .A2(new_n292), .A3(new_n817), .A4(new_n1096), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(new_n833), .A2(G97), .B1(new_n797), .B2(G68), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n1121), .A2(new_n1124), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1113), .B1(new_n1129), .B2(new_n836), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n921), .A2(new_n930), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1130), .B1(new_n1131), .B2(new_n777), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n932), .B1(new_n929), .B2(new_n950), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n735), .A2(new_n744), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1136), .A2(new_n707), .A3(new_n853), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n851), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1135), .B1(new_n1139), .B2(new_n938), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n938), .B1(new_n849), .B2(new_n851), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n1141), .A2(new_n931), .B1(new_n921), .B2(new_n930), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n766), .A2(new_n938), .A3(G330), .A4(new_n853), .ZN(new_n1143));
  INV_X1    g0943(.A(KEYINPUT116), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1145), .ZN(new_n1146));
  NOR3_X1   g0946(.A1(new_n1140), .A2(new_n1142), .A3(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1141), .A2(new_n931), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1148), .A2(new_n1131), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n851), .B1(new_n745), .B2(new_n853), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n938), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1134), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1145), .B1(new_n1149), .B2(new_n1152), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n1147), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n772), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1133), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1146), .B1(new_n1140), .B2(new_n1142), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1149), .A2(new_n1152), .A3(new_n1145), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  OR2_X1    g0959(.A1(new_n767), .A2(new_n458), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n853), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1151), .B1(new_n767), .B2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1162), .A2(new_n1143), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n850), .A2(new_n1138), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1162), .A2(new_n1150), .A3(new_n1143), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  NAND4_X1  g0967(.A1(new_n1159), .A2(new_n894), .A3(new_n1160), .A4(new_n1167), .ZN(new_n1168));
  NOR3_X1   g0968(.A1(new_n749), .A2(new_n750), .A3(KEYINPUT29), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n459), .B1(new_n1169), .B2(new_n747), .ZN(new_n1170));
  NAND4_X1  g0970(.A1(new_n1167), .A2(new_n698), .A3(new_n1170), .A4(new_n1160), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n724), .B1(new_n1154), .B2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1156), .B1(new_n1168), .B2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(G378));
  OAI211_X1 g0974(.A(new_n698), .B(new_n1160), .C1(new_n752), .C2(new_n458), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1175), .A2(KEYINPUT120), .ZN(new_n1176));
  INV_X1    g0976(.A(KEYINPUT120), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n894), .A2(new_n1177), .A3(new_n1160), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n1176), .B(new_n1178), .C1(new_n1154), .C2(new_n1171), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n842), .B1(new_n944), .B2(new_n951), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n927), .A2(new_n915), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(new_n1182), .A2(new_n922), .B1(new_n927), .B2(new_n928), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n766), .A2(new_n938), .A3(new_n853), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n946), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n314), .A2(new_n315), .A3(new_n457), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n270), .A2(new_n898), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1186), .A2(new_n1188), .ZN(new_n1189));
  NAND4_X1  g0989(.A1(new_n314), .A2(new_n315), .A3(new_n457), .A4(new_n1187), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1191));
  AND3_X1   g0991(.A1(new_n1189), .A2(new_n1190), .A3(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1191), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  AND3_X1   g0994(.A1(new_n1181), .A2(new_n1185), .A3(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1194), .B1(new_n1181), .B2(new_n1185), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n942), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(KEYINPUT121), .ZN(new_n1198));
  OAI21_X1  g0998(.A(KEYINPUT40), .B1(new_n917), .B2(new_n920), .ZN(new_n1199));
  OAI21_X1  g0999(.A(G330), .B1(new_n1199), .B2(new_n1184), .ZN(new_n1200));
  OAI22_X1  g1000(.A1(new_n1200), .A2(new_n945), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1181), .A2(new_n1185), .A3(new_n1194), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1201), .A2(new_n941), .A3(new_n1202), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1197), .A2(new_n1198), .A3(new_n1203), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n942), .B(KEYINPUT121), .C1(new_n1195), .C2(new_n1196), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1204), .A2(KEYINPUT57), .A3(new_n1205), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n725), .B1(new_n1180), .B2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1197), .A2(new_n1203), .ZN(new_n1208));
  AOI21_X1  g1008(.A(KEYINPUT57), .B1(new_n1179), .B2(new_n1208), .ZN(new_n1209));
  OR2_X1    g1009(.A1(new_n1207), .A2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1194), .A2(new_n777), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n796), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1212), .A2(G58), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n298), .A2(new_n462), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1214), .B1(new_n857), .B2(G77), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n1213), .B(new_n1215), .C1(new_n859), .C2(new_n1087), .ZN(new_n1216));
  XNOR2_X1  g1016(.A(new_n1216), .B(KEYINPUT118), .ZN(new_n1217));
  OAI22_X1  g1017(.A1(new_n808), .A2(new_n215), .B1(new_n813), .B2(new_n614), .ZN(new_n1218));
  XNOR2_X1  g1018(.A(new_n1218), .B(KEYINPUT119), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n819), .A2(G97), .B1(G107), .B2(new_n810), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1219), .B(new_n1220), .C1(new_n360), .C2(new_n803), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n1217), .A2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1222), .A2(KEYINPUT58), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n1214), .B(new_n257), .C1(G33), .C2(G41), .ZN(new_n1224));
  AND2_X1   g1024(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(new_n810), .A2(G128), .B1(new_n807), .B2(G150), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1226), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1227), .B1(G132), .B2(new_n819), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(new_n829), .A2(G125), .B1(new_n857), .B2(new_n1120), .ZN(new_n1229));
  OAI211_X1 g1029(.A(new_n1228), .B(new_n1229), .C1(new_n1114), .C2(new_n803), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1230), .A2(KEYINPUT59), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1230), .A2(KEYINPUT59), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1212), .A2(G159), .ZN(new_n1233));
  AOI211_X1 g1033(.A(G33), .B(G41), .C1(new_n822), .C2(G124), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1232), .A2(new_n1233), .A3(new_n1234), .ZN(new_n1235));
  OAI221_X1 g1035(.A(new_n1225), .B1(KEYINPUT58), .B2(new_n1222), .C1(new_n1231), .C2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(new_n780), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n875), .A2(new_n257), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1211), .A2(new_n846), .A3(new_n1237), .A4(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1240), .B1(new_n1208), .B2(new_n772), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1210), .A2(new_n1241), .ZN(G375));
  AND2_X1   g1042(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1175), .A2(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n983), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1244), .A2(new_n1245), .A3(new_n1171), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1151), .A2(new_n777), .ZN(new_n1247));
  NOR3_X1   g1047(.A1(new_n780), .A2(G68), .A3(new_n777), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n811), .A2(new_n1114), .ZN(new_n1249));
  OAI211_X1 g1049(.A(new_n1213), .B(new_n292), .C1(new_n864), .C2(new_n816), .ZN(new_n1250));
  AOI211_X1 g1050(.A(new_n1249), .B(new_n1250), .C1(new_n819), .C2(new_n1120), .ZN(new_n1251));
  OAI22_X1  g1051(.A1(new_n859), .A2(new_n1118), .B1(new_n860), .B2(new_n813), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1252), .B1(G50), .B2(new_n807), .ZN(new_n1253));
  OAI211_X1 g1053(.A(new_n1251), .B(new_n1253), .C1(new_n863), .C2(new_n803), .ZN(new_n1254));
  OAI221_X1 g1054(.A(new_n298), .B1(new_n550), .B2(new_n816), .C1(new_n859), .C2(new_n632), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1255), .B1(G294), .B2(new_n829), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1050), .B1(new_n811), .B2(new_n1087), .ZN(new_n1257));
  XNOR2_X1  g1057(.A(new_n1257), .B(KEYINPUT123), .ZN(new_n1258));
  OAI211_X1 g1058(.A(new_n1256), .B(new_n1258), .C1(new_n204), .C2(new_n798), .ZN(new_n1259));
  OAI22_X1  g1059(.A1(new_n803), .A2(new_n222), .B1(new_n614), .B2(new_n818), .ZN(new_n1260));
  XNOR2_X1  g1060(.A(new_n1260), .B(KEYINPUT122), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1254), .B1(new_n1259), .B2(new_n1261), .ZN(new_n1262));
  AOI211_X1 g1062(.A(new_n775), .B(new_n1248), .C1(new_n1262), .C2(new_n780), .ZN(new_n1263));
  AOI22_X1  g1063(.A1(new_n1167), .A2(new_n772), .B1(new_n1247), .B2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1246), .A2(new_n1264), .ZN(G381));
  INV_X1    g1065(.A(G387), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1077), .A2(new_n844), .A3(new_n1079), .ZN(new_n1267));
  NOR3_X1   g1067(.A1(new_n1267), .A2(G384), .A3(G381), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1266), .A2(new_n1111), .A3(new_n1173), .A4(new_n1268), .ZN(new_n1269));
  OR2_X1    g1069(.A1(new_n1269), .A2(G375), .ZN(G407));
  NAND2_X1  g1070(.A1(new_n705), .A2(G213), .ZN(new_n1271));
  OR3_X1    g1071(.A1(G375), .A2(G378), .A3(new_n1271), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1272), .A2(G407), .A3(G213), .ZN(G409));
  NAND2_X1  g1073(.A1(G387), .A2(new_n1111), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(KEYINPUT127), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(G393), .A2(G396), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(new_n1267), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1275), .A2(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1266), .A2(G390), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1279), .A2(new_n1274), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1278), .A2(new_n1280), .ZN(new_n1281));
  NAND4_X1  g1081(.A1(new_n1275), .A2(new_n1277), .A3(new_n1279), .A4(new_n1274), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1171), .A2(KEYINPUT60), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1285), .A2(new_n1244), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1175), .A2(KEYINPUT60), .A3(new_n1243), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1286), .A2(new_n725), .A3(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1288), .A2(new_n1264), .ZN(new_n1289));
  INV_X1    g1089(.A(G384), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1288), .A2(G384), .A3(new_n1264), .ZN(new_n1292));
  AND2_X1   g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT125), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1204), .A2(new_n772), .A3(new_n1205), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1295), .A2(KEYINPUT124), .A3(new_n1239), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1179), .A2(new_n1245), .A3(new_n1208), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  AOI21_X1  g1098(.A(KEYINPUT124), .B1(new_n1295), .B2(new_n1239), .ZN(new_n1299));
  OAI211_X1 g1099(.A(new_n1294), .B(new_n1173), .C1(new_n1298), .C2(new_n1299), .ZN(new_n1300));
  OAI211_X1 g1100(.A(G378), .B(new_n1241), .C1(new_n1207), .C2(new_n1209), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1295), .A2(new_n1239), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT124), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1305), .A2(new_n1297), .A3(new_n1296), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1294), .B1(new_n1306), .B2(new_n1173), .ZN(new_n1307));
  OAI211_X1 g1107(.A(new_n1271), .B(new_n1293), .C1(new_n1302), .C2(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1308), .A2(KEYINPUT126), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1173), .B1(new_n1298), .B2(new_n1299), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1310), .A2(KEYINPUT125), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1311), .A2(new_n1300), .A3(new_n1301), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT126), .ZN(new_n1313));
  NAND4_X1  g1113(.A1(new_n1312), .A2(new_n1313), .A3(new_n1271), .A4(new_n1293), .ZN(new_n1314));
  AOI21_X1  g1114(.A(KEYINPUT62), .B1(new_n1309), .B2(new_n1314), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1271), .B1(new_n1302), .B2(new_n1307), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n705), .A2(G213), .A3(G2897), .ZN(new_n1317));
  AND3_X1   g1117(.A1(new_n1291), .A2(new_n1292), .A3(new_n1317), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1317), .B1(new_n1291), .B2(new_n1292), .ZN(new_n1319));
  NOR2_X1   g1119(.A1(new_n1318), .A2(new_n1319), .ZN(new_n1320));
  AOI21_X1  g1120(.A(KEYINPUT61), .B1(new_n1316), .B2(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1308), .A2(KEYINPUT62), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1321), .A2(new_n1322), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1284), .B1(new_n1315), .B2(new_n1323), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT63), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1309), .A2(new_n1325), .A3(new_n1314), .ZN(new_n1326));
  OR2_X1    g1126(.A1(new_n1308), .A2(new_n1325), .ZN(new_n1327));
  NAND4_X1  g1127(.A1(new_n1326), .A2(new_n1283), .A3(new_n1321), .A4(new_n1327), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1324), .A2(new_n1328), .ZN(G405));
  AOI21_X1  g1129(.A(G378), .B1(new_n1210), .B2(new_n1241), .ZN(new_n1330));
  INV_X1    g1130(.A(new_n1301), .ZN(new_n1331));
  NOR2_X1   g1131(.A1(new_n1330), .A2(new_n1331), .ZN(new_n1332));
  NOR2_X1   g1132(.A1(new_n1278), .A2(new_n1280), .ZN(new_n1333));
  AOI22_X1  g1133(.A1(new_n1275), .A2(new_n1277), .B1(new_n1279), .B2(new_n1274), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n1332), .B1(new_n1333), .B2(new_n1334), .ZN(new_n1335));
  OAI211_X1 g1135(.A(new_n1281), .B(new_n1282), .C1(new_n1331), .C2(new_n1330), .ZN(new_n1336));
  AND3_X1   g1136(.A1(new_n1335), .A2(new_n1336), .A3(new_n1293), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n1293), .B1(new_n1335), .B2(new_n1336), .ZN(new_n1338));
  NOR2_X1   g1138(.A1(new_n1337), .A2(new_n1338), .ZN(G402));
endmodule


