

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596;

  XNOR2_X1 U328 ( .A(n435), .B(n434), .ZN(n439) );
  XNOR2_X1 U329 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U330 ( .A(n442), .B(n441), .ZN(n443) );
  INV_X1 U331 ( .A(n440), .ZN(n441) );
  XOR2_X1 U332 ( .A(n422), .B(n421), .Z(n574) );
  XOR2_X1 U333 ( .A(n346), .B(n345), .Z(n538) );
  XOR2_X1 U334 ( .A(n339), .B(n338), .Z(n296) );
  XOR2_X1 U335 ( .A(KEYINPUT94), .B(n436), .Z(n297) );
  XNOR2_X1 U336 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U337 ( .A(G99GAT), .B(G85GAT), .ZN(n440) );
  XNOR2_X1 U338 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U339 ( .A(n340), .B(n296), .ZN(n341) );
  XOR2_X1 U340 ( .A(KEYINPUT36), .B(n574), .Z(n592) );
  XNOR2_X1 U341 ( .A(n342), .B(n341), .ZN(n343) );
  NOR2_X1 U342 ( .A1(n536), .A2(n481), .ZN(n580) );
  NOR2_X1 U343 ( .A1(n534), .A2(n505), .ZN(n462) );
  XNOR2_X1 U344 ( .A(n444), .B(n443), .ZN(n585) );
  XNOR2_X1 U345 ( .A(n462), .B(n461), .ZN(n520) );
  XNOR2_X1 U346 ( .A(G169GAT), .B(KEYINPUT123), .ZN(n486) );
  XNOR2_X1 U347 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U348 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U349 ( .A(n487), .B(n486), .ZN(G1348GAT) );
  XNOR2_X1 U350 ( .A(n466), .B(n465), .ZN(G1330GAT) );
  XOR2_X1 U351 ( .A(G22GAT), .B(G155GAT), .Z(n387) );
  XOR2_X1 U352 ( .A(G78GAT), .B(G148GAT), .Z(n299) );
  XNOR2_X1 U353 ( .A(G106GAT), .B(KEYINPUT71), .ZN(n298) );
  XNOR2_X1 U354 ( .A(n299), .B(n298), .ZN(n425) );
  XOR2_X1 U355 ( .A(n387), .B(n425), .Z(n301) );
  NAND2_X1 U356 ( .A1(G228GAT), .A2(G233GAT), .ZN(n300) );
  XNOR2_X1 U357 ( .A(n301), .B(n300), .ZN(n305) );
  XOR2_X1 U358 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n303) );
  XNOR2_X1 U359 ( .A(KEYINPUT88), .B(KEYINPUT22), .ZN(n302) );
  XNOR2_X1 U360 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U361 ( .A(n305), .B(n304), .Z(n310) );
  XNOR2_X1 U362 ( .A(G50GAT), .B(KEYINPUT73), .ZN(n306) );
  XNOR2_X1 U363 ( .A(n306), .B(G162GAT), .ZN(n420) );
  XOR2_X1 U364 ( .A(KEYINPUT2), .B(KEYINPUT90), .Z(n308) );
  XNOR2_X1 U365 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n307) );
  XNOR2_X1 U366 ( .A(n308), .B(n307), .ZN(n368) );
  XNOR2_X1 U367 ( .A(n420), .B(n368), .ZN(n309) );
  XNOR2_X1 U368 ( .A(n310), .B(n309), .ZN(n315) );
  XOR2_X1 U369 ( .A(KEYINPUT21), .B(G204GAT), .Z(n312) );
  XNOR2_X1 U370 ( .A(G197GAT), .B(G211GAT), .ZN(n311) );
  XNOR2_X1 U371 ( .A(n312), .B(n311), .ZN(n314) );
  XOR2_X1 U372 ( .A(G218GAT), .B(KEYINPUT89), .Z(n313) );
  XNOR2_X1 U373 ( .A(n314), .B(n313), .ZN(n345) );
  XNOR2_X1 U374 ( .A(n315), .B(n345), .ZN(n482) );
  XOR2_X1 U375 ( .A(KEYINPUT17), .B(KEYINPUT85), .Z(n317) );
  XNOR2_X1 U376 ( .A(KEYINPUT19), .B(G183GAT), .ZN(n316) );
  XNOR2_X1 U377 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U378 ( .A(KEYINPUT18), .B(n318), .Z(n335) );
  XOR2_X1 U379 ( .A(G176GAT), .B(KEYINPUT86), .Z(n320) );
  XNOR2_X1 U380 ( .A(G113GAT), .B(KEYINPUT87), .ZN(n319) );
  XNOR2_X1 U381 ( .A(n320), .B(n319), .ZN(n333) );
  XOR2_X1 U382 ( .A(G190GAT), .B(G99GAT), .Z(n322) );
  XNOR2_X1 U383 ( .A(G43GAT), .B(G134GAT), .ZN(n321) );
  XNOR2_X1 U384 ( .A(n322), .B(n321), .ZN(n326) );
  XOR2_X1 U385 ( .A(KEYINPUT84), .B(KEYINPUT20), .Z(n324) );
  XNOR2_X1 U386 ( .A(G169GAT), .B(KEYINPUT83), .ZN(n323) );
  XNOR2_X1 U387 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U388 ( .A(n326), .B(n325), .Z(n331) );
  XOR2_X1 U389 ( .A(KEYINPUT0), .B(KEYINPUT82), .Z(n361) );
  XOR2_X1 U390 ( .A(G120GAT), .B(G71GAT), .Z(n442) );
  XOR2_X1 U391 ( .A(G15GAT), .B(G127GAT), .Z(n388) );
  XOR2_X1 U392 ( .A(n442), .B(n388), .Z(n328) );
  NAND2_X1 U393 ( .A1(G227GAT), .A2(G233GAT), .ZN(n327) );
  XNOR2_X1 U394 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U395 ( .A(n361), .B(n329), .ZN(n330) );
  XNOR2_X1 U396 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U397 ( .A(n333), .B(n332), .Z(n334) );
  XOR2_X1 U398 ( .A(n335), .B(n334), .Z(n541) );
  INV_X1 U399 ( .A(n335), .ZN(n344) );
  XNOR2_X1 U400 ( .A(G176GAT), .B(G92GAT), .ZN(n336) );
  XNOR2_X1 U401 ( .A(n336), .B(G64GAT), .ZN(n436) );
  NAND2_X1 U402 ( .A1(G226GAT), .A2(G233GAT), .ZN(n337) );
  XNOR2_X1 U403 ( .A(n297), .B(n337), .ZN(n342) );
  XOR2_X1 U404 ( .A(G169GAT), .B(G8GAT), .Z(n451) );
  XOR2_X1 U405 ( .A(G36GAT), .B(G190GAT), .Z(n407) );
  XNOR2_X1 U406 ( .A(n451), .B(n407), .ZN(n340) );
  XOR2_X1 U407 ( .A(KEYINPUT93), .B(KEYINPUT95), .Z(n339) );
  XNOR2_X1 U408 ( .A(KEYINPUT78), .B(KEYINPUT96), .ZN(n338) );
  XOR2_X1 U409 ( .A(n344), .B(n343), .Z(n346) );
  NAND2_X1 U410 ( .A1(n541), .A2(n538), .ZN(n347) );
  NAND2_X1 U411 ( .A1(n482), .A2(n347), .ZN(n348) );
  XOR2_X1 U412 ( .A(KEYINPUT25), .B(n348), .Z(n351) );
  XNOR2_X1 U413 ( .A(KEYINPUT27), .B(n538), .ZN(n376) );
  NOR2_X1 U414 ( .A1(n482), .A2(n541), .ZN(n349) );
  XNOR2_X1 U415 ( .A(n349), .B(KEYINPUT26), .ZN(n579) );
  NAND2_X1 U416 ( .A1(n376), .A2(n579), .ZN(n350) );
  NAND2_X1 U417 ( .A1(n351), .A2(n350), .ZN(n352) );
  XOR2_X1 U418 ( .A(KEYINPUT97), .B(n352), .Z(n373) );
  XOR2_X1 U419 ( .A(KEYINPUT6), .B(KEYINPUT92), .Z(n354) );
  XNOR2_X1 U420 ( .A(KEYINPUT91), .B(KEYINPUT5), .ZN(n353) );
  XNOR2_X1 U421 ( .A(n354), .B(n353), .ZN(n372) );
  XOR2_X1 U422 ( .A(G85GAT), .B(G162GAT), .Z(n356) );
  XNOR2_X1 U423 ( .A(G29GAT), .B(G127GAT), .ZN(n355) );
  XNOR2_X1 U424 ( .A(n356), .B(n355), .ZN(n360) );
  XOR2_X1 U425 ( .A(G57GAT), .B(G148GAT), .Z(n358) );
  XNOR2_X1 U426 ( .A(G120GAT), .B(G155GAT), .ZN(n357) );
  XNOR2_X1 U427 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U428 ( .A(n360), .B(n359), .Z(n366) );
  XOR2_X1 U429 ( .A(G113GAT), .B(G1GAT), .Z(n455) );
  XOR2_X1 U430 ( .A(G134GAT), .B(KEYINPUT77), .Z(n409) );
  XOR2_X1 U431 ( .A(n409), .B(n361), .Z(n363) );
  NAND2_X1 U432 ( .A1(G225GAT), .A2(G233GAT), .ZN(n362) );
  XNOR2_X1 U433 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U434 ( .A(n455), .B(n364), .ZN(n365) );
  XNOR2_X1 U435 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U436 ( .A(n367), .B(KEYINPUT1), .Z(n370) );
  XNOR2_X1 U437 ( .A(n368), .B(KEYINPUT4), .ZN(n369) );
  XNOR2_X1 U438 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U439 ( .A(n372), .B(n371), .Z(n375) );
  NAND2_X1 U440 ( .A1(n373), .A2(n375), .ZN(n380) );
  XNOR2_X1 U441 ( .A(n482), .B(KEYINPUT28), .ZN(n374) );
  XNOR2_X1 U442 ( .A(n374), .B(KEYINPUT67), .ZN(n544) );
  INV_X1 U443 ( .A(n375), .ZN(n536) );
  NAND2_X1 U444 ( .A1(n536), .A2(n376), .ZN(n488) );
  NOR2_X1 U445 ( .A1(n544), .A2(n488), .ZN(n378) );
  INV_X1 U446 ( .A(n541), .ZN(n377) );
  NAND2_X1 U447 ( .A1(n378), .A2(n377), .ZN(n379) );
  NAND2_X1 U448 ( .A1(n380), .A2(n379), .ZN(n502) );
  XOR2_X1 U449 ( .A(KEYINPUT78), .B(G64GAT), .Z(n382) );
  XNOR2_X1 U450 ( .A(G1GAT), .B(G8GAT), .ZN(n381) );
  XNOR2_X1 U451 ( .A(n382), .B(n381), .ZN(n386) );
  XOR2_X1 U452 ( .A(KEYINPUT15), .B(KEYINPUT80), .Z(n384) );
  XNOR2_X1 U453 ( .A(KEYINPUT79), .B(KEYINPUT14), .ZN(n383) );
  XNOR2_X1 U454 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U455 ( .A(n386), .B(n385), .ZN(n399) );
  XOR2_X1 U456 ( .A(G78GAT), .B(n387), .Z(n390) );
  XNOR2_X1 U457 ( .A(n388), .B(G211GAT), .ZN(n389) );
  XNOR2_X1 U458 ( .A(n390), .B(n389), .ZN(n395) );
  XNOR2_X1 U459 ( .A(G57GAT), .B(KEYINPUT70), .ZN(n391) );
  XNOR2_X1 U460 ( .A(n391), .B(KEYINPUT13), .ZN(n437) );
  XOR2_X1 U461 ( .A(KEYINPUT12), .B(n437), .Z(n393) );
  NAND2_X1 U462 ( .A1(G231GAT), .A2(G233GAT), .ZN(n392) );
  XNOR2_X1 U463 ( .A(n393), .B(n392), .ZN(n394) );
  XOR2_X1 U464 ( .A(n395), .B(n394), .Z(n397) );
  XNOR2_X1 U465 ( .A(G183GAT), .B(G71GAT), .ZN(n396) );
  XNOR2_X1 U466 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U467 ( .A(n399), .B(n398), .Z(n555) );
  INV_X1 U468 ( .A(n555), .ZN(n588) );
  NAND2_X1 U469 ( .A1(n502), .A2(n588), .ZN(n400) );
  XNOR2_X1 U470 ( .A(n400), .B(KEYINPUT103), .ZN(n423) );
  XOR2_X1 U471 ( .A(KEYINPUT9), .B(KEYINPUT75), .Z(n402) );
  XNOR2_X1 U472 ( .A(G218GAT), .B(KEYINPUT65), .ZN(n401) );
  XNOR2_X1 U473 ( .A(n402), .B(n401), .ZN(n406) );
  XOR2_X1 U474 ( .A(KEYINPUT64), .B(KEYINPUT11), .Z(n404) );
  XNOR2_X1 U475 ( .A(G106GAT), .B(G92GAT), .ZN(n403) );
  XNOR2_X1 U476 ( .A(n404), .B(n403), .ZN(n405) );
  XOR2_X1 U477 ( .A(n406), .B(n405), .Z(n413) );
  XNOR2_X1 U478 ( .A(n440), .B(n407), .ZN(n411) );
  NAND2_X1 U479 ( .A1(G232GAT), .A2(G233GAT), .ZN(n408) );
  XNOR2_X1 U480 ( .A(n413), .B(n412), .ZN(n417) );
  XOR2_X1 U481 ( .A(KEYINPUT74), .B(KEYINPUT76), .Z(n415) );
  XNOR2_X1 U482 ( .A(KEYINPUT10), .B(KEYINPUT66), .ZN(n414) );
  XNOR2_X1 U483 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U484 ( .A(n417), .B(n416), .Z(n422) );
  XOR2_X1 U485 ( .A(G29GAT), .B(G43GAT), .Z(n419) );
  XNOR2_X1 U486 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n418) );
  XNOR2_X1 U487 ( .A(n419), .B(n418), .ZN(n452) );
  XNOR2_X1 U488 ( .A(n452), .B(n420), .ZN(n421) );
  NAND2_X1 U489 ( .A1(n423), .A2(n592), .ZN(n424) );
  XOR2_X1 U490 ( .A(KEYINPUT37), .B(n424), .Z(n534) );
  NAND2_X1 U491 ( .A1(KEYINPUT72), .A2(n425), .ZN(n429) );
  INV_X1 U492 ( .A(KEYINPUT72), .ZN(n427) );
  INV_X1 U493 ( .A(n425), .ZN(n426) );
  NAND2_X1 U494 ( .A1(n427), .A2(n426), .ZN(n428) );
  NAND2_X1 U495 ( .A1(n429), .A2(n428), .ZN(n435) );
  XOR2_X1 U496 ( .A(KEYINPUT31), .B(KEYINPUT32), .Z(n431) );
  XNOR2_X1 U497 ( .A(G204GAT), .B(KEYINPUT33), .ZN(n430) );
  XNOR2_X1 U498 ( .A(n431), .B(n430), .ZN(n433) );
  AND2_X1 U499 ( .A1(G230GAT), .A2(G233GAT), .ZN(n432) );
  XOR2_X1 U500 ( .A(n437), .B(n436), .Z(n438) );
  XNOR2_X1 U501 ( .A(n439), .B(n438), .ZN(n444) );
  XOR2_X1 U502 ( .A(G197GAT), .B(G141GAT), .Z(n446) );
  XNOR2_X1 U503 ( .A(G15GAT), .B(G22GAT), .ZN(n445) );
  XNOR2_X1 U504 ( .A(n446), .B(n445), .ZN(n450) );
  XOR2_X1 U505 ( .A(KEYINPUT68), .B(KEYINPUT30), .Z(n448) );
  XNOR2_X1 U506 ( .A(KEYINPUT69), .B(KEYINPUT29), .ZN(n447) );
  XNOR2_X1 U507 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U508 ( .A(n450), .B(n449), .ZN(n460) );
  XOR2_X1 U509 ( .A(n452), .B(n451), .Z(n454) );
  NAND2_X1 U510 ( .A1(G229GAT), .A2(G233GAT), .ZN(n453) );
  XNOR2_X1 U511 ( .A(n454), .B(n453), .ZN(n456) );
  XOR2_X1 U512 ( .A(n456), .B(n455), .Z(n458) );
  XNOR2_X1 U513 ( .A(G50GAT), .B(G36GAT), .ZN(n457) );
  XNOR2_X1 U514 ( .A(n458), .B(n457), .ZN(n459) );
  XOR2_X1 U515 ( .A(n460), .B(n459), .Z(n548) );
  NAND2_X1 U516 ( .A1(n585), .A2(n548), .ZN(n505) );
  XNOR2_X1 U517 ( .A(KEYINPUT38), .B(KEYINPUT104), .ZN(n461) );
  NAND2_X1 U518 ( .A1(n520), .A2(n541), .ZN(n466) );
  XOR2_X1 U519 ( .A(KEYINPUT106), .B(KEYINPUT40), .Z(n464) );
  XNOR2_X1 U520 ( .A(G43GAT), .B(KEYINPUT105), .ZN(n463) );
  INV_X1 U521 ( .A(n548), .ZN(n581) );
  INV_X1 U522 ( .A(KEYINPUT54), .ZN(n480) );
  XOR2_X1 U523 ( .A(KEYINPUT41), .B(n585), .Z(n570) );
  NOR2_X1 U524 ( .A1(n581), .A2(n570), .ZN(n467) );
  XOR2_X1 U525 ( .A(n467), .B(KEYINPUT46), .Z(n469) );
  INV_X1 U526 ( .A(n574), .ZN(n495) );
  NOR2_X1 U527 ( .A1(n495), .A2(n555), .ZN(n468) );
  NAND2_X1 U528 ( .A1(n469), .A2(n468), .ZN(n470) );
  XNOR2_X1 U529 ( .A(n470), .B(KEYINPUT47), .ZN(n476) );
  NAND2_X1 U530 ( .A1(n555), .A2(n592), .ZN(n472) );
  XNOR2_X1 U531 ( .A(KEYINPUT45), .B(KEYINPUT113), .ZN(n471) );
  XNOR2_X1 U532 ( .A(n472), .B(n471), .ZN(n473) );
  NAND2_X1 U533 ( .A1(n473), .A2(n585), .ZN(n474) );
  NOR2_X1 U534 ( .A1(n548), .A2(n474), .ZN(n475) );
  NOR2_X1 U535 ( .A1(n476), .A2(n475), .ZN(n477) );
  XNOR2_X1 U536 ( .A(n477), .B(KEYINPUT48), .ZN(n489) );
  INV_X1 U537 ( .A(n538), .ZN(n478) );
  NOR2_X1 U538 ( .A1(n489), .A2(n478), .ZN(n479) );
  XNOR2_X1 U539 ( .A(n480), .B(n479), .ZN(n481) );
  NAND2_X1 U540 ( .A1(n482), .A2(n580), .ZN(n483) );
  XNOR2_X1 U541 ( .A(n483), .B(KEYINPUT55), .ZN(n484) );
  NAND2_X1 U542 ( .A1(n484), .A2(n541), .ZN(n485) );
  XNOR2_X1 U543 ( .A(n485), .B(KEYINPUT122), .ZN(n575) );
  NOR2_X1 U544 ( .A1(n581), .A2(n575), .ZN(n487) );
  NOR2_X1 U545 ( .A1(n489), .A2(n488), .ZN(n490) );
  XNOR2_X1 U546 ( .A(n490), .B(KEYINPUT114), .ZN(n559) );
  NAND2_X1 U547 ( .A1(n559), .A2(n541), .ZN(n492) );
  INV_X1 U548 ( .A(KEYINPUT115), .ZN(n491) );
  XNOR2_X1 U549 ( .A(n492), .B(n491), .ZN(n493) );
  NOR2_X1 U550 ( .A1(n544), .A2(n493), .ZN(n494) );
  XNOR2_X1 U551 ( .A(KEYINPUT116), .B(n494), .ZN(n556) );
  NAND2_X1 U552 ( .A1(n495), .A2(n556), .ZN(n499) );
  XOR2_X1 U553 ( .A(KEYINPUT119), .B(KEYINPUT51), .Z(n497) );
  XOR2_X1 U554 ( .A(G134GAT), .B(KEYINPUT120), .Z(n496) );
  XNOR2_X1 U555 ( .A(n499), .B(n498), .ZN(G1343GAT) );
  XOR2_X1 U556 ( .A(KEYINPUT34), .B(KEYINPUT100), .Z(n508) );
  NAND2_X1 U557 ( .A1(n555), .A2(n574), .ZN(n500) );
  XNOR2_X1 U558 ( .A(n500), .B(KEYINPUT81), .ZN(n501) );
  XNOR2_X1 U559 ( .A(KEYINPUT16), .B(n501), .ZN(n503) );
  NAND2_X1 U560 ( .A1(n503), .A2(n502), .ZN(n504) );
  XNOR2_X1 U561 ( .A(n504), .B(KEYINPUT98), .ZN(n526) );
  NOR2_X1 U562 ( .A1(n526), .A2(n505), .ZN(n506) );
  XOR2_X1 U563 ( .A(KEYINPUT99), .B(n506), .Z(n515) );
  NAND2_X1 U564 ( .A1(n515), .A2(n536), .ZN(n507) );
  XNOR2_X1 U565 ( .A(n508), .B(n507), .ZN(n509) );
  XOR2_X1 U566 ( .A(G1GAT), .B(n509), .Z(G1324GAT) );
  NAND2_X1 U567 ( .A1(n515), .A2(n538), .ZN(n510) );
  XNOR2_X1 U568 ( .A(n510), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U569 ( .A(KEYINPUT35), .B(KEYINPUT102), .Z(n512) );
  NAND2_X1 U570 ( .A1(n515), .A2(n541), .ZN(n511) );
  XNOR2_X1 U571 ( .A(n512), .B(n511), .ZN(n514) );
  XOR2_X1 U572 ( .A(G15GAT), .B(KEYINPUT101), .Z(n513) );
  XNOR2_X1 U573 ( .A(n514), .B(n513), .ZN(G1326GAT) );
  NAND2_X1 U574 ( .A1(n515), .A2(n544), .ZN(n516) );
  XNOR2_X1 U575 ( .A(n516), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U576 ( .A1(n520), .A2(n536), .ZN(n518) );
  XOR2_X1 U577 ( .A(G29GAT), .B(KEYINPUT39), .Z(n517) );
  XNOR2_X1 U578 ( .A(n518), .B(n517), .ZN(G1328GAT) );
  NAND2_X1 U579 ( .A1(n520), .A2(n538), .ZN(n519) );
  XNOR2_X1 U580 ( .A(n519), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U581 ( .A(G50GAT), .B(KEYINPUT107), .Z(n522) );
  NAND2_X1 U582 ( .A1(n520), .A2(n544), .ZN(n521) );
  XNOR2_X1 U583 ( .A(n522), .B(n521), .ZN(G1331GAT) );
  XNOR2_X1 U584 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n523) );
  XNOR2_X1 U585 ( .A(n523), .B(KEYINPUT110), .ZN(n524) );
  XOR2_X1 U586 ( .A(KEYINPUT109), .B(n524), .Z(n528) );
  INV_X1 U587 ( .A(n570), .ZN(n550) );
  NAND2_X1 U588 ( .A1(n550), .A2(n581), .ZN(n525) );
  XNOR2_X1 U589 ( .A(n525), .B(KEYINPUT108), .ZN(n535) );
  NOR2_X1 U590 ( .A1(n535), .A2(n526), .ZN(n531) );
  NAND2_X1 U591 ( .A1(n531), .A2(n536), .ZN(n527) );
  XNOR2_X1 U592 ( .A(n528), .B(n527), .ZN(G1332GAT) );
  NAND2_X1 U593 ( .A1(n531), .A2(n538), .ZN(n529) );
  XNOR2_X1 U594 ( .A(n529), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U595 ( .A1(n531), .A2(n541), .ZN(n530) );
  XNOR2_X1 U596 ( .A(n530), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U597 ( .A(G78GAT), .B(KEYINPUT43), .Z(n533) );
  NAND2_X1 U598 ( .A1(n531), .A2(n544), .ZN(n532) );
  XNOR2_X1 U599 ( .A(n533), .B(n532), .ZN(G1335GAT) );
  NOR2_X1 U600 ( .A1(n535), .A2(n534), .ZN(n545) );
  NAND2_X1 U601 ( .A1(n545), .A2(n536), .ZN(n537) );
  XNOR2_X1 U602 ( .A(G85GAT), .B(n537), .ZN(G1336GAT) );
  XOR2_X1 U603 ( .A(G92GAT), .B(KEYINPUT111), .Z(n540) );
  NAND2_X1 U604 ( .A1(n545), .A2(n538), .ZN(n539) );
  XNOR2_X1 U605 ( .A(n540), .B(n539), .ZN(G1337GAT) );
  NAND2_X1 U606 ( .A1(n545), .A2(n541), .ZN(n542) );
  XNOR2_X1 U607 ( .A(n542), .B(KEYINPUT112), .ZN(n543) );
  XNOR2_X1 U608 ( .A(G99GAT), .B(n543), .ZN(G1338GAT) );
  NAND2_X1 U609 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U610 ( .A(n546), .B(KEYINPUT44), .ZN(n547) );
  XNOR2_X1 U611 ( .A(G106GAT), .B(n547), .ZN(G1339GAT) );
  NAND2_X1 U612 ( .A1(n548), .A2(n556), .ZN(n549) );
  XNOR2_X1 U613 ( .A(G113GAT), .B(n549), .ZN(G1340GAT) );
  XOR2_X1 U614 ( .A(G120GAT), .B(KEYINPUT117), .Z(n552) );
  NAND2_X1 U615 ( .A1(n556), .A2(n550), .ZN(n551) );
  XNOR2_X1 U616 ( .A(n552), .B(n551), .ZN(n554) );
  XOR2_X1 U617 ( .A(KEYINPUT49), .B(KEYINPUT118), .Z(n553) );
  XNOR2_X1 U618 ( .A(n554), .B(n553), .ZN(G1341GAT) );
  NAND2_X1 U619 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U620 ( .A(n557), .B(KEYINPUT50), .ZN(n558) );
  XNOR2_X1 U621 ( .A(G127GAT), .B(n558), .ZN(G1342GAT) );
  NAND2_X1 U622 ( .A1(n559), .A2(n579), .ZN(n566) );
  NOR2_X1 U623 ( .A1(n581), .A2(n566), .ZN(n561) );
  XNOR2_X1 U624 ( .A(G141GAT), .B(KEYINPUT121), .ZN(n560) );
  XNOR2_X1 U625 ( .A(n561), .B(n560), .ZN(G1344GAT) );
  NOR2_X1 U626 ( .A1(n570), .A2(n566), .ZN(n563) );
  XNOR2_X1 U627 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n563), .B(n562), .ZN(n564) );
  XNOR2_X1 U629 ( .A(G148GAT), .B(n564), .ZN(G1345GAT) );
  NOR2_X1 U630 ( .A1(n588), .A2(n566), .ZN(n565) );
  XOR2_X1 U631 ( .A(G155GAT), .B(n565), .Z(G1346GAT) );
  NOR2_X1 U632 ( .A1(n574), .A2(n566), .ZN(n567) );
  XOR2_X1 U633 ( .A(G162GAT), .B(n567), .Z(G1347GAT) );
  XOR2_X1 U634 ( .A(KEYINPUT56), .B(KEYINPUT124), .Z(n569) );
  XNOR2_X1 U635 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n568) );
  XNOR2_X1 U636 ( .A(n569), .B(n568), .ZN(n572) );
  NOR2_X1 U637 ( .A1(n570), .A2(n575), .ZN(n571) );
  XOR2_X1 U638 ( .A(n572), .B(n571), .Z(G1349GAT) );
  NOR2_X1 U639 ( .A1(n588), .A2(n575), .ZN(n573) );
  XOR2_X1 U640 ( .A(G183GAT), .B(n573), .Z(G1350GAT) );
  NOR2_X1 U641 ( .A1(n575), .A2(n574), .ZN(n577) );
  XNOR2_X1 U642 ( .A(KEYINPUT58), .B(KEYINPUT125), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U644 ( .A(G190GAT), .B(n578), .ZN(G1351GAT) );
  NAND2_X1 U645 ( .A1(n580), .A2(n579), .ZN(n590) );
  NOR2_X1 U646 ( .A1(n581), .A2(n590), .ZN(n583) );
  XNOR2_X1 U647 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U649 ( .A(G197GAT), .B(n584), .ZN(G1352GAT) );
  NOR2_X1 U650 ( .A1(n585), .A2(n590), .ZN(n587) );
  XNOR2_X1 U651 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n586) );
  XNOR2_X1 U652 ( .A(n587), .B(n586), .ZN(G1353GAT) );
  NOR2_X1 U653 ( .A1(n588), .A2(n590), .ZN(n589) );
  XOR2_X1 U654 ( .A(G211GAT), .B(n589), .Z(G1354GAT) );
  INV_X1 U655 ( .A(n590), .ZN(n591) );
  NAND2_X1 U656 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U657 ( .A(n593), .B(KEYINPUT62), .ZN(n594) );
  XOR2_X1 U658 ( .A(n594), .B(KEYINPUT126), .Z(n596) );
  XNOR2_X1 U659 ( .A(G218GAT), .B(KEYINPUT127), .ZN(n595) );
  XNOR2_X1 U660 ( .A(n596), .B(n595), .ZN(G1355GAT) );
endmodule

