

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593;

  NOR2_X2 U322 ( .A1(n584), .A2(n517), .ZN(n518) );
  XNOR2_X2 U323 ( .A(n340), .B(n521), .ZN(n472) );
  XOR2_X2 U324 ( .A(n339), .B(n338), .Z(n521) );
  NOR2_X2 U325 ( .A1(n579), .A2(n578), .ZN(n589) );
  NOR2_X2 U326 ( .A1(n565), .A2(n564), .ZN(n573) );
  INV_X1 U327 ( .A(KEYINPUT27), .ZN(n355) );
  XNOR2_X1 U328 ( .A(KEYINPUT38), .B(n464), .ZN(n492) );
  XOR2_X1 U329 ( .A(n562), .B(KEYINPUT28), .Z(n529) );
  XNOR2_X1 U330 ( .A(n392), .B(n391), .ZN(n565) );
  XOR2_X1 U331 ( .A(n373), .B(n372), .Z(n290) );
  XOR2_X1 U332 ( .A(G204GAT), .B(G92GAT), .Z(n291) );
  XNOR2_X1 U333 ( .A(n318), .B(n317), .ZN(n319) );
  INV_X1 U334 ( .A(G22GAT), .ZN(n365) );
  XNOR2_X1 U335 ( .A(n320), .B(n319), .ZN(n323) );
  XNOR2_X1 U336 ( .A(n366), .B(n365), .ZN(n367) );
  XNOR2_X1 U337 ( .A(n355), .B(KEYINPUT100), .ZN(n356) );
  XNOR2_X1 U338 ( .A(n368), .B(n367), .ZN(n369) );
  XNOR2_X1 U339 ( .A(n556), .B(n356), .ZN(n396) );
  XNOR2_X1 U340 ( .A(KEYINPUT125), .B(KEYINPUT54), .ZN(n558) );
  XNOR2_X1 U341 ( .A(n559), .B(n558), .ZN(n561) );
  XNOR2_X1 U342 ( .A(n446), .B(n291), .ZN(n351) );
  XNOR2_X1 U343 ( .A(n352), .B(n351), .ZN(n353) );
  INV_X1 U344 ( .A(KEYINPUT114), .ZN(n469) );
  INV_X1 U345 ( .A(G29GAT), .ZN(n465) );
  XNOR2_X1 U346 ( .A(n469), .B(G50GAT), .ZN(n470) );
  XNOR2_X1 U347 ( .A(n466), .B(n465), .ZN(n467) );
  XNOR2_X1 U348 ( .A(n471), .B(n470), .ZN(G1331GAT) );
  XOR2_X1 U349 ( .A(KEYINPUT91), .B(KEYINPUT3), .Z(n293) );
  XNOR2_X1 U350 ( .A(KEYINPUT2), .B(G155GAT), .ZN(n292) );
  XNOR2_X1 U351 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U352 ( .A(G141GAT), .B(n294), .Z(n374) );
  XOR2_X1 U353 ( .A(G29GAT), .B(G134GAT), .Z(n312) );
  XOR2_X1 U354 ( .A(G1GAT), .B(G127GAT), .Z(n408) );
  XOR2_X1 U355 ( .A(n312), .B(n408), .Z(n296) );
  XNOR2_X1 U356 ( .A(G162GAT), .B(G85GAT), .ZN(n295) );
  XNOR2_X1 U357 ( .A(n296), .B(n295), .ZN(n308) );
  XOR2_X1 U358 ( .A(KEYINPUT94), .B(KEYINPUT1), .Z(n298) );
  XNOR2_X1 U359 ( .A(KEYINPUT4), .B(KEYINPUT92), .ZN(n297) );
  XNOR2_X1 U360 ( .A(n298), .B(n297), .ZN(n302) );
  XOR2_X1 U361 ( .A(KEYINPUT5), .B(KEYINPUT93), .Z(n300) );
  XNOR2_X1 U362 ( .A(KEYINPUT6), .B(KEYINPUT95), .ZN(n299) );
  XNOR2_X1 U363 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U364 ( .A(n302), .B(n301), .Z(n306) );
  XNOR2_X1 U365 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n303) );
  XNOR2_X1 U366 ( .A(n303), .B(KEYINPUT87), .ZN(n383) );
  XNOR2_X1 U367 ( .A(G120GAT), .B(G148GAT), .ZN(n304) );
  XNOR2_X1 U368 ( .A(n304), .B(G57GAT), .ZN(n455) );
  XNOR2_X1 U369 ( .A(n383), .B(n455), .ZN(n305) );
  XNOR2_X1 U370 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X1 U371 ( .A(n308), .B(n307), .Z(n310) );
  NAND2_X1 U372 ( .A1(G225GAT), .A2(G233GAT), .ZN(n309) );
  XNOR2_X1 U373 ( .A(n310), .B(n309), .ZN(n311) );
  XNOR2_X1 U374 ( .A(n374), .B(n311), .ZN(n402) );
  XNOR2_X1 U375 ( .A(KEYINPUT96), .B(n402), .ZN(n560) );
  INV_X1 U376 ( .A(KEYINPUT82), .ZN(n340) );
  XOR2_X1 U377 ( .A(KEYINPUT79), .B(KEYINPUT67), .Z(n314) );
  XOR2_X1 U378 ( .A(G50GAT), .B(G162GAT), .Z(n361) );
  XNOR2_X1 U379 ( .A(n361), .B(n312), .ZN(n313) );
  XNOR2_X1 U380 ( .A(n314), .B(n313), .ZN(n320) );
  XOR2_X1 U381 ( .A(KEYINPUT9), .B(KEYINPUT68), .Z(n316) );
  XNOR2_X1 U382 ( .A(KEYINPUT80), .B(KEYINPUT11), .ZN(n315) );
  XNOR2_X1 U383 ( .A(n316), .B(n315), .ZN(n318) );
  AND2_X1 U384 ( .A1(G232GAT), .A2(G233GAT), .ZN(n317) );
  INV_X1 U385 ( .A(n323), .ZN(n321) );
  NAND2_X1 U386 ( .A1(n321), .A2(KEYINPUT10), .ZN(n325) );
  INV_X1 U387 ( .A(KEYINPUT10), .ZN(n322) );
  NAND2_X1 U388 ( .A1(n323), .A2(n322), .ZN(n324) );
  NAND2_X1 U389 ( .A1(n325), .A2(n324), .ZN(n329) );
  XOR2_X1 U390 ( .A(KEYINPUT81), .B(G218GAT), .Z(n327) );
  XNOR2_X1 U391 ( .A(G36GAT), .B(G190GAT), .ZN(n326) );
  XNOR2_X1 U392 ( .A(n327), .B(n326), .ZN(n343) );
  XNOR2_X1 U393 ( .A(n343), .B(KEYINPUT65), .ZN(n328) );
  XNOR2_X1 U394 ( .A(n329), .B(n328), .ZN(n339) );
  XOR2_X1 U395 ( .A(G43GAT), .B(KEYINPUT8), .Z(n331) );
  XNOR2_X1 U396 ( .A(KEYINPUT74), .B(KEYINPUT7), .ZN(n330) );
  XNOR2_X1 U397 ( .A(n331), .B(n330), .ZN(n437) );
  INV_X1 U398 ( .A(G92GAT), .ZN(n332) );
  NAND2_X1 U399 ( .A1(G85GAT), .A2(n332), .ZN(n335) );
  INV_X1 U400 ( .A(G85GAT), .ZN(n333) );
  NAND2_X1 U401 ( .A1(n333), .A2(G92GAT), .ZN(n334) );
  NAND2_X1 U402 ( .A1(n335), .A2(n334), .ZN(n337) );
  XNOR2_X1 U403 ( .A(G99GAT), .B(G106GAT), .ZN(n336) );
  XNOR2_X1 U404 ( .A(n337), .B(n336), .ZN(n448) );
  XOR2_X1 U405 ( .A(n437), .B(n448), .Z(n338) );
  XOR2_X1 U406 ( .A(n472), .B(KEYINPUT36), .Z(n591) );
  XOR2_X1 U407 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n342) );
  XNOR2_X1 U408 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n341) );
  XNOR2_X1 U409 ( .A(n342), .B(n341), .ZN(n385) );
  XOR2_X1 U410 ( .A(n385), .B(n343), .Z(n354) );
  XOR2_X1 U411 ( .A(KEYINPUT97), .B(KEYINPUT98), .Z(n345) );
  NAND2_X1 U412 ( .A1(G226GAT), .A2(G233GAT), .ZN(n344) );
  XNOR2_X1 U413 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U414 ( .A(n346), .B(KEYINPUT99), .Z(n350) );
  XNOR2_X1 U415 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n347) );
  XNOR2_X1 U416 ( .A(n347), .B(G211GAT), .ZN(n368) );
  XNOR2_X1 U417 ( .A(G8GAT), .B(G183GAT), .ZN(n348) );
  XNOR2_X1 U418 ( .A(n348), .B(KEYINPUT83), .ZN(n420) );
  XNOR2_X1 U419 ( .A(n368), .B(n420), .ZN(n349) );
  XNOR2_X1 U420 ( .A(n350), .B(n349), .ZN(n352) );
  XOR2_X1 U421 ( .A(G176GAT), .B(G64GAT), .Z(n446) );
  XNOR2_X1 U422 ( .A(n354), .B(n353), .ZN(n556) );
  INV_X1 U423 ( .A(n396), .ZN(n357) );
  NOR2_X1 U424 ( .A1(n357), .A2(n560), .ZN(n358) );
  XNOR2_X1 U425 ( .A(n358), .B(KEYINPUT101), .ZN(n528) );
  XOR2_X1 U426 ( .A(KEYINPUT89), .B(KEYINPUT24), .Z(n360) );
  XNOR2_X1 U427 ( .A(KEYINPUT22), .B(KEYINPUT23), .ZN(n359) );
  XNOR2_X1 U428 ( .A(n360), .B(n359), .ZN(n373) );
  XOR2_X1 U429 ( .A(KEYINPUT90), .B(G148GAT), .Z(n363) );
  XOR2_X1 U430 ( .A(G204GAT), .B(G78GAT), .Z(n447) );
  XNOR2_X1 U431 ( .A(n361), .B(n447), .ZN(n362) );
  XNOR2_X1 U432 ( .A(n363), .B(n362), .ZN(n364) );
  XOR2_X1 U433 ( .A(n364), .B(G106GAT), .Z(n371) );
  NAND2_X1 U434 ( .A1(G228GAT), .A2(G233GAT), .ZN(n366) );
  XNOR2_X1 U435 ( .A(n369), .B(G218GAT), .ZN(n370) );
  XNOR2_X1 U436 ( .A(n371), .B(n370), .ZN(n372) );
  XOR2_X1 U437 ( .A(n374), .B(n290), .Z(n562) );
  INV_X1 U438 ( .A(n529), .ZN(n375) );
  NOR2_X1 U439 ( .A1(n528), .A2(n375), .ZN(n393) );
  XOR2_X1 U440 ( .A(G183GAT), .B(G120GAT), .Z(n377) );
  XNOR2_X1 U441 ( .A(G15GAT), .B(G127GAT), .ZN(n376) );
  XNOR2_X1 U442 ( .A(n377), .B(n376), .ZN(n381) );
  XOR2_X1 U443 ( .A(KEYINPUT88), .B(KEYINPUT66), .Z(n379) );
  XNOR2_X1 U444 ( .A(G176GAT), .B(KEYINPUT20), .ZN(n378) );
  XNOR2_X1 U445 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U446 ( .A(n381), .B(n380), .ZN(n392) );
  XNOR2_X1 U447 ( .A(G99GAT), .B(G190GAT), .ZN(n382) );
  XNOR2_X1 U448 ( .A(n382), .B(G134GAT), .ZN(n384) );
  XOR2_X1 U449 ( .A(n384), .B(n383), .Z(n390) );
  XOR2_X1 U450 ( .A(n385), .B(G71GAT), .Z(n387) );
  NAND2_X1 U451 ( .A1(G227GAT), .A2(G233GAT), .ZN(n386) );
  XNOR2_X1 U452 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U453 ( .A(G43GAT), .B(n388), .ZN(n389) );
  XNOR2_X1 U454 ( .A(n390), .B(n389), .ZN(n391) );
  NAND2_X1 U455 ( .A1(n393), .A2(n565), .ZN(n394) );
  XNOR2_X1 U456 ( .A(n394), .B(KEYINPUT102), .ZN(n405) );
  NAND2_X1 U457 ( .A1(n562), .A2(n565), .ZN(n395) );
  XOR2_X1 U458 ( .A(KEYINPUT26), .B(n395), .Z(n577) );
  NAND2_X1 U459 ( .A1(n577), .A2(n396), .ZN(n401) );
  NOR2_X1 U460 ( .A1(n565), .A2(n556), .ZN(n397) );
  NOR2_X1 U461 ( .A1(n562), .A2(n397), .ZN(n398) );
  XOR2_X1 U462 ( .A(n398), .B(KEYINPUT25), .Z(n399) );
  XNOR2_X1 U463 ( .A(KEYINPUT103), .B(n399), .ZN(n400) );
  NAND2_X1 U464 ( .A1(n401), .A2(n400), .ZN(n403) );
  NAND2_X1 U465 ( .A1(n403), .A2(n402), .ZN(n404) );
  NAND2_X1 U466 ( .A1(n405), .A2(n404), .ZN(n476) );
  XOR2_X1 U467 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n407) );
  XNOR2_X1 U468 ( .A(KEYINPUT12), .B(KEYINPUT84), .ZN(n406) );
  XNOR2_X1 U469 ( .A(n407), .B(n406), .ZN(n412) );
  XOR2_X1 U470 ( .A(n408), .B(G78GAT), .Z(n410) );
  XOR2_X1 U471 ( .A(G15GAT), .B(G22GAT), .Z(n436) );
  XNOR2_X1 U472 ( .A(n436), .B(G155GAT), .ZN(n409) );
  XNOR2_X1 U473 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U474 ( .A(n412), .B(n411), .Z(n414) );
  NAND2_X1 U475 ( .A1(G231GAT), .A2(G233GAT), .ZN(n413) );
  XNOR2_X1 U476 ( .A(n414), .B(n413), .ZN(n418) );
  XOR2_X1 U477 ( .A(KEYINPUT85), .B(G57GAT), .Z(n416) );
  XNOR2_X1 U478 ( .A(G211GAT), .B(G64GAT), .ZN(n415) );
  XNOR2_X1 U479 ( .A(n416), .B(n415), .ZN(n417) );
  XOR2_X1 U480 ( .A(n418), .B(n417), .Z(n422) );
  XNOR2_X1 U481 ( .A(G71GAT), .B(KEYINPUT13), .ZN(n419) );
  XNOR2_X1 U482 ( .A(n419), .B(KEYINPUT75), .ZN(n456) );
  XNOR2_X1 U483 ( .A(n420), .B(n456), .ZN(n421) );
  XOR2_X1 U484 ( .A(n422), .B(n421), .Z(n587) );
  INV_X1 U485 ( .A(n587), .ZN(n551) );
  NAND2_X1 U486 ( .A1(n476), .A2(n551), .ZN(n423) );
  XNOR2_X1 U487 ( .A(n423), .B(KEYINPUT108), .ZN(n424) );
  NOR2_X1 U488 ( .A1(n591), .A2(n424), .ZN(n425) );
  XNOR2_X1 U489 ( .A(n425), .B(KEYINPUT37), .ZN(n508) );
  XOR2_X1 U490 ( .A(KEYINPUT30), .B(KEYINPUT71), .Z(n427) );
  XNOR2_X1 U491 ( .A(KEYINPUT72), .B(KEYINPUT70), .ZN(n426) );
  XNOR2_X1 U492 ( .A(n427), .B(n426), .ZN(n445) );
  XOR2_X1 U493 ( .A(G50GAT), .B(G29GAT), .Z(n429) );
  XNOR2_X1 U494 ( .A(G169GAT), .B(G36GAT), .ZN(n428) );
  XNOR2_X1 U495 ( .A(n429), .B(n428), .ZN(n433) );
  XOR2_X1 U496 ( .A(G8GAT), .B(G197GAT), .Z(n431) );
  XNOR2_X1 U497 ( .A(G113GAT), .B(G141GAT), .ZN(n430) );
  XNOR2_X1 U498 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U499 ( .A(n433), .B(n432), .Z(n443) );
  XOR2_X1 U500 ( .A(G1GAT), .B(KEYINPUT73), .Z(n435) );
  XNOR2_X1 U501 ( .A(KEYINPUT69), .B(KEYINPUT29), .ZN(n434) );
  XNOR2_X1 U502 ( .A(n435), .B(n434), .ZN(n441) );
  XOR2_X1 U503 ( .A(n437), .B(n436), .Z(n439) );
  NAND2_X1 U504 ( .A1(G229GAT), .A2(G233GAT), .ZN(n438) );
  XNOR2_X1 U505 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U506 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U507 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U508 ( .A(n445), .B(n444), .ZN(n580) );
  INV_X1 U509 ( .A(n580), .ZN(n544) );
  XNOR2_X1 U510 ( .A(n447), .B(n446), .ZN(n460) );
  XOR2_X1 U511 ( .A(n448), .B(KEYINPUT33), .Z(n450) );
  NAND2_X1 U512 ( .A1(G230GAT), .A2(G233GAT), .ZN(n449) );
  XNOR2_X1 U513 ( .A(n450), .B(n449), .ZN(n454) );
  XOR2_X1 U514 ( .A(KEYINPUT31), .B(KEYINPUT76), .Z(n452) );
  XNOR2_X1 U515 ( .A(KEYINPUT77), .B(KEYINPUT32), .ZN(n451) );
  XNOR2_X1 U516 ( .A(n452), .B(n451), .ZN(n453) );
  XOR2_X1 U517 ( .A(n454), .B(n453), .Z(n458) );
  XNOR2_X1 U518 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U519 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U520 ( .A(n460), .B(n459), .ZN(n495) );
  BUF_X1 U521 ( .A(n495), .Z(n584) );
  NOR2_X1 U522 ( .A1(n544), .A2(n584), .ZN(n461) );
  XOR2_X1 U523 ( .A(KEYINPUT78), .B(n461), .Z(n478) );
  NOR2_X1 U524 ( .A1(n508), .A2(n478), .ZN(n463) );
  XNOR2_X1 U525 ( .A(KEYINPUT109), .B(KEYINPUT110), .ZN(n462) );
  XNOR2_X1 U526 ( .A(n463), .B(n462), .ZN(n464) );
  NOR2_X1 U527 ( .A1(n560), .A2(n492), .ZN(n468) );
  XNOR2_X1 U528 ( .A(KEYINPUT111), .B(KEYINPUT39), .ZN(n466) );
  XNOR2_X1 U529 ( .A(n468), .B(n467), .ZN(G1328GAT) );
  NOR2_X1 U530 ( .A1(n529), .A2(n492), .ZN(n471) );
  XOR2_X1 U531 ( .A(KEYINPUT16), .B(KEYINPUT86), .Z(n474) );
  INV_X1 U532 ( .A(n472), .ZN(n538) );
  NAND2_X1 U533 ( .A1(n587), .A2(n538), .ZN(n473) );
  XNOR2_X1 U534 ( .A(n474), .B(n473), .ZN(n475) );
  NAND2_X1 U535 ( .A1(n476), .A2(n475), .ZN(n477) );
  XNOR2_X1 U536 ( .A(n477), .B(KEYINPUT104), .ZN(n497) );
  OR2_X1 U537 ( .A1(n478), .A2(n497), .ZN(n486) );
  NOR2_X1 U538 ( .A1(n560), .A2(n486), .ZN(n480) );
  XNOR2_X1 U539 ( .A(KEYINPUT34), .B(KEYINPUT105), .ZN(n479) );
  XNOR2_X1 U540 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U541 ( .A(G1GAT), .B(n481), .ZN(G1324GAT) );
  NOR2_X1 U542 ( .A1(n556), .A2(n486), .ZN(n482) );
  XOR2_X1 U543 ( .A(G8GAT), .B(n482), .Z(G1325GAT) );
  NOR2_X1 U544 ( .A1(n565), .A2(n486), .ZN(n484) );
  XNOR2_X1 U545 ( .A(KEYINPUT106), .B(KEYINPUT35), .ZN(n483) );
  XNOR2_X1 U546 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U547 ( .A(G15GAT), .B(n485), .ZN(G1326GAT) );
  NOR2_X1 U548 ( .A1(n529), .A2(n486), .ZN(n488) );
  XNOR2_X1 U549 ( .A(G22GAT), .B(KEYINPUT107), .ZN(n487) );
  XNOR2_X1 U550 ( .A(n488), .B(n487), .ZN(G1327GAT) );
  NOR2_X1 U551 ( .A1(n556), .A2(n492), .ZN(n489) );
  XOR2_X1 U552 ( .A(G36GAT), .B(n489), .Z(G1329GAT) );
  XOR2_X1 U553 ( .A(KEYINPUT112), .B(KEYINPUT113), .Z(n491) );
  XNOR2_X1 U554 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n490) );
  XNOR2_X1 U555 ( .A(n491), .B(n490), .ZN(n494) );
  NOR2_X1 U556 ( .A1(n565), .A2(n492), .ZN(n493) );
  XOR2_X1 U557 ( .A(n494), .B(n493), .Z(G1330GAT) );
  XNOR2_X1 U558 ( .A(n495), .B(KEYINPUT41), .ZN(n496) );
  XNOR2_X1 U559 ( .A(n496), .B(KEYINPUT64), .ZN(n546) );
  XNOR2_X1 U560 ( .A(n546), .B(KEYINPUT115), .ZN(n567) );
  NAND2_X1 U561 ( .A1(n544), .A2(n567), .ZN(n507) );
  OR2_X1 U562 ( .A1(n497), .A2(n507), .ZN(n504) );
  NOR2_X1 U563 ( .A1(n560), .A2(n504), .ZN(n498) );
  XOR2_X1 U564 ( .A(n498), .B(KEYINPUT42), .Z(n499) );
  XNOR2_X1 U565 ( .A(G57GAT), .B(n499), .ZN(G1332GAT) );
  NOR2_X1 U566 ( .A1(n556), .A2(n504), .ZN(n500) );
  XOR2_X1 U567 ( .A(KEYINPUT116), .B(n500), .Z(n501) );
  XNOR2_X1 U568 ( .A(G64GAT), .B(n501), .ZN(G1333GAT) );
  NOR2_X1 U569 ( .A1(n565), .A2(n504), .ZN(n503) );
  XNOR2_X1 U570 ( .A(G71GAT), .B(KEYINPUT117), .ZN(n502) );
  XNOR2_X1 U571 ( .A(n503), .B(n502), .ZN(G1334GAT) );
  NOR2_X1 U572 ( .A1(n529), .A2(n504), .ZN(n506) );
  XNOR2_X1 U573 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n505) );
  XNOR2_X1 U574 ( .A(n506), .B(n505), .ZN(G1335GAT) );
  OR2_X1 U575 ( .A1(n508), .A2(n507), .ZN(n512) );
  NOR2_X1 U576 ( .A1(n560), .A2(n512), .ZN(n509) );
  XOR2_X1 U577 ( .A(G85GAT), .B(n509), .Z(G1336GAT) );
  NOR2_X1 U578 ( .A1(n556), .A2(n512), .ZN(n510) );
  XOR2_X1 U579 ( .A(G92GAT), .B(n510), .Z(G1337GAT) );
  NOR2_X1 U580 ( .A1(n565), .A2(n512), .ZN(n511) );
  XOR2_X1 U581 ( .A(G99GAT), .B(n511), .Z(G1338GAT) );
  NOR2_X1 U582 ( .A1(n529), .A2(n512), .ZN(n514) );
  XNOR2_X1 U583 ( .A(KEYINPUT44), .B(KEYINPUT118), .ZN(n513) );
  XNOR2_X1 U584 ( .A(n514), .B(n513), .ZN(n515) );
  XOR2_X1 U585 ( .A(G106GAT), .B(n515), .Z(G1339GAT) );
  NOR2_X1 U586 ( .A1(n591), .A2(n551), .ZN(n516) );
  XOR2_X1 U587 ( .A(KEYINPUT45), .B(n516), .Z(n517) );
  NAND2_X1 U588 ( .A1(n518), .A2(n544), .ZN(n526) );
  NOR2_X1 U589 ( .A1(n546), .A2(n544), .ZN(n519) );
  XNOR2_X1 U590 ( .A(n519), .B(KEYINPUT119), .ZN(n520) );
  XNOR2_X1 U591 ( .A(KEYINPUT46), .B(n520), .ZN(n523) );
  AND2_X1 U592 ( .A1(n551), .A2(n521), .ZN(n522) );
  AND2_X1 U593 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U594 ( .A(n524), .B(KEYINPUT47), .ZN(n525) );
  NAND2_X1 U595 ( .A1(n526), .A2(n525), .ZN(n527) );
  XOR2_X1 U596 ( .A(KEYINPUT48), .B(n527), .Z(n557) );
  NOR2_X1 U597 ( .A1(n557), .A2(n528), .ZN(n543) );
  NAND2_X1 U598 ( .A1(n529), .A2(n543), .ZN(n530) );
  NOR2_X1 U599 ( .A1(n565), .A2(n530), .ZN(n539) );
  NAND2_X1 U600 ( .A1(n539), .A2(n580), .ZN(n531) );
  XNOR2_X1 U601 ( .A(G113GAT), .B(n531), .ZN(G1340GAT) );
  XOR2_X1 U602 ( .A(KEYINPUT120), .B(KEYINPUT49), .Z(n533) );
  NAND2_X1 U603 ( .A1(n539), .A2(n567), .ZN(n532) );
  XNOR2_X1 U604 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U605 ( .A(G120GAT), .B(n534), .ZN(G1341GAT) );
  XOR2_X1 U606 ( .A(KEYINPUT50), .B(KEYINPUT121), .Z(n536) );
  NAND2_X1 U607 ( .A1(n539), .A2(n587), .ZN(n535) );
  XNOR2_X1 U608 ( .A(n536), .B(n535), .ZN(n537) );
  XNOR2_X1 U609 ( .A(G127GAT), .B(n537), .ZN(G1342GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT122), .B(KEYINPUT51), .Z(n541) );
  NAND2_X1 U611 ( .A1(n539), .A2(n472), .ZN(n540) );
  XNOR2_X1 U612 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U613 ( .A(G134GAT), .B(n542), .ZN(G1343GAT) );
  NAND2_X1 U614 ( .A1(n543), .A2(n577), .ZN(n553) );
  NOR2_X1 U615 ( .A1(n544), .A2(n553), .ZN(n545) );
  XOR2_X1 U616 ( .A(G141GAT), .B(n545), .Z(G1344GAT) );
  NOR2_X1 U617 ( .A1(n553), .A2(n546), .ZN(n550) );
  XOR2_X1 U618 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n548) );
  XNOR2_X1 U619 ( .A(G148GAT), .B(KEYINPUT123), .ZN(n547) );
  XNOR2_X1 U620 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U621 ( .A(n550), .B(n549), .ZN(G1345GAT) );
  NOR2_X1 U622 ( .A1(n551), .A2(n553), .ZN(n552) );
  XOR2_X1 U623 ( .A(G155GAT), .B(n552), .Z(G1346GAT) );
  NOR2_X1 U624 ( .A1(n521), .A2(n553), .ZN(n554) );
  XOR2_X1 U625 ( .A(KEYINPUT124), .B(n554), .Z(n555) );
  XNOR2_X1 U626 ( .A(G162GAT), .B(n555), .ZN(G1347GAT) );
  OR2_X1 U627 ( .A1(n557), .A2(n556), .ZN(n559) );
  NAND2_X1 U628 ( .A1(n561), .A2(n560), .ZN(n578) );
  NOR2_X1 U629 ( .A1(n562), .A2(n578), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n563), .B(KEYINPUT55), .ZN(n564) );
  NAND2_X1 U631 ( .A1(n573), .A2(n580), .ZN(n566) );
  XNOR2_X1 U632 ( .A(G169GAT), .B(n566), .ZN(G1348GAT) );
  XNOR2_X1 U633 ( .A(KEYINPUT126), .B(KEYINPUT57), .ZN(n571) );
  NAND2_X1 U634 ( .A1(n573), .A2(n567), .ZN(n569) );
  XOR2_X1 U635 ( .A(G176GAT), .B(KEYINPUT56), .Z(n568) );
  XNOR2_X1 U636 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(G1349GAT) );
  NAND2_X1 U638 ( .A1(n587), .A2(n573), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n572), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U640 ( .A1(n573), .A2(n472), .ZN(n575) );
  XOR2_X1 U641 ( .A(KEYINPUT58), .B(KEYINPUT127), .Z(n574) );
  XNOR2_X1 U642 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n576), .B(G190GAT), .ZN(G1351GAT) );
  XOR2_X1 U644 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n582) );
  INV_X1 U645 ( .A(n577), .ZN(n579) );
  NAND2_X1 U646 ( .A1(n589), .A2(n580), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U648 ( .A(G197GAT), .B(n583), .ZN(G1352GAT) );
  XOR2_X1 U649 ( .A(G204GAT), .B(KEYINPUT61), .Z(n586) );
  NAND2_X1 U650 ( .A1(n589), .A2(n584), .ZN(n585) );
  XNOR2_X1 U651 ( .A(n586), .B(n585), .ZN(G1353GAT) );
  NAND2_X1 U652 ( .A1(n587), .A2(n589), .ZN(n588) );
  XNOR2_X1 U653 ( .A(n588), .B(G211GAT), .ZN(G1354GAT) );
  INV_X1 U654 ( .A(n589), .ZN(n590) );
  NOR2_X1 U655 ( .A1(n591), .A2(n590), .ZN(n592) );
  XOR2_X1 U656 ( .A(KEYINPUT62), .B(n592), .Z(n593) );
  XNOR2_X1 U657 ( .A(G218GAT), .B(n593), .ZN(G1355GAT) );
endmodule

