//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 1 0 0 0 0 1 0 1 1 1 0 0 0 1 0 0 1 0 1 0 0 0 0 1 1 0 1 0 1 0 1 0 1 0 0 0 0 0 0 1 1 1 1 0 1 1 1 0 1 1 0 0 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:24 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n449, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n546, new_n547, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n604, new_n605, new_n608, new_n609, new_n611, new_n612,
    new_n613, new_n615, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1201;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT64), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT65), .B(G2066), .ZN(G384));
  XNOR2_X1  g008(.A(KEYINPUT66), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT67), .B(G69), .Z(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  OR4_X1    g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n454), .A2(new_n455), .ZN(G325));
  XOR2_X1   g031(.A(G325), .B(KEYINPUT68), .Z(G261));
  AOI22_X1  g032(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  NAND3_X1  g034(.A1(new_n459), .A2(G101), .A3(G2104), .ZN(new_n460));
  OR2_X1    g035(.A1(new_n460), .A2(KEYINPUT69), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(KEYINPUT69), .ZN(new_n462));
  OR2_X1    g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(G2105), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  AOI22_X1  g040(.A1(new_n461), .A2(new_n462), .B1(new_n465), .B2(G137), .ZN(new_n466));
  INV_X1    g041(.A(new_n466), .ZN(new_n467));
  XNOR2_X1  g042(.A(KEYINPUT3), .B(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G125), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n459), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n467), .A2(new_n471), .ZN(G160));
  NAND2_X1  g047(.A1(new_n468), .A2(G2105), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G124), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n465), .A2(G136), .ZN(new_n476));
  OR2_X1    g051(.A1(G100), .A2(G2105), .ZN(new_n477));
  OAI211_X1 g052(.A(new_n477), .B(G2104), .C1(G112), .C2(new_n459), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n475), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G162));
  NAND2_X1  g055(.A1(G126), .A2(G2105), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n481), .B1(new_n463), .B2(new_n464), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n459), .A2(G114), .ZN(new_n483));
  OAI21_X1  g058(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  OAI21_X1  g060(.A(KEYINPUT70), .B1(new_n482), .B2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n481), .ZN(new_n487));
  AND2_X1   g062(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n488));
  NOR2_X1   g063(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(G102), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(new_n459), .ZN(new_n492));
  INV_X1    g067(.A(G114), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(G2105), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n492), .A2(new_n494), .A3(G2104), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT70), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n490), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  OAI211_X1 g072(.A(G138), .B(new_n459), .C1(new_n488), .C2(new_n489), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT4), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n468), .A2(new_n500), .A3(G138), .A4(new_n459), .ZN(new_n501));
  AOI22_X1  g076(.A1(new_n486), .A2(new_n497), .B1(new_n499), .B2(new_n501), .ZN(G164));
  INV_X1    g077(.A(G651), .ZN(new_n503));
  NAND2_X1  g078(.A1(G75), .A2(G543), .ZN(new_n504));
  XOR2_X1   g079(.A(new_n504), .B(KEYINPUT71), .Z(new_n505));
  XNOR2_X1  g080(.A(KEYINPUT5), .B(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(G62), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n503), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  XNOR2_X1  g083(.A(KEYINPUT6), .B(G651), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G88), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n509), .A2(G543), .ZN(new_n512));
  INV_X1    g087(.A(G50), .ZN(new_n513));
  OAI22_X1  g088(.A1(new_n510), .A2(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  OR2_X1    g089(.A1(new_n508), .A2(new_n514), .ZN(G303));
  INV_X1    g090(.A(G303), .ZN(G166));
  NAND3_X1  g091(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n517));
  XNOR2_X1  g092(.A(new_n517), .B(KEYINPUT7), .ZN(new_n518));
  INV_X1    g093(.A(G51), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n518), .B1(new_n512), .B2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(new_n506), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n509), .A2(G89), .ZN(new_n522));
  NAND2_X1  g097(.A1(G63), .A2(G651), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n520), .A2(new_n524), .ZN(G168));
  AOI22_X1  g100(.A1(new_n506), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n526));
  OR2_X1    g101(.A1(new_n526), .A2(new_n503), .ZN(new_n527));
  OR2_X1    g102(.A1(new_n527), .A2(KEYINPUT72), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n527), .A2(KEYINPUT72), .ZN(new_n529));
  INV_X1    g104(.A(new_n510), .ZN(new_n530));
  AND2_X1   g105(.A1(new_n509), .A2(G543), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n530), .A2(G90), .B1(new_n531), .B2(G52), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n528), .A2(new_n529), .A3(new_n532), .ZN(G301));
  INV_X1    g108(.A(G301), .ZN(G171));
  NAND2_X1  g109(.A1(new_n506), .A2(G56), .ZN(new_n535));
  NAND2_X1  g110(.A1(G68), .A2(G543), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G651), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(KEYINPUT73), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT73), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n537), .A2(new_n540), .A3(G651), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n530), .A2(G81), .B1(new_n531), .B2(G43), .ZN(new_n542));
  AND3_X1   g117(.A1(new_n539), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G860), .ZN(G153));
  NAND4_X1  g119(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g120(.A1(G1), .A2(G3), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT8), .ZN(new_n547));
  NAND4_X1  g122(.A1(G319), .A2(G483), .A3(G661), .A4(new_n547), .ZN(G188));
  INV_X1    g123(.A(KEYINPUT75), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n510), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n506), .A2(new_n509), .A3(KEYINPUT75), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G91), .ZN(new_n554));
  NAND2_X1  g129(.A1(KEYINPUT74), .A2(G53), .ZN(new_n555));
  OR3_X1    g130(.A1(new_n512), .A2(KEYINPUT9), .A3(new_n555), .ZN(new_n556));
  OAI21_X1  g131(.A(KEYINPUT9), .B1(new_n512), .B2(new_n555), .ZN(new_n557));
  NAND2_X1  g132(.A1(G78), .A2(G543), .ZN(new_n558));
  INV_X1    g133(.A(G65), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n558), .B1(new_n521), .B2(new_n559), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n556), .A2(new_n557), .B1(G651), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n554), .A2(new_n561), .ZN(G299));
  INV_X1    g137(.A(G168), .ZN(G286));
  INV_X1    g138(.A(G87), .ZN(new_n564));
  OAI21_X1  g139(.A(KEYINPUT76), .B1(new_n552), .B2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT76), .ZN(new_n566));
  NAND4_X1  g141(.A1(new_n550), .A2(new_n566), .A3(G87), .A4(new_n551), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  OR2_X1    g143(.A1(new_n506), .A2(G74), .ZN(new_n569));
  AOI22_X1  g144(.A1(G651), .A2(new_n569), .B1(new_n531), .B2(G49), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n568), .A2(new_n570), .ZN(G288));
  INV_X1    g146(.A(G48), .ZN(new_n572));
  OAI21_X1  g147(.A(KEYINPUT77), .B1(new_n512), .B2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT77), .ZN(new_n574));
  NAND4_X1  g149(.A1(new_n509), .A2(new_n574), .A3(G48), .A4(G543), .ZN(new_n575));
  NAND2_X1  g150(.A1(G73), .A2(G543), .ZN(new_n576));
  INV_X1    g151(.A(G61), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n576), .B1(new_n521), .B2(new_n577), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n573), .A2(new_n575), .B1(new_n578), .B2(G651), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n550), .A2(G86), .A3(new_n551), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(G305));
  INV_X1    g156(.A(G85), .ZN(new_n582));
  INV_X1    g157(.A(G47), .ZN(new_n583));
  OAI22_X1  g158(.A1(new_n510), .A2(new_n582), .B1(new_n512), .B2(new_n583), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n506), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n585), .A2(new_n503), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(G290));
  NAND2_X1  g163(.A1(G301), .A2(G868), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n589), .A2(KEYINPUT78), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n553), .A2(G92), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT10), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n591), .B(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(G79), .A2(G543), .ZN(new_n594));
  INV_X1    g169(.A(G66), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n521), .B2(new_n595), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n596), .A2(G651), .B1(new_n531), .B2(G54), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(G868), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AND2_X1   g175(.A1(new_n589), .A2(KEYINPUT78), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n590), .B1(new_n600), .B2(new_n601), .ZN(G284));
  AOI21_X1  g177(.A(new_n590), .B1(new_n600), .B2(new_n601), .ZN(G321));
  NAND2_X1  g178(.A1(G286), .A2(G868), .ZN(new_n604));
  INV_X1    g179(.A(G299), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n605), .B2(G868), .ZN(G297));
  OAI21_X1  g181(.A(new_n604), .B1(new_n605), .B2(G868), .ZN(G280));
  INV_X1    g182(.A(new_n598), .ZN(new_n608));
  INV_X1    g183(.A(G559), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n609), .B2(G860), .ZN(G148));
  NOR2_X1   g185(.A1(new_n598), .A2(G559), .ZN(new_n611));
  INV_X1    g186(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(G868), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n613), .B1(G868), .B2(new_n543), .ZN(G323));
  XOR2_X1   g189(.A(KEYINPUT79), .B(KEYINPUT11), .Z(new_n615));
  XNOR2_X1  g190(.A(G323), .B(new_n615), .ZN(G282));
  AND2_X1   g191(.A1(new_n459), .A2(G2104), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n468), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT12), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT13), .ZN(new_n620));
  INV_X1    g195(.A(G2100), .ZN(new_n621));
  OR2_X1    g196(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  AOI22_X1  g197(.A1(new_n474), .A2(G123), .B1(G135), .B2(new_n465), .ZN(new_n623));
  NOR3_X1   g198(.A1(new_n459), .A2(KEYINPUT80), .A3(G111), .ZN(new_n624));
  OAI21_X1  g199(.A(KEYINPUT80), .B1(new_n459), .B2(G111), .ZN(new_n625));
  OAI211_X1 g200(.A(new_n625), .B(G2104), .C1(G99), .C2(G2105), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n623), .B1(new_n624), .B2(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(G2096), .Z(new_n628));
  NAND2_X1  g203(.A1(new_n620), .A2(new_n621), .ZN(new_n629));
  NAND3_X1  g204(.A1(new_n622), .A2(new_n628), .A3(new_n629), .ZN(G156));
  XNOR2_X1  g205(.A(G2427), .B(G2438), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2430), .ZN(new_n632));
  XNOR2_X1  g207(.A(KEYINPUT15), .B(G2435), .ZN(new_n633));
  OR2_X1    g208(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n632), .A2(new_n633), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n634), .A2(KEYINPUT14), .A3(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(G1341), .B(G1348), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n636), .B(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(G2451), .B(G2454), .Z(new_n641));
  XNOR2_X1  g216(.A(G2443), .B(G2446), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n644), .A2(G14), .ZN(new_n645));
  NOR2_X1   g220(.A1(new_n640), .A2(new_n643), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(G401));
  INV_X1    g223(.A(KEYINPUT18), .ZN(new_n649));
  XOR2_X1   g224(.A(G2084), .B(G2090), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT82), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2067), .B(G2678), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n653), .A2(KEYINPUT17), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n651), .A2(new_n652), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n649), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(new_n621), .ZN(new_n657));
  XOR2_X1   g232(.A(G2072), .B(G2078), .Z(new_n658));
  AOI21_X1  g233(.A(new_n658), .B1(new_n653), .B2(KEYINPUT18), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n659), .B(G2096), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n657), .B(new_n660), .ZN(G227));
  XNOR2_X1  g236(.A(G1956), .B(G2474), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1961), .B(G1966), .ZN(new_n663));
  OR2_X1    g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g239(.A(KEYINPUT83), .ZN(new_n665));
  OR2_X1    g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(G1971), .B(G1976), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT19), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n664), .A2(new_n665), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n666), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT20), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n662), .A2(new_n663), .ZN(new_n672));
  OAI21_X1  g247(.A(new_n672), .B1(new_n668), .B2(new_n664), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n668), .A2(KEYINPUT84), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT85), .ZN(new_n677));
  AND3_X1   g252(.A1(new_n671), .A2(new_n675), .A3(new_n677), .ZN(new_n678));
  AOI21_X1  g253(.A(new_n677), .B1(new_n671), .B2(new_n675), .ZN(new_n679));
  XOR2_X1   g254(.A(G1991), .B(G1996), .Z(new_n680));
  OR3_X1    g255(.A1(new_n678), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  OAI21_X1  g256(.A(new_n680), .B1(new_n678), .B2(new_n679), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1981), .B(G1986), .ZN(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n681), .A2(new_n684), .A3(new_n682), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n686), .A2(new_n687), .ZN(G229));
  NAND3_X1  g263(.A1(new_n459), .A2(G103), .A3(G2104), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT25), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n468), .A2(G127), .ZN(new_n691));
  NAND2_X1  g266(.A1(G115), .A2(G2104), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n459), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  AOI211_X1 g268(.A(new_n690), .B(new_n693), .C1(G139), .C2(new_n465), .ZN(new_n694));
  INV_X1    g269(.A(G29), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(new_n695), .B2(G33), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n697), .A2(new_n442), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT94), .ZN(new_n699));
  NAND2_X1  g274(.A1(G171), .A2(G16), .ZN(new_n700));
  NOR2_X1   g275(.A1(G5), .A2(G16), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT96), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n699), .B1(G1961), .B2(new_n704), .ZN(new_n705));
  NOR2_X1   g280(.A1(G16), .A2(G19), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n706), .B1(new_n543), .B2(G16), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n707), .A2(G1341), .ZN(new_n708));
  INV_X1    g283(.A(G1961), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n708), .B1(new_n703), .B2(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n695), .A2(G26), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT28), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n474), .A2(G128), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n465), .A2(G140), .ZN(new_n714));
  OR2_X1    g289(.A1(G104), .A2(G2105), .ZN(new_n715));
  OAI211_X1 g290(.A(new_n715), .B(G2104), .C1(G116), .C2(new_n459), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n713), .A2(new_n714), .A3(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(new_n717), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n712), .B1(new_n718), .B2(new_n695), .ZN(new_n719));
  XNOR2_X1  g294(.A(KEYINPUT93), .B(G2067), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n695), .A2(G27), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(G164), .B2(new_n695), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(G2078), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n721), .A2(new_n724), .ZN(new_n725));
  XOR2_X1   g300(.A(KEYINPUT31), .B(G11), .Z(new_n726));
  INV_X1    g301(.A(G28), .ZN(new_n727));
  OR2_X1    g302(.A1(new_n727), .A2(KEYINPUT30), .ZN(new_n728));
  AOI21_X1  g303(.A(G29), .B1(new_n727), .B2(KEYINPUT30), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n726), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(new_n627), .B2(new_n695), .ZN(new_n731));
  INV_X1    g306(.A(G16), .ZN(new_n732));
  NOR2_X1   g307(.A1(G168), .A2(new_n732), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(new_n732), .B2(G21), .ZN(new_n734));
  INV_X1    g309(.A(G1966), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n731), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(KEYINPUT24), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n695), .B1(new_n737), .B2(G34), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(new_n737), .B2(G34), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(G160), .B2(G29), .ZN(new_n740));
  NAND3_X1  g315(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n741));
  XOR2_X1   g316(.A(new_n741), .B(KEYINPUT26), .Z(new_n742));
  INV_X1    g317(.A(G129), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n742), .B1(new_n473), .B2(new_n743), .ZN(new_n744));
  AOI22_X1  g319(.A1(new_n465), .A2(G141), .B1(G105), .B2(new_n617), .ZN(new_n745));
  INV_X1    g320(.A(new_n745), .ZN(new_n746));
  OR2_X1    g321(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n748), .A2(new_n695), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(new_n695), .B2(G32), .ZN(new_n750));
  XNOR2_X1  g325(.A(KEYINPUT27), .B(G1996), .ZN(new_n751));
  OAI221_X1 g326(.A(new_n736), .B1(G2084), .B2(new_n740), .C1(new_n750), .C2(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n740), .A2(G2084), .ZN(new_n753));
  OAI221_X1 g328(.A(new_n753), .B1(new_n735), .B2(new_n734), .C1(new_n697), .C2(new_n442), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  NAND4_X1  g330(.A1(new_n705), .A2(new_n710), .A3(new_n725), .A4(new_n755), .ZN(new_n756));
  NOR2_X1   g331(.A1(G162), .A2(new_n695), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(new_n695), .B2(G35), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT29), .ZN(new_n759));
  INV_X1    g334(.A(G2090), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT97), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n750), .A2(new_n751), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT95), .ZN(new_n764));
  INV_X1    g339(.A(new_n759), .ZN(new_n765));
  AOI22_X1  g340(.A1(new_n765), .A2(G2090), .B1(G1341), .B2(new_n707), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n762), .A2(new_n764), .A3(new_n766), .ZN(new_n767));
  NOR2_X1   g342(.A1(G4), .A2(G16), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(new_n608), .B2(G16), .ZN(new_n769));
  XNOR2_X1  g344(.A(KEYINPUT92), .B(G1348), .ZN(new_n770));
  NOR2_X1   g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n769), .A2(new_n770), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n732), .A2(G20), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(KEYINPUT23), .Z(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(G299), .B2(G16), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(G1956), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n772), .A2(new_n776), .ZN(new_n777));
  NOR4_X1   g352(.A1(new_n756), .A2(new_n767), .A3(new_n771), .A4(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n695), .A2(G25), .ZN(new_n779));
  OR2_X1    g354(.A1(G95), .A2(G2105), .ZN(new_n780));
  OAI211_X1 g355(.A(new_n780), .B(G2104), .C1(G107), .C2(new_n459), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT86), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n465), .A2(G131), .ZN(new_n783));
  INV_X1    g358(.A(G119), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n783), .B1(new_n784), .B2(new_n473), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n782), .A2(new_n785), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n779), .B1(new_n786), .B2(new_n695), .ZN(new_n787));
  XOR2_X1   g362(.A(KEYINPUT35), .B(G1991), .Z(new_n788));
  XOR2_X1   g363(.A(new_n787), .B(new_n788), .Z(new_n789));
  NOR2_X1   g364(.A1(G16), .A2(G24), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(new_n587), .B2(G16), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT88), .ZN(new_n792));
  XOR2_X1   g367(.A(KEYINPUT87), .B(G1986), .Z(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  AOI211_X1 g369(.A(new_n789), .B(new_n794), .C1(KEYINPUT91), .C2(KEYINPUT36), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n732), .A2(G22), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(G166), .B2(new_n732), .ZN(new_n797));
  XOR2_X1   g372(.A(new_n797), .B(G1971), .Z(new_n798));
  AND2_X1   g373(.A1(new_n732), .A2(G6), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n799), .B1(G305), .B2(G16), .ZN(new_n800));
  XNOR2_X1  g375(.A(KEYINPUT32), .B(G1981), .ZN(new_n801));
  INV_X1    g376(.A(new_n801), .ZN(new_n802));
  OR2_X1    g377(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n800), .A2(new_n802), .ZN(new_n804));
  NAND3_X1  g379(.A1(new_n798), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  NOR2_X1   g380(.A1(G16), .A2(G23), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT89), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(G288), .B2(new_n732), .ZN(new_n808));
  XOR2_X1   g383(.A(KEYINPUT33), .B(G1976), .Z(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT90), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n808), .B(new_n810), .ZN(new_n811));
  OAI21_X1  g386(.A(KEYINPUT34), .B1(new_n805), .B2(new_n811), .ZN(new_n812));
  OR3_X1    g387(.A1(new_n805), .A2(KEYINPUT34), .A3(new_n811), .ZN(new_n813));
  AND3_X1   g388(.A1(new_n795), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  OR2_X1    g389(.A1(KEYINPUT91), .A2(KEYINPUT36), .ZN(new_n815));
  OR2_X1    g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n814), .A2(new_n815), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n778), .A2(new_n816), .A3(new_n817), .ZN(G150));
  INV_X1    g393(.A(G150), .ZN(G311));
  XNOR2_X1  g394(.A(KEYINPUT100), .B(G860), .ZN(new_n820));
  INV_X1    g395(.A(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(G93), .ZN(new_n822));
  INV_X1    g397(.A(G55), .ZN(new_n823));
  OAI22_X1  g398(.A1(new_n510), .A2(new_n822), .B1(new_n512), .B2(new_n823), .ZN(new_n824));
  AND2_X1   g399(.A1(new_n824), .A2(KEYINPUT98), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n824), .A2(KEYINPUT98), .ZN(new_n826));
  AOI22_X1  g401(.A1(new_n506), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n827));
  OAI22_X1  g402(.A1(new_n825), .A2(new_n826), .B1(new_n503), .B2(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT99), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n543), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n830), .B1(new_n829), .B2(new_n828), .ZN(new_n831));
  INV_X1    g406(.A(new_n828), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n832), .A2(KEYINPUT99), .A3(new_n543), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT38), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n608), .A2(G559), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n835), .B(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT39), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n821), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n839), .B1(new_n838), .B2(new_n837), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n828), .A2(new_n821), .ZN(new_n841));
  XOR2_X1   g416(.A(new_n841), .B(KEYINPUT37), .Z(new_n842));
  NAND2_X1  g417(.A1(new_n840), .A2(new_n842), .ZN(G145));
  XNOR2_X1  g418(.A(new_n786), .B(new_n619), .ZN(new_n844));
  OR2_X1    g419(.A1(G106), .A2(G2105), .ZN(new_n845));
  OAI211_X1 g420(.A(new_n845), .B(G2104), .C1(G118), .C2(new_n459), .ZN(new_n846));
  INV_X1    g421(.A(G130), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n846), .B1(new_n473), .B2(new_n847), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n848), .B1(G142), .B2(new_n465), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n844), .B(new_n849), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n850), .B(KEYINPUT102), .Z(new_n851));
  OAI21_X1  g426(.A(KEYINPUT101), .B1(new_n482), .B2(new_n485), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT101), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n490), .A2(new_n495), .A3(new_n853), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n500), .B1(new_n465), .B2(G138), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n498), .A2(KEYINPUT4), .ZN(new_n856));
  OAI211_X1 g431(.A(new_n852), .B(new_n854), .C1(new_n855), .C2(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n717), .B(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(new_n748), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(new_n694), .ZN(new_n860));
  OR2_X1    g435(.A1(new_n851), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n627), .B(new_n479), .ZN(new_n862));
  XOR2_X1   g437(.A(new_n862), .B(G160), .Z(new_n863));
  AOI21_X1  g438(.A(new_n863), .B1(new_n860), .B2(new_n850), .ZN(new_n864));
  AOI21_X1  g439(.A(G37), .B1(new_n861), .B2(new_n864), .ZN(new_n865));
  AND2_X1   g440(.A1(new_n851), .A2(new_n860), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n851), .A2(new_n860), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n863), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n865), .A2(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g445(.A1(new_n612), .A2(new_n834), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n611), .A2(new_n833), .A3(new_n831), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n598), .A2(G299), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n593), .A2(new_n605), .A3(new_n597), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n873), .A2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT41), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n874), .A2(new_n879), .A3(new_n875), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n879), .B1(new_n874), .B2(new_n875), .ZN(new_n882));
  OAI211_X1 g457(.A(new_n872), .B(new_n871), .C1(new_n881), .C2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n878), .A2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT104), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n884), .A2(new_n885), .A3(KEYINPUT42), .ZN(new_n886));
  XNOR2_X1  g461(.A(G166), .B(G305), .ZN(new_n887));
  INV_X1    g462(.A(new_n570), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n888), .B1(new_n565), .B2(new_n567), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(G290), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT103), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n887), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n890), .A2(new_n891), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n892), .B(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT42), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n895), .B1(KEYINPUT104), .B2(new_n896), .ZN(new_n897));
  OAI211_X1 g472(.A(new_n878), .B(new_n883), .C1(KEYINPUT104), .C2(new_n896), .ZN(new_n898));
  AND3_X1   g473(.A1(new_n886), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n897), .B1(new_n886), .B2(new_n898), .ZN(new_n900));
  OAI21_X1  g475(.A(G868), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n901), .B1(G868), .B2(new_n832), .ZN(G295));
  OAI21_X1  g477(.A(new_n901), .B1(G868), .B2(new_n832), .ZN(G331));
  XNOR2_X1  g478(.A(G301), .B(G168), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n904), .A2(new_n831), .A3(new_n833), .ZN(new_n905));
  INV_X1    g480(.A(new_n904), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n834), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n877), .A2(new_n905), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n905), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT106), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n909), .B1(new_n910), .B2(new_n880), .ZN(new_n911));
  INV_X1    g486(.A(new_n875), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n605), .B1(new_n593), .B2(new_n597), .ZN(new_n913));
  OAI21_X1  g488(.A(KEYINPUT41), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n914), .A2(new_n910), .A3(new_n880), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n908), .B1(new_n911), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(new_n895), .ZN(new_n918));
  INV_X1    g493(.A(G37), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n909), .B1(new_n881), .B2(new_n882), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n920), .A2(new_n894), .A3(new_n908), .ZN(new_n921));
  XNOR2_X1  g496(.A(KEYINPUT105), .B(KEYINPUT43), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n918), .A2(new_n919), .A3(new_n921), .A4(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(new_n908), .ZN(new_n924));
  AOI22_X1  g499(.A1(new_n880), .A2(new_n914), .B1(new_n907), .B2(new_n905), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n895), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n926), .A2(new_n921), .A3(new_n919), .ZN(new_n927));
  INV_X1    g502(.A(new_n922), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT44), .ZN(new_n930));
  AND3_X1   g505(.A1(new_n923), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n921), .A2(new_n919), .ZN(new_n932));
  OAI211_X1 g507(.A(new_n915), .B(new_n909), .C1(new_n910), .C2(new_n880), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n894), .B1(new_n933), .B2(new_n908), .ZN(new_n934));
  OAI21_X1  g509(.A(KEYINPUT43), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n926), .A2(new_n921), .A3(new_n919), .A4(new_n922), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n930), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n931), .A2(new_n937), .ZN(G397));
  AND3_X1   g513(.A1(new_n490), .A2(new_n495), .A3(new_n853), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n853), .B1(new_n490), .B2(new_n495), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n499), .A2(new_n501), .ZN(new_n942));
  AOI21_X1  g517(.A(G1384), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  AND2_X1   g518(.A1(new_n469), .A2(new_n470), .ZN(new_n944));
  OAI211_X1 g519(.A(new_n466), .B(G40), .C1(new_n944), .C2(new_n459), .ZN(new_n945));
  NOR3_X1   g520(.A1(new_n943), .A2(KEYINPUT45), .A3(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(G1996), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n747), .B(new_n947), .ZN(new_n948));
  XOR2_X1   g523(.A(new_n717), .B(G2067), .Z(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  XNOR2_X1  g525(.A(new_n786), .B(new_n788), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n946), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(new_n946), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n587), .B(G1986), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n952), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n955), .B(KEYINPUT107), .ZN(new_n956));
  INV_X1    g531(.A(G1976), .ZN(new_n957));
  NAND2_X1  g532(.A1(G288), .A2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(G1384), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n857), .A2(new_n959), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n960), .A2(new_n945), .ZN(new_n961));
  INV_X1    g536(.A(G8), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT52), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n889), .A2(G1976), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n958), .A2(new_n963), .A3(new_n964), .A4(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n573), .A2(new_n575), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n578), .A2(G651), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n530), .A2(G86), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n967), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(G1981), .ZN(new_n971));
  INV_X1    g546(.A(G1981), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n579), .A2(new_n972), .A3(new_n580), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT114), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n975), .A2(KEYINPUT49), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  OAI211_X1 g552(.A(new_n971), .B(new_n973), .C1(new_n975), .C2(KEYINPUT49), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n977), .A2(new_n963), .A3(new_n978), .ZN(new_n979));
  AOI211_X1 g554(.A(new_n957), .B(new_n888), .C1(new_n565), .C2(new_n567), .ZN(new_n980));
  INV_X1    g555(.A(new_n945), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(new_n943), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(G8), .ZN(new_n983));
  OAI21_X1  g558(.A(KEYINPUT52), .B1(new_n980), .B2(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n966), .A2(new_n979), .A3(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT115), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n966), .A2(new_n979), .A3(new_n984), .A4(KEYINPUT115), .ZN(new_n988));
  AND2_X1   g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  XNOR2_X1  g564(.A(KEYINPUT110), .B(G1971), .ZN(new_n990));
  INV_X1    g565(.A(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT109), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT45), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n993), .A2(G1384), .ZN(new_n994));
  AND3_X1   g569(.A1(new_n857), .A2(new_n992), .A3(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n992), .B1(new_n857), .B2(new_n994), .ZN(new_n996));
  NOR3_X1   g571(.A1(new_n482), .A2(new_n485), .A3(KEYINPUT70), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n496), .B1(new_n490), .B2(new_n495), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n942), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(KEYINPUT45), .B1(new_n999), .B2(new_n959), .ZN(new_n1000));
  OAI22_X1  g575(.A1(new_n995), .A2(new_n996), .B1(new_n1000), .B2(KEYINPUT108), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n993), .B1(G164), .B2(G1384), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT108), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n981), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n991), .B1(new_n1001), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT111), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT112), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1008), .B1(new_n960), .B2(KEYINPUT50), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT50), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n857), .A2(KEYINPUT112), .A3(new_n1010), .A4(new_n959), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n999), .A2(new_n959), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n945), .B1(new_n1013), .B2(KEYINPUT50), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1012), .A2(new_n760), .A3(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT113), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n945), .B1(new_n1000), .B2(KEYINPUT108), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n857), .A2(new_n994), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(KEYINPUT109), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n857), .A2(new_n992), .A3(new_n994), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1018), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1024), .A2(KEYINPUT111), .A3(new_n991), .ZN(new_n1025));
  NOR2_X1   g600(.A1(G164), .A2(G1384), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n981), .B1(new_n1026), .B2(new_n1010), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1027), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1028), .A2(KEYINPUT113), .A3(new_n760), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1007), .A2(new_n1017), .A3(new_n1025), .A4(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(G303), .A2(G8), .ZN(new_n1031));
  XNOR2_X1  g606(.A(new_n1031), .B(KEYINPUT55), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1030), .A2(G8), .A3(new_n1033), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n979), .A2(new_n957), .A3(new_n889), .ZN(new_n1035));
  AND2_X1   g610(.A1(new_n1035), .A2(new_n973), .ZN(new_n1036));
  OAI22_X1  g611(.A1(new_n989), .A2(new_n1034), .B1(new_n983), .B2(new_n1036), .ZN(new_n1037));
  AOI22_X1  g612(.A1(new_n1020), .A2(new_n1021), .B1(new_n1003), .B2(new_n1002), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n990), .B1(new_n1038), .B2(new_n1018), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n960), .A2(KEYINPUT50), .ZN(new_n1040));
  OAI211_X1 g615(.A(new_n1040), .B(new_n981), .C1(KEYINPUT50), .C2(new_n1013), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1041), .A2(G2090), .ZN(new_n1042));
  OAI21_X1  g617(.A(G8), .B1(new_n1039), .B2(new_n1042), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n985), .B1(new_n1032), .B2(new_n1043), .ZN(new_n1044));
  XOR2_X1   g619(.A(KEYINPUT117), .B(G2084), .Z(new_n1045));
  AOI21_X1  g620(.A(KEYINPUT112), .B1(new_n943), .B2(new_n1010), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1011), .ZN(new_n1047));
  OAI211_X1 g622(.A(new_n1014), .B(new_n1045), .C1(new_n1046), .C2(new_n1047), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n981), .B1(new_n943), .B2(KEYINPUT45), .ZN(new_n1049));
  INV_X1    g624(.A(new_n994), .ZN(new_n1050));
  OAI21_X1  g625(.A(KEYINPUT116), .B1(G164), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT116), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n999), .A2(new_n1052), .A3(new_n994), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n735), .B1(new_n1049), .B2(new_n1054), .ZN(new_n1055));
  AOI211_X1 g630(.A(new_n962), .B(G286), .C1(new_n1048), .C2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1034), .A2(new_n1044), .A3(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT63), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1030), .A2(G8), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(new_n1032), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n987), .A2(new_n988), .ZN(new_n1062));
  AND2_X1   g637(.A1(new_n1056), .A2(KEYINPUT63), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1061), .A2(new_n1034), .A3(new_n1062), .A4(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1037), .B1(new_n1059), .B2(new_n1064), .ZN(new_n1065));
  NOR2_X1   g640(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT57), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1067), .B1(new_n554), .B2(new_n561), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1066), .A2(new_n1068), .ZN(new_n1069));
  XNOR2_X1  g644(.A(KEYINPUT56), .B(G2072), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1018), .A2(new_n1022), .A3(new_n1023), .A4(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(G1956), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1041), .A2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1069), .B1(new_n1071), .B2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(G1348), .B1(new_n1012), .B2(new_n1014), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n982), .A2(G2067), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1077), .A2(new_n598), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1071), .A2(new_n1073), .A3(new_n1069), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1074), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  AND3_X1   g655(.A1(new_n1071), .A2(new_n1073), .A3(new_n1069), .ZN(new_n1081));
  NOR3_X1   g656(.A1(new_n1081), .A2(new_n1074), .A3(KEYINPUT61), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT61), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1071), .A2(new_n1073), .ZN(new_n1084));
  INV_X1    g659(.A(new_n1069), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1083), .B1(new_n1086), .B2(new_n1079), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1082), .A2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT60), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1089), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1076), .ZN(new_n1091));
  OAI211_X1 g666(.A(KEYINPUT60), .B(new_n1091), .C1(new_n1028), .C2(G1348), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1090), .A2(new_n608), .A3(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1077), .A2(KEYINPUT60), .A3(new_n598), .ZN(new_n1094));
  XOR2_X1   g669(.A(KEYINPUT58), .B(G1341), .Z(new_n1095));
  NAND2_X1  g670(.A1(new_n982), .A2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1096), .B1(new_n1024), .B2(G1996), .ZN(new_n1097));
  AND2_X1   g672(.A1(new_n543), .A2(KEYINPUT118), .ZN(new_n1098));
  XNOR2_X1  g673(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n1099));
  AND3_X1   g674(.A1(new_n1097), .A2(new_n1098), .A3(new_n1099), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1099), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1101));
  OAI211_X1 g676(.A(new_n1093), .B(new_n1094), .C1(new_n1100), .C2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1080), .B1(new_n1088), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT54), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1049), .A2(new_n1054), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT53), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1107), .A2(G2078), .ZN(new_n1108));
  AOI22_X1  g683(.A1(new_n1105), .A2(new_n709), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1038), .A2(new_n443), .A3(new_n1018), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(new_n1107), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1109), .A2(G301), .A3(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT122), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1109), .A2(new_n1111), .A3(KEYINPUT122), .A4(G301), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1104), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  OAI21_X1  g691(.A(KEYINPUT120), .B1(new_n1028), .B2(G1961), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT120), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1105), .A2(new_n1118), .A3(new_n709), .ZN(new_n1119));
  AND2_X1   g694(.A1(new_n1022), .A2(new_n1108), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1049), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1117), .A2(new_n1111), .A3(new_n1119), .A4(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(KEYINPUT123), .ZN(new_n1124));
  AOI22_X1  g699(.A1(new_n1110), .A2(new_n1107), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT123), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1125), .A2(new_n1126), .A3(new_n1117), .A4(new_n1119), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1124), .A2(G171), .A3(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1116), .A2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1048), .A2(new_n1055), .A3(G168), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(G8), .ZN(new_n1131));
  AOI21_X1  g706(.A(G168), .B1(new_n1048), .B2(new_n1055), .ZN(new_n1132));
  OAI21_X1  g707(.A(KEYINPUT51), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT51), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1130), .A2(new_n1134), .A3(G8), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1133), .A2(new_n1135), .ZN(new_n1136));
  AND3_X1   g711(.A1(new_n1136), .A2(new_n1034), .A3(new_n1044), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1103), .A2(new_n1129), .A3(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT121), .ZN(new_n1139));
  AOI21_X1  g714(.A(G301), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1140), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1125), .A2(G301), .A3(new_n1117), .A4(new_n1119), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1139), .B1(new_n1143), .B2(new_n1104), .ZN(new_n1144));
  AOI211_X1 g719(.A(KEYINPUT121), .B(KEYINPUT54), .C1(new_n1141), .C2(new_n1142), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1065), .B1(new_n1138), .B2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT125), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1148), .B1(new_n1136), .B2(KEYINPUT62), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT62), .ZN(new_n1150));
  AOI211_X1 g725(.A(KEYINPUT125), .B(new_n1150), .C1(new_n1133), .C2(new_n1135), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1149), .A2(new_n1151), .ZN(new_n1152));
  AND3_X1   g727(.A1(new_n966), .A2(new_n979), .A3(new_n984), .ZN(new_n1153));
  OR2_X1    g728(.A1(new_n1041), .A2(G2090), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n962), .B1(new_n1154), .B2(new_n1005), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1153), .B1(new_n1155), .B2(new_n1033), .ZN(new_n1156));
  AOI211_X1 g731(.A(new_n1006), .B(new_n990), .C1(new_n1038), .C2(new_n1018), .ZN(new_n1157));
  AOI21_X1  g732(.A(KEYINPUT111), .B1(new_n1024), .B2(new_n991), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g734(.A(KEYINPUT113), .B1(new_n1028), .B2(new_n760), .ZN(new_n1160));
  AND4_X1   g735(.A1(KEYINPUT113), .A2(new_n1012), .A3(new_n760), .A4(new_n1014), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n962), .B1(new_n1159), .B2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1156), .B1(new_n1163), .B2(new_n1033), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT124), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1133), .A2(new_n1150), .A3(new_n1135), .ZN(new_n1166));
  NAND4_X1  g741(.A1(new_n1164), .A2(new_n1165), .A3(new_n1166), .A4(new_n1140), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1034), .A2(new_n1140), .A3(new_n1044), .ZN(new_n1168));
  AND3_X1   g743(.A1(new_n1133), .A2(new_n1150), .A3(new_n1135), .ZN(new_n1169));
  OAI21_X1  g744(.A(KEYINPUT124), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  AND3_X1   g745(.A1(new_n1152), .A2(new_n1167), .A3(new_n1170), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n956), .B1(new_n1147), .B2(new_n1171), .ZN(new_n1172));
  NOR2_X1   g747(.A1(G290), .A2(G1986), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n946), .A2(KEYINPUT48), .A3(new_n1173), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT48), .ZN(new_n1175));
  INV_X1    g750(.A(new_n1173), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1175), .B1(new_n953), .B2(new_n1176), .ZN(new_n1177));
  AND3_X1   g752(.A1(new_n952), .A2(new_n1174), .A3(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n946), .A2(new_n947), .ZN(new_n1179));
  XNOR2_X1  g754(.A(new_n1179), .B(KEYINPUT46), .ZN(new_n1180));
  AND2_X1   g755(.A1(new_n949), .A2(new_n748), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1180), .B1(new_n953), .B2(new_n1181), .ZN(new_n1182));
  XOR2_X1   g757(.A(new_n1182), .B(KEYINPUT47), .Z(new_n1183));
  NAND2_X1  g758(.A1(new_n786), .A2(new_n788), .ZN(new_n1184));
  OAI22_X1  g759(.A1(new_n950), .A2(new_n1184), .B1(G2067), .B2(new_n717), .ZN(new_n1185));
  AOI211_X1 g760(.A(new_n1178), .B(new_n1183), .C1(new_n946), .C2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1172), .A2(new_n1186), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g762(.A(G229), .ZN(new_n1189));
  INV_X1    g763(.A(KEYINPUT127), .ZN(new_n1190));
  OAI21_X1  g764(.A(G319), .B1(new_n645), .B2(new_n646), .ZN(new_n1191));
  NOR2_X1   g765(.A1(G227), .A2(new_n1191), .ZN(new_n1192));
  INV_X1    g766(.A(KEYINPUT126), .ZN(new_n1193));
  NAND2_X1  g767(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  OAI21_X1  g768(.A(KEYINPUT126), .B1(G227), .B2(new_n1191), .ZN(new_n1195));
  NAND2_X1  g769(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  AND3_X1   g770(.A1(new_n1189), .A2(new_n1190), .A3(new_n1196), .ZN(new_n1197));
  AOI21_X1  g771(.A(new_n1190), .B1(new_n1189), .B2(new_n1196), .ZN(new_n1198));
  OAI21_X1  g772(.A(new_n869), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  AOI21_X1  g773(.A(new_n1199), .B1(new_n929), .B2(new_n923), .ZN(G308));
  NAND2_X1  g774(.A1(new_n923), .A2(new_n929), .ZN(new_n1201));
  OAI211_X1 g775(.A(new_n1201), .B(new_n869), .C1(new_n1198), .C2(new_n1197), .ZN(G225));
endmodule


