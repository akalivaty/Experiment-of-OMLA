//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 0 1 0 1 0 1 0 1 1 0 1 1 0 0 1 0 1 0 0 1 1 1 1 0 0 1 1 0 0 0 1 0 0 1 0 0 0 1 1 1 0 0 1 0 0 0 1 0 0 1 1 1 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:51 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n697, new_n698, new_n699, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n756, new_n757, new_n758, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n965, new_n966, new_n967, new_n968, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019;
  INV_X1    g000(.A(KEYINPUT89), .ZN(new_n187));
  XNOR2_X1  g001(.A(G113), .B(G122), .ZN(new_n188));
  INV_X1    g002(.A(G104), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n188), .B(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G237), .ZN(new_n191));
  INV_X1    g005(.A(G953), .ZN(new_n192));
  AND4_X1   g006(.A1(G143), .A2(new_n191), .A3(new_n192), .A4(G214), .ZN(new_n193));
  NOR2_X1   g007(.A1(G237), .A2(G953), .ZN(new_n194));
  AOI21_X1  g008(.A(G143), .B1(new_n194), .B2(G214), .ZN(new_n195));
  OAI21_X1  g009(.A(G131), .B1(new_n193), .B2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT17), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n191), .A2(new_n192), .A3(G214), .ZN(new_n198));
  INV_X1    g012(.A(G143), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G131), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n194), .A2(G143), .A3(G214), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n200), .A2(new_n201), .A3(new_n202), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n196), .A2(new_n197), .A3(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G140), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G125), .ZN(new_n206));
  INV_X1    g020(.A(G125), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G140), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n206), .A2(new_n208), .A3(KEYINPUT16), .ZN(new_n209));
  OR3_X1    g023(.A1(new_n207), .A2(KEYINPUT16), .A3(G140), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G146), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n209), .A2(new_n210), .A3(G146), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n200), .A2(new_n202), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n215), .A2(KEYINPUT17), .A3(G131), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n204), .A2(new_n213), .A3(new_n214), .A4(new_n216), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n193), .A2(new_n195), .ZN(new_n218));
  NAND2_X1  g032(.A1(KEYINPUT18), .A2(G131), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n206), .A2(new_n208), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G146), .ZN(new_n221));
  XNOR2_X1  g035(.A(G125), .B(G140), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(new_n212), .ZN(new_n223));
  AOI22_X1  g037(.A1(new_n218), .A2(new_n219), .B1(new_n221), .B2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(new_n219), .ZN(new_n225));
  AOI21_X1  g039(.A(KEYINPUT86), .B1(new_n215), .B2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT86), .ZN(new_n227));
  AOI211_X1 g041(.A(new_n227), .B(new_n219), .C1(new_n200), .C2(new_n202), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n224), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n190), .B1(new_n217), .B2(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n217), .A2(new_n229), .A3(new_n190), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(KEYINPUT88), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT88), .ZN(new_n233));
  NAND4_X1  g047(.A1(new_n217), .A2(new_n229), .A3(new_n233), .A4(new_n190), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n230), .B1(new_n232), .B2(new_n234), .ZN(new_n235));
  OAI21_X1  g049(.A(G475), .B1(new_n235), .B2(G902), .ZN(new_n236));
  XOR2_X1   g050(.A(KEYINPUT85), .B(KEYINPUT20), .Z(new_n237));
  NAND2_X1  g051(.A1(new_n232), .A2(new_n234), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n196), .A2(new_n203), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT87), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n222), .A2(new_n240), .ZN(new_n241));
  XNOR2_X1  g055(.A(new_n241), .B(KEYINPUT19), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n239), .B1(new_n242), .B2(G146), .ZN(new_n243));
  OR2_X1    g057(.A1(new_n214), .A2(KEYINPUT73), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n214), .A2(KEYINPUT73), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n229), .B1(new_n243), .B2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n190), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n238), .A2(new_n249), .ZN(new_n250));
  NOR2_X1   g064(.A1(G475), .A2(G902), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n237), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  AOI22_X1  g066(.A1(new_n232), .A2(new_n234), .B1(new_n247), .B2(new_n248), .ZN(new_n253));
  INV_X1    g067(.A(new_n251), .ZN(new_n254));
  NOR3_X1   g068(.A1(new_n253), .A2(KEYINPUT20), .A3(new_n254), .ZN(new_n255));
  OAI211_X1 g069(.A(new_n187), .B(new_n236), .C1(new_n252), .C2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT20), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n250), .A2(new_n258), .A3(new_n251), .ZN(new_n259));
  INV_X1    g073(.A(new_n237), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n260), .B1(new_n253), .B2(new_n254), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n187), .B1(new_n262), .B2(new_n236), .ZN(new_n263));
  NAND2_X1  g077(.A1(G234), .A2(G237), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n264), .A2(G952), .A3(new_n192), .ZN(new_n265));
  XOR2_X1   g079(.A(new_n265), .B(KEYINPUT92), .Z(new_n266));
  AND3_X1   g080(.A1(new_n264), .A2(G902), .A3(G953), .ZN(new_n267));
  XNOR2_X1  g081(.A(KEYINPUT21), .B(G898), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  AND2_X1   g083(.A1(new_n266), .A2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(G128), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n272), .A2(G143), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(G143), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n273), .B1(KEYINPUT13), .B2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT90), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n199), .A2(G128), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT13), .ZN(new_n279));
  OAI21_X1  g093(.A(KEYINPUT90), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  OAI211_X1 g094(.A(new_n277), .B(G134), .C1(new_n275), .C2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(G134), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n278), .A2(new_n274), .A3(new_n282), .ZN(new_n283));
  XNOR2_X1  g097(.A(G116), .B(G122), .ZN(new_n284));
  INV_X1    g098(.A(G107), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(G122), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(G116), .ZN(new_n288));
  INV_X1    g102(.A(G116), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(G122), .ZN(new_n290));
  AND3_X1   g104(.A1(new_n288), .A2(new_n290), .A3(new_n285), .ZN(new_n291));
  OR2_X1    g105(.A1(new_n286), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n281), .A2(new_n283), .A3(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(new_n291), .ZN(new_n294));
  INV_X1    g108(.A(new_n283), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n282), .B1(new_n278), .B2(new_n274), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n294), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT14), .ZN(new_n298));
  OAI21_X1  g112(.A(G107), .B1(new_n290), .B2(new_n298), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n299), .B1(new_n298), .B2(new_n284), .ZN(new_n300));
  OR2_X1    g114(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  XNOR2_X1  g115(.A(KEYINPUT9), .B(G234), .ZN(new_n302));
  INV_X1    g116(.A(G217), .ZN(new_n303));
  NOR3_X1   g117(.A1(new_n302), .A2(new_n303), .A3(G953), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n293), .A2(new_n301), .A3(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(new_n304), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n283), .B1(new_n286), .B2(new_n291), .ZN(new_n307));
  OR2_X1    g121(.A1(new_n275), .A2(new_n280), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n282), .B1(new_n275), .B2(new_n276), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n307), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n297), .A2(new_n300), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n306), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n305), .A2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(G902), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(G478), .ZN(new_n316));
  NOR2_X1   g130(.A1(new_n316), .A2(KEYINPUT15), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  OAI211_X1 g132(.A(new_n313), .B(new_n314), .C1(KEYINPUT15), .C2(new_n316), .ZN(new_n319));
  AND3_X1   g133(.A1(new_n318), .A2(new_n319), .A3(KEYINPUT91), .ZN(new_n320));
  AOI21_X1  g134(.A(KEYINPUT91), .B1(new_n318), .B2(new_n319), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n271), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NOR3_X1   g136(.A1(new_n257), .A2(new_n263), .A3(new_n322), .ZN(new_n323));
  OAI21_X1  g137(.A(G214), .B1(G237), .B2(G902), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n192), .A2(G224), .ZN(new_n326));
  XOR2_X1   g140(.A(new_n326), .B(KEYINPUT83), .Z(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT65), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n329), .B1(new_n212), .B2(G143), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n199), .A2(KEYINPUT65), .A3(G146), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  AOI21_X1  g146(.A(KEYINPUT64), .B1(new_n212), .B2(G143), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n212), .A2(KEYINPUT64), .A3(G143), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n272), .A2(KEYINPUT1), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n332), .A2(new_n334), .A3(new_n335), .A4(new_n336), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n199), .A2(G146), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT1), .ZN(new_n339));
  OAI21_X1  g153(.A(G128), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n199), .A2(G146), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n212), .A2(G143), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n340), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n337), .A2(new_n344), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n345), .A2(G125), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT0), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n347), .A2(new_n272), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n332), .A2(new_n334), .A3(new_n335), .A4(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n348), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n347), .A2(new_n272), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n350), .A2(new_n343), .A3(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n207), .B1(new_n349), .B2(new_n352), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n328), .B1(new_n346), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n349), .A2(new_n352), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(G125), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n356), .B(new_n327), .C1(G125), .C2(new_n345), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n354), .A2(new_n357), .ZN(new_n358));
  XNOR2_X1  g172(.A(G110), .B(G122), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT2), .ZN(new_n360));
  INV_X1    g174(.A(G113), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n360), .A2(new_n361), .A3(KEYINPUT67), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT67), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n363), .B1(KEYINPUT2), .B2(G113), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(KEYINPUT2), .A2(G113), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  XNOR2_X1  g181(.A(G116), .B(G119), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n365), .A2(new_n366), .A3(new_n368), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  OAI21_X1  g186(.A(KEYINPUT3), .B1(new_n189), .B2(G107), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT3), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n374), .A2(new_n285), .A3(G104), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n189), .A2(G107), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n373), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT4), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n377), .A2(new_n378), .A3(G101), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n377), .A2(KEYINPUT77), .A3(G101), .ZN(new_n380));
  INV_X1    g194(.A(G101), .ZN(new_n381));
  NAND4_X1  g195(.A1(new_n373), .A2(new_n375), .A3(new_n381), .A4(new_n376), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n380), .A2(KEYINPUT4), .A3(new_n382), .ZN(new_n383));
  AOI21_X1  g197(.A(KEYINPUT77), .B1(new_n377), .B2(G101), .ZN(new_n384));
  OAI211_X1 g198(.A(new_n372), .B(new_n379), .C1(new_n383), .C2(new_n384), .ZN(new_n385));
  XNOR2_X1  g199(.A(KEYINPUT81), .B(KEYINPUT5), .ZN(new_n386));
  INV_X1    g200(.A(G119), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n386), .A2(G116), .A3(new_n387), .ZN(new_n388));
  OAI211_X1 g202(.A(new_n388), .B(G113), .C1(new_n369), .C2(new_n386), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n189), .A2(G107), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n285), .A2(G104), .ZN(new_n391));
  OAI21_X1  g205(.A(G101), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  AND2_X1   g206(.A1(new_n382), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n389), .A2(new_n371), .A3(new_n393), .ZN(new_n394));
  AOI211_X1 g208(.A(KEYINPUT6), .B(new_n359), .C1(new_n385), .C2(new_n394), .ZN(new_n395));
  AND3_X1   g209(.A1(new_n377), .A2(KEYINPUT77), .A3(G101), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n382), .A2(KEYINPUT4), .ZN(new_n397));
  NOR3_X1   g211(.A1(new_n396), .A2(new_n384), .A3(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(new_n371), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n368), .B1(new_n365), .B2(new_n366), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n379), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  OAI211_X1 g215(.A(new_n359), .B(new_n394), .C1(new_n398), .C2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT82), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n385), .A2(KEYINPUT82), .A3(new_n359), .A4(new_n394), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n359), .B1(new_n385), .B2(new_n394), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT6), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  AOI211_X1 g223(.A(new_n358), .B(new_n395), .C1(new_n406), .C2(new_n409), .ZN(new_n410));
  XNOR2_X1  g224(.A(new_n359), .B(KEYINPUT8), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n368), .A2(KEYINPUT5), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n388), .A2(new_n412), .A3(G113), .ZN(new_n413));
  AND3_X1   g227(.A1(new_n393), .A2(new_n413), .A3(new_n371), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n393), .B1(new_n389), .B2(new_n371), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n411), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n326), .A2(KEYINPUT7), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n417), .B1(new_n346), .B2(new_n353), .ZN(new_n418));
  INV_X1    g232(.A(new_n417), .ZN(new_n419));
  OAI211_X1 g233(.A(new_n356), .B(new_n419), .C1(G125), .C2(new_n345), .ZN(new_n420));
  AND3_X1   g234(.A1(new_n416), .A2(new_n418), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n406), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(new_n314), .ZN(new_n423));
  OAI21_X1  g237(.A(KEYINPUT84), .B1(new_n410), .B2(new_n423), .ZN(new_n424));
  OAI21_X1  g238(.A(G210), .B1(G237), .B2(G902), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n406), .A2(new_n409), .ZN(new_n427));
  INV_X1    g241(.A(new_n395), .ZN(new_n428));
  INV_X1    g242(.A(new_n358), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n427), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT84), .ZN(new_n431));
  AOI21_X1  g245(.A(G902), .B1(new_n406), .B2(new_n421), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n430), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n424), .A2(new_n426), .A3(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n430), .A2(new_n432), .A3(new_n425), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n325), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(G469), .ZN(new_n437));
  INV_X1    g251(.A(new_n355), .ZN(new_n438));
  OAI211_X1 g252(.A(new_n438), .B(new_n379), .C1(new_n383), .C2(new_n384), .ZN(new_n439));
  INV_X1    g253(.A(new_n337), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n272), .B1(new_n342), .B2(KEYINPUT1), .ZN(new_n441));
  AND3_X1   g255(.A1(new_n212), .A2(KEYINPUT64), .A3(G143), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n442), .A2(new_n333), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n441), .B1(new_n443), .B2(new_n332), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n393), .B1(new_n440), .B2(new_n444), .ZN(new_n445));
  XOR2_X1   g259(.A(KEYINPUT78), .B(KEYINPUT10), .Z(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(G137), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n449), .A2(KEYINPUT11), .A3(G134), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n282), .A2(G137), .ZN(new_n451));
  AND2_X1   g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT66), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT11), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n454), .B1(new_n282), .B2(G137), .ZN(new_n455));
  NAND4_X1  g269(.A1(new_n452), .A2(new_n453), .A3(new_n201), .A4(new_n455), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n455), .A2(new_n450), .A3(new_n201), .A4(new_n451), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(KEYINPUT66), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n455), .A2(new_n450), .A3(new_n451), .ZN(new_n459));
  AOI22_X1  g273(.A1(new_n456), .A2(new_n458), .B1(G131), .B2(new_n459), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n345), .A2(KEYINPUT10), .A3(new_n393), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n439), .A2(new_n448), .A3(new_n460), .A4(new_n461), .ZN(new_n462));
  XNOR2_X1  g276(.A(G110), .B(G140), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n192), .A2(G227), .ZN(new_n464));
  XNOR2_X1  g278(.A(new_n463), .B(new_n464), .ZN(new_n465));
  XNOR2_X1  g279(.A(KEYINPUT75), .B(KEYINPUT76), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n465), .B(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n462), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n382), .A2(new_n392), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n470), .A2(new_n337), .A3(new_n344), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n460), .B1(new_n445), .B2(new_n471), .ZN(new_n472));
  OAI21_X1  g286(.A(KEYINPUT80), .B1(new_n472), .B2(KEYINPUT12), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n459), .A2(G131), .ZN(new_n474));
  AND2_X1   g288(.A1(new_n457), .A2(KEYINPUT66), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n457), .A2(KEYINPUT66), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n332), .A2(new_n334), .A3(new_n335), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(new_n340), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n470), .B1(new_n479), .B2(new_n337), .ZN(new_n480));
  INV_X1    g294(.A(new_n471), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n477), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT80), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT12), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n482), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n473), .A2(new_n485), .ZN(new_n486));
  OAI211_X1 g300(.A(KEYINPUT12), .B(new_n477), .C1(new_n480), .C2(new_n481), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(KEYINPUT79), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT79), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n472), .A2(new_n489), .A3(KEYINPUT12), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n469), .B1(new_n486), .B2(new_n491), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n461), .B1(new_n480), .B2(new_n446), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n379), .A2(new_n349), .A3(new_n352), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n398), .A2(new_n494), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n477), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n468), .B1(new_n496), .B2(new_n462), .ZN(new_n497));
  OAI211_X1 g311(.A(new_n437), .B(new_n314), .C1(new_n492), .C2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(new_n469), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(new_n496), .ZN(new_n500));
  INV_X1    g314(.A(new_n462), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n501), .B1(new_n486), .B2(new_n491), .ZN(new_n502));
  OAI211_X1 g316(.A(G469), .B(new_n500), .C1(new_n502), .C2(new_n468), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n437), .A2(new_n314), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n498), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  OAI21_X1  g320(.A(G221), .B1(new_n302), .B2(G902), .ZN(new_n507));
  AND2_X1   g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n323), .A2(new_n436), .A3(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT93), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT74), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n512), .A2(KEYINPUT25), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n272), .A2(G119), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT23), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n514), .B1(KEYINPUT71), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n387), .A2(G128), .ZN(new_n517));
  XNOR2_X1  g331(.A(KEYINPUT71), .B(KEYINPUT23), .ZN(new_n518));
  OAI211_X1 g332(.A(new_n516), .B(new_n517), .C1(new_n518), .C2(new_n514), .ZN(new_n519));
  XNOR2_X1  g333(.A(KEYINPUT72), .B(G110), .ZN(new_n520));
  AND2_X1   g334(.A1(new_n514), .A2(new_n517), .ZN(new_n521));
  XOR2_X1   g335(.A(KEYINPUT24), .B(G110), .Z(new_n522));
  OAI22_X1  g336(.A1(new_n519), .A2(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n523), .A2(new_n244), .A3(new_n245), .A4(new_n223), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n213), .A2(new_n214), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n521), .A2(new_n522), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n519), .A2(G110), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n525), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n524), .A2(new_n528), .ZN(new_n529));
  XNOR2_X1  g343(.A(KEYINPUT22), .B(G137), .ZN(new_n530));
  AND3_X1   g344(.A1(new_n192), .A2(G221), .A3(G234), .ZN(new_n531));
  XNOR2_X1  g345(.A(new_n530), .B(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n529), .A2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(new_n532), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n524), .A2(new_n528), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n513), .B1(new_n536), .B2(G902), .ZN(new_n537));
  INV_X1    g351(.A(new_n513), .ZN(new_n538));
  NAND4_X1  g352(.A1(new_n533), .A2(new_n314), .A3(new_n535), .A4(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n303), .B1(G234), .B2(new_n314), .ZN(new_n541));
  AND2_X1   g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NOR3_X1   g356(.A1(new_n536), .A2(G902), .A3(new_n541), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT31), .ZN(new_n546));
  INV_X1    g360(.A(new_n372), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n477), .A2(new_n438), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n449), .A2(G134), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n201), .B1(new_n549), .B2(new_n451), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n550), .B1(new_n337), .B2(new_n344), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n456), .A2(new_n458), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n551), .A2(new_n552), .A3(KEYINPUT68), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n548), .A2(new_n553), .ZN(new_n554));
  AOI21_X1  g368(.A(KEYINPUT68), .B1(new_n551), .B2(new_n552), .ZN(new_n555));
  OAI21_X1  g369(.A(KEYINPUT30), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT30), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n551), .A2(new_n552), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n548), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n547), .B1(new_n556), .B2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT68), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  NAND4_X1  g376(.A1(new_n562), .A2(new_n547), .A3(new_n548), .A4(new_n553), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n194), .A2(G210), .ZN(new_n564));
  XNOR2_X1  g378(.A(new_n564), .B(KEYINPUT27), .ZN(new_n565));
  XNOR2_X1  g379(.A(KEYINPUT26), .B(G101), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n565), .B(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n563), .A2(new_n567), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n546), .B1(new_n560), .B2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n568), .ZN(new_n570));
  AND3_X1   g384(.A1(new_n548), .A2(new_n557), .A3(new_n558), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n562), .A2(new_n548), .A3(new_n553), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n571), .B1(KEYINPUT30), .B2(new_n572), .ZN(new_n573));
  OAI211_X1 g387(.A(new_n570), .B(KEYINPUT31), .C1(new_n573), .C2(new_n547), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n548), .A2(new_n547), .A3(new_n558), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT28), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT70), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n575), .A2(KEYINPUT70), .A3(new_n576), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n460), .A2(new_n355), .ZN(new_n581));
  AND2_X1   g395(.A1(new_n551), .A2(new_n552), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n372), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  AND2_X1   g397(.A1(new_n563), .A2(new_n583), .ZN(new_n584));
  OAI211_X1 g398(.A(new_n579), .B(new_n580), .C1(new_n584), .C2(new_n576), .ZN(new_n585));
  XOR2_X1   g399(.A(new_n567), .B(KEYINPUT69), .Z(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  AOI22_X1  g401(.A1(new_n569), .A2(new_n574), .B1(new_n585), .B2(new_n587), .ZN(new_n588));
  NOR2_X1   g402(.A1(G472), .A2(G902), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  OAI21_X1  g404(.A(KEYINPUT32), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n569), .A2(new_n574), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n585), .A2(new_n587), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT32), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n594), .A2(new_n595), .A3(new_n589), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n591), .A2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT29), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n586), .A2(new_n598), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n585), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n579), .A2(new_n580), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n372), .B1(new_n554), .B2(new_n555), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n576), .B1(new_n602), .B2(new_n563), .ZN(new_n603));
  OAI21_X1  g417(.A(KEYINPUT29), .B1(new_n601), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(new_n567), .ZN(new_n605));
  INV_X1    g419(.A(new_n563), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n560), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(new_n598), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n600), .B1(new_n605), .B2(new_n608), .ZN(new_n609));
  OAI21_X1  g423(.A(G472), .B1(new_n609), .B2(G902), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n545), .B1(new_n597), .B2(new_n610), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n323), .A2(new_n436), .A3(new_n508), .A4(KEYINPUT93), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n511), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n613), .B(G101), .ZN(G3));
  OAI21_X1  g428(.A(new_n236), .B1(new_n252), .B2(new_n255), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(KEYINPUT89), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(new_n256), .ZN(new_n617));
  NAND2_X1  g431(.A1(G478), .A2(G902), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n618), .B1(new_n315), .B2(G478), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT33), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n313), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(KEYINPUT94), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT94), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n313), .A2(new_n624), .A3(new_n621), .ZN(new_n625));
  OAI21_X1  g439(.A(KEYINPUT95), .B1(new_n313), .B2(new_n621), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT95), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n305), .A2(new_n312), .A3(new_n627), .A4(KEYINPUT33), .ZN(new_n628));
  AOI22_X1  g442(.A1(new_n623), .A2(new_n625), .B1(new_n626), .B2(new_n628), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n620), .B1(new_n629), .B2(new_n316), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n617), .A2(new_n631), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n426), .B1(new_n410), .B2(new_n423), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n325), .B1(new_n633), .B2(new_n435), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  NOR3_X1   g449(.A1(new_n632), .A2(new_n270), .A3(new_n635), .ZN(new_n636));
  OAI21_X1  g450(.A(G472), .B1(new_n588), .B2(G902), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n594), .A2(new_n589), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n544), .A2(new_n507), .A3(new_n506), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n636), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT34), .B(G104), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G6));
  NOR2_X1   g458(.A1(new_n320), .A2(new_n321), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n250), .A2(new_n251), .A3(new_n237), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(new_n261), .ZN(new_n647));
  AND2_X1   g461(.A1(new_n647), .A2(new_n236), .ZN(new_n648));
  AND4_X1   g462(.A1(new_n271), .A2(new_n634), .A3(new_n645), .A4(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n641), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(KEYINPUT96), .ZN(new_n651));
  XNOR2_X1  g465(.A(KEYINPUT35), .B(G107), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G9));
  NAND2_X1  g467(.A1(new_n540), .A2(new_n541), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n532), .A2(KEYINPUT36), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n529), .B(new_n655), .ZN(new_n656));
  OAI211_X1 g470(.A(new_n656), .B(new_n314), .C1(new_n303), .C2(G234), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n654), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(KEYINPUT97), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT97), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n654), .A2(new_n660), .A3(new_n657), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n639), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n511), .A2(new_n612), .A3(new_n663), .ZN(new_n664));
  XOR2_X1   g478(.A(KEYINPUT37), .B(G110), .Z(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G12));
  NAND2_X1  g480(.A1(new_n597), .A2(new_n610), .ZN(new_n667));
  INV_X1    g481(.A(G900), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n267), .A2(new_n668), .ZN(new_n669));
  AND2_X1   g483(.A1(new_n266), .A2(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n648), .A2(new_n645), .A3(new_n671), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n662), .A2(new_n672), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n667), .A2(new_n673), .A3(new_n508), .A4(new_n634), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G128), .ZN(G30));
  XNOR2_X1  g489(.A(KEYINPUT100), .B(KEYINPUT39), .ZN(new_n676));
  XOR2_X1   g490(.A(new_n670), .B(new_n676), .Z(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n508), .A2(new_n678), .ZN(new_n679));
  OR2_X1    g493(.A1(new_n679), .A2(KEYINPUT40), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n679), .A2(KEYINPUT40), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n257), .A2(new_n263), .ZN(new_n682));
  INV_X1    g496(.A(new_n645), .ZN(new_n683));
  NOR4_X1   g497(.A1(new_n682), .A2(new_n325), .A3(new_n683), .A4(new_n658), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n586), .B1(new_n563), .B2(new_n602), .ZN(new_n685));
  OAI22_X1  g499(.A1(new_n685), .A2(KEYINPUT99), .B1(new_n560), .B2(new_n568), .ZN(new_n686));
  AND2_X1   g500(.A1(new_n685), .A2(KEYINPUT99), .ZN(new_n687));
  OAI21_X1  g501(.A(new_n314), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(G472), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n597), .A2(new_n689), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n680), .A2(new_n681), .A3(new_n684), .A4(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n434), .A2(new_n435), .ZN(new_n692));
  XNOR2_X1  g506(.A(KEYINPUT98), .B(KEYINPUT38), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(new_n199), .ZN(G45));
  OAI211_X1 g510(.A(new_n631), .B(new_n671), .C1(new_n257), .C2(new_n263), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n697), .A2(new_n662), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n698), .A2(new_n667), .A3(new_n508), .A4(new_n634), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G146), .ZN(G48));
  NAND2_X1  g514(.A1(new_n486), .A2(new_n491), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n497), .B1(new_n701), .B2(new_n499), .ZN(new_n702));
  OAI21_X1  g516(.A(G469), .B1(new_n702), .B2(G902), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n703), .A2(new_n507), .A3(new_n498), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT101), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n703), .A2(KEYINPUT101), .A3(new_n507), .A4(new_n498), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n636), .A2(new_n611), .A3(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(KEYINPUT41), .B(G113), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n710), .B(new_n711), .ZN(G15));
  NAND3_X1  g526(.A1(new_n611), .A2(new_n709), .A3(new_n649), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G116), .ZN(G18));
  NAND3_X1  g528(.A1(new_n706), .A2(new_n634), .A3(new_n707), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT102), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n706), .A2(KEYINPUT102), .A3(new_n634), .A4(new_n707), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  AOI22_X1  g533(.A1(new_n604), .A2(new_n567), .B1(new_n607), .B2(new_n598), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n314), .B1(new_n720), .B2(new_n600), .ZN(new_n721));
  AOI22_X1  g535(.A1(new_n591), .A2(new_n596), .B1(new_n721), .B2(G472), .ZN(new_n722));
  INV_X1    g536(.A(new_n323), .ZN(new_n723));
  NOR3_X1   g537(.A1(new_n722), .A2(new_n723), .A3(new_n662), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n719), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G119), .ZN(G21));
  OAI21_X1  g540(.A(new_n587), .B1(new_n601), .B2(new_n603), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n592), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(new_n589), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n637), .A2(new_n544), .A3(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(KEYINPUT103), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n617), .A2(new_n645), .A3(new_n634), .ZN(new_n732));
  NOR3_X1   g546(.A1(new_n708), .A2(new_n732), .A3(new_n270), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G122), .ZN(G24));
  NAND2_X1  g549(.A1(new_n594), .A2(new_n314), .ZN(new_n736));
  AOI22_X1  g550(.A1(new_n736), .A2(G472), .B1(new_n589), .B2(new_n728), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n630), .B1(new_n616), .B2(new_n256), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n737), .A2(new_n738), .A3(new_n658), .A4(new_n671), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n739), .B1(new_n717), .B2(new_n718), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(new_n207), .ZN(G27));
  AND2_X1   g555(.A1(new_n435), .A2(new_n324), .ZN(new_n742));
  AND3_X1   g556(.A1(new_n434), .A2(new_n742), .A3(KEYINPUT104), .ZN(new_n743));
  AOI21_X1  g557(.A(KEYINPUT104), .B1(new_n434), .B2(new_n742), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n697), .A2(KEYINPUT42), .ZN(new_n746));
  AND4_X1   g560(.A1(new_n611), .A2(new_n745), .A3(new_n508), .A4(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n506), .A2(new_n507), .ZN(new_n748));
  NOR4_X1   g562(.A1(new_n697), .A2(new_n743), .A3(new_n744), .A4(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT105), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n750), .B1(new_n722), .B2(new_n545), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n611), .A2(KEYINPUT105), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n749), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n747), .B1(new_n753), .B2(KEYINPUT42), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G131), .ZN(G33));
  INV_X1    g569(.A(new_n672), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n611), .A2(new_n745), .A3(new_n508), .A4(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(KEYINPUT106), .B(G134), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n757), .B(new_n758), .ZN(G36));
  INV_X1    g573(.A(new_n498), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n500), .B1(new_n502), .B2(new_n468), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT45), .ZN(new_n762));
  OR2_X1    g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n437), .B1(new_n761), .B2(new_n762), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n504), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT46), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n760), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NOR3_X1   g582(.A1(new_n766), .A2(KEYINPUT107), .A3(new_n767), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT107), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n770), .B1(new_n765), .B2(KEYINPUT46), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n768), .B1(new_n769), .B2(new_n771), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n772), .A2(new_n507), .A3(new_n678), .A4(new_n745), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n639), .A2(new_n658), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(KEYINPUT108), .ZN(new_n775));
  INV_X1    g589(.A(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n682), .A2(new_n631), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(KEYINPUT43), .ZN(new_n778));
  OR3_X1    g592(.A1(new_n617), .A2(KEYINPUT43), .A3(new_n630), .ZN(new_n779));
  AND2_X1   g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT44), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n776), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(new_n780), .ZN(new_n783));
  OAI21_X1  g597(.A(KEYINPUT44), .B1(new_n783), .B2(new_n775), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n773), .B1(new_n782), .B2(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(new_n449), .ZN(G39));
  INV_X1    g600(.A(new_n745), .ZN(new_n787));
  OR4_X1    g601(.A1(new_n667), .A2(new_n787), .A3(new_n544), .A4(new_n697), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n772), .A2(new_n507), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT47), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n772), .A2(KEYINPUT47), .A3(new_n507), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n788), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(new_n205), .ZN(G42));
  INV_X1    g608(.A(KEYINPUT51), .ZN(new_n795));
  NOR3_X1   g609(.A1(new_n690), .A2(new_n545), .A3(new_n266), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n796), .A2(new_n709), .A3(new_n745), .ZN(new_n797));
  NOR3_X1   g611(.A1(new_n797), .A2(new_n617), .A3(new_n631), .ZN(new_n798));
  NOR4_X1   g612(.A1(new_n783), .A2(new_n266), .A3(new_n708), .A4(new_n787), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n637), .A2(new_n658), .A3(new_n729), .ZN(new_n800));
  INV_X1    g614(.A(new_n800), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n798), .B1(new_n799), .B2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(new_n266), .ZN(new_n803));
  AND3_X1   g617(.A1(new_n780), .A2(new_n803), .A3(new_n731), .ZN(new_n804));
  INV_X1    g618(.A(new_n694), .ZN(new_n805));
  OR3_X1    g619(.A1(new_n708), .A2(KEYINPUT112), .A3(new_n324), .ZN(new_n806));
  OAI21_X1  g620(.A(KEYINPUT112), .B1(new_n708), .B2(new_n324), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n805), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n804), .A2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT50), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n804), .A2(KEYINPUT50), .A3(new_n808), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n811), .A2(KEYINPUT113), .A3(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(new_n813), .ZN(new_n814));
  AOI21_X1  g628(.A(KEYINPUT113), .B1(new_n811), .B2(new_n812), .ZN(new_n815));
  OAI211_X1 g629(.A(KEYINPUT114), .B(new_n802), .C1(new_n814), .C2(new_n815), .ZN(new_n816));
  AND2_X1   g630(.A1(new_n791), .A2(new_n792), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n703), .A2(new_n498), .ZN(new_n818));
  OR2_X1    g632(.A1(new_n818), .A2(new_n507), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n804), .A2(new_n745), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n816), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n811), .A2(new_n812), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT113), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(new_n813), .ZN(new_n827));
  AOI21_X1  g641(.A(KEYINPUT114), .B1(new_n827), .B2(new_n802), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n795), .B1(new_n823), .B2(new_n828), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n751), .A2(new_n752), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n799), .A2(new_n830), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n831), .B(KEYINPUT48), .ZN(new_n832));
  INV_X1    g646(.A(G952), .ZN(new_n833));
  AOI211_X1 g647(.A(new_n833), .B(G953), .C1(new_n804), .C2(new_n719), .ZN(new_n834));
  OAI211_X1 g648(.A(new_n832), .B(new_n834), .C1(new_n632), .C2(new_n797), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT115), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n820), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n817), .A2(KEYINPUT115), .A3(new_n819), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n837), .A2(new_n821), .A3(new_n838), .ZN(new_n839));
  AND3_X1   g653(.A1(new_n824), .A2(KEYINPUT51), .A3(new_n802), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n835), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n692), .A2(new_n324), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n842), .A2(new_n270), .ZN(new_n843));
  OR2_X1    g657(.A1(new_n738), .A2(KEYINPUT109), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n738), .A2(KEYINPUT109), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n843), .A2(new_n844), .A3(new_n641), .A4(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n613), .A2(new_n710), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n318), .A2(new_n319), .ZN(new_n848));
  INV_X1    g662(.A(new_n848), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n617), .A2(new_n849), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n850), .A2(KEYINPUT110), .A3(new_n436), .A4(new_n271), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT110), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n616), .A2(new_n256), .A3(new_n271), .A4(new_n848), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n852), .B1(new_n842), .B2(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n851), .A2(new_n854), .A3(new_n641), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n664), .A2(new_n855), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n847), .A2(new_n856), .ZN(new_n857));
  AND3_X1   g671(.A1(new_n725), .A2(new_n734), .A3(new_n713), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n800), .A2(new_n697), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n745), .A2(new_n859), .A3(new_n508), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n748), .B1(new_n597), .B2(new_n610), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n648), .A2(new_n671), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n662), .A2(new_n848), .A3(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n861), .A2(new_n745), .A3(new_n863), .ZN(new_n864));
  AND3_X1   g678(.A1(new_n757), .A2(new_n860), .A3(new_n864), .ZN(new_n865));
  AND4_X1   g679(.A1(new_n754), .A2(new_n857), .A3(new_n858), .A4(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n719), .A2(new_n859), .ZN(new_n867));
  OAI211_X1 g681(.A(new_n861), .B(new_n634), .C1(new_n673), .C2(new_n698), .ZN(new_n868));
  INV_X1    g682(.A(new_n732), .ZN(new_n869));
  NOR3_X1   g683(.A1(new_n748), .A2(new_n658), .A3(new_n670), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n869), .A2(new_n690), .A3(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n867), .A2(new_n868), .A3(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT52), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n867), .A2(KEYINPUT52), .A3(new_n868), .A4(new_n871), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n866), .A2(KEYINPUT53), .A3(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n753), .A2(KEYINPUT42), .ZN(new_n878));
  INV_X1    g692(.A(new_n747), .ZN(new_n879));
  AND3_X1   g693(.A1(new_n878), .A2(new_n865), .A3(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n725), .A2(new_n734), .A3(new_n713), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n881), .A2(new_n847), .A3(new_n856), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n876), .A2(new_n880), .A3(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT53), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n877), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n699), .A2(new_n674), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n887), .A2(new_n740), .ZN(new_n888));
  AOI21_X1  g702(.A(KEYINPUT52), .B1(new_n888), .B2(new_n871), .ZN(new_n889));
  INV_X1    g703(.A(new_n875), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  AND4_X1   g705(.A1(KEYINPUT53), .A2(new_n757), .A3(new_n860), .A4(new_n864), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n857), .A2(new_n858), .A3(new_n754), .A4(new_n892), .ZN(new_n893));
  OAI21_X1  g707(.A(KEYINPUT111), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  AND2_X1   g708(.A1(new_n754), .A2(new_n892), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT111), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n895), .A2(new_n876), .A3(new_n896), .A4(new_n882), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n894), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g712(.A(KEYINPUT54), .B1(new_n883), .B2(new_n884), .ZN(new_n899));
  AOI22_X1  g713(.A1(new_n886), .A2(KEYINPUT54), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n829), .A2(new_n841), .A3(new_n900), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n901), .B1(G952), .B2(G953), .ZN(new_n902));
  AND3_X1   g716(.A1(new_n544), .A2(new_n324), .A3(new_n507), .ZN(new_n903));
  OR2_X1    g717(.A1(new_n818), .A2(KEYINPUT49), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n818), .A2(KEYINPUT49), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n903), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  OR4_X1    g720(.A1(new_n805), .A2(new_n906), .A3(new_n690), .A4(new_n777), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n902), .A2(new_n907), .ZN(G75));
  NAND2_X1  g722(.A1(new_n833), .A2(G953), .ZN(new_n909));
  XOR2_X1   g723(.A(new_n909), .B(KEYINPUT116), .Z(new_n910));
  INV_X1    g724(.A(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT56), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n898), .A2(new_n885), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(G902), .ZN(new_n914));
  INV_X1    g728(.A(G210), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n912), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n427), .A2(new_n428), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(new_n358), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n918), .A2(new_n430), .ZN(new_n919));
  XOR2_X1   g733(.A(new_n919), .B(KEYINPUT55), .Z(new_n920));
  NAND2_X1  g734(.A1(new_n916), .A2(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(new_n920), .ZN(new_n922));
  OAI211_X1 g736(.A(new_n912), .B(new_n922), .C1(new_n914), .C2(new_n915), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n911), .B1(new_n921), .B2(new_n923), .ZN(G51));
  XNOR2_X1  g738(.A(new_n504), .B(KEYINPUT57), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT117), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n898), .A2(new_n926), .A3(new_n899), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT54), .ZN(new_n928));
  AOI22_X1  g742(.A1(new_n894), .A2(new_n897), .B1(new_n884), .B2(new_n883), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n927), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n926), .B1(new_n898), .B2(new_n899), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n925), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(new_n702), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(new_n914), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n935), .A2(new_n763), .A3(new_n764), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n911), .B1(new_n934), .B2(new_n936), .ZN(G54));
  NAND2_X1  g751(.A1(KEYINPUT58), .A2(G475), .ZN(new_n938));
  OR3_X1    g752(.A1(new_n914), .A2(new_n250), .A3(new_n938), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n250), .B1(new_n914), .B2(new_n938), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n911), .B1(new_n939), .B2(new_n940), .ZN(G60));
  INV_X1    g755(.A(KEYINPUT118), .ZN(new_n942));
  XOR2_X1   g756(.A(new_n618), .B(KEYINPUT59), .Z(new_n943));
  AOI21_X1  g757(.A(KEYINPUT53), .B1(new_n866), .B2(new_n876), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n883), .A2(new_n884), .ZN(new_n945));
  OAI21_X1  g759(.A(KEYINPUT54), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n898), .A2(new_n899), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n943), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n942), .B1(new_n948), .B2(new_n629), .ZN(new_n949));
  INV_X1    g763(.A(new_n629), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n950), .A2(new_n943), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n951), .B1(new_n930), .B2(new_n931), .ZN(new_n952));
  OAI211_X1 g766(.A(KEYINPUT118), .B(new_n950), .C1(new_n900), .C2(new_n943), .ZN(new_n953));
  AND4_X1   g767(.A1(new_n910), .A2(new_n949), .A3(new_n952), .A4(new_n953), .ZN(G63));
  XNOR2_X1  g768(.A(KEYINPUT120), .B(KEYINPUT60), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n303), .A2(new_n314), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n955), .B(new_n956), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n913), .A2(new_n656), .A3(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(new_n957), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n536), .B1(new_n929), .B2(new_n959), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n958), .A2(new_n960), .A3(new_n910), .ZN(new_n961));
  AND3_X1   g775(.A1(new_n961), .A2(KEYINPUT119), .A3(KEYINPUT61), .ZN(new_n962));
  AOI21_X1  g776(.A(KEYINPUT61), .B1(new_n961), .B2(KEYINPUT119), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n962), .A2(new_n963), .ZN(G66));
  INV_X1    g778(.A(G224), .ZN(new_n965));
  OAI21_X1  g779(.A(G953), .B1(new_n268), .B2(new_n965), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n966), .B1(new_n882), .B2(G953), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n917), .B1(G898), .B2(new_n192), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n967), .B(new_n968), .ZN(G69));
  AND3_X1   g783(.A1(new_n611), .A2(new_n745), .A3(new_n508), .ZN(new_n970));
  AND2_X1   g784(.A1(new_n844), .A2(new_n845), .ZN(new_n971));
  OAI211_X1 g785(.A(new_n970), .B(new_n678), .C1(new_n971), .C2(new_n850), .ZN(new_n972));
  INV_X1    g786(.A(KEYINPUT123), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n972), .B(new_n973), .ZN(new_n974));
  NOR3_X1   g788(.A1(new_n974), .A2(new_n785), .A3(new_n793), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n888), .A2(KEYINPUT122), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT122), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n977), .B1(new_n887), .B2(new_n740), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(new_n695), .ZN(new_n980));
  AOI21_X1  g794(.A(KEYINPUT62), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  AND3_X1   g795(.A1(new_n979), .A2(KEYINPUT62), .A3(new_n980), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n975), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n983), .A2(new_n192), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n242), .B(KEYINPUT121), .ZN(new_n985));
  XOR2_X1   g799(.A(new_n573), .B(new_n985), .Z(new_n986));
  NAND2_X1  g800(.A1(new_n830), .A2(new_n869), .ZN(new_n987));
  NOR3_X1   g801(.A1(new_n987), .A2(new_n677), .A3(new_n789), .ZN(new_n988));
  INV_X1    g802(.A(new_n754), .ZN(new_n989));
  INV_X1    g803(.A(new_n757), .ZN(new_n990));
  NOR3_X1   g804(.A1(new_n988), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n793), .A2(new_n785), .ZN(new_n992));
  NAND4_X1  g806(.A1(new_n991), .A2(new_n992), .A3(new_n192), .A4(new_n979), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n986), .B1(G900), .B2(G953), .ZN(new_n994));
  AOI22_X1  g808(.A1(new_n984), .A2(new_n986), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n192), .B1(G227), .B2(G900), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n993), .A2(new_n994), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n996), .B1(new_n997), .B2(KEYINPUT124), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n995), .B(new_n998), .ZN(G72));
  INV_X1    g813(.A(new_n567), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n607), .A2(new_n1000), .ZN(new_n1001));
  XOR2_X1   g815(.A(new_n1001), .B(KEYINPUT126), .Z(new_n1002));
  NAND4_X1  g816(.A1(new_n991), .A2(new_n992), .A3(new_n882), .A4(new_n979), .ZN(new_n1003));
  NAND2_X1  g817(.A1(G472), .A2(G902), .ZN(new_n1004));
  XOR2_X1   g818(.A(new_n1004), .B(KEYINPUT63), .Z(new_n1005));
  AOI21_X1  g819(.A(new_n1002), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g820(.A1(new_n607), .A2(new_n1000), .ZN(new_n1007));
  INV_X1    g821(.A(new_n1007), .ZN(new_n1008));
  NAND3_X1  g822(.A1(new_n1008), .A2(new_n1005), .A3(new_n1001), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n1009), .B1(new_n877), .B2(new_n885), .ZN(new_n1010));
  NOR3_X1   g824(.A1(new_n1006), .A2(new_n1010), .A3(new_n911), .ZN(new_n1011));
  OAI211_X1 g825(.A(new_n975), .B(new_n882), .C1(new_n981), .C2(new_n982), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n1012), .A2(KEYINPUT125), .A3(new_n1005), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1013), .A2(new_n1007), .ZN(new_n1014));
  AOI21_X1  g828(.A(KEYINPUT125), .B1(new_n1012), .B2(new_n1005), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n1011), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1016), .A2(KEYINPUT127), .ZN(new_n1017));
  INV_X1    g831(.A(KEYINPUT127), .ZN(new_n1018));
  OAI211_X1 g832(.A(new_n1018), .B(new_n1011), .C1(new_n1014), .C2(new_n1015), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1017), .A2(new_n1019), .ZN(G57));
endmodule


