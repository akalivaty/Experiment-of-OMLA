//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 1 0 1 0 1 0 0 0 0 1 0 1 0 1 1 1 0 0 1 1 1 1 1 1 0 1 0 1 1 0 1 0 1 1 1 1 1 0 1 0 1 1 1 0 1 1 1 1 1 1 1 0 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:59 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n728, new_n729, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n741, new_n742, new_n743,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001;
  INV_X1    g000(.A(G472), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(G101), .ZN(new_n189));
  INV_X1    g003(.A(G237), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(KEYINPUT73), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT73), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G237), .ZN(new_n193));
  AOI21_X1  g007(.A(G953), .B1(new_n191), .B2(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G210), .ZN(new_n195));
  XNOR2_X1  g009(.A(new_n189), .B(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT28), .ZN(new_n197));
  INV_X1    g011(.A(G134), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G137), .ZN(new_n199));
  INV_X1    g013(.A(G137), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G134), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n199), .A2(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G131), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT11), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n204), .B1(new_n198), .B2(G137), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n200), .A2(KEYINPUT11), .A3(G134), .ZN(new_n206));
  INV_X1    g020(.A(G131), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n205), .A2(new_n206), .A3(new_n207), .A4(new_n199), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT68), .ZN(new_n209));
  AND2_X1   g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n208), .A2(new_n209), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n203), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT70), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT64), .ZN(new_n215));
  INV_X1    g029(.A(G146), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n215), .B1(new_n216), .B2(G143), .ZN(new_n217));
  INV_X1    g031(.A(G143), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n218), .A2(KEYINPUT64), .A3(G146), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n216), .A2(G143), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  AOI21_X1  g036(.A(KEYINPUT69), .B1(new_n221), .B2(KEYINPUT1), .ZN(new_n223));
  OAI211_X1 g037(.A(KEYINPUT69), .B(KEYINPUT1), .C1(new_n218), .C2(G146), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(G128), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n222), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  OAI21_X1  g040(.A(KEYINPUT65), .B1(new_n218), .B2(G146), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT65), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n228), .A2(new_n216), .A3(G143), .ZN(new_n229));
  AND2_X1   g043(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  OAI21_X1  g044(.A(KEYINPUT66), .B1(new_n216), .B2(G143), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT66), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n232), .A2(new_n218), .A3(G146), .ZN(new_n233));
  INV_X1    g047(.A(G128), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n234), .A2(KEYINPUT1), .ZN(new_n235));
  NAND4_X1  g049(.A1(new_n230), .A2(new_n231), .A3(new_n233), .A4(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n226), .A2(new_n236), .ZN(new_n237));
  XNOR2_X1  g051(.A(new_n208), .B(new_n209), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n238), .A2(KEYINPUT70), .A3(new_n203), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n214), .A2(new_n237), .A3(new_n239), .ZN(new_n240));
  XOR2_X1   g054(.A(G116), .B(G119), .Z(new_n241));
  XNOR2_X1  g055(.A(KEYINPUT2), .B(G113), .ZN(new_n242));
  XNOR2_X1  g056(.A(new_n241), .B(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(KEYINPUT0), .A2(G128), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  NOR2_X1   g060(.A1(KEYINPUT0), .A2(G128), .ZN(new_n247));
  AOI211_X1 g061(.A(new_n246), .B(new_n247), .C1(new_n220), .C2(new_n221), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n231), .A2(new_n227), .A3(new_n233), .A4(new_n229), .ZN(new_n249));
  OR3_X1    g063(.A1(new_n249), .A2(KEYINPUT67), .A3(new_n245), .ZN(new_n250));
  OAI21_X1  g064(.A(KEYINPUT67), .B1(new_n249), .B2(new_n245), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n248), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n205), .A2(new_n199), .A3(new_n206), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G131), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n238), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n252), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n240), .A2(new_n244), .A3(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT72), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n240), .A2(KEYINPUT72), .A3(new_n244), .A4(new_n256), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(new_n211), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n208), .A2(new_n209), .ZN(new_n263));
  AOI22_X1  g077(.A1(new_n262), .A2(new_n263), .B1(G131), .B2(new_n202), .ZN(new_n264));
  AOI22_X1  g078(.A1(new_n252), .A2(new_n255), .B1(new_n264), .B2(new_n237), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(new_n243), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n197), .B1(new_n261), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n257), .A2(new_n197), .ZN(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n196), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n240), .A2(KEYINPUT30), .A3(new_n256), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(KEYINPUT71), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT71), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n240), .A2(new_n274), .A3(KEYINPUT30), .A4(new_n256), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n243), .B1(new_n265), .B2(KEYINPUT30), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(new_n196), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n279), .A2(new_n261), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n271), .A2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT29), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n280), .A2(new_n283), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n244), .B1(new_n240), .B2(new_n256), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n286), .B1(new_n259), .B2(new_n260), .ZN(new_n287));
  OAI211_X1 g101(.A(new_n269), .B(new_n285), .C1(new_n287), .C2(new_n197), .ZN(new_n288));
  INV_X1    g102(.A(G902), .ZN(new_n289));
  AND2_X1   g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n187), .B1(new_n284), .B2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT32), .ZN(new_n292));
  NOR2_X1   g106(.A1(G472), .A2(G902), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n261), .A2(new_n196), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n277), .B1(new_n273), .B2(new_n275), .ZN(new_n296));
  NOR3_X1   g110(.A1(new_n295), .A2(KEYINPUT31), .A3(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT31), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n280), .B1(new_n259), .B2(new_n260), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n298), .B1(new_n279), .B2(new_n299), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n280), .B1(new_n268), .B2(new_n270), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n294), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n292), .B1(new_n303), .B2(KEYINPUT74), .ZN(new_n304));
  OAI21_X1  g118(.A(KEYINPUT31), .B1(new_n295), .B2(new_n296), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n279), .A2(new_n298), .A3(new_n299), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n302), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(new_n293), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT74), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n308), .A2(new_n309), .A3(KEYINPUT32), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n291), .B1(new_n304), .B2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT23), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n312), .A2(new_n234), .A3(G119), .ZN(new_n313));
  INV_X1    g127(.A(G119), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(G128), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n234), .A2(G119), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n313), .B1(new_n317), .B2(new_n312), .ZN(new_n318));
  INV_X1    g132(.A(G110), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  OR2_X1    g134(.A1(KEYINPUT24), .A2(G110), .ZN(new_n321));
  NAND2_X1  g135(.A1(KEYINPUT24), .A2(G110), .ZN(new_n322));
  AND3_X1   g136(.A1(new_n321), .A2(KEYINPUT75), .A3(new_n322), .ZN(new_n323));
  AOI21_X1  g137(.A(KEYINPUT75), .B1(new_n321), .B2(new_n322), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n317), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n320), .A2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(G140), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(G125), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n328), .A2(KEYINPUT16), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n327), .A2(KEYINPUT77), .A3(G125), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT77), .ZN(new_n333));
  XNOR2_X1  g147(.A(G125), .B(G140), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n332), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT16), .ZN(new_n336));
  OAI211_X1 g150(.A(G146), .B(new_n330), .C1(new_n335), .C2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n334), .A2(new_n216), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n326), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(KEYINPUT78), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT78), .ZN(new_n341));
  NAND4_X1  g155(.A1(new_n326), .A2(new_n337), .A3(new_n341), .A4(new_n338), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  OAI211_X1 g157(.A(new_n313), .B(G110), .C1(new_n317), .C2(new_n312), .ZN(new_n344));
  XOR2_X1   g158(.A(new_n344), .B(KEYINPUT76), .Z(new_n345));
  INV_X1    g159(.A(G125), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(G140), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n328), .A2(new_n347), .A3(new_n333), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n336), .B1(new_n348), .B2(new_n331), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n216), .B1(new_n349), .B2(new_n329), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n337), .A2(new_n350), .ZN(new_n351));
  OR2_X1    g165(.A1(new_n323), .A2(new_n324), .ZN(new_n352));
  OAI211_X1 g166(.A(new_n345), .B(new_n351), .C1(new_n317), .C2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(G953), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n354), .A2(G221), .A3(G234), .ZN(new_n355));
  XNOR2_X1  g169(.A(new_n355), .B(KEYINPUT22), .ZN(new_n356));
  XNOR2_X1  g170(.A(new_n356), .B(G137), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n343), .A2(new_n353), .A3(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  AOI21_X1  g173(.A(KEYINPUT79), .B1(new_n343), .B2(new_n353), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n343), .A2(KEYINPUT79), .A3(new_n353), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n357), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n359), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(G217), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n366), .B1(G234), .B2(new_n289), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n367), .A2(G902), .ZN(new_n368));
  AND3_X1   g182(.A1(new_n365), .A2(KEYINPUT80), .A3(new_n368), .ZN(new_n369));
  AOI21_X1  g183(.A(KEYINPUT80), .B1(new_n365), .B2(new_n368), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  AND3_X1   g185(.A1(new_n343), .A2(KEYINPUT79), .A3(new_n353), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n364), .B1(new_n372), .B2(new_n360), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n373), .A2(new_n289), .A3(new_n358), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(KEYINPUT25), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT25), .ZN(new_n376));
  NAND4_X1  g190(.A1(new_n373), .A2(new_n376), .A3(new_n289), .A4(new_n358), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n375), .A2(new_n367), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n371), .A2(new_n378), .ZN(new_n379));
  OAI21_X1  g193(.A(KEYINPUT81), .B1(new_n311), .B2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(new_n291), .ZN(new_n381));
  AOI21_X1  g195(.A(KEYINPUT32), .B1(new_n308), .B2(new_n309), .ZN(new_n382));
  AOI211_X1 g196(.A(KEYINPUT74), .B(new_n292), .C1(new_n307), .C2(new_n293), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n381), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT81), .ZN(new_n385));
  INV_X1    g199(.A(new_n379), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n384), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n380), .A2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT12), .ZN(new_n389));
  INV_X1    g203(.A(G104), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(G107), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n390), .A2(G107), .ZN(new_n393));
  OAI21_X1  g207(.A(G101), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  OAI21_X1  g208(.A(KEYINPUT3), .B1(new_n390), .B2(G107), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT3), .ZN(new_n396));
  INV_X1    g210(.A(G107), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n396), .A2(new_n397), .A3(G104), .ZN(new_n398));
  INV_X1    g212(.A(G101), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n395), .A2(new_n398), .A3(new_n399), .A4(new_n391), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n394), .A2(new_n400), .ZN(new_n401));
  AND3_X1   g215(.A1(new_n226), .A2(new_n236), .A3(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(new_n401), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n221), .A2(KEYINPUT1), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(G128), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n249), .A2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT84), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n249), .A2(KEYINPUT84), .A3(new_n405), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n408), .A2(new_n236), .A3(new_n409), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n402), .B1(new_n403), .B2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(new_n255), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n389), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n226), .A2(new_n236), .A3(new_n401), .ZN(new_n414));
  AND3_X1   g228(.A1(new_n249), .A2(KEYINPUT84), .A3(new_n405), .ZN(new_n415));
  AOI21_X1  g229(.A(KEYINPUT84), .B1(new_n249), .B2(new_n405), .ZN(new_n416));
  INV_X1    g230(.A(new_n235), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n249), .A2(new_n417), .ZN(new_n418));
  NOR3_X1   g232(.A1(new_n415), .A2(new_n416), .A3(new_n418), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n414), .B1(new_n419), .B2(new_n401), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n420), .A2(KEYINPUT12), .A3(new_n255), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n413), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n410), .A2(new_n403), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT10), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n395), .A2(new_n398), .A3(new_n391), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT4), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n425), .A2(new_n426), .A3(G101), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(KEYINPUT83), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT83), .ZN(new_n429));
  NAND4_X1  g243(.A1(new_n425), .A2(new_n429), .A3(new_n426), .A4(G101), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n426), .B1(new_n425), .B2(G101), .ZN(new_n431));
  AOI22_X1  g245(.A1(new_n428), .A2(new_n430), .B1(new_n400), .B2(new_n431), .ZN(new_n432));
  AOI22_X1  g246(.A1(new_n423), .A2(new_n424), .B1(new_n252), .B2(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n237), .A2(KEYINPUT10), .A3(new_n403), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n433), .A2(new_n412), .A3(new_n434), .ZN(new_n435));
  AOI21_X1  g249(.A(KEYINPUT82), .B1(new_n422), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n423), .A2(new_n424), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n252), .A2(new_n432), .ZN(new_n438));
  AND4_X1   g252(.A1(new_n412), .A2(new_n437), .A3(new_n438), .A4(new_n434), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n412), .B1(new_n433), .B2(new_n434), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  XNOR2_X1  g255(.A(G110), .B(G140), .ZN(new_n442));
  AND2_X1   g256(.A1(new_n354), .A2(G227), .ZN(new_n443));
  XOR2_X1   g257(.A(new_n442), .B(new_n443), .Z(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  NOR3_X1   g259(.A1(new_n436), .A2(new_n441), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n422), .A2(new_n435), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n444), .B1(new_n447), .B2(KEYINPUT82), .ZN(new_n448));
  OAI21_X1  g262(.A(G469), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  NOR3_X1   g263(.A1(new_n411), .A2(new_n389), .A3(new_n412), .ZN(new_n450));
  AOI21_X1  g264(.A(KEYINPUT12), .B1(new_n420), .B2(new_n255), .ZN(new_n451));
  OAI21_X1  g265(.A(KEYINPUT85), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT85), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n413), .A2(new_n453), .A3(new_n421), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n452), .A2(new_n435), .A3(new_n444), .A4(new_n454), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n445), .B1(new_n439), .B2(new_n440), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(G469), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n457), .A2(new_n458), .A3(new_n289), .ZN(new_n459));
  NAND2_X1  g273(.A1(G469), .A2(G902), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n449), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  XOR2_X1   g275(.A(KEYINPUT9), .B(G234), .Z(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  OAI21_X1  g277(.A(G221), .B1(new_n463), .B2(G902), .ZN(new_n464));
  AND2_X1   g278(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  OAI21_X1  g279(.A(G214), .B1(G237), .B2(G902), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n432), .A2(new_n243), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT5), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n469), .A2(new_n314), .A3(G116), .ZN(new_n470));
  OAI211_X1 g284(.A(G113), .B(new_n470), .C1(new_n241), .C2(new_n469), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n471), .B1(new_n241), .B2(new_n242), .ZN(new_n472));
  OR2_X1    g286(.A1(new_n472), .A2(new_n401), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n468), .A2(new_n473), .ZN(new_n474));
  XOR2_X1   g288(.A(G110), .B(G122), .Z(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(new_n475), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n468), .A2(new_n473), .A3(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n476), .A2(KEYINPUT6), .A3(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(G224), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n480), .A2(G953), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n252), .A2(new_n346), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n237), .A2(G125), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(new_n237), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(new_n346), .ZN(new_n486));
  INV_X1    g300(.A(new_n481), .ZN(new_n487));
  OAI211_X1 g301(.A(new_n486), .B(new_n487), .C1(new_n346), .C2(new_n252), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n484), .A2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT6), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n474), .A2(new_n490), .A3(new_n475), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n479), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n486), .B1(new_n346), .B2(new_n252), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n487), .A2(KEYINPUT7), .ZN(new_n494));
  OAI211_X1 g308(.A(new_n493), .B(new_n494), .C1(KEYINPUT87), .C2(new_n482), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n401), .A2(KEYINPUT86), .ZN(new_n496));
  XOR2_X1   g310(.A(new_n472), .B(new_n496), .Z(new_n497));
  XOR2_X1   g311(.A(new_n475), .B(KEYINPUT8), .Z(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n494), .A2(KEYINPUT87), .ZN(new_n500));
  OAI211_X1 g314(.A(new_n486), .B(new_n500), .C1(new_n346), .C2(new_n252), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n495), .A2(new_n499), .A3(new_n478), .A4(new_n501), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n492), .A2(new_n502), .A3(new_n289), .ZN(new_n503));
  OAI21_X1  g317(.A(G210), .B1(G237), .B2(G902), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n492), .A2(new_n502), .A3(new_n289), .A4(new_n504), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n467), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  AND2_X1   g322(.A1(new_n465), .A2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(G475), .ZN(new_n510));
  AND3_X1   g324(.A1(new_n194), .A2(G143), .A3(G214), .ZN(new_n511));
  AOI21_X1  g325(.A(G143), .B1(new_n194), .B2(G214), .ZN(new_n512));
  OAI211_X1 g326(.A(KEYINPUT18), .B(G131), .C1(new_n511), .C2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(KEYINPUT88), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n194), .A2(G214), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(new_n218), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n194), .A2(G143), .A3(G214), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT88), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n518), .A2(new_n519), .A3(KEYINPUT18), .A4(G131), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n514), .A2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT90), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n348), .A2(G146), .A3(new_n331), .ZN(new_n523));
  AND3_X1   g337(.A1(new_n523), .A2(KEYINPUT89), .A3(new_n338), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n523), .A2(KEYINPUT89), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n522), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n523), .A2(KEYINPUT89), .A3(new_n338), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n527), .B(KEYINPUT90), .C1(KEYINPUT89), .C2(new_n523), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n511), .A2(new_n512), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT18), .ZN(new_n531));
  OAI211_X1 g345(.A(new_n530), .B(KEYINPUT91), .C1(new_n531), .C2(new_n207), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n516), .A2(new_n207), .A3(new_n517), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT91), .ZN(new_n534));
  OAI211_X1 g348(.A(new_n533), .B(new_n534), .C1(new_n518), .C2(KEYINPUT18), .ZN(new_n535));
  NAND4_X1  g349(.A1(new_n521), .A2(new_n529), .A3(new_n532), .A4(new_n535), .ZN(new_n536));
  XNOR2_X1  g350(.A(G113), .B(G122), .ZN(new_n537));
  XNOR2_X1  g351(.A(new_n537), .B(new_n390), .ZN(new_n538));
  INV_X1    g352(.A(new_n351), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n518), .A2(KEYINPUT17), .A3(G131), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n518), .A2(G131), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(new_n533), .ZN(new_n542));
  OAI211_X1 g356(.A(new_n539), .B(new_n540), .C1(new_n542), .C2(KEYINPUT17), .ZN(new_n543));
  AND3_X1   g357(.A1(new_n536), .A2(new_n538), .A3(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n334), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT92), .ZN(new_n546));
  NOR3_X1   g360(.A1(new_n545), .A2(new_n546), .A3(KEYINPUT19), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n348), .A2(new_n331), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n548), .B1(KEYINPUT92), .B2(new_n545), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n547), .B1(new_n549), .B2(KEYINPUT19), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(new_n216), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n542), .A2(new_n337), .A3(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n538), .B1(new_n536), .B2(new_n552), .ZN(new_n553));
  OAI211_X1 g367(.A(new_n510), .B(new_n289), .C1(new_n544), .C2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(KEYINPUT20), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(KEYINPUT93), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT93), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n554), .A2(new_n557), .A3(KEYINPUT20), .ZN(new_n558));
  INV_X1    g372(.A(new_n553), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n536), .A2(new_n543), .A3(new_n538), .ZN(new_n560));
  AOI21_X1  g374(.A(G475), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT20), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n561), .A2(new_n562), .A3(new_n289), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n556), .A2(new_n558), .A3(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n538), .B1(new_n536), .B2(new_n543), .ZN(new_n565));
  OR2_X1    g379(.A1(new_n544), .A2(new_n565), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n510), .B1(new_n566), .B2(new_n289), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n564), .A2(new_n568), .ZN(new_n569));
  NOR3_X1   g383(.A1(new_n463), .A2(new_n366), .A3(G953), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  XNOR2_X1  g385(.A(G128), .B(G143), .ZN(new_n572));
  XNOR2_X1  g386(.A(new_n572), .B(G134), .ZN(new_n573));
  INV_X1    g387(.A(G116), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(G122), .ZN(new_n575));
  INV_X1    g389(.A(G122), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(G116), .ZN(new_n577));
  AND2_X1   g391(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  AND2_X1   g392(.A1(new_n578), .A2(new_n397), .ZN(new_n579));
  OAI21_X1  g393(.A(KEYINPUT14), .B1(new_n576), .B2(G116), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT96), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n575), .A2(KEYINPUT96), .A3(KEYINPUT14), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n582), .A2(new_n577), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(KEYINPUT97), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT97), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n582), .A2(new_n583), .A3(new_n586), .A4(new_n577), .ZN(new_n587));
  OAI211_X1 g401(.A(new_n585), .B(new_n587), .C1(KEYINPUT14), .C2(new_n575), .ZN(new_n588));
  AOI211_X1 g402(.A(new_n573), .B(new_n579), .C1(new_n588), .C2(G107), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n578), .B(G107), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n572), .A2(new_n198), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n591), .B(KEYINPUT95), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n572), .A2(KEYINPUT13), .ZN(new_n593));
  OR3_X1    g407(.A1(new_n234), .A2(KEYINPUT13), .A3(G143), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n593), .A2(G134), .A3(new_n594), .ZN(new_n595));
  OR2_X1    g409(.A1(new_n595), .A2(KEYINPUT94), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(KEYINPUT94), .ZN(new_n597));
  AOI211_X1 g411(.A(new_n590), .B(new_n592), .C1(new_n596), .C2(new_n597), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n571), .B1(new_n589), .B2(new_n598), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n579), .B1(new_n588), .B2(G107), .ZN(new_n600));
  INV_X1    g414(.A(new_n573), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n590), .B1(new_n596), .B2(new_n597), .ZN(new_n603));
  INV_X1    g417(.A(new_n592), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n602), .A2(new_n605), .A3(new_n570), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n599), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(new_n289), .ZN(new_n608));
  INV_X1    g422(.A(G478), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n609), .A2(KEYINPUT15), .ZN(new_n610));
  XOR2_X1   g424(.A(new_n608), .B(new_n610), .Z(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  AND2_X1   g426(.A1(new_n354), .A2(G952), .ZN(new_n613));
  NAND2_X1  g427(.A1(G234), .A2(G237), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  XOR2_X1   g430(.A(KEYINPUT21), .B(G898), .Z(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n614), .A2(G902), .A3(G953), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n616), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  NOR3_X1   g435(.A1(new_n569), .A2(new_n612), .A3(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n388), .A2(new_n509), .A3(new_n622), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n623), .B(KEYINPUT98), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(new_n399), .ZN(G3));
  AOI21_X1  g439(.A(G902), .B1(new_n301), .B2(new_n302), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n308), .B1(new_n626), .B2(new_n187), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n371), .A2(new_n464), .A3(new_n378), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  AOI211_X1 g443(.A(new_n467), .B(new_n621), .C1(new_n506), .C2(new_n507), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n608), .A2(G478), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n609), .A2(new_n289), .ZN(new_n632));
  XNOR2_X1  g446(.A(KEYINPUT99), .B(KEYINPUT33), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n607), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(KEYINPUT100), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n599), .A2(new_n606), .A3(KEYINPUT33), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT100), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n607), .A2(new_n638), .A3(new_n634), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n636), .A2(new_n637), .A3(new_n639), .ZN(new_n640));
  AOI211_X1 g454(.A(new_n631), .B(new_n632), .C1(new_n640), .C2(G478), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n569), .A2(new_n630), .A3(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n629), .A2(new_n643), .A3(new_n461), .ZN(new_n644));
  XOR2_X1   g458(.A(KEYINPUT34), .B(G104), .Z(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G6));
  NAND4_X1  g460(.A1(new_n561), .A2(KEYINPUT101), .A3(new_n562), .A4(new_n289), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT101), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n648), .B1(new_n554), .B2(KEYINPUT20), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n556), .A2(new_n558), .A3(new_n647), .A4(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(new_n568), .ZN(new_n651));
  INV_X1    g465(.A(new_n508), .ZN(new_n652));
  NOR4_X1   g466(.A1(new_n651), .A2(new_n652), .A3(new_n611), .A4(new_n621), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n653), .A2(new_n629), .A3(new_n461), .ZN(new_n654));
  XOR2_X1   g468(.A(KEYINPUT35), .B(G107), .Z(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G9));
  NOR2_X1   g470(.A1(new_n364), .A2(KEYINPUT36), .ZN(new_n657));
  AND2_X1   g471(.A1(new_n363), .A2(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n363), .A2(new_n657), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n368), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n378), .A2(new_n660), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n461), .A2(new_n661), .A3(new_n464), .A4(new_n508), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n627), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(new_n622), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(KEYINPUT37), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(new_n319), .ZN(G12));
  XOR2_X1   g480(.A(KEYINPUT102), .B(G900), .Z(new_n667));
  AOI21_X1  g481(.A(new_n616), .B1(new_n620), .B2(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n650), .A2(new_n612), .A3(new_n568), .A4(new_n669), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n662), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n384), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G128), .ZN(G30));
  NAND2_X1  g487(.A1(new_n506), .A2(new_n507), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(KEYINPUT38), .ZN(new_n675));
  XOR2_X1   g489(.A(new_n668), .B(KEYINPUT39), .Z(new_n676));
  NAND2_X1  g490(.A1(new_n465), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(KEYINPUT104), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT40), .ZN(new_n679));
  AND2_X1   g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n678), .A2(new_n679), .ZN(new_n681));
  OAI211_X1 g495(.A(new_n466), .B(new_n675), .C1(new_n680), .C2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n287), .A2(new_n280), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(new_n289), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n280), .B1(new_n279), .B2(new_n261), .ZN(new_n685));
  OAI21_X1  g499(.A(G472), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n686), .B1(new_n382), .B2(new_n383), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(KEYINPUT103), .ZN(new_n688));
  INV_X1    g502(.A(new_n661), .ZN(new_n689));
  AND3_X1   g503(.A1(new_n554), .A2(new_n557), .A3(KEYINPUT20), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n557), .B1(new_n554), .B2(KEYINPUT20), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n554), .A2(KEYINPUT20), .ZN(new_n692));
  NOR3_X1   g506(.A1(new_n690), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n693), .A2(new_n567), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n694), .A2(new_n611), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n688), .A2(new_n689), .A3(new_n695), .ZN(new_n696));
  OR2_X1    g510(.A1(new_n682), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G143), .ZN(G45));
  OAI211_X1 g512(.A(new_n641), .B(new_n669), .C1(new_n693), .C2(new_n567), .ZN(new_n699));
  NOR3_X1   g513(.A1(new_n311), .A2(new_n662), .A3(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(new_n216), .ZN(G48));
  NOR2_X1   g515(.A1(new_n311), .A2(new_n379), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT107), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT105), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n704), .A2(new_n458), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n706), .B1(new_n457), .B2(new_n289), .ZN(new_n707));
  AOI211_X1 g521(.A(G902), .B(new_n705), .C1(new_n455), .C2(new_n456), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  AOI21_X1  g523(.A(KEYINPUT106), .B1(new_n709), .B2(new_n464), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT106), .ZN(new_n711));
  INV_X1    g525(.A(new_n464), .ZN(new_n712));
  NOR4_X1   g526(.A1(new_n707), .A2(new_n708), .A3(new_n711), .A4(new_n712), .ZN(new_n713));
  OAI21_X1  g527(.A(new_n703), .B1(new_n710), .B2(new_n713), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n457), .A2(new_n289), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(new_n705), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n457), .A2(new_n289), .A3(new_n706), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n716), .A2(new_n464), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(new_n711), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n709), .A2(KEYINPUT106), .A3(new_n464), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n719), .A2(new_n720), .A3(KEYINPUT107), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n714), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n702), .A2(new_n643), .A3(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(KEYINPUT41), .B(G113), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n723), .B(new_n724), .ZN(G15));
  NAND3_X1  g539(.A1(new_n702), .A2(new_n653), .A3(new_n722), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G116), .ZN(G18));
  NOR3_X1   g541(.A1(new_n710), .A2(new_n713), .A3(new_n652), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n384), .A2(new_n728), .A3(new_n622), .A4(new_n661), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G119), .ZN(G21));
  OAI21_X1  g544(.A(new_n269), .B1(new_n287), .B2(new_n197), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(new_n280), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n294), .B1(new_n301), .B2(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT108), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n734), .B1(new_n626), .B2(new_n187), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n307), .A2(new_n289), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n736), .A2(KEYINPUT108), .A3(G472), .ZN(new_n737));
  AOI211_X1 g551(.A(new_n379), .B(new_n733), .C1(new_n735), .C2(new_n737), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n722), .A2(new_n738), .A3(new_n630), .A4(new_n695), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G122), .ZN(G24));
  AOI21_X1  g554(.A(new_n733), .B1(new_n735), .B2(new_n737), .ZN(new_n741));
  INV_X1    g555(.A(new_n699), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n728), .A2(new_n741), .A3(new_n661), .A4(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G125), .ZN(G27));
  INV_X1    g558(.A(KEYINPUT42), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n506), .A2(new_n466), .A3(new_n507), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT109), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n746), .B(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n465), .A2(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(new_n749), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n750), .A2(new_n384), .A3(new_n742), .A4(new_n386), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n308), .B(KEYINPUT32), .ZN(new_n752));
  AOI211_X1 g566(.A(new_n745), .B(new_n379), .C1(new_n752), .C2(new_n381), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n749), .A2(new_n699), .ZN(new_n754));
  AOI22_X1  g568(.A1(new_n745), .A2(new_n751), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(new_n207), .ZN(G33));
  NOR4_X1   g570(.A1(new_n311), .A2(new_n749), .A3(new_n379), .A4(new_n670), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(new_n198), .ZN(G36));
  INV_X1    g572(.A(new_n748), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT111), .ZN(new_n760));
  OAI211_X1 g574(.A(new_n694), .B(new_n641), .C1(new_n760), .C2(KEYINPUT43), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n641), .A2(new_n564), .A3(new_n568), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT43), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n564), .A2(new_n760), .A3(new_n568), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n762), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n761), .A2(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n766), .A2(new_n627), .A3(new_n661), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT44), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  OR2_X1    g583(.A1(new_n769), .A2(KEYINPUT112), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(KEYINPUT112), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n759), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT110), .ZN(new_n773));
  OAI21_X1  g587(.A(KEYINPUT45), .B1(new_n446), .B2(new_n448), .ZN(new_n774));
  OR2_X1    g588(.A1(new_n439), .A2(new_n440), .ZN(new_n775));
  AND2_X1   g589(.A1(new_n422), .A2(new_n435), .ZN(new_n776));
  OAI211_X1 g590(.A(new_n775), .B(new_n444), .C1(new_n776), .C2(KEYINPUT82), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT45), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT82), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n445), .B1(new_n776), .B2(new_n779), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n777), .A2(new_n778), .A3(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n774), .A2(new_n781), .A3(G469), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n782), .A2(new_n460), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT46), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n773), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n783), .A2(new_n784), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n782), .A2(KEYINPUT110), .A3(KEYINPUT46), .A4(new_n460), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n785), .A2(new_n786), .A3(new_n459), .A4(new_n787), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n788), .A2(new_n464), .A3(new_n676), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n789), .B1(new_n768), .B2(new_n767), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n772), .A2(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(G137), .ZN(G39));
  NAND2_X1  g606(.A1(new_n788), .A2(new_n464), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT47), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n788), .A2(KEYINPUT47), .A3(new_n464), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n797), .A2(new_n742), .A3(new_n748), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n311), .A2(new_n379), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(new_n327), .ZN(G42));
  NOR2_X1   g615(.A1(new_n628), .A2(new_n467), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(KEYINPUT113), .ZN(new_n803));
  INV_X1    g617(.A(new_n762), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT49), .ZN(new_n805));
  OAI211_X1 g619(.A(new_n803), .B(new_n804), .C1(new_n805), .C2(new_n709), .ZN(new_n806));
  XOR2_X1   g620(.A(new_n806), .B(KEYINPUT114), .Z(new_n807));
  INV_X1    g621(.A(new_n675), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n688), .B1(new_n805), .B2(new_n709), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n807), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n709), .A2(new_n712), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n795), .A2(new_n796), .A3(new_n811), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n615), .B1(new_n761), .B2(new_n765), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n813), .A2(new_n738), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n812), .A2(new_n748), .A3(new_n814), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n688), .A2(new_n379), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n710), .A2(new_n713), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT118), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n817), .A2(new_n818), .A3(new_n748), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n748), .A2(new_n719), .A3(new_n720), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n615), .B1(new_n820), .B2(KEYINPUT118), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n569), .A2(new_n641), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n816), .A2(new_n819), .A3(new_n821), .A4(new_n822), .ZN(new_n823));
  AND2_X1   g637(.A1(new_n815), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n821), .A2(new_n766), .A3(new_n819), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT119), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n821), .A2(KEYINPUT119), .A3(new_n766), .A4(new_n819), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n829), .A2(new_n661), .A3(new_n741), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n675), .A2(new_n466), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n813), .A2(new_n817), .A3(new_n738), .A4(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT50), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n832), .B(new_n833), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n824), .A2(KEYINPUT51), .A3(new_n830), .A4(new_n834), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n830), .A2(new_n834), .A3(new_n815), .A4(new_n823), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT51), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n835), .A2(new_n613), .A3(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n814), .A2(new_n728), .ZN(new_n840));
  AND2_X1   g654(.A1(new_n739), .A2(new_n723), .ZN(new_n841));
  AND2_X1   g655(.A1(new_n726), .A2(new_n729), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n751), .A2(new_n745), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n753), .A2(new_n754), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n841), .A2(new_n842), .A3(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n741), .A2(new_n742), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n650), .A2(new_n611), .A3(new_n568), .A4(new_n669), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n847), .B1(new_n848), .B2(new_n311), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n749), .A2(new_n689), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n757), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n630), .A2(new_n564), .A3(new_n612), .A4(new_n568), .ZN(new_n852));
  OR2_X1    g666(.A1(new_n852), .A2(KEYINPUT115), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(KEYINPUT115), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n853), .A2(new_n854), .A3(new_n461), .A4(new_n629), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n855), .A2(new_n644), .A3(new_n664), .ZN(new_n856));
  INV_X1    g670(.A(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n851), .A2(new_n623), .A3(new_n857), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n846), .A2(new_n858), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n699), .A2(new_n662), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n384), .B1(new_n860), .B2(new_n671), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n661), .A2(new_n668), .ZN(new_n862));
  AND3_X1   g676(.A1(new_n569), .A2(new_n508), .A3(new_n612), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n687), .A2(new_n465), .A3(new_n862), .A4(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n743), .A2(new_n861), .A3(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT52), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n743), .A2(new_n861), .A3(new_n864), .A4(KEYINPUT52), .ZN(new_n868));
  AOI21_X1  g682(.A(KEYINPUT53), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n859), .A2(new_n869), .ZN(new_n870));
  AND4_X1   g684(.A1(new_n723), .A2(new_n739), .A3(new_n726), .A4(new_n729), .ZN(new_n871));
  INV_X1    g685(.A(new_n622), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n872), .B1(new_n380), .B2(new_n387), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n856), .B1(new_n873), .B2(new_n509), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n871), .A2(new_n874), .A3(new_n845), .A4(new_n851), .ZN(new_n875));
  AOI21_X1  g689(.A(KEYINPUT116), .B1(new_n867), .B2(new_n868), .ZN(new_n876));
  AND3_X1   g690(.A1(new_n867), .A2(KEYINPUT116), .A3(new_n868), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT53), .ZN(new_n879));
  OAI211_X1 g693(.A(KEYINPUT54), .B(new_n870), .C1(new_n878), .C2(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT54), .ZN(new_n881));
  INV_X1    g695(.A(new_n858), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n723), .A2(new_n739), .A3(new_n726), .A4(new_n729), .ZN(new_n883));
  OAI21_X1  g697(.A(KEYINPUT117), .B1(new_n883), .B2(new_n755), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT117), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n841), .A2(new_n842), .A3(new_n845), .A4(new_n885), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n879), .B1(new_n867), .B2(new_n868), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n882), .A2(new_n884), .A3(new_n886), .A4(new_n887), .ZN(new_n888));
  OAI211_X1 g702(.A(new_n881), .B(new_n888), .C1(new_n878), .C2(KEYINPUT53), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n839), .A2(new_n840), .A3(new_n880), .A4(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n816), .A2(new_n819), .A3(new_n821), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n569), .A2(new_n641), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n752), .A2(new_n381), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n894), .A2(new_n386), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n895), .B1(new_n827), .B2(new_n828), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n896), .B(KEYINPUT48), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n890), .A2(new_n893), .A3(new_n897), .ZN(new_n898));
  NOR2_X1   g712(.A1(G952), .A2(G953), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n810), .B1(new_n898), .B2(new_n899), .ZN(G75));
  NOR2_X1   g714(.A1(new_n354), .A2(G952), .ZN(new_n901));
  INV_X1    g715(.A(new_n901), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n877), .A2(new_n876), .ZN(new_n903));
  AOI21_X1  g717(.A(KEYINPUT53), .B1(new_n903), .B2(new_n859), .ZN(new_n904));
  AND4_X1   g718(.A1(new_n882), .A2(new_n884), .A3(new_n886), .A4(new_n887), .ZN(new_n905));
  OAI211_X1 g719(.A(G210), .B(G902), .C1(new_n904), .C2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT56), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT120), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n902), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n479), .A2(new_n491), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n911), .B(new_n489), .ZN(new_n912));
  XOR2_X1   g726(.A(new_n912), .B(KEYINPUT55), .Z(new_n913));
  AOI21_X1  g727(.A(new_n913), .B1(new_n908), .B2(new_n909), .ZN(new_n914));
  INV_X1    g728(.A(new_n913), .ZN(new_n915));
  AOI211_X1 g729(.A(KEYINPUT120), .B(new_n915), .C1(new_n906), .C2(new_n907), .ZN(new_n916));
  NOR3_X1   g730(.A1(new_n910), .A2(new_n914), .A3(new_n916), .ZN(G51));
  OAI21_X1  g731(.A(KEYINPUT54), .B1(new_n904), .B2(new_n905), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT121), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n918), .A2(new_n919), .A3(new_n889), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n904), .A2(new_n905), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n921), .A2(KEYINPUT121), .A3(new_n881), .ZN(new_n922));
  XOR2_X1   g736(.A(new_n460), .B(KEYINPUT57), .Z(new_n923));
  NAND3_X1  g737(.A1(new_n920), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n924), .A2(new_n457), .ZN(new_n925));
  OR3_X1    g739(.A1(new_n921), .A2(new_n289), .A3(new_n782), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n901), .B1(new_n925), .B2(new_n926), .ZN(G54));
  OAI21_X1  g741(.A(new_n888), .B1(new_n878), .B2(KEYINPUT53), .ZN(new_n928));
  AND3_X1   g742(.A1(new_n928), .A2(KEYINPUT58), .A3(G902), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT122), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n544), .A2(new_n553), .ZN(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n929), .A2(new_n930), .A3(G475), .A4(new_n932), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n928), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n901), .B1(new_n934), .B2(new_n931), .ZN(new_n935));
  OAI21_X1  g749(.A(KEYINPUT122), .B1(new_n934), .B2(new_n931), .ZN(new_n936));
  AND3_X1   g750(.A1(new_n933), .A2(new_n935), .A3(new_n936), .ZN(G60));
  XNOR2_X1  g751(.A(new_n632), .B(KEYINPUT59), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n938), .B1(new_n880), .B2(new_n889), .ZN(new_n939));
  INV_X1    g753(.A(new_n640), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n902), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n920), .A2(new_n922), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n942), .A2(new_n938), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n941), .B1(new_n943), .B2(new_n940), .ZN(G63));
  INV_X1    g758(.A(new_n365), .ZN(new_n945));
  XNOR2_X1  g759(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n366), .A2(new_n289), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n946), .B(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(new_n948), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n945), .B1(new_n921), .B2(new_n949), .ZN(new_n950));
  OAI211_X1 g764(.A(new_n928), .B(new_n948), .C1(new_n658), .C2(new_n659), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n950), .A2(new_n951), .A3(new_n902), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT61), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n950), .A2(new_n951), .A3(KEYINPUT61), .A4(new_n902), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(new_n955), .ZN(G66));
  NAND2_X1  g770(.A1(new_n871), .A2(new_n874), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n957), .A2(new_n354), .ZN(new_n958));
  OAI21_X1  g772(.A(G953), .B1(new_n618), .B2(new_n480), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n911), .B1(G898), .B2(new_n354), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n960), .B(new_n961), .ZN(G69));
  AOI21_X1  g776(.A(new_n800), .B1(new_n772), .B2(new_n790), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n789), .A2(new_n895), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(new_n863), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n743), .A2(new_n861), .ZN(new_n966));
  NOR3_X1   g780(.A1(new_n755), .A2(new_n757), .A3(new_n966), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n963), .A2(new_n354), .A3(new_n965), .A4(new_n967), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n276), .B1(KEYINPUT30), .B2(new_n265), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n969), .B(new_n550), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n970), .B1(G900), .B2(G953), .ZN(new_n971));
  AOI21_X1  g785(.A(KEYINPUT126), .B1(new_n968), .B2(new_n971), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n354), .B1(G227), .B2(G900), .ZN(new_n973));
  XOR2_X1   g787(.A(new_n973), .B(KEYINPUT127), .Z(new_n974));
  NOR2_X1   g788(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(new_n800), .ZN(new_n976));
  INV_X1    g790(.A(new_n966), .ZN(new_n977));
  NAND2_X1  g791(.A1(KEYINPUT124), .A2(KEYINPUT62), .ZN(new_n978));
  OAI211_X1 g792(.A(new_n977), .B(new_n978), .C1(new_n682), .C2(new_n696), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n892), .B1(new_n611), .B2(new_n569), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n980), .A2(new_n748), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n678), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n982), .A2(new_n388), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n983), .B(KEYINPUT125), .ZN(new_n984));
  NAND4_X1  g798(.A1(new_n791), .A2(new_n976), .A3(new_n979), .A4(new_n984), .ZN(new_n985));
  OR2_X1    g799(.A1(KEYINPUT124), .A2(KEYINPUT62), .ZN(new_n986));
  AOI22_X1  g800(.A1(new_n697), .A2(new_n977), .B1(new_n978), .B2(new_n986), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n354), .B1(new_n985), .B2(new_n987), .ZN(new_n988));
  AOI22_X1  g802(.A1(new_n988), .A2(new_n970), .B1(new_n968), .B2(new_n971), .ZN(new_n989));
  XNOR2_X1  g803(.A(new_n975), .B(new_n989), .ZN(G72));
  NOR3_X1   g804(.A1(new_n985), .A2(new_n987), .A3(new_n957), .ZN(new_n991));
  NAND2_X1  g805(.A1(G472), .A2(G902), .ZN(new_n992));
  XOR2_X1   g806(.A(new_n992), .B(KEYINPUT63), .Z(new_n993));
  INV_X1    g807(.A(new_n993), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n685), .B1(new_n991), .B2(new_n994), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n963), .A2(new_n965), .A3(new_n967), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n993), .B1(new_n996), .B2(new_n957), .ZN(new_n997));
  INV_X1    g811(.A(new_n281), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NOR3_X1   g813(.A1(new_n998), .A2(new_n685), .A3(new_n994), .ZN(new_n1000));
  OAI211_X1 g814(.A(new_n870), .B(new_n1000), .C1(new_n878), .C2(new_n879), .ZN(new_n1001));
  AND4_X1   g815(.A1(new_n902), .A2(new_n995), .A3(new_n999), .A4(new_n1001), .ZN(G57));
endmodule


