//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 0 0 0 0 1 1 0 1 1 1 1 0 1 0 0 1 1 0 1 1 0 1 1 1 0 0 0 1 0 1 0 0 0 1 0 1 1 1 1 0 1 1 1 1 1 1 0 0 1 0 0 1 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:40 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n446, new_n448, new_n449, new_n451, new_n454, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n560, new_n561, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n576,
    new_n577, new_n578, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n609,
    new_n612, new_n613, new_n615, new_n616, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n897, new_n898, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1148,
    new_n1149;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT64), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT65), .Z(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  NAND2_X1  g020(.A1(G94), .A2(G452), .ZN(new_n446));
  XNOR2_X1  g021(.A(new_n446), .B(KEYINPUT66), .ZN(G173));
  XNOR2_X1  g022(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n448));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n448), .B(new_n449), .ZN(G223));
  INV_X1    g025(.A(new_n449), .ZN(new_n451));
  NAND2_X1  g026(.A1(new_n451), .A2(G567), .ZN(G234));
  NAND2_X1  g027(.A1(new_n451), .A2(G2106), .ZN(G217));
  NOR4_X1   g028(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT2), .Z(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AOI22_X1  g034(.A1(new_n455), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  OAI211_X1 g037(.A(KEYINPUT68), .B(new_n461), .C1(new_n462), .C2(KEYINPUT69), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT68), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT69), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n464), .B1(new_n465), .B2(G2104), .ZN(new_n466));
  OAI21_X1  g041(.A(KEYINPUT3), .B1(new_n462), .B2(KEYINPUT68), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n463), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  AND2_X1   g044(.A1(new_n469), .A2(G137), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n462), .A2(G2105), .ZN(new_n471));
  AOI22_X1  g046(.A1(new_n468), .A2(new_n470), .B1(G101), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n461), .A2(G2104), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n473), .A2(new_n474), .A3(G125), .ZN(new_n475));
  NAND2_X1  g050(.A1(G113), .A2(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n472), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G160));
  AOI21_X1  g055(.A(new_n461), .B1(new_n464), .B2(G2104), .ZN(new_n481));
  OAI21_X1  g056(.A(KEYINPUT68), .B1(new_n462), .B2(KEYINPUT69), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g058(.A(G2105), .B1(new_n483), .B2(new_n463), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G136), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n469), .B1(new_n483), .B2(new_n463), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G124), .ZN(new_n487));
  INV_X1    g062(.A(G100), .ZN(new_n488));
  AND3_X1   g063(.A1(new_n488), .A2(new_n469), .A3(KEYINPUT70), .ZN(new_n489));
  AOI21_X1  g064(.A(KEYINPUT70), .B1(new_n488), .B2(new_n469), .ZN(new_n490));
  OAI221_X1 g065(.A(G2104), .B1(G112), .B2(new_n469), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n485), .A2(new_n487), .A3(new_n491), .ZN(new_n492));
  XNOR2_X1  g067(.A(new_n492), .B(KEYINPUT71), .ZN(G162));
  NAND3_X1  g068(.A1(new_n468), .A2(G126), .A3(G2105), .ZN(new_n494));
  OAI21_X1  g069(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n495));
  INV_X1    g070(.A(G114), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n495), .B1(new_n496), .B2(G2105), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n469), .A2(G138), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n499), .B1(new_n468), .B2(new_n501), .ZN(new_n502));
  XNOR2_X1  g077(.A(KEYINPUT3), .B(G2104), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n503), .A2(new_n499), .A3(new_n501), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(new_n505));
  OAI211_X1 g080(.A(new_n494), .B(new_n498), .C1(new_n502), .C2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(G164));
  NAND2_X1  g082(.A1(G75), .A2(G543), .ZN(new_n508));
  XNOR2_X1  g083(.A(new_n508), .B(KEYINPUT74), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT72), .ZN(new_n510));
  INV_X1    g085(.A(G543), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n510), .B1(new_n511), .B2(KEYINPUT5), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT5), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n513), .A2(KEYINPUT72), .A3(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n511), .A2(KEYINPUT5), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(G62), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n509), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  AND2_X1   g094(.A1(KEYINPUT6), .A2(G651), .ZN(new_n520));
  NOR2_X1   g095(.A1(KEYINPUT6), .A2(G651), .ZN(new_n521));
  OAI21_X1  g096(.A(G543), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(new_n522), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n519), .A2(G651), .B1(G50), .B2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(G88), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n520), .A2(new_n521), .ZN(new_n526));
  OAI21_X1  g101(.A(KEYINPUT73), .B1(new_n517), .B2(new_n526), .ZN(new_n527));
  AOI22_X1  g102(.A1(new_n512), .A2(new_n514), .B1(KEYINPUT5), .B2(new_n511), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT73), .ZN(new_n529));
  OAI211_X1 g104(.A(new_n528), .B(new_n529), .C1(new_n521), .C2(new_n520), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n527), .A2(new_n530), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n524), .B1(new_n525), .B2(new_n531), .ZN(G303));
  INV_X1    g107(.A(G303), .ZN(G166));
  NAND3_X1  g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  XOR2_X1   g109(.A(new_n534), .B(KEYINPUT7), .Z(new_n535));
  AND3_X1   g110(.A1(new_n528), .A2(G63), .A3(G651), .ZN(new_n536));
  AOI211_X1 g111(.A(new_n535), .B(new_n536), .C1(G51), .C2(new_n523), .ZN(new_n537));
  INV_X1    g112(.A(new_n531), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G89), .ZN(new_n539));
  AND2_X1   g114(.A1(new_n537), .A2(new_n539), .ZN(G168));
  NAND3_X1  g115(.A1(new_n527), .A2(new_n530), .A3(G90), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n523), .A2(G52), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(KEYINPUT75), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT75), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n541), .A2(new_n545), .A3(new_n542), .ZN(new_n546));
  NAND2_X1  g121(.A1(G77), .A2(G543), .ZN(new_n547));
  INV_X1    g122(.A(G64), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n547), .B1(new_n517), .B2(new_n548), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n544), .A2(new_n546), .B1(G651), .B2(new_n549), .ZN(G171));
  NAND2_X1  g125(.A1(new_n538), .A2(G81), .ZN(new_n551));
  NAND2_X1  g126(.A1(G68), .A2(G543), .ZN(new_n552));
  INV_X1    g127(.A(G56), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n552), .B1(new_n517), .B2(new_n553), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n554), .A2(G651), .B1(G43), .B2(new_n523), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n551), .A2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G860), .ZN(G153));
  NAND4_X1  g133(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND4_X1  g136(.A1(G319), .A2(G483), .A3(G661), .A4(new_n561), .ZN(G188));
  NAND2_X1  g137(.A1(G78), .A2(G543), .ZN(new_n563));
  INV_X1    g138(.A(G65), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n563), .B1(new_n517), .B2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT9), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(KEYINPUT76), .ZN(new_n567));
  OAI21_X1  g142(.A(G53), .B1(new_n566), .B2(KEYINPUT76), .ZN(new_n568));
  OR3_X1    g143(.A1(new_n522), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n567), .B1(new_n522), .B2(new_n568), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n565), .A2(G651), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n527), .A2(new_n530), .A3(G91), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n571), .A2(new_n572), .ZN(G299));
  INV_X1    g148(.A(G171), .ZN(G301));
  INV_X1    g149(.A(G168), .ZN(G286));
  OR2_X1    g150(.A1(new_n528), .A2(G74), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n576), .A2(G651), .B1(G49), .B2(new_n523), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n527), .A2(new_n530), .A3(G87), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(G288));
  NAND2_X1  g154(.A1(G73), .A2(G543), .ZN(new_n580));
  INV_X1    g155(.A(G61), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n517), .B2(new_n581), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n582), .A2(G651), .B1(G48), .B2(new_n523), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n527), .A2(new_n530), .A3(G86), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n583), .A2(KEYINPUT77), .A3(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(new_n586));
  AOI21_X1  g161(.A(KEYINPUT77), .B1(new_n583), .B2(new_n584), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n586), .A2(new_n587), .ZN(G305));
  NAND2_X1  g163(.A1(G72), .A2(G543), .ZN(new_n589));
  INV_X1    g164(.A(G60), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n517), .B2(new_n590), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n591), .A2(G651), .B1(G47), .B2(new_n523), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n527), .A2(new_n530), .A3(G85), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(new_n593), .ZN(G290));
  NAND2_X1  g169(.A1(new_n523), .A2(G54), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n528), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n596));
  INV_X1    g171(.A(G651), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n595), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT78), .ZN(new_n599));
  XNOR2_X1  g174(.A(new_n598), .B(new_n599), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n527), .A2(new_n530), .A3(G92), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT10), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n601), .B(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(G868), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n606), .B1(new_n605), .B2(G171), .ZN(G321));
  XNOR2_X1  g182(.A(G321), .B(KEYINPUT79), .ZN(G284));
  XOR2_X1   g183(.A(G299), .B(KEYINPUT80), .Z(new_n609));
  MUX2_X1   g184(.A(G286), .B(new_n609), .S(new_n605), .Z(G297));
  MUX2_X1   g185(.A(G286), .B(new_n609), .S(new_n605), .Z(G280));
  INV_X1    g186(.A(new_n604), .ZN(new_n612));
  INV_X1    g187(.A(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n613), .B2(G860), .ZN(G148));
  NAND2_X1  g189(.A1(new_n612), .A2(new_n613), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n615), .A2(G868), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n616), .B1(G868), .B2(new_n557), .ZN(G323));
  XNOR2_X1  g192(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g193(.A1(new_n503), .A2(new_n471), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT12), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT13), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(G2100), .ZN(new_n622));
  INV_X1    g197(.A(KEYINPUT81), .ZN(new_n623));
  AND3_X1   g198(.A1(new_n486), .A2(new_n623), .A3(G123), .ZN(new_n624));
  AOI21_X1  g199(.A(new_n623), .B1(new_n486), .B2(G123), .ZN(new_n625));
  OR2_X1    g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  OAI21_X1  g201(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n627));
  INV_X1    g202(.A(G111), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n627), .B1(new_n628), .B2(G2105), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n629), .B1(new_n484), .B2(G135), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n626), .A2(new_n630), .ZN(new_n631));
  OR2_X1    g206(.A1(new_n631), .A2(G2096), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n631), .A2(G2096), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n622), .A2(new_n632), .A3(new_n633), .ZN(G156));
  XOR2_X1   g209(.A(G1341), .B(G1348), .Z(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT83), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT82), .B(KEYINPUT16), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  INV_X1    g213(.A(KEYINPUT14), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2427), .B(G2438), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2430), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT15), .B(G2435), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n639), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n643), .B1(new_n642), .B2(new_n641), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n638), .B(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(G2451), .B(G2454), .Z(new_n646));
  XNOR2_X1  g221(.A(G2443), .B(G2446), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  OR2_X1    g223(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n645), .A2(new_n648), .ZN(new_n650));
  AND3_X1   g225(.A1(new_n649), .A2(G14), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT84), .ZN(G401));
  XOR2_X1   g227(.A(G2072), .B(G2078), .Z(new_n653));
  XOR2_X1   g228(.A(new_n653), .B(KEYINPUT17), .Z(new_n654));
  XNOR2_X1  g229(.A(G2067), .B(G2678), .ZN(new_n655));
  XOR2_X1   g230(.A(G2084), .B(G2090), .Z(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  NOR3_X1   g232(.A1(new_n654), .A2(new_n655), .A3(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT86), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n654), .A2(new_n655), .ZN(new_n660));
  INV_X1    g235(.A(new_n653), .ZN(new_n661));
  OAI211_X1 g236(.A(new_n660), .B(new_n657), .C1(new_n661), .C2(new_n655), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n661), .A2(new_n655), .A3(new_n656), .ZN(new_n663));
  XOR2_X1   g238(.A(KEYINPUT85), .B(KEYINPUT18), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n659), .A2(new_n662), .A3(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(G2096), .B(G2100), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(G227));
  XOR2_X1   g243(.A(G1961), .B(G1966), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT87), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1956), .B(G2474), .ZN(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1971), .B(G1976), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT19), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n676), .B(KEYINPUT20), .Z(new_n677));
  NOR2_X1   g252(.A1(new_n670), .A2(new_n672), .ZN(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n679), .A2(new_n675), .A3(new_n673), .ZN(new_n680));
  OAI211_X1 g255(.A(new_n677), .B(new_n680), .C1(new_n675), .C2(new_n679), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1991), .B(G1996), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1981), .B(G1986), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(G229));
  NAND2_X1  g262(.A1(G305), .A2(G16), .ZN(new_n688));
  INV_X1    g263(.A(G16), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n689), .A2(G6), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT32), .B(G1981), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  XOR2_X1   g268(.A(KEYINPUT90), .B(G16), .Z(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n695), .A2(G22), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(G166), .B2(new_n695), .ZN(new_n697));
  INV_X1    g272(.A(G1971), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  OR2_X1    g274(.A1(new_n691), .A2(new_n692), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n689), .A2(G23), .ZN(new_n701));
  INV_X1    g276(.A(G288), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n701), .B1(new_n702), .B2(new_n689), .ZN(new_n703));
  XNOR2_X1  g278(.A(KEYINPUT33), .B(G1976), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  AND4_X1   g280(.A1(new_n693), .A2(new_n699), .A3(new_n700), .A4(new_n705), .ZN(new_n706));
  XOR2_X1   g281(.A(KEYINPUT91), .B(KEYINPUT34), .Z(new_n707));
  OR2_X1    g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n706), .A2(new_n707), .ZN(new_n709));
  INV_X1    g284(.A(G29), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(G25), .ZN(new_n711));
  OR2_X1    g286(.A1(G95), .A2(G2105), .ZN(new_n712));
  OAI211_X1 g287(.A(new_n712), .B(G2104), .C1(G107), .C2(new_n469), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT88), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n484), .A2(G131), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n486), .A2(G119), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n714), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(KEYINPUT89), .Z(new_n718));
  INV_X1    g293(.A(new_n718), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n711), .B1(new_n719), .B2(new_n710), .ZN(new_n720));
  XOR2_X1   g295(.A(KEYINPUT35), .B(G1991), .Z(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n695), .A2(G24), .ZN(new_n723));
  INV_X1    g298(.A(G290), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n723), .B1(new_n724), .B2(new_n695), .ZN(new_n725));
  INV_X1    g300(.A(G1986), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n725), .B(new_n726), .ZN(new_n727));
  NAND4_X1  g302(.A1(new_n708), .A2(new_n709), .A3(new_n722), .A4(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(KEYINPUT36), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n728), .B(new_n729), .ZN(new_n730));
  NOR2_X1   g305(.A1(G5), .A2(G16), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(KEYINPUT97), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(G301), .B2(new_n689), .ZN(new_n733));
  INV_X1    g308(.A(G1961), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT98), .ZN(new_n736));
  NAND3_X1  g311(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT95), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT26), .ZN(new_n739));
  AOI22_X1  g314(.A1(new_n484), .A2(G141), .B1(G105), .B2(new_n471), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n486), .A2(G129), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n739), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n743), .A2(new_n710), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(new_n710), .B2(G32), .ZN(new_n745));
  XNOR2_X1  g320(.A(KEYINPUT27), .B(G1996), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n710), .A2(G27), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(KEYINPUT99), .Z(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G164), .B2(new_n710), .ZN(new_n749));
  XOR2_X1   g324(.A(KEYINPUT100), .B(G2078), .Z(new_n750));
  AOI22_X1  g325(.A1(new_n745), .A2(new_n746), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(KEYINPUT30), .ZN(new_n752));
  AND2_X1   g327(.A1(new_n752), .A2(G28), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n710), .B1(new_n752), .B2(G28), .ZN(new_n754));
  AND2_X1   g329(.A1(KEYINPUT31), .A2(G11), .ZN(new_n755));
  NOR2_X1   g330(.A1(KEYINPUT31), .A2(G11), .ZN(new_n756));
  OAI22_X1  g331(.A1(new_n753), .A2(new_n754), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(new_n631), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n757), .B1(new_n758), .B2(G29), .ZN(new_n759));
  OAI211_X1 g334(.A(new_n751), .B(new_n759), .C1(new_n749), .C2(new_n750), .ZN(new_n760));
  INV_X1    g335(.A(G34), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n761), .A2(KEYINPUT24), .ZN(new_n762));
  AOI21_X1  g337(.A(G29), .B1(new_n761), .B2(KEYINPUT24), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n762), .B1(new_n763), .B2(KEYINPUT93), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(KEYINPUT93), .B2(new_n763), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(new_n479), .B2(new_n710), .ZN(new_n766));
  INV_X1    g341(.A(G2084), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT94), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(new_n745), .B2(new_n746), .ZN(new_n770));
  NOR2_X1   g345(.A1(new_n760), .A2(new_n770), .ZN(new_n771));
  AND2_X1   g346(.A1(new_n710), .A2(G33), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n484), .A2(G139), .ZN(new_n773));
  NAND3_X1  g348(.A1(new_n469), .A2(G103), .A3(G2104), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(KEYINPUT25), .Z(new_n775));
  AOI22_X1  g350(.A1(new_n503), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n776));
  OAI211_X1 g351(.A(new_n773), .B(new_n775), .C1(new_n469), .C2(new_n776), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n772), .B1(new_n777), .B2(G29), .ZN(new_n778));
  INV_X1    g353(.A(G2072), .ZN(new_n779));
  AOI22_X1  g354(.A1(new_n778), .A2(new_n779), .B1(new_n767), .B2(new_n766), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(new_n779), .B2(new_n778), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n710), .A2(G26), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(KEYINPUT28), .Z(new_n783));
  NAND2_X1  g358(.A1(new_n484), .A2(G140), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n486), .A2(G128), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n469), .A2(G116), .ZN(new_n786));
  OAI21_X1  g361(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n787));
  OAI211_X1 g362(.A(new_n784), .B(new_n785), .C1(new_n786), .C2(new_n787), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n783), .B1(new_n788), .B2(G29), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(G2067), .ZN(new_n790));
  XNOR2_X1  g365(.A(KEYINPUT101), .B(G1956), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n694), .A2(G20), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(KEYINPUT23), .Z(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(G299), .B2(G16), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n790), .B1(new_n791), .B2(new_n794), .ZN(new_n795));
  AOI211_X1 g370(.A(new_n781), .B(new_n795), .C1(new_n791), .C2(new_n794), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n694), .A2(G19), .ZN(new_n797));
  XOR2_X1   g372(.A(new_n797), .B(KEYINPUT92), .Z(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(new_n556), .B2(new_n695), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(G1341), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n689), .A2(G21), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(G168), .B2(new_n689), .ZN(new_n802));
  XOR2_X1   g377(.A(KEYINPUT96), .B(G1966), .Z(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NAND4_X1  g379(.A1(new_n771), .A2(new_n796), .A3(new_n800), .A4(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n710), .A2(G35), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(G162), .B2(new_n710), .ZN(new_n807));
  XOR2_X1   g382(.A(new_n807), .B(KEYINPUT29), .Z(new_n808));
  INV_X1    g383(.A(G2090), .ZN(new_n809));
  AOI22_X1  g384(.A1(new_n808), .A2(new_n809), .B1(new_n734), .B2(new_n733), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n689), .A2(G4), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(new_n612), .B2(new_n689), .ZN(new_n812));
  XOR2_X1   g387(.A(new_n812), .B(G1348), .Z(new_n813));
  OAI211_X1 g388(.A(new_n810), .B(new_n813), .C1(new_n809), .C2(new_n808), .ZN(new_n814));
  NOR4_X1   g389(.A1(new_n730), .A2(new_n736), .A3(new_n805), .A4(new_n814), .ZN(G311));
  OR4_X1    g390(.A1(new_n730), .A2(new_n736), .A3(new_n805), .A4(new_n814), .ZN(G150));
  NOR2_X1   g391(.A1(new_n604), .A2(new_n613), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT38), .ZN(new_n818));
  NAND2_X1  g393(.A1(G80), .A2(G543), .ZN(new_n819));
  INV_X1    g394(.A(G67), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n819), .B1(new_n517), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n821), .A2(G651), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT102), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n821), .A2(KEYINPUT102), .A3(G651), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n523), .A2(G55), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n527), .A2(new_n530), .A3(G93), .ZN(new_n827));
  NAND4_X1  g402(.A1(new_n824), .A2(new_n825), .A3(new_n826), .A4(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n557), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n556), .A2(new_n828), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n818), .B(new_n832), .ZN(new_n833));
  AND2_X1   g408(.A1(new_n833), .A2(KEYINPUT39), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n833), .A2(KEYINPUT39), .ZN(new_n835));
  NOR3_X1   g410(.A1(new_n834), .A2(new_n835), .A3(G860), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n828), .A2(G860), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT37), .ZN(new_n838));
  OR2_X1    g413(.A1(new_n836), .A2(new_n838), .ZN(G145));
  XNOR2_X1  g414(.A(new_n788), .B(new_n506), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(new_n743), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(new_n777), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n717), .B(new_n620), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n486), .A2(G130), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n469), .A2(G118), .ZN(new_n845));
  OAI21_X1  g420(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n844), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n847), .B1(G142), .B2(new_n484), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n843), .B(new_n848), .ZN(new_n849));
  OR2_X1    g424(.A1(new_n842), .A2(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n631), .B(new_n479), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(G162), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n842), .A2(new_n849), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n850), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(KEYINPUT104), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT103), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n853), .A2(new_n856), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n857), .A2(new_n852), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n850), .A2(new_n856), .A3(new_n853), .ZN(new_n859));
  AOI21_X1  g434(.A(G37), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n855), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g437(.A(new_n702), .B(G303), .ZN(new_n863));
  NOR3_X1   g438(.A1(new_n586), .A2(new_n724), .A3(new_n587), .ZN(new_n864));
  INV_X1    g439(.A(new_n587), .ZN(new_n865));
  AOI21_X1  g440(.A(G290), .B1(new_n865), .B2(new_n585), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n863), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  NOR3_X1   g443(.A1(new_n863), .A2(new_n864), .A3(new_n866), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n870), .B1(KEYINPUT105), .B2(KEYINPUT42), .ZN(new_n871));
  NAND2_X1  g446(.A1(KEYINPUT105), .A2(KEYINPUT42), .ZN(new_n872));
  XOR2_X1   g447(.A(new_n872), .B(KEYINPUT106), .Z(new_n873));
  OR2_X1    g448(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n871), .A2(new_n873), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n615), .B(new_n832), .ZN(new_n877));
  INV_X1    g452(.A(G299), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n600), .A2(new_n603), .A3(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n878), .B1(new_n600), .B2(new_n603), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  AND2_X1   g458(.A1(new_n877), .A2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n881), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n885), .A2(KEYINPUT41), .A3(new_n879), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT41), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n887), .B1(new_n880), .B2(new_n881), .ZN(new_n888));
  AND2_X1   g463(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n877), .A2(new_n889), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n884), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n876), .A2(new_n891), .ZN(new_n892));
  OAI211_X1 g467(.A(new_n874), .B(new_n875), .C1(new_n884), .C2(new_n890), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n605), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n829), .A2(G868), .ZN(new_n895));
  OR2_X1    g470(.A1(new_n894), .A2(new_n895), .ZN(G295));
  NAND2_X1  g471(.A1(G295), .A2(KEYINPUT107), .ZN(new_n897));
  OR3_X1    g472(.A1(new_n894), .A2(KEYINPUT107), .A3(new_n895), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(G331));
  INV_X1    g474(.A(KEYINPUT44), .ZN(new_n900));
  INV_X1    g475(.A(new_n831), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n556), .A2(new_n828), .ZN(new_n902));
  OAI21_X1  g477(.A(G171), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND3_X1  g478(.A1(G301), .A2(new_n830), .A3(new_n831), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(G286), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n903), .A2(new_n904), .A3(G168), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n889), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  AND3_X1   g483(.A1(new_n903), .A2(new_n904), .A3(G168), .ZN(new_n909));
  AOI21_X1  g484(.A(G168), .B1(new_n903), .B2(new_n904), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n882), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n908), .A2(new_n911), .A3(new_n870), .ZN(new_n912));
  INV_X1    g487(.A(G37), .ZN(new_n913));
  AND2_X1   g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n908), .A2(new_n911), .ZN(new_n915));
  INV_X1    g490(.A(new_n869), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT108), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n916), .A2(new_n917), .A3(new_n867), .ZN(new_n918));
  OAI21_X1  g493(.A(KEYINPUT108), .B1(new_n868), .B2(new_n869), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT109), .ZN(new_n922));
  AND3_X1   g497(.A1(new_n915), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n922), .B1(new_n915), .B2(new_n921), .ZN(new_n924));
  OAI211_X1 g499(.A(new_n914), .B(KEYINPUT43), .C1(new_n923), .C2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT43), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n912), .A2(new_n913), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n920), .B1(new_n911), .B2(new_n908), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n926), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n900), .B1(new_n925), .B2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  OAI211_X1 g506(.A(new_n914), .B(new_n926), .C1(new_n923), .C2(new_n924), .ZN(new_n932));
  OAI21_X1  g507(.A(KEYINPUT43), .B1(new_n927), .B2(new_n928), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(new_n900), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT110), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n931), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  AOI21_X1  g512(.A(KEYINPUT44), .B1(new_n932), .B2(new_n933), .ZN(new_n938));
  OAI21_X1  g513(.A(KEYINPUT110), .B1(new_n930), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n937), .A2(new_n939), .ZN(G397));
  INV_X1    g515(.A(G1384), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n468), .A2(new_n501), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n505), .B1(new_n942), .B2(KEYINPUT4), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n494), .A2(new_n498), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n941), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT45), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n468), .A2(new_n470), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n471), .A2(G101), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n476), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n952), .B1(new_n503), .B2(G125), .ZN(new_n953));
  OAI21_X1  g528(.A(G40), .B1(new_n953), .B2(new_n469), .ZN(new_n954));
  OAI21_X1  g529(.A(KEYINPUT111), .B1(new_n951), .B2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(G40), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n956), .B1(new_n477), .B2(G2105), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT111), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n957), .A2(new_n472), .A3(new_n958), .ZN(new_n959));
  AND2_X1   g534(.A1(new_n955), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n948), .A2(new_n960), .ZN(new_n961));
  XOR2_X1   g536(.A(new_n788), .B(G2067), .Z(new_n962));
  AOI21_X1  g537(.A(new_n961), .B1(new_n962), .B2(new_n743), .ZN(new_n963));
  OR3_X1    g538(.A1(new_n961), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n964));
  OAI21_X1  g539(.A(KEYINPUT46), .B1(new_n961), .B2(G1996), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n963), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  XNOR2_X1  g541(.A(new_n966), .B(KEYINPUT47), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n962), .A2(new_n961), .ZN(new_n968));
  XNOR2_X1  g543(.A(new_n968), .B(KEYINPUT113), .ZN(new_n969));
  INV_X1    g544(.A(G1996), .ZN(new_n970));
  NOR3_X1   g545(.A1(new_n961), .A2(new_n970), .A3(new_n743), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(new_n961), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n973), .A2(new_n970), .A3(new_n743), .ZN(new_n974));
  XNOR2_X1  g549(.A(new_n974), .B(KEYINPUT112), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n972), .A2(new_n719), .A3(new_n721), .A4(new_n975), .ZN(new_n976));
  OR2_X1    g551(.A1(new_n788), .A2(G2067), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n961), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n972), .A2(new_n975), .ZN(new_n979));
  XOR2_X1   g554(.A(new_n717), .B(new_n721), .Z(new_n980));
  AOI21_X1  g555(.A(new_n979), .B1(new_n973), .B2(new_n980), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n973), .A2(new_n726), .A3(new_n724), .ZN(new_n982));
  XNOR2_X1  g557(.A(new_n982), .B(KEYINPUT48), .ZN(new_n983));
  AOI211_X1 g558(.A(new_n967), .B(new_n978), .C1(new_n981), .C2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n583), .A2(new_n584), .ZN(new_n985));
  OR2_X1    g560(.A1(new_n985), .A2(G1981), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(G1981), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT49), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n986), .A2(KEYINPUT49), .A3(new_n987), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n955), .A2(new_n506), .A3(new_n941), .A4(new_n959), .ZN(new_n992));
  AND2_X1   g567(.A1(new_n992), .A2(G8), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n990), .A2(new_n991), .A3(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n702), .A2(G1976), .ZN(new_n995));
  INV_X1    g570(.A(G1976), .ZN(new_n996));
  AOI21_X1  g571(.A(KEYINPUT52), .B1(G288), .B2(new_n996), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n993), .A2(new_n995), .A3(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n993), .A2(new_n995), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(KEYINPUT52), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n994), .A2(new_n998), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT114), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n994), .A2(new_n998), .A3(KEYINPUT114), .A4(new_n1000), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(G8), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n500), .B1(new_n483), .B2(new_n463), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n504), .B1(new_n1007), .B2(new_n499), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n497), .B1(new_n486), .B2(G126), .ZN(new_n1009));
  AOI21_X1  g584(.A(G1384), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT50), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n945), .A2(KEYINPUT50), .ZN(new_n1013));
  AND3_X1   g588(.A1(new_n1012), .A2(new_n960), .A3(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(new_n809), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n506), .A2(KEYINPUT45), .A3(new_n941), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n960), .A2(new_n947), .A3(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(new_n698), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1006), .B1(new_n1015), .B2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(G303), .A2(G8), .ZN(new_n1020));
  XOR2_X1   g595(.A(new_n1020), .B(KEYINPUT55), .Z(new_n1021));
  AND2_X1   g596(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1005), .A2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g598(.A1(G288), .A2(G1976), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n994), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(new_n986), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(KEYINPUT115), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(new_n993), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n1026), .A2(KEYINPUT115), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1023), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT63), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1032));
  OR3_X1    g607(.A1(new_n1022), .A2(new_n1032), .A3(new_n1001), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1012), .A2(new_n960), .A3(new_n1013), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1034), .A2(G2084), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT116), .ZN(new_n1036));
  AOI22_X1  g611(.A1(new_n1035), .A2(new_n1036), .B1(new_n803), .B2(new_n1017), .ZN(new_n1037));
  OAI21_X1  g612(.A(KEYINPUT116), .B1(new_n1034), .B2(G2084), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1039), .A2(G8), .A3(G168), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1031), .B1(new_n1033), .B2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1040), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1042));
  NOR3_X1   g617(.A1(new_n1022), .A2(new_n1032), .A3(new_n1031), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1030), .B1(new_n1041), .B2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(G168), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1014), .A2(new_n1036), .A3(new_n767), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1017), .A2(new_n803), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1047), .A2(new_n1038), .A3(G168), .A4(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(G8), .ZN(new_n1050));
  OAI21_X1  g625(.A(KEYINPUT51), .B1(new_n1046), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT62), .ZN(new_n1052));
  OAI211_X1 g627(.A(new_n1051), .B(new_n1052), .C1(KEYINPUT51), .C2(new_n1050), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT53), .ZN(new_n1054));
  OR3_X1    g629(.A1(new_n1017), .A2(new_n1054), .A3(G2078), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1054), .B1(new_n1017), .B2(G2078), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1034), .A2(new_n734), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1055), .A2(new_n1056), .A3(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(G171), .ZN(new_n1059));
  NOR4_X1   g634(.A1(new_n1022), .A2(new_n1059), .A3(new_n1032), .A4(new_n1001), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1053), .A2(KEYINPUT127), .A3(new_n1060), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1051), .B1(KEYINPUT51), .B2(new_n1050), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(KEYINPUT62), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(KEYINPUT127), .B1(new_n1053), .B2(new_n1060), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1045), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n947), .A2(new_n1016), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n957), .A2(new_n472), .ZN(new_n1068));
  AOI211_X1 g643(.A(new_n1054), .B(G2078), .C1(new_n1068), .C2(KEYINPUT124), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1069), .B1(KEYINPUT124), .B2(new_n1068), .ZN(new_n1070));
  OAI211_X1 g645(.A(new_n1056), .B(new_n1057), .C1(new_n1067), .C2(new_n1070), .ZN(new_n1071));
  OR2_X1    g646(.A1(new_n1071), .A2(G171), .ZN(new_n1072));
  AOI21_X1  g647(.A(KEYINPUT54), .B1(new_n1072), .B2(new_n1059), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1033), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1071), .A2(G171), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT125), .ZN(new_n1076));
  XNOR2_X1  g651(.A(new_n1075), .B(new_n1076), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1055), .A2(G301), .A3(new_n1056), .A4(new_n1057), .ZN(new_n1078));
  AND2_X1   g653(.A1(new_n1078), .A2(KEYINPUT54), .ZN(new_n1079));
  AOI21_X1  g654(.A(KEYINPUT126), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1081));
  AOI21_X1  g656(.A(KEYINPUT125), .B1(new_n1071), .B2(G171), .ZN(new_n1082));
  OAI211_X1 g657(.A(KEYINPUT126), .B(new_n1079), .C1(new_n1081), .C2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1083), .ZN(new_n1084));
  OAI211_X1 g659(.A(new_n1062), .B(new_n1074), .C1(new_n1080), .C2(new_n1084), .ZN(new_n1085));
  NOR2_X1   g660(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT57), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1087), .B1(new_n571), .B2(new_n572), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1011), .B1(new_n506), .B2(new_n941), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n955), .A2(new_n959), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(G1956), .B1(new_n1093), .B2(new_n1012), .ZN(new_n1094));
  XNOR2_X1  g669(.A(KEYINPUT56), .B(G2072), .ZN(new_n1095));
  AND4_X1   g670(.A1(new_n960), .A2(new_n947), .A3(new_n1016), .A4(new_n1095), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1090), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT117), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n992), .A2(new_n1098), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1010), .A2(KEYINPUT117), .A3(new_n955), .A4(new_n959), .ZN(new_n1100));
  AOI21_X1  g675(.A(G2067), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT118), .ZN(new_n1102));
  OAI22_X1  g677(.A1(new_n1101), .A2(new_n1102), .B1(new_n1014), .B2(G1348), .ZN(new_n1103));
  AND2_X1   g678(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1097), .B1(new_n1105), .B2(new_n604), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n960), .A2(new_n947), .A3(new_n1016), .A4(new_n1095), .ZN(new_n1107));
  OAI211_X1 g682(.A(new_n1089), .B(new_n1107), .C1(new_n1014), .C2(G1956), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1106), .A2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n604), .B1(new_n1105), .B2(KEYINPUT60), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT60), .ZN(new_n1111));
  NOR4_X1   g686(.A1(new_n1103), .A2(new_n1104), .A3(new_n1111), .A4(new_n612), .ZN(new_n1112));
  OAI22_X1  g687(.A1(new_n1110), .A2(new_n1112), .B1(KEYINPUT60), .B2(new_n1105), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT61), .ZN(new_n1114));
  AND3_X1   g689(.A1(new_n1097), .A2(new_n1114), .A3(new_n1108), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1114), .B1(new_n1097), .B2(new_n1108), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  XOR2_X1   g692(.A(KEYINPUT58), .B(G1341), .Z(new_n1118));
  NAND3_X1  g693(.A1(new_n1099), .A2(new_n1100), .A3(new_n1118), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n960), .A2(new_n947), .A3(new_n970), .A4(new_n1016), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT119), .ZN(new_n1122));
  AND3_X1   g697(.A1(new_n1122), .A2(KEYINPUT120), .A3(KEYINPUT59), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1121), .A2(new_n557), .A3(new_n1123), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n556), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1124), .B1(new_n1122), .B2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g701(.A(KEYINPUT59), .B1(new_n1125), .B2(KEYINPUT120), .ZN(new_n1127));
  OAI21_X1  g702(.A(KEYINPUT121), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1121), .A2(KEYINPUT120), .A3(new_n557), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT59), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  OR2_X1    g706(.A1(new_n1125), .A2(new_n1122), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT121), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1131), .A2(new_n1132), .A3(new_n1133), .A4(new_n1124), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1117), .B1(new_n1128), .B2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT122), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1113), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  AOI211_X1 g712(.A(KEYINPUT122), .B(new_n1117), .C1(new_n1134), .C2(new_n1128), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1109), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1085), .B1(new_n1139), .B2(KEYINPUT123), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT123), .ZN(new_n1141));
  OAI211_X1 g716(.A(new_n1141), .B(new_n1109), .C1(new_n1137), .C2(new_n1138), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1066), .B1(new_n1140), .B2(new_n1142), .ZN(new_n1143));
  XNOR2_X1  g718(.A(G290), .B(new_n726), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n981), .B1(new_n961), .B2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n984), .B1(new_n1143), .B2(new_n1145), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g721(.A(G319), .ZN(new_n1148));
  NOR4_X1   g722(.A1(G229), .A2(new_n1148), .A3(new_n651), .A4(G227), .ZN(new_n1149));
  NAND3_X1  g723(.A1(new_n1149), .A2(new_n861), .A3(new_n934), .ZN(G225));
  INV_X1    g724(.A(G225), .ZN(G308));
endmodule


