//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 0 0 0 1 1 1 1 1 0 1 0 1 1 1 1 1 1 1 1 0 0 1 0 0 0 0 0 0 1 0 1 0 1 1 0 0 1 1 0 0 0 1 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:59 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n450, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n533, new_n534,
    new_n535, new_n536, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n550, new_n552,
    new_n553, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n578, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n610, new_n611, new_n612, new_n615, new_n617, new_n618, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1171, new_n1172,
    new_n1173;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT64), .Z(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  XNOR2_X1  g039(.A(new_n464), .B(KEYINPUT65), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  AOI22_X1  g046(.A1(G101), .A2(new_n465), .B1(new_n471), .B2(G137), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  INV_X1    g048(.A(G125), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n473), .B1(new_n470), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n472), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G160));
  XNOR2_X1  g053(.A(KEYINPUT3), .B(G2104), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G2105), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n471), .A2(G136), .ZN(new_n483));
  OR2_X1    g058(.A1(G100), .A2(G2105), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n484), .B(G2104), .C1(G112), .C2(new_n463), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n482), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G162));
  NAND4_X1  g062(.A1(new_n467), .A2(new_n469), .A3(KEYINPUT4), .A4(G138), .ZN(new_n488));
  NAND2_X1  g063(.A1(G102), .A2(G2104), .ZN(new_n489));
  AOI21_X1  g064(.A(G2105), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(G114), .A2(G2104), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n492), .B1(new_n479), .B2(G126), .ZN(new_n493));
  OAI21_X1  g068(.A(KEYINPUT4), .B1(new_n493), .B2(new_n463), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n479), .A2(G138), .A3(new_n463), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n490), .B1(new_n494), .B2(new_n495), .ZN(G164));
  INV_X1    g071(.A(KEYINPUT66), .ZN(new_n497));
  INV_X1    g072(.A(G543), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n497), .B1(new_n498), .B2(KEYINPUT5), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT5), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n500), .A2(KEYINPUT66), .A3(G543), .ZN(new_n501));
  AOI22_X1  g076(.A1(new_n499), .A2(new_n501), .B1(KEYINPUT5), .B2(new_n498), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G62), .ZN(new_n503));
  NAND2_X1  g078(.A1(G75), .A2(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G651), .ZN(new_n506));
  AND2_X1   g081(.A1(KEYINPUT6), .A2(G651), .ZN(new_n507));
  NOR2_X1   g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(new_n510));
  AND2_X1   g085(.A1(new_n502), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G88), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n509), .A2(new_n498), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G50), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n506), .A2(new_n512), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(KEYINPUT67), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n502), .A2(new_n510), .ZN(new_n517));
  INV_X1    g092(.A(G88), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n514), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(G651), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n520), .B1(new_n503), .B2(new_n504), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT67), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n516), .A2(new_n524), .ZN(G166));
  NAND2_X1  g100(.A1(new_n511), .A2(G89), .ZN(new_n526));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n527), .B(KEYINPUT7), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n502), .A2(G63), .A3(G651), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n513), .A2(G51), .ZN(new_n530));
  NAND4_X1  g105(.A1(new_n526), .A2(new_n528), .A3(new_n529), .A4(new_n530), .ZN(G286));
  INV_X1    g106(.A(G286), .ZN(G168));
  AOI22_X1  g107(.A1(new_n502), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n533));
  OR2_X1    g108(.A1(new_n533), .A2(new_n520), .ZN(new_n534));
  XOR2_X1   g109(.A(KEYINPUT68), .B(G90), .Z(new_n535));
  AOI22_X1  g110(.A1(new_n511), .A2(new_n535), .B1(G52), .B2(new_n513), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n534), .A2(new_n536), .ZN(G301));
  INV_X1    g112(.A(G301), .ZN(G171));
  XOR2_X1   g113(.A(KEYINPUT70), .B(G81), .Z(new_n539));
  NAND2_X1  g114(.A1(new_n511), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n513), .A2(G43), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n502), .A2(G56), .ZN(new_n542));
  INV_X1    g117(.A(G68), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n542), .B1(new_n543), .B2(new_n498), .ZN(new_n544));
  AND3_X1   g119(.A1(new_n544), .A2(KEYINPUT69), .A3(G651), .ZN(new_n545));
  AOI21_X1  g120(.A(KEYINPUT69), .B1(new_n544), .B2(G651), .ZN(new_n546));
  OAI211_X1 g121(.A(new_n540), .B(new_n541), .C1(new_n545), .C2(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  AND3_X1   g124(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G36), .ZN(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n550), .A2(new_n553), .ZN(G188));
  OAI211_X1 g129(.A(G53), .B(G543), .C1(new_n507), .C2(new_n508), .ZN(new_n555));
  XOR2_X1   g130(.A(KEYINPUT71), .B(KEYINPUT9), .Z(new_n556));
  OR2_X1    g131(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT72), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n555), .A2(KEYINPUT9), .ZN(new_n560));
  AND2_X1   g135(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  OAI211_X1 g136(.A(KEYINPUT73), .B(new_n559), .C1(new_n561), .C2(new_n558), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT73), .ZN(new_n563));
  INV_X1    g138(.A(new_n559), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n558), .B1(new_n557), .B2(new_n560), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n563), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n562), .A2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(new_n567), .ZN(new_n568));
  AOI22_X1  g143(.A1(new_n502), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n569));
  OR2_X1    g144(.A1(new_n569), .A2(new_n520), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT74), .ZN(new_n571));
  INV_X1    g146(.A(G91), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n571), .B1(new_n517), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n511), .A2(KEYINPUT74), .A3(G91), .ZN(new_n574));
  AND3_X1   g149(.A1(new_n570), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n568), .A2(new_n575), .ZN(G299));
  INV_X1    g151(.A(G166), .ZN(G303));
  NAND2_X1  g152(.A1(new_n511), .A2(G87), .ZN(new_n578));
  OAI21_X1  g153(.A(G651), .B1(new_n502), .B2(G74), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n513), .A2(G49), .ZN(new_n580));
  AND3_X1   g155(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(G288));
  NAND2_X1  g157(.A1(new_n513), .A2(G48), .ZN(new_n583));
  INV_X1    g158(.A(G86), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n517), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n502), .A2(G61), .ZN(new_n586));
  NAND2_X1  g161(.A1(G73), .A2(G543), .ZN(new_n587));
  XNOR2_X1  g162(.A(new_n587), .B(KEYINPUT75), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n520), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n585), .A2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(G305));
  XNOR2_X1  g166(.A(KEYINPUT76), .B(G47), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n511), .A2(G85), .B1(new_n513), .B2(new_n592), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n502), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n520), .B2(new_n594), .ZN(G290));
  NAND2_X1  g170(.A1(G301), .A2(G868), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n511), .A2(G92), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT10), .ZN(new_n598));
  XNOR2_X1  g173(.A(new_n597), .B(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n513), .A2(G54), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n502), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n601));
  OR2_X1    g176(.A1(new_n601), .A2(new_n520), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n599), .A2(new_n600), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n603), .A2(KEYINPUT77), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT77), .ZN(new_n605));
  NAND4_X1  g180(.A1(new_n599), .A2(new_n605), .A3(new_n600), .A4(new_n602), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n596), .B1(new_n607), .B2(G868), .ZN(G284));
  OAI21_X1  g183(.A(new_n596), .B1(new_n607), .B2(G868), .ZN(G321));
  NAND2_X1  g184(.A1(G286), .A2(G868), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n570), .A2(new_n573), .A3(new_n574), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n567), .A2(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n610), .B1(new_n612), .B2(G868), .ZN(G297));
  XNOR2_X1  g188(.A(G297), .B(KEYINPUT78), .ZN(G280));
  INV_X1    g189(.A(G559), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n607), .B1(new_n615), .B2(G860), .ZN(G148));
  NAND2_X1  g191(.A1(new_n607), .A2(new_n615), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n617), .A2(G868), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n618), .B1(G868), .B2(new_n548), .ZN(G323));
  XNOR2_X1  g194(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g195(.A1(new_n465), .A2(new_n479), .ZN(new_n621));
  XNOR2_X1  g196(.A(KEYINPUT79), .B(KEYINPUT12), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n621), .B(new_n622), .ZN(new_n623));
  XOR2_X1   g198(.A(KEYINPUT13), .B(G2100), .Z(new_n624));
  XNOR2_X1  g199(.A(new_n623), .B(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n481), .A2(G123), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n471), .A2(G135), .ZN(new_n627));
  NOR2_X1   g202(.A1(G99), .A2(G2105), .ZN(new_n628));
  OAI21_X1  g203(.A(G2104), .B1(new_n463), .B2(G111), .ZN(new_n629));
  OAI211_X1 g204(.A(new_n626), .B(new_n627), .C1(new_n628), .C2(new_n629), .ZN(new_n630));
  XOR2_X1   g205(.A(new_n630), .B(G2096), .Z(new_n631));
  NAND2_X1  g206(.A1(new_n625), .A2(new_n631), .ZN(G156));
  XNOR2_X1  g207(.A(G2427), .B(G2438), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2430), .ZN(new_n634));
  XOR2_X1   g209(.A(KEYINPUT15), .B(G2435), .Z(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n636), .A2(KEYINPUT14), .ZN(new_n637));
  XOR2_X1   g212(.A(G2451), .B(G2454), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2443), .B(G2446), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(KEYINPUT16), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n639), .B(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(G1341), .B(G1348), .Z(new_n643));
  INV_X1    g218(.A(new_n643), .ZN(new_n644));
  AND2_X1   g219(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n645), .A2(KEYINPUT80), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n642), .A2(new_n644), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n645), .A2(KEYINPUT80), .ZN(new_n648));
  NAND4_X1  g223(.A1(new_n646), .A2(G14), .A3(new_n647), .A4(new_n648), .ZN(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(G401));
  XOR2_X1   g225(.A(G2084), .B(G2090), .Z(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(G2067), .B(G2678), .Z(new_n653));
  OR2_X1    g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n652), .A2(new_n653), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n654), .A2(new_n655), .A3(KEYINPUT17), .ZN(new_n656));
  INV_X1    g231(.A(KEYINPUT18), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(G2096), .B(G2100), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(G2072), .B(G2078), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT81), .ZN(new_n662));
  AOI21_X1  g237(.A(new_n662), .B1(KEYINPUT18), .B2(new_n654), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n660), .B(new_n663), .Z(G227));
  XOR2_X1   g239(.A(G1956), .B(G2474), .Z(new_n665));
  XOR2_X1   g240(.A(G1961), .B(G1966), .Z(new_n666));
  NOR2_X1   g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1971), .B(G1976), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT19), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n671), .B(KEYINPUT82), .Z(new_n672));
  NAND2_X1  g247(.A1(new_n665), .A2(new_n666), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(new_n674), .B(KEYINPUT20), .Z(new_n675));
  NAND3_X1  g250(.A1(new_n668), .A2(new_n670), .A3(new_n673), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n672), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1991), .B(G1996), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1981), .B(G1986), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n677), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT83), .ZN(new_n683));
  XOR2_X1   g258(.A(new_n681), .B(new_n683), .Z(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(G229));
  OR2_X1    g260(.A1(G5), .A2(G16), .ZN(new_n686));
  INV_X1    g261(.A(G16), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n686), .B1(G301), .B2(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(G1961), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT93), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n688), .A2(new_n689), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT92), .B(G2067), .ZN(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT91), .B(KEYINPUT28), .ZN(new_n694));
  INV_X1    g269(.A(G29), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n695), .A2(G26), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n694), .B(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n471), .A2(G140), .ZN(new_n698));
  OR2_X1    g273(.A1(G104), .A2(G2105), .ZN(new_n699));
  OAI211_X1 g274(.A(new_n699), .B(G2104), .C1(G116), .C2(new_n463), .ZN(new_n700));
  INV_X1    g275(.A(G128), .ZN(new_n701));
  OAI211_X1 g276(.A(new_n698), .B(new_n700), .C1(new_n701), .C2(new_n480), .ZN(new_n702));
  OR2_X1    g277(.A1(new_n702), .A2(KEYINPUT90), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n702), .A2(KEYINPUT90), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n697), .B1(new_n705), .B2(G29), .ZN(new_n706));
  OAI211_X1 g281(.A(new_n691), .B(new_n692), .C1(new_n693), .C2(new_n706), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n708));
  XOR2_X1   g283(.A(new_n708), .B(KEYINPUT25), .Z(new_n709));
  NAND2_X1  g284(.A1(new_n471), .A2(G139), .ZN(new_n710));
  AOI22_X1  g285(.A1(new_n479), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n711));
  OAI211_X1 g286(.A(new_n709), .B(new_n710), .C1(new_n463), .C2(new_n711), .ZN(new_n712));
  MUX2_X1   g287(.A(G33), .B(new_n712), .S(G29), .Z(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(G2072), .ZN(new_n714));
  INV_X1    g289(.A(G28), .ZN(new_n715));
  AOI21_X1  g290(.A(G29), .B1(new_n715), .B2(KEYINPUT30), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(KEYINPUT30), .B2(new_n715), .ZN(new_n717));
  AND2_X1   g292(.A1(KEYINPUT24), .A2(G34), .ZN(new_n718));
  NOR2_X1   g293(.A1(KEYINPUT24), .A2(G34), .ZN(new_n719));
  NOR3_X1   g294(.A1(new_n718), .A2(new_n719), .A3(G29), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(new_n477), .B2(G29), .ZN(new_n721));
  INV_X1    g296(.A(G2084), .ZN(new_n722));
  OAI221_X1 g297(.A(new_n717), .B1(new_n695), .B2(new_n630), .C1(new_n721), .C2(new_n722), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n714), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n687), .A2(G21), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(G168), .B2(new_n687), .ZN(new_n726));
  INV_X1    g301(.A(G1966), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  XNOR2_X1  g303(.A(KEYINPUT31), .B(G11), .ZN(new_n729));
  AOI22_X1  g304(.A1(new_n706), .A2(new_n693), .B1(new_n722), .B2(new_n721), .ZN(new_n730));
  NAND4_X1  g305(.A1(new_n724), .A2(new_n728), .A3(new_n729), .A4(new_n730), .ZN(new_n731));
  NOR2_X1   g306(.A1(G29), .A2(G32), .ZN(new_n732));
  AOI22_X1  g307(.A1(G105), .A2(new_n465), .B1(new_n471), .B2(G141), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n481), .A2(G129), .ZN(new_n734));
  NAND3_X1  g309(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(KEYINPUT26), .Z(new_n736));
  NAND3_X1  g311(.A1(new_n733), .A2(new_n734), .A3(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(new_n737), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n732), .B1(new_n738), .B2(G29), .ZN(new_n739));
  XOR2_X1   g314(.A(KEYINPUT27), .B(G1996), .Z(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n695), .A2(G27), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G164), .B2(new_n695), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(G2078), .ZN(new_n744));
  NOR4_X1   g319(.A1(new_n707), .A2(new_n731), .A3(new_n741), .A4(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n695), .A2(G35), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(G162), .B2(new_n695), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(KEYINPUT29), .Z(new_n748));
  INV_X1    g323(.A(G2090), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g325(.A1(G4), .A2(G16), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(new_n607), .B2(G16), .ZN(new_n752));
  XOR2_X1   g327(.A(KEYINPUT87), .B(G1348), .Z(new_n753));
  XNOR2_X1  g328(.A(new_n752), .B(new_n753), .ZN(new_n754));
  AND3_X1   g329(.A1(new_n745), .A2(new_n750), .A3(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(KEYINPUT94), .ZN(new_n756));
  INV_X1    g331(.A(KEYINPUT23), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(G299), .B2(G16), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n687), .A2(G20), .ZN(new_n759));
  MUX2_X1   g334(.A(new_n757), .B(new_n758), .S(new_n759), .Z(new_n760));
  INV_X1    g335(.A(G1956), .ZN(new_n761));
  OR2_X1    g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n760), .A2(new_n761), .ZN(new_n763));
  OAI211_X1 g338(.A(new_n762), .B(new_n763), .C1(new_n749), .C2(new_n748), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n755), .B1(new_n756), .B2(new_n764), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(new_n756), .B2(new_n764), .ZN(new_n766));
  INV_X1    g341(.A(G19), .ZN(new_n767));
  OAI21_X1  g342(.A(KEYINPUT88), .B1(new_n767), .B2(G16), .ZN(new_n768));
  OR3_X1    g343(.A1(new_n767), .A2(KEYINPUT88), .A3(G16), .ZN(new_n769));
  OAI211_X1 g344(.A(new_n768), .B(new_n769), .C1(new_n548), .C2(new_n687), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT89), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(G1341), .ZN(new_n772));
  NAND2_X1  g347(.A1(G166), .A2(G16), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G16), .B2(G22), .ZN(new_n774));
  XNOR2_X1  g349(.A(KEYINPUT86), .B(G1971), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n687), .A2(G23), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(new_n581), .B2(new_n687), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT33), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(G1976), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n687), .A2(G6), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(new_n590), .B2(new_n687), .ZN(new_n782));
  XNOR2_X1  g357(.A(KEYINPUT32), .B(G1981), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  INV_X1    g359(.A(new_n784), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n776), .A2(new_n780), .A3(new_n785), .ZN(new_n786));
  OR2_X1    g361(.A1(new_n786), .A2(KEYINPUT34), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n481), .A2(G119), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n471), .A2(G131), .ZN(new_n789));
  NOR2_X1   g364(.A1(G95), .A2(G2105), .ZN(new_n790));
  OAI21_X1  g365(.A(G2104), .B1(new_n463), .B2(G107), .ZN(new_n791));
  OAI211_X1 g366(.A(new_n788), .B(new_n789), .C1(new_n790), .C2(new_n791), .ZN(new_n792));
  MUX2_X1   g367(.A(G25), .B(new_n792), .S(G29), .Z(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT84), .ZN(new_n794));
  XNOR2_X1  g369(.A(KEYINPUT35), .B(G1991), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n794), .B(new_n795), .Z(new_n796));
  NOR2_X1   g371(.A1(G16), .A2(G24), .ZN(new_n797));
  XOR2_X1   g372(.A(G290), .B(KEYINPUT85), .Z(new_n798));
  AOI21_X1  g373(.A(new_n797), .B1(new_n798), .B2(G16), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(G1986), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n800), .B1(new_n786), .B2(KEYINPUT34), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n787), .A2(new_n796), .A3(new_n801), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT36), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n766), .A2(new_n772), .A3(new_n803), .ZN(G150));
  INV_X1    g379(.A(G150), .ZN(G311));
  AOI22_X1  g380(.A1(new_n511), .A2(G93), .B1(G55), .B2(new_n513), .ZN(new_n806));
  INV_X1    g381(.A(KEYINPUT95), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  AOI22_X1  g383(.A1(new_n502), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n809));
  OR2_X1    g384(.A1(new_n809), .A2(new_n520), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  XOR2_X1   g386(.A(KEYINPUT96), .B(G860), .Z(new_n812));
  NAND2_X1  g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n813), .B(KEYINPUT37), .Z(new_n814));
  INV_X1    g389(.A(KEYINPUT39), .ZN(new_n815));
  AND2_X1   g390(.A1(new_n604), .A2(new_n606), .ZN(new_n816));
  OAI21_X1  g391(.A(KEYINPUT38), .B1(new_n816), .B2(new_n615), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT38), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n607), .A2(new_n818), .A3(G559), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(new_n811), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n821), .A2(new_n547), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n811), .A2(new_n548), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n820), .A2(new_n824), .ZN(new_n825));
  NAND4_X1  g400(.A1(new_n817), .A2(new_n823), .A3(new_n822), .A4(new_n819), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n815), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  AND2_X1   g402(.A1(new_n827), .A2(KEYINPUT97), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n825), .A2(new_n815), .A3(new_n826), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n829), .B1(new_n827), .B2(KEYINPUT97), .ZN(new_n830));
  NOR3_X1   g405(.A1(new_n828), .A2(new_n830), .A3(new_n812), .ZN(new_n831));
  AND2_X1   g406(.A1(new_n831), .A2(KEYINPUT98), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n831), .A2(KEYINPUT98), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n814), .B1(new_n832), .B2(new_n833), .ZN(G145));
  XNOR2_X1  g409(.A(new_n623), .B(KEYINPUT102), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n792), .B(KEYINPUT101), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n835), .B(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n481), .A2(G130), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n471), .A2(G142), .ZN(new_n839));
  OR2_X1    g414(.A1(G106), .A2(G2105), .ZN(new_n840));
  OAI211_X1 g415(.A(new_n840), .B(G2104), .C1(G118), .C2(new_n463), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n838), .A2(new_n839), .A3(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n837), .B(new_n843), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n467), .A2(new_n469), .A3(G126), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n463), .B1(new_n845), .B2(new_n491), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT4), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n495), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(new_n490), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n705), .B(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT100), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n712), .A2(new_n852), .ZN(new_n853));
  XOR2_X1   g428(.A(new_n853), .B(KEYINPUT99), .Z(new_n854));
  OR2_X1    g429(.A1(new_n851), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n851), .A2(new_n854), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n855), .A2(new_n738), .A3(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n738), .B1(new_n855), .B2(new_n856), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n844), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n630), .B(new_n477), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(new_n486), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n851), .B(new_n854), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n864), .A2(new_n737), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n837), .B(new_n842), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n865), .A2(new_n866), .A3(new_n857), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n860), .A2(new_n863), .A3(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT104), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND4_X1  g445(.A1(new_n860), .A2(new_n867), .A3(KEYINPUT104), .A4(new_n863), .ZN(new_n871));
  AOI21_X1  g446(.A(G37), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT103), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n860), .A2(new_n873), .A3(new_n867), .ZN(new_n874));
  OAI211_X1 g449(.A(new_n874), .B(new_n862), .C1(new_n873), .C2(new_n860), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g452(.A(KEYINPUT107), .ZN(new_n878));
  XNOR2_X1  g453(.A(G290), .B(new_n590), .ZN(new_n879));
  OR2_X1    g454(.A1(new_n879), .A2(G303), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(G303), .ZN(new_n881));
  AND3_X1   g456(.A1(new_n880), .A2(new_n581), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n581), .B1(new_n880), .B2(new_n881), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n824), .A2(new_n617), .ZN(new_n885));
  NAND4_X1  g460(.A1(new_n822), .A2(new_n607), .A3(new_n615), .A4(new_n823), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NOR2_X1   g462(.A1(G299), .A2(new_n603), .ZN(new_n888));
  INV_X1    g463(.A(new_n603), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n889), .A2(new_n612), .ZN(new_n890));
  OAI21_X1  g465(.A(KEYINPUT41), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(G299), .A2(new_n603), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n889), .A2(new_n612), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT41), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n891), .A2(KEYINPUT105), .A3(new_n895), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n888), .A2(new_n890), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT105), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n897), .A2(new_n898), .A3(new_n894), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n887), .A2(new_n896), .A3(new_n899), .ZN(new_n900));
  XOR2_X1   g475(.A(KEYINPUT106), .B(KEYINPUT42), .Z(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n885), .A2(new_n897), .A3(new_n886), .ZN(new_n903));
  AND3_X1   g478(.A1(new_n900), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n902), .B1(new_n900), .B2(new_n903), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n884), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n900), .A2(new_n903), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(new_n901), .ZN(new_n908));
  INV_X1    g483(.A(new_n884), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n900), .A2(new_n902), .A3(new_n903), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n908), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n906), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(G868), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n821), .A2(G868), .ZN(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n878), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  AOI211_X1 g491(.A(KEYINPUT107), .B(new_n914), .C1(new_n912), .C2(G868), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n916), .A2(new_n917), .ZN(G295));
  NAND2_X1  g493(.A1(new_n913), .A2(new_n915), .ZN(G331));
  XNOR2_X1  g494(.A(G301), .B(G286), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n824), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n822), .A2(new_n823), .A3(new_n920), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n924), .A2(new_n896), .A3(new_n899), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n922), .A2(new_n897), .A3(new_n923), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g502(.A(KEYINPUT108), .B1(new_n927), .B2(new_n909), .ZN(new_n928));
  INV_X1    g503(.A(G37), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n927), .A2(new_n909), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT108), .ZN(new_n931));
  NAND4_X1  g506(.A1(new_n925), .A2(new_n884), .A3(new_n931), .A4(new_n926), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n928), .A2(new_n929), .A3(new_n930), .A4(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT43), .ZN(new_n934));
  AND2_X1   g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT109), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n891), .A2(new_n936), .A3(new_n895), .ZN(new_n937));
  OAI211_X1 g512(.A(new_n924), .B(new_n937), .C1(new_n936), .C2(new_n891), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n938), .A2(new_n926), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n939), .A2(new_n909), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n928), .A2(new_n940), .A3(new_n929), .A4(new_n932), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n941), .A2(new_n934), .ZN(new_n942));
  OAI21_X1  g517(.A(KEYINPUT44), .B1(new_n935), .B2(new_n942), .ZN(new_n943));
  OR2_X1    g518(.A1(new_n933), .A2(new_n934), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT44), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n941), .A2(new_n934), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n943), .A2(new_n947), .ZN(G397));
  AOI21_X1  g523(.A(G1384), .B1(new_n848), .B2(new_n849), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n949), .A2(KEYINPUT45), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n465), .A2(G101), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n471), .A2(G137), .ZN(new_n952));
  AND4_X1   g527(.A1(G40), .A2(new_n476), .A3(new_n951), .A4(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n950), .A2(new_n953), .ZN(new_n954));
  OR2_X1    g529(.A1(new_n792), .A2(new_n795), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n792), .A2(new_n795), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n954), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n705), .A2(G2067), .ZN(new_n958));
  INV_X1    g533(.A(G2067), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n703), .A2(new_n959), .A3(new_n704), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(new_n954), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  XOR2_X1   g538(.A(new_n963), .B(KEYINPUT111), .Z(new_n964));
  NOR2_X1   g539(.A1(new_n954), .A2(G1996), .ZN(new_n965));
  XNOR2_X1  g540(.A(new_n965), .B(KEYINPUT110), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(new_n738), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n962), .A2(G1996), .A3(new_n737), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n964), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  XNOR2_X1  g544(.A(G290), .B(G1986), .ZN(new_n970));
  AOI211_X1 g545(.A(new_n957), .B(new_n969), .C1(new_n962), .C2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT52), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n949), .A2(new_n953), .ZN(new_n973));
  INV_X1    g548(.A(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(G8), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n581), .A2(G1976), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n972), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n977), .A2(new_n972), .A3(G8), .A4(new_n973), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n581), .A2(G1976), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  OAI21_X1  g556(.A(KEYINPUT115), .B1(new_n978), .B2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(G1981), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n590), .B(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT49), .ZN(new_n985));
  OR2_X1    g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n984), .A2(new_n985), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n986), .A2(new_n987), .A3(new_n976), .ZN(new_n988));
  OAI211_X1 g563(.A(new_n982), .B(new_n988), .C1(KEYINPUT115), .C2(new_n981), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n516), .A2(G8), .A3(new_n524), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT113), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(KEYINPUT114), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT55), .ZN(new_n994));
  NAND4_X1  g569(.A1(new_n516), .A2(new_n524), .A3(KEYINPUT113), .A4(G8), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT114), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n990), .A2(new_n991), .A3(new_n996), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n993), .A2(new_n994), .A3(new_n995), .A4(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n995), .A2(new_n994), .ZN(new_n999));
  AND3_X1   g574(.A1(new_n990), .A2(new_n991), .A3(new_n996), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n996), .B1(new_n990), .B2(new_n991), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n999), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  AND2_X1   g577(.A1(new_n998), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n472), .A2(G40), .A3(new_n476), .ZN(new_n1004));
  INV_X1    g579(.A(G1384), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n850), .A2(KEYINPUT45), .A3(new_n1005), .ZN(new_n1006));
  OR2_X1    g581(.A1(new_n1006), .A2(KEYINPUT112), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT45), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1008), .B1(G164), .B2(G1384), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1009), .A2(KEYINPUT112), .A3(new_n1006), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1004), .B1(new_n1007), .B2(new_n1010), .ZN(new_n1011));
  OR2_X1    g586(.A1(new_n1011), .A2(G1971), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT50), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n953), .B1(new_n949), .B2(new_n1013), .ZN(new_n1014));
  NOR3_X1   g589(.A1(G164), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(new_n749), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n975), .B1(new_n1012), .B2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n989), .B1(new_n1003), .B2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n998), .A2(new_n1002), .ZN(new_n1020));
  INV_X1    g595(.A(new_n495), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n845), .A2(new_n491), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(G2105), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1021), .B1(new_n1023), .B2(KEYINPUT4), .ZN(new_n1024));
  OAI211_X1 g599(.A(new_n1013), .B(new_n1005), .C1(new_n1024), .C2(new_n490), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(KEYINPUT118), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT118), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n949), .A2(new_n1027), .A3(new_n1013), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT117), .ZN(new_n1030));
  OAI211_X1 g605(.A(new_n1030), .B(new_n953), .C1(new_n949), .C2(new_n1013), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1014), .A2(KEYINPUT117), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1029), .A2(new_n1031), .A3(new_n1032), .ZN(new_n1033));
  OR2_X1    g608(.A1(new_n1033), .A2(G2090), .ZN(new_n1034));
  AND2_X1   g609(.A1(new_n1012), .A2(new_n1034), .ZN(new_n1035));
  OAI211_X1 g610(.A(KEYINPUT119), .B(new_n1020), .C1(new_n1035), .C2(new_n975), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT119), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n975), .B1(new_n1012), .B2(new_n1034), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1037), .B1(new_n1003), .B2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1019), .A2(new_n1036), .A3(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT61), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n568), .A2(KEYINPUT123), .A3(KEYINPUT57), .A4(new_n575), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n575), .A2(new_n562), .A3(KEYINPUT57), .A4(new_n566), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT123), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT57), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n564), .A2(new_n565), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1045), .B1(new_n611), .B2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1043), .A2(new_n1044), .A3(new_n1047), .ZN(new_n1048));
  AND2_X1   g623(.A1(new_n1042), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1033), .A2(new_n761), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(KEYINPUT122), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT122), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1033), .A2(new_n1052), .A3(new_n761), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1054));
  XNOR2_X1  g629(.A(KEYINPUT56), .B(G2072), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1011), .A2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1049), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1057));
  AND3_X1   g632(.A1(new_n1033), .A2(new_n1052), .A3(new_n761), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1052), .B1(new_n1033), .B2(new_n761), .ZN(new_n1059));
  OAI211_X1 g634(.A(new_n1049), .B(new_n1056), .C1(new_n1058), .C2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1060), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1041), .B1(new_n1057), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT59), .ZN(new_n1063));
  XNOR2_X1  g638(.A(KEYINPUT58), .B(G1341), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n974), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(G1996), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1065), .B1(new_n1011), .B2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1063), .B1(new_n1067), .B2(new_n547), .ZN(new_n1068));
  AOI211_X1 g643(.A(G1996), .B(new_n1004), .C1(new_n1007), .C2(new_n1010), .ZN(new_n1069));
  OAI211_X1 g644(.A(KEYINPUT59), .B(new_n548), .C1(new_n1069), .C2(new_n1065), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1068), .A2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(G1348), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1072), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n974), .A2(new_n959), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT60), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1077), .A2(KEYINPUT124), .A3(new_n889), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT124), .ZN(new_n1079));
  AOI21_X1  g654(.A(KEYINPUT60), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1079), .B1(new_n1080), .B2(new_n603), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1078), .A2(new_n1081), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  OAI211_X1 g659(.A(new_n1078), .B(new_n1081), .C1(new_n1076), .C2(new_n1075), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1071), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1056), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1049), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1089), .A2(KEYINPUT61), .A3(new_n1060), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1062), .A2(new_n1086), .A3(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n603), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1060), .B1(new_n1057), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n951), .A2(new_n952), .ZN(new_n1095));
  INV_X1    g670(.A(G2078), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(KEYINPUT53), .ZN(new_n1097));
  AOI211_X1 g672(.A(new_n1095), .B(new_n1097), .C1(new_n1007), .C2(new_n1010), .ZN(new_n1098));
  XNOR2_X1  g673(.A(new_n475), .B(KEYINPUT127), .ZN(new_n1099));
  OAI211_X1 g674(.A(new_n1098), .B(G40), .C1(new_n463), .C2(new_n1099), .ZN(new_n1100));
  XNOR2_X1  g675(.A(G301), .B(KEYINPUT54), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(KEYINPUT53), .B1(new_n1011), .B2(new_n1096), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1103), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n689), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1100), .A2(new_n1102), .A3(new_n1104), .A4(new_n1105), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1009), .A2(new_n953), .A3(new_n1006), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1105), .B1(new_n1097), .B2(new_n1107), .ZN(new_n1108));
  XNOR2_X1  g683(.A(new_n1108), .B(KEYINPUT126), .ZN(new_n1109));
  OR2_X1    g684(.A1(new_n1109), .A2(new_n1103), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(new_n1101), .ZN(new_n1111));
  AND3_X1   g686(.A1(new_n1107), .A2(KEYINPUT120), .A3(new_n727), .ZN(new_n1112));
  AOI21_X1  g687(.A(KEYINPUT120), .B1(new_n1107), .B2(new_n727), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1016), .A2(new_n722), .ZN(new_n1115));
  AOI21_X1  g690(.A(KEYINPUT125), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1107), .A2(new_n727), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT120), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1107), .A2(KEYINPUT120), .A3(new_n727), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1119), .A2(KEYINPUT125), .A3(new_n1115), .A4(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1121), .ZN(new_n1122));
  OAI211_X1 g697(.A(G8), .B(G286), .C1(new_n1116), .C2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT51), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1119), .A2(new_n1115), .A3(new_n1120), .ZN(new_n1125));
  OAI211_X1 g700(.A(new_n1124), .B(G8), .C1(new_n1125), .C2(G286), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1123), .A2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT125), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1125), .A2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1129), .A2(G168), .A3(new_n1121), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1124), .B1(new_n1130), .B2(G8), .ZN(new_n1131));
  OAI211_X1 g706(.A(new_n1106), .B(new_n1111), .C1(new_n1127), .C2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1094), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1131), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT62), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1135), .A2(new_n1136), .A3(new_n1126), .A4(new_n1123), .ZN(new_n1137));
  OAI21_X1  g712(.A(KEYINPUT62), .B1(new_n1127), .B2(new_n1131), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1137), .A2(new_n1138), .A3(G171), .A4(new_n1110), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1040), .B1(new_n1134), .B2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT63), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1125), .A2(G8), .A3(G168), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1141), .B1(new_n1040), .B2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT121), .ZN(new_n1144));
  NOR3_X1   g719(.A1(new_n1003), .A2(new_n1018), .A3(new_n1144), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1145), .A2(new_n1141), .ZN(new_n1146));
  INV_X1    g721(.A(new_n989), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1142), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1018), .B1(new_n1003), .B2(new_n1144), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n1146), .A2(new_n1147), .A3(new_n1148), .A4(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1143), .A2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1147), .A2(new_n1018), .A3(new_n1003), .ZN(new_n1152));
  INV_X1    g727(.A(G1976), .ZN(new_n1153));
  AND3_X1   g728(.A1(new_n988), .A2(new_n1153), .A3(new_n581), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n590), .A2(new_n983), .ZN(new_n1155));
  XOR2_X1   g730(.A(new_n1155), .B(KEYINPUT116), .Z(new_n1156));
  OAI21_X1  g731(.A(new_n976), .B1(new_n1154), .B2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1151), .A2(new_n1152), .A3(new_n1157), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n971), .B1(new_n1140), .B2(new_n1158), .ZN(new_n1159));
  XOR2_X1   g734(.A(new_n966), .B(KEYINPUT46), .Z(new_n1160));
  OAI211_X1 g735(.A(new_n1160), .B(new_n963), .C1(new_n738), .C2(new_n954), .ZN(new_n1161));
  XOR2_X1   g736(.A(new_n1161), .B(KEYINPUT47), .Z(new_n1162));
  NOR3_X1   g737(.A1(new_n954), .A2(G1986), .A3(G290), .ZN(new_n1163));
  XNOR2_X1  g738(.A(new_n1163), .B(KEYINPUT48), .ZN(new_n1164));
  NOR3_X1   g739(.A1(new_n969), .A2(new_n957), .A3(new_n1164), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n960), .B1(new_n969), .B2(new_n955), .ZN(new_n1166));
  AND2_X1   g741(.A1(new_n1166), .A2(new_n962), .ZN(new_n1167));
  NOR3_X1   g742(.A1(new_n1162), .A2(new_n1165), .A3(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1159), .A2(new_n1168), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g744(.A1(new_n649), .A2(new_n684), .ZN(new_n1171));
  AOI21_X1  g745(.A(new_n1171), .B1(new_n872), .B2(new_n875), .ZN(new_n1172));
  NOR2_X1   g746(.A1(G227), .A2(new_n461), .ZN(new_n1173));
  NAND4_X1  g747(.A1(new_n1172), .A2(new_n944), .A3(new_n946), .A4(new_n1173), .ZN(G225));
  INV_X1    g748(.A(G225), .ZN(G308));
endmodule


