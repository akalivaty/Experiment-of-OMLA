//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 1 1 0 0 1 0 1 1 0 1 1 1 1 1 0 1 0 1 0 1 1 1 1 1 0 1 1 1 0 0 0 1 0 1 1 0 1 1 1 0 1 0 0 1 1 0 1 0 0 1 0 1 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:45 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n210));
  INV_X1    g0010(.A(G87), .ZN(new_n211));
  INV_X1    g0011(.A(G250), .ZN(new_n212));
  OAI21_X1  g0012(.A(new_n210), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  AOI21_X1  g0013(.A(new_n213), .B1(G116), .B2(G270), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G58), .A2(G232), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G107), .A2(G264), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G50), .A2(G226), .ZN(new_n217));
  NAND4_X1  g0017(.A1(new_n214), .A2(new_n215), .A3(new_n216), .A4(new_n217), .ZN(new_n218));
  INV_X1    g0018(.A(G68), .ZN(new_n219));
  INV_X1    g0019(.A(G238), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n209), .B1(new_n218), .B2(new_n221), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT1), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n209), .A2(G13), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n224), .B(G250), .C1(G257), .C2(G264), .ZN(new_n225));
  INV_X1    g0025(.A(KEYINPUT0), .ZN(new_n226));
  OR2_X1    g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(G50), .B1(G58), .B2(G68), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  INV_X1    g0030(.A(G20), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n229), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n225), .A2(new_n226), .ZN(new_n234));
  NAND3_X1  g0034(.A1(new_n227), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n235), .B(KEYINPUT64), .Z(new_n236));
  NOR2_X1   g0036(.A1(new_n223), .A2(new_n236), .ZN(G361));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT2), .B(G226), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G250), .B(G257), .Z(new_n242));
  XNOR2_X1  g0042(.A(G264), .B(G270), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G358));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(G68), .B(G77), .Z(new_n249));
  XNOR2_X1  g0049(.A(G50), .B(G58), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n248), .B(new_n251), .ZN(G351));
  INV_X1    g0052(.A(KEYINPUT17), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT74), .ZN(new_n254));
  INV_X1    g0054(.A(G1), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n255), .B1(G41), .B2(G45), .ZN(new_n256));
  INV_X1    g0056(.A(G274), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(KEYINPUT3), .ZN(new_n260));
  OR2_X1    g0060(.A1(G223), .A2(G1698), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT3), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G33), .ZN(new_n263));
  INV_X1    g0063(.A(G226), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G1698), .ZN(new_n265));
  NAND4_X1  g0065(.A1(new_n260), .A2(new_n261), .A3(new_n263), .A4(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(G33), .A2(G87), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(G33), .A2(G41), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n269), .A2(G1), .A3(G13), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n258), .B1(new_n268), .B2(new_n271), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n270), .A2(G232), .A3(new_n256), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n254), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n270), .B1(new_n266), .B2(new_n267), .ZN(new_n275));
  INV_X1    g0075(.A(new_n273), .ZN(new_n276));
  NOR4_X1   g0076(.A1(new_n275), .A2(new_n276), .A3(KEYINPUT74), .A4(new_n258), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n274), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G200), .ZN(new_n279));
  INV_X1    g0079(.A(G190), .ZN(new_n280));
  NOR3_X1   g0080(.A1(new_n275), .A2(new_n258), .A3(new_n276), .ZN(new_n281));
  AOI22_X1  g0081(.A1(new_n278), .A2(new_n279), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  XOR2_X1   g0082(.A(KEYINPUT8), .B(G58), .Z(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n255), .A2(G13), .A3(G20), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g0087(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(new_n230), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n255), .A2(G20), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n287), .B1(new_n292), .B2(new_n284), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT16), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT7), .ZN(new_n296));
  XNOR2_X1  g0096(.A(KEYINPUT3), .B(G33), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n296), .B1(new_n297), .B2(G20), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n260), .A2(new_n263), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n296), .A2(G20), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n219), .B1(new_n298), .B2(new_n301), .ZN(new_n302));
  AND2_X1   g0102(.A1(G58), .A2(G68), .ZN(new_n303));
  OAI21_X1  g0103(.A(G20), .B1(new_n303), .B2(new_n201), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(KEYINPUT71), .ZN(new_n305));
  NOR2_X1   g0105(.A1(G20), .A2(G33), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(G159), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT71), .ZN(new_n308));
  OAI211_X1 g0108(.A(new_n308), .B(G20), .C1(new_n303), .C2(new_n201), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n305), .A2(new_n307), .A3(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(KEYINPUT72), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT72), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n305), .A2(new_n312), .A3(new_n307), .A4(new_n309), .ZN(new_n313));
  AOI211_X1 g0113(.A(new_n295), .B(new_n302), .C1(new_n311), .C2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT73), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n315), .B1(new_n262), .B2(G33), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n259), .A2(KEYINPUT73), .A3(KEYINPUT3), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n316), .A2(new_n263), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(new_n300), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n219), .B1(new_n319), .B2(new_n298), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n295), .B1(new_n320), .B2(new_n310), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(new_n289), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n294), .B1(new_n314), .B2(new_n322), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n253), .B1(new_n282), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n268), .A2(new_n271), .ZN(new_n325));
  INV_X1    g0125(.A(new_n258), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n325), .A2(new_n326), .A3(new_n273), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(KEYINPUT74), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n281), .A2(new_n254), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n328), .A2(new_n329), .A3(new_n279), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n330), .B1(G190), .B2(new_n327), .ZN(new_n331));
  AND2_X1   g0131(.A1(new_n305), .A2(new_n309), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n262), .A2(G33), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n259), .A2(KEYINPUT3), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n231), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  AOI22_X1  g0135(.A1(new_n296), .A2(new_n335), .B1(new_n318), .B2(new_n300), .ZN(new_n336));
  OAI211_X1 g0136(.A(new_n332), .B(new_n307), .C1(new_n336), .C2(new_n219), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n290), .B1(new_n337), .B2(new_n295), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n311), .A2(new_n313), .ZN(new_n339));
  INV_X1    g0139(.A(new_n302), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n339), .A2(KEYINPUT16), .A3(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n293), .B1(new_n338), .B2(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n331), .A2(new_n342), .A3(KEYINPUT17), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n324), .A2(new_n343), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n327), .A2(G179), .ZN(new_n345));
  INV_X1    g0145(.A(G169), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n345), .B1(new_n278), .B2(new_n346), .ZN(new_n347));
  NAND4_X1  g0147(.A1(new_n347), .A2(new_n323), .A3(KEYINPUT75), .A4(KEYINPUT18), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT18), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n328), .A2(new_n329), .A3(new_n346), .ZN(new_n350));
  INV_X1    g0150(.A(new_n345), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n349), .B1(new_n342), .B2(new_n352), .ZN(new_n353));
  AND2_X1   g0153(.A1(new_n348), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n347), .A2(new_n323), .A3(KEYINPUT18), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT75), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n344), .B1(new_n354), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n203), .A2(G20), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n259), .A2(G20), .ZN(new_n360));
  AOI22_X1  g0160(.A1(new_n359), .A2(KEYINPUT66), .B1(new_n283), .B2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(G150), .ZN(new_n362));
  INV_X1    g0162(.A(new_n306), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n361), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n359), .A2(KEYINPUT66), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n289), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n286), .A2(new_n202), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n291), .A2(G50), .ZN(new_n368));
  XOR2_X1   g0168(.A(new_n368), .B(KEYINPUT67), .Z(new_n369));
  NAND3_X1  g0169(.A1(new_n369), .A2(new_n285), .A3(new_n290), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n366), .A2(new_n367), .A3(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT9), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n366), .A2(KEYINPUT9), .A3(new_n367), .A4(new_n370), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n270), .A2(new_n256), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT65), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n270), .A2(KEYINPUT65), .A3(new_n256), .ZN(new_n378));
  AND2_X1   g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(G226), .ZN(new_n380));
  NOR2_X1   g0180(.A1(G222), .A2(G1698), .ZN(new_n381));
  INV_X1    g0181(.A(G1698), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n382), .A2(G223), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n297), .B1(new_n381), .B2(new_n383), .ZN(new_n384));
  OAI211_X1 g0184(.A(new_n384), .B(new_n271), .C1(G77), .C2(new_n297), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n380), .A2(new_n326), .A3(new_n385), .ZN(new_n386));
  AOI22_X1  g0186(.A1(new_n386), .A2(G200), .B1(KEYINPUT68), .B2(KEYINPUT10), .ZN(new_n387));
  INV_X1    g0187(.A(new_n386), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(G190), .ZN(new_n389));
  NAND4_X1  g0189(.A1(new_n373), .A2(new_n374), .A3(new_n387), .A4(new_n389), .ZN(new_n390));
  NOR2_X1   g0190(.A1(KEYINPUT68), .A2(KEYINPUT10), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  AOI22_X1  g0192(.A1(new_n371), .A2(new_n372), .B1(new_n388), .B2(G190), .ZN(new_n393));
  INV_X1    g0193(.A(new_n391), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n393), .A2(new_n394), .A3(new_n374), .A4(new_n387), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n386), .A2(new_n346), .ZN(new_n396));
  OAI211_X1 g0196(.A(new_n371), .B(new_n396), .C1(G179), .C2(new_n386), .ZN(new_n397));
  AND3_X1   g0197(.A1(new_n392), .A2(new_n395), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n379), .A2(G244), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n297), .A2(G232), .A3(new_n382), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n297), .A2(G238), .A3(G1698), .ZN(new_n401));
  OAI211_X1 g0201(.A(new_n400), .B(new_n401), .C1(new_n206), .C2(new_n297), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(new_n271), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n399), .A2(new_n403), .A3(new_n326), .ZN(new_n404));
  OR2_X1    g0204(.A1(new_n404), .A2(G179), .ZN(new_n405));
  AOI22_X1  g0205(.A1(new_n283), .A2(new_n306), .B1(G20), .B2(G77), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n231), .A2(G33), .ZN(new_n407));
  XOR2_X1   g0207(.A(KEYINPUT15), .B(G87), .Z(new_n408));
  INV_X1    g0208(.A(new_n408), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n406), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n292), .ZN(new_n411));
  AOI22_X1  g0211(.A1(new_n410), .A2(new_n289), .B1(G77), .B2(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n412), .B1(G77), .B2(new_n285), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n404), .A2(new_n346), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n405), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  AND3_X1   g0215(.A1(new_n358), .A2(new_n398), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n264), .A2(new_n382), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n417), .B1(G232), .B2(new_n382), .ZN(new_n418));
  OAI22_X1  g0218(.A1(new_n418), .A2(new_n299), .B1(new_n259), .B2(new_n205), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(new_n271), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n377), .A2(G238), .A3(new_n378), .ZN(new_n421));
  AND3_X1   g0221(.A1(new_n421), .A2(KEYINPUT69), .A3(new_n326), .ZN(new_n422));
  AOI21_X1  g0222(.A(KEYINPUT69), .B1(new_n421), .B2(new_n326), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n420), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(KEYINPUT13), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT13), .ZN(new_n426));
  OAI211_X1 g0226(.A(new_n426), .B(new_n420), .C1(new_n422), .C2(new_n423), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n425), .A2(KEYINPUT70), .A3(new_n427), .ZN(new_n428));
  OR3_X1    g0228(.A1(new_n424), .A2(KEYINPUT70), .A3(KEYINPUT13), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n428), .A2(new_n429), .A3(G200), .ZN(new_n430));
  OAI22_X1  g0230(.A1(new_n363), .A2(new_n202), .B1(new_n231), .B2(G68), .ZN(new_n431));
  INV_X1    g0231(.A(G77), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n407), .A2(new_n432), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n289), .B1(new_n431), .B2(new_n433), .ZN(new_n434));
  XNOR2_X1  g0234(.A(new_n434), .B(KEYINPUT11), .ZN(new_n435));
  OAI21_X1  g0235(.A(KEYINPUT12), .B1(new_n285), .B2(G68), .ZN(new_n436));
  OR3_X1    g0236(.A1(new_n285), .A2(KEYINPUT12), .A3(G68), .ZN(new_n437));
  AOI22_X1  g0237(.A1(new_n411), .A2(G68), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n435), .A2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n425), .A2(G190), .A3(new_n427), .ZN(new_n441));
  AND3_X1   g0241(.A1(new_n430), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n428), .A2(new_n429), .A3(G169), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(KEYINPUT14), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT14), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n428), .A2(new_n429), .A3(new_n445), .A4(G169), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n425), .A2(G179), .A3(new_n427), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n444), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n442), .B1(new_n448), .B2(new_n439), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n413), .B1(G200), .B2(new_n404), .ZN(new_n450));
  OR2_X1    g0250(.A1(new_n404), .A2(new_n280), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  AND3_X1   g0252(.A1(new_n416), .A2(new_n449), .A3(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n297), .A2(G257), .A3(G1698), .ZN(new_n455));
  NAND2_X1  g0255(.A1(G33), .A2(G294), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n260), .A2(new_n263), .A3(G250), .A4(new_n382), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n455), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(new_n271), .ZN(new_n459));
  INV_X1    g0259(.A(G41), .ZN(new_n460));
  OAI211_X1 g0260(.A(new_n255), .B(G45), .C1(new_n460), .C2(KEYINPUT5), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT77), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT5), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n463), .B1(new_n464), .B2(G41), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n460), .A2(KEYINPUT77), .A3(KEYINPUT5), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n462), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n468), .A2(G264), .A3(new_n270), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n461), .B1(new_n465), .B2(new_n466), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(G274), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n459), .A2(new_n469), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(G169), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT86), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(new_n472), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(G179), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n472), .A2(KEYINPUT86), .A3(G169), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n475), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT24), .ZN(new_n480));
  OAI21_X1  g0280(.A(KEYINPUT23), .B1(new_n231), .B2(G107), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT23), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n482), .A2(new_n206), .A3(G20), .ZN(new_n483));
  INV_X1    g0283(.A(G116), .ZN(new_n484));
  OAI211_X1 g0284(.A(new_n481), .B(new_n483), .C1(new_n484), .C2(new_n407), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT84), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n360), .A2(G116), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n488), .A2(KEYINPUT84), .A3(new_n481), .A4(new_n483), .ZN(new_n489));
  AND2_X1   g0289(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  XOR2_X1   g0290(.A(KEYINPUT83), .B(KEYINPUT22), .Z(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n297), .A2(new_n231), .A3(G87), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n491), .A2(new_n231), .A3(G87), .A4(new_n297), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n480), .B1(new_n490), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n487), .A2(new_n489), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n498), .A2(KEYINPUT24), .A3(new_n495), .A4(new_n494), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n497), .A2(new_n289), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n255), .A2(G33), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n285), .A2(new_n501), .A3(new_n230), .A4(new_n288), .ZN(new_n502));
  INV_X1    g0302(.A(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(G107), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n286), .B(new_n206), .C1(KEYINPUT85), .C2(KEYINPUT25), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT85), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT25), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n506), .B(new_n507), .C1(new_n285), .C2(G107), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n505), .B(new_n508), .C1(new_n506), .C2(new_n507), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n500), .A2(new_n504), .A3(new_n509), .ZN(new_n510));
  AND2_X1   g0310(.A1(new_n479), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n472), .A2(G200), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n500), .A2(new_n504), .A3(new_n509), .A4(new_n512), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n472), .A2(new_n280), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n220), .A2(new_n382), .ZN(new_n516));
  INV_X1    g0316(.A(G244), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(G1698), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n260), .A2(new_n516), .A3(new_n263), .A4(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(G33), .A2(G116), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(new_n271), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n255), .A2(G45), .ZN(new_n523));
  AND2_X1   g0323(.A1(G33), .A2(G41), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n523), .B(G250), .C1(new_n524), .C2(new_n230), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n255), .A2(G45), .A3(G274), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n525), .A2(KEYINPUT78), .A3(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(KEYINPUT78), .B1(new_n525), .B2(new_n526), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n522), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(new_n346), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n525), .A2(new_n526), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT78), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(new_n527), .ZN(new_n535));
  INV_X1    g0335(.A(G179), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n535), .A2(new_n536), .A3(new_n522), .ZN(new_n537));
  NAND3_X1  g0337(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(new_n231), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n211), .A2(new_n205), .A3(new_n206), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n260), .A2(new_n263), .A3(new_n231), .A4(G68), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT19), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n543), .B1(new_n407), .B2(new_n205), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n541), .A2(new_n542), .A3(new_n544), .ZN(new_n545));
  AOI22_X1  g0345(.A1(new_n545), .A2(new_n289), .B1(new_n286), .B2(new_n409), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT79), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n503), .A2(new_n408), .ZN(new_n548));
  AND3_X1   g0348(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n547), .B1(new_n546), .B2(new_n548), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n531), .B(new_n537), .C1(new_n549), .C2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(new_n530), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(G190), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n530), .A2(G200), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT80), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n503), .A2(new_n555), .A3(G87), .ZN(new_n556));
  OAI21_X1  g0356(.A(KEYINPUT80), .B1(new_n502), .B2(new_n211), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  AND2_X1   g0358(.A1(new_n558), .A2(new_n546), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n553), .A2(new_n554), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n551), .A2(new_n560), .ZN(new_n561));
  NOR3_X1   g0361(.A1(new_n511), .A2(new_n515), .A3(new_n561), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n285), .A2(G97), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n502), .A2(new_n205), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n306), .A2(G77), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT76), .ZN(new_n566));
  NAND2_X1  g0366(.A1(KEYINPUT6), .A2(G97), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n566), .B1(new_n567), .B2(G107), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n206), .A2(KEYINPUT76), .A3(KEYINPUT6), .A4(G97), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(G97), .A2(G107), .ZN(new_n571));
  AOI21_X1  g0371(.A(KEYINPUT6), .B1(new_n207), .B2(new_n571), .ZN(new_n572));
  OAI21_X1  g0372(.A(G20), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n565), .B(new_n573), .C1(new_n336), .C2(new_n206), .ZN(new_n574));
  AOI211_X1 g0374(.A(new_n563), .B(new_n564), .C1(new_n574), .C2(new_n289), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n260), .A2(new_n263), .A3(G244), .A4(new_n382), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT4), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n297), .A2(KEYINPUT4), .A3(G244), .A4(new_n382), .ZN(new_n579));
  NAND2_X1  g0379(.A1(G33), .A2(G283), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n297), .A2(G250), .A3(G1698), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n578), .A2(new_n579), .A3(new_n580), .A4(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n271), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n470), .A2(new_n271), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(G257), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n583), .A2(new_n471), .A3(new_n585), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n586), .A2(G190), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n582), .A2(new_n271), .B1(new_n584), .B2(G257), .ZN(new_n588));
  AOI21_X1  g0388(.A(G200), .B1(new_n588), .B2(new_n471), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n575), .B1(new_n587), .B2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(new_n563), .ZN(new_n591));
  INV_X1    g0391(.A(new_n564), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n206), .B1(new_n319), .B2(new_n298), .ZN(new_n593));
  AND2_X1   g0393(.A1(new_n568), .A2(new_n569), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n207), .A2(new_n571), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT6), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n231), .B1(new_n594), .B2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(new_n565), .ZN(new_n599));
  NOR3_X1   g0399(.A1(new_n593), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n591), .B(new_n592), .C1(new_n600), .C2(new_n290), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n588), .A2(new_n536), .A3(new_n471), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n586), .A2(new_n346), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  AND2_X1   g0404(.A1(new_n590), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n468), .A2(G270), .A3(new_n270), .ZN(new_n606));
  AND2_X1   g0406(.A1(new_n606), .A2(new_n471), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n297), .A2(G257), .A3(new_n382), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n299), .A2(G303), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n260), .A2(new_n263), .A3(G264), .A4(G1698), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT81), .ZN(new_n612));
  AND3_X1   g0412(.A1(new_n611), .A2(new_n612), .A3(new_n271), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n612), .B1(new_n611), .B2(new_n271), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n607), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n286), .A2(new_n484), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n503), .A2(G116), .ZN(new_n617));
  OAI211_X1 g0417(.A(new_n580), .B(new_n231), .C1(G33), .C2(new_n205), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n618), .B(new_n289), .C1(new_n231), .C2(G116), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT20), .ZN(new_n620));
  AND2_X1   g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n619), .A2(new_n620), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n616), .B(new_n617), .C1(new_n621), .C2(new_n622), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n615), .A2(G169), .A3(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT21), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  OAI211_X1 g0426(.A(new_n607), .B(G190), .C1(new_n613), .C2(new_n614), .ZN(new_n627));
  INV_X1    g0427(.A(new_n623), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n606), .A2(new_n471), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n611), .A2(new_n271), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(KEYINPUT81), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n611), .A2(new_n612), .A3(new_n271), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n629), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  OAI211_X1 g0433(.A(new_n627), .B(new_n628), .C1(new_n633), .C2(new_n279), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n633), .A2(G179), .A3(new_n623), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n615), .A2(KEYINPUT21), .A3(G169), .A4(new_n623), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n626), .A2(new_n634), .A3(new_n635), .A4(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT82), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n637), .A2(new_n638), .ZN(new_n640));
  OAI211_X1 g0440(.A(new_n562), .B(new_n605), .C1(new_n639), .C2(new_n640), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n454), .A2(new_n641), .ZN(G372));
  NAND2_X1  g0442(.A1(new_n448), .A2(new_n439), .ZN(new_n643));
  AOI211_X1 g0443(.A(new_n344), .B(new_n442), .C1(new_n643), .C2(new_n415), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n353), .A2(new_n355), .ZN(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  OAI211_X1 g0446(.A(new_n392), .B(new_n395), .C1(new_n644), .C2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT87), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n279), .B1(new_n535), .B2(new_n522), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n558), .A2(new_n546), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n648), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n559), .A2(new_n554), .A3(KEYINPUT87), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n651), .A2(new_n652), .A3(new_n553), .ZN(new_n653));
  AND2_X1   g0453(.A1(new_n653), .A2(new_n551), .ZN(new_n654));
  AND2_X1   g0454(.A1(new_n500), .A2(new_n509), .ZN(new_n655));
  INV_X1    g0455(.A(new_n514), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n655), .A2(new_n504), .A3(new_n656), .A4(new_n512), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT88), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n605), .A2(new_n654), .A3(new_n657), .A4(new_n658), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n590), .A2(new_n653), .A3(new_n604), .A4(new_n551), .ZN(new_n660));
  OAI21_X1  g0460(.A(KEYINPUT88), .B1(new_n660), .B2(new_n515), .ZN(new_n661));
  AND2_X1   g0461(.A1(new_n626), .A2(new_n636), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n479), .A2(new_n510), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n662), .A2(new_n663), .A3(new_n635), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n659), .A2(new_n661), .A3(new_n664), .ZN(new_n665));
  AND3_X1   g0465(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT26), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n666), .A2(new_n667), .A3(new_n551), .A4(new_n653), .ZN(new_n668));
  OAI21_X1  g0468(.A(KEYINPUT26), .B1(new_n561), .B2(new_n604), .ZN(new_n669));
  AND3_X1   g0469(.A1(new_n668), .A2(new_n669), .A3(new_n551), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n665), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n453), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n647), .A2(new_n672), .A3(new_n397), .ZN(G369));
  INV_X1    g0473(.A(G330), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n662), .A2(new_n635), .ZN(new_n675));
  INV_X1    g0475(.A(G13), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n676), .A2(G20), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  OR3_X1    g0478(.A1(new_n678), .A2(KEYINPUT27), .A3(G1), .ZN(new_n679));
  OAI21_X1  g0479(.A(KEYINPUT27), .B1(new_n678), .B2(G1), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n679), .A2(G213), .A3(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(G343), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n628), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n675), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g0486(.A(new_n637), .B(KEYINPUT82), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n686), .B1(new_n687), .B2(new_n685), .ZN(new_n688));
  OR2_X1    g0488(.A1(new_n688), .A2(KEYINPUT89), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(KEYINPUT89), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n674), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n510), .A2(new_n683), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n657), .A2(new_n663), .A3(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n693), .B1(new_n663), .B2(new_n684), .ZN(new_n694));
  AND2_X1   g0494(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n675), .A2(new_n684), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT90), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  AOI21_X1  g0498(.A(KEYINPUT90), .B1(new_n675), .B2(new_n684), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n694), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n663), .A2(new_n683), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  OR2_X1    g0503(.A1(new_n695), .A2(new_n703), .ZN(G399));
  INV_X1    g0504(.A(new_n224), .ZN(new_n705));
  OR3_X1    g0505(.A1(new_n705), .A2(KEYINPUT91), .A3(G41), .ZN(new_n706));
  OAI21_X1  g0506(.A(KEYINPUT91), .B1(new_n705), .B2(G41), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n709), .A2(new_n255), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n540), .A2(G116), .ZN(new_n711));
  AOI22_X1  g0511(.A1(new_n710), .A2(new_n711), .B1(new_n229), .B2(new_n709), .ZN(new_n712));
  XOR2_X1   g0512(.A(new_n712), .B(KEYINPUT28), .Z(new_n713));
  AOI21_X1  g0513(.A(new_n683), .B1(new_n665), .B2(new_n670), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  XOR2_X1   g0515(.A(KEYINPUT92), .B(KEYINPUT29), .Z(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT29), .ZN(new_n718));
  INV_X1    g0518(.A(new_n664), .ZN(new_n719));
  NOR3_X1   g0519(.A1(new_n719), .A2(new_n515), .A3(new_n660), .ZN(new_n720));
  INV_X1    g0520(.A(new_n654), .ZN(new_n721));
  OAI21_X1  g0521(.A(KEYINPUT26), .B1(new_n721), .B2(new_n604), .ZN(new_n722));
  INV_X1    g0522(.A(new_n551), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n561), .A2(new_n604), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n723), .B1(new_n724), .B2(new_n667), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n722), .A2(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n684), .B1(new_n720), .B2(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n717), .B1(new_n718), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n633), .A2(G179), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  AND3_X1   g0530(.A1(new_n476), .A2(new_n552), .A3(new_n588), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT30), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n730), .A2(KEYINPUT30), .A3(new_n731), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n552), .B1(new_n471), .B2(new_n588), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n736), .A2(new_n536), .A3(new_n472), .A4(new_n615), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n734), .A2(new_n735), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(new_n683), .ZN(new_n739));
  OAI211_X1 g0539(.A(KEYINPUT31), .B(new_n739), .C1(new_n641), .C2(new_n683), .ZN(new_n740));
  OR2_X1    g0540(.A1(new_n739), .A2(KEYINPUT31), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n740), .A2(G330), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n728), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n713), .B1(new_n744), .B2(G1), .ZN(G364));
  AOI21_X1  g0545(.A(new_n255), .B1(new_n677), .B2(G45), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n709), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n691), .A2(new_n748), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n689), .A2(new_n674), .A3(new_n690), .ZN(new_n750));
  NOR2_X1   g0550(.A1(G13), .A2(G33), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(G20), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  OR2_X1    g0554(.A1(new_n688), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(G45), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n229), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n705), .A2(new_n297), .ZN(new_n758));
  OAI211_X1 g0558(.A(new_n757), .B(new_n758), .C1(new_n251), .C2(new_n756), .ZN(new_n759));
  INV_X1    g0559(.A(G355), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n297), .A2(new_n224), .ZN(new_n761));
  OAI221_X1 g0561(.A(new_n759), .B1(G116), .B2(new_n224), .C1(new_n760), .C2(new_n761), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n230), .B1(G20), .B2(new_n346), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n753), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  XOR2_X1   g0565(.A(KEYINPUT33), .B(G317), .Z(new_n766));
  NOR2_X1   g0566(.A1(new_n536), .A2(new_n279), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n231), .A2(G190), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n766), .A2(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n231), .A2(new_n280), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n279), .A2(G179), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n768), .A2(new_n772), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  AOI22_X1  g0576(.A1(G303), .A2(new_n774), .B1(new_n776), .B2(G283), .ZN(new_n777));
  NOR2_X1   g0577(.A1(G179), .A2(G200), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n768), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(G329), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n777), .A2(new_n299), .A3(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n536), .A2(G200), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(new_n768), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  AOI211_X1 g0585(.A(new_n770), .B(new_n782), .C1(G311), .C2(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n771), .A2(new_n767), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n231), .B1(new_n778), .B2(G190), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  AOI22_X1  g0590(.A1(new_n788), .A2(G326), .B1(new_n790), .B2(G294), .ZN(new_n791));
  XNOR2_X1  g0591(.A(new_n791), .B(KEYINPUT95), .ZN(new_n792));
  INV_X1    g0592(.A(G322), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n771), .A2(new_n783), .ZN(new_n794));
  OAI211_X1 g0594(.A(new_n786), .B(new_n792), .C1(new_n793), .C2(new_n794), .ZN(new_n795));
  OAI22_X1  g0595(.A1(new_n787), .A2(new_n202), .B1(new_n784), .B2(new_n432), .ZN(new_n796));
  INV_X1    g0596(.A(new_n794), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n796), .B1(G58), .B2(new_n797), .ZN(new_n798));
  XNOR2_X1  g0598(.A(new_n798), .B(KEYINPUT93), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n799), .B1(G107), .B2(new_n776), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n299), .B1(new_n774), .B2(G87), .ZN(new_n801));
  INV_X1    g0601(.A(new_n769), .ZN(new_n802));
  AOI22_X1  g0602(.A1(new_n802), .A2(G68), .B1(new_n790), .B2(G97), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n800), .A2(new_n801), .A3(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(G159), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n779), .A2(new_n805), .ZN(new_n806));
  XOR2_X1   g0606(.A(KEYINPUT94), .B(KEYINPUT32), .Z(new_n807));
  XNOR2_X1  g0607(.A(new_n806), .B(new_n807), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n795), .B1(new_n804), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(new_n763), .ZN(new_n810));
  AND3_X1   g0610(.A1(new_n755), .A2(new_n765), .A3(new_n810), .ZN(new_n811));
  AOI22_X1  g0611(.A1(new_n749), .A2(new_n750), .B1(new_n748), .B2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(G396));
  INV_X1    g0613(.A(KEYINPUT100), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n415), .A2(new_n683), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  AOI22_X1  g0616(.A1(new_n450), .A2(new_n451), .B1(new_n413), .B2(new_n683), .ZN(new_n817));
  INV_X1    g0617(.A(new_n415), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n816), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  XOR2_X1   g0619(.A(new_n819), .B(KEYINPUT98), .Z(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(new_n715), .ZN(new_n821));
  XOR2_X1   g0621(.A(new_n821), .B(KEYINPUT99), .Z(new_n822));
  INV_X1    g0622(.A(new_n819), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n671), .A2(new_n684), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n814), .B1(new_n825), .B2(new_n742), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n748), .B1(new_n825), .B2(new_n742), .ZN(new_n827));
  INV_X1    g0627(.A(new_n742), .ZN(new_n828));
  NAND4_X1  g0628(.A1(new_n822), .A2(KEYINPUT100), .A3(new_n828), .A4(new_n824), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n826), .A2(new_n827), .A3(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(G137), .ZN(new_n831));
  OAI22_X1  g0631(.A1(new_n787), .A2(new_n831), .B1(new_n769), .B2(new_n362), .ZN(new_n832));
  XNOR2_X1  g0632(.A(new_n832), .B(KEYINPUT97), .ZN(new_n833));
  INV_X1    g0633(.A(G143), .ZN(new_n834));
  OAI221_X1 g0634(.A(new_n833), .B1(new_n834), .B2(new_n794), .C1(new_n805), .C2(new_n784), .ZN(new_n835));
  XNOR2_X1  g0635(.A(new_n835), .B(KEYINPUT34), .ZN(new_n836));
  INV_X1    g0636(.A(G58), .ZN(new_n837));
  OAI221_X1 g0637(.A(new_n836), .B1(new_n202), .B2(new_n773), .C1(new_n837), .C2(new_n789), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n775), .A2(new_n219), .ZN(new_n839));
  INV_X1    g0639(.A(G132), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n779), .A2(new_n840), .ZN(new_n841));
  NOR4_X1   g0641(.A1(new_n838), .A2(new_n299), .A3(new_n839), .A4(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(G294), .ZN(new_n843));
  OAI22_X1  g0643(.A1(new_n794), .A2(new_n843), .B1(new_n789), .B2(new_n205), .ZN(new_n844));
  XNOR2_X1  g0644(.A(new_n844), .B(KEYINPUT96), .ZN(new_n845));
  INV_X1    g0645(.A(G303), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n787), .A2(new_n846), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n775), .A2(new_n211), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n299), .B1(new_n784), .B2(new_n484), .ZN(new_n849));
  NOR4_X1   g0649(.A1(new_n845), .A2(new_n847), .A3(new_n848), .A4(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(G283), .ZN(new_n851));
  OAI221_X1 g0651(.A(new_n850), .B1(new_n206), .B2(new_n773), .C1(new_n851), .C2(new_n769), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n852), .B1(G311), .B2(new_n780), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n763), .B1(new_n842), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n819), .A2(new_n751), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n763), .A2(new_n751), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(new_n432), .ZN(new_n857));
  NAND4_X1  g0657(.A1(new_n854), .A2(new_n748), .A3(new_n855), .A4(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n830), .A2(new_n858), .ZN(G384));
  AND2_X1   g0659(.A1(new_n740), .A2(new_n741), .ZN(new_n860));
  AND2_X1   g0660(.A1(new_n448), .A2(new_n439), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(new_n683), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n440), .A2(new_n684), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n449), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n819), .B1(new_n862), .B2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT102), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT38), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n341), .A2(new_n289), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n302), .B1(new_n311), .B2(new_n313), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n870), .A2(KEYINPUT16), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n294), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n681), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n357), .A2(new_n353), .A3(new_n348), .ZN(new_n875));
  INV_X1    g0675(.A(new_n344), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n874), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n323), .B1(new_n347), .B2(new_n873), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT37), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n331), .A2(new_n342), .ZN(new_n880));
  AND3_X1   g0680(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n872), .A2(new_n347), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n874), .A2(new_n882), .A3(new_n880), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n881), .B1(KEYINPUT37), .B2(new_n883), .ZN(new_n884));
  OAI211_X1 g0684(.A(new_n867), .B(new_n868), .C1(new_n877), .C2(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n868), .B1(new_n877), .B2(new_n884), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n339), .A2(new_n340), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(new_n295), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n290), .B1(new_n870), .B2(KEYINPUT16), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n293), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  OAI22_X1  g0690(.A1(new_n890), .A2(new_n352), .B1(new_n323), .B2(new_n282), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n890), .A2(new_n681), .ZN(new_n892));
  OAI21_X1  g0692(.A(KEYINPUT37), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n895), .B(KEYINPUT38), .C1(new_n358), .C2(new_n874), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n886), .A2(KEYINPUT102), .A3(new_n896), .ZN(new_n897));
  NAND4_X1  g0697(.A1(new_n860), .A2(new_n866), .A3(new_n885), .A4(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT40), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(KEYINPUT103), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT103), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n898), .A2(new_n902), .A3(new_n899), .ZN(new_n903));
  AND2_X1   g0703(.A1(new_n860), .A2(new_n866), .ZN(new_n904));
  AOI211_X1 g0704(.A(new_n342), .B(new_n681), .C1(new_n876), .C2(new_n645), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n879), .B1(new_n878), .B2(new_n880), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n881), .A2(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n868), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n899), .B1(new_n908), .B2(new_n896), .ZN(new_n909));
  AOI22_X1  g0709(.A1(new_n901), .A2(new_n903), .B1(new_n904), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n860), .A2(new_n453), .ZN(new_n911));
  XOR2_X1   g0711(.A(new_n911), .B(KEYINPUT104), .Z(new_n912));
  XNOR2_X1  g0712(.A(new_n910), .B(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(G330), .ZN(new_n914));
  AOI211_X1 g0714(.A(new_n863), .B(new_n442), .C1(new_n448), .C2(new_n439), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n643), .A2(new_n684), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT101), .ZN(new_n918));
  AOI211_X1 g0718(.A(new_n683), .B(new_n819), .C1(new_n665), .C2(new_n670), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n918), .B1(new_n919), .B2(new_n815), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n824), .A2(KEYINPUT101), .A3(new_n816), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n917), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  AND2_X1   g0722(.A1(new_n897), .A2(new_n885), .ZN(new_n923));
  AOI22_X1  g0723(.A1(new_n922), .A2(new_n923), .B1(new_n646), .B2(new_n681), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n897), .A2(KEYINPUT39), .A3(new_n885), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT39), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n908), .A2(new_n926), .A3(new_n896), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n643), .A2(new_n683), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n924), .A2(new_n930), .ZN(new_n931));
  OAI211_X1 g0731(.A(new_n453), .B(new_n717), .C1(new_n718), .C2(new_n727), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n932), .A2(new_n397), .A3(new_n647), .ZN(new_n933));
  INV_X1    g0733(.A(new_n933), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n931), .B(new_n934), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n914), .B(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n936), .B1(new_n255), .B2(new_n677), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n594), .A2(new_n597), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n484), .B1(new_n938), .B2(KEYINPUT35), .ZN(new_n939));
  OAI211_X1 g0739(.A(new_n939), .B(new_n232), .C1(KEYINPUT35), .C2(new_n938), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n940), .B(KEYINPUT36), .ZN(new_n941));
  OAI21_X1  g0741(.A(G77), .B1(new_n837), .B2(new_n219), .ZN(new_n942));
  OAI22_X1  g0742(.A1(new_n942), .A2(new_n228), .B1(G50), .B2(new_n219), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n943), .A2(G1), .A3(new_n676), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n937), .A2(new_n941), .A3(new_n944), .ZN(G367));
  XNOR2_X1  g0745(.A(new_n696), .B(new_n697), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n605), .B1(new_n575), .B2(new_n684), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n666), .A2(new_n683), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n946), .A2(new_n694), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(KEYINPUT42), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n604), .B1(new_n947), .B2(new_n663), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(new_n684), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(KEYINPUT105), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT105), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n951), .A2(new_n956), .A3(new_n953), .ZN(new_n957));
  AND2_X1   g0757(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT43), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n654), .B1(new_n559), .B2(new_n684), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n723), .A2(new_n650), .A3(new_n683), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  OR2_X1    g0763(.A1(new_n950), .A2(KEYINPUT42), .ZN(new_n964));
  NAND4_X1  g0764(.A1(new_n958), .A2(new_n959), .A3(new_n963), .A4(new_n964), .ZN(new_n965));
  AND2_X1   g0765(.A1(new_n695), .A2(new_n949), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n955), .A2(new_n964), .A3(new_n957), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n963), .A2(new_n959), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n962), .A2(KEYINPUT43), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n967), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  AND3_X1   g0770(.A1(new_n965), .A2(new_n966), .A3(new_n970), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n966), .B1(new_n965), .B2(new_n970), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n708), .B(KEYINPUT41), .ZN(new_n974));
  INV_X1    g0774(.A(new_n949), .ZN(new_n975));
  XOR2_X1   g0775(.A(KEYINPUT106), .B(KEYINPUT44), .Z(new_n976));
  NAND3_X1  g0776(.A1(new_n703), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(new_n976), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n701), .B1(new_n946), .B2(new_n694), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n978), .B1(new_n979), .B2(new_n949), .ZN(new_n980));
  AOI21_X1  g0780(.A(KEYINPUT45), .B1(new_n979), .B2(new_n949), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT45), .ZN(new_n982));
  NOR3_X1   g0782(.A1(new_n703), .A2(new_n982), .A3(new_n975), .ZN(new_n983));
  OAI211_X1 g0783(.A(new_n977), .B(new_n980), .C1(new_n981), .C2(new_n983), .ZN(new_n984));
  OAI21_X1  g0784(.A(KEYINPUT107), .B1(new_n984), .B2(new_n695), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n695), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n691), .A2(KEYINPUT108), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n946), .B(new_n694), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(new_n989), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n991), .B1(KEYINPUT108), .B2(new_n691), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n990), .A2(new_n744), .A3(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n993), .A2(KEYINPUT109), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT109), .ZN(new_n995));
  NAND4_X1  g0795(.A1(new_n990), .A2(new_n744), .A3(new_n992), .A4(new_n995), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n984), .A2(KEYINPUT107), .A3(new_n695), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n987), .A2(new_n994), .A3(new_n996), .A4(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n974), .B1(new_n998), .B2(new_n744), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n973), .B1(new_n999), .B2(new_n747), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n764), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n758), .ZN(new_n1002));
  OAI22_X1  g0802(.A1(new_n244), .A2(new_n1002), .B1(new_n224), .B2(new_n409), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n748), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT110), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n299), .B1(new_n789), .B2(new_n206), .ZN(new_n1006));
  INV_X1    g0806(.A(G317), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n794), .A2(new_n846), .B1(new_n779), .B2(new_n1007), .ZN(new_n1008));
  AOI211_X1 g0808(.A(new_n1006), .B(new_n1008), .C1(G294), .C2(new_n802), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n773), .A2(new_n484), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1010), .A2(KEYINPUT46), .ZN(new_n1011));
  INV_X1    g0811(.A(G311), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n1010), .A2(KEYINPUT46), .B1(new_n1012), .B2(new_n787), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n205), .A2(new_n775), .B1(new_n784), .B2(new_n851), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1009), .A2(new_n1011), .A3(new_n1015), .ZN(new_n1016));
  OAI22_X1  g0816(.A1(new_n794), .A2(new_n362), .B1(new_n789), .B2(new_n219), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1017), .B(KEYINPUT111), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n299), .B1(new_n774), .B2(G58), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n776), .A2(G77), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n769), .A2(new_n805), .B1(new_n784), .B2(new_n202), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1021), .B1(G137), .B2(new_n780), .ZN(new_n1022));
  NAND4_X1  g0822(.A1(new_n1018), .A2(new_n1019), .A3(new_n1020), .A4(new_n1022), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n787), .A2(new_n834), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1016), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  XOR2_X1   g0825(.A(new_n1025), .B(KEYINPUT47), .Z(new_n1026));
  INV_X1    g0826(.A(new_n763), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n1005), .B1(new_n1026), .B2(new_n1027), .C1(new_n962), .C2(new_n754), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1000), .A2(new_n1028), .ZN(G387));
  NAND2_X1  g0829(.A1(new_n990), .A2(new_n992), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1030), .A2(new_n743), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1031), .A2(new_n709), .A3(new_n993), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n758), .B1(new_n241), .B2(new_n756), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n711), .B2(new_n761), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n283), .A2(new_n202), .ZN(new_n1035));
  XOR2_X1   g0835(.A(KEYINPUT112), .B(KEYINPUT50), .Z(new_n1036));
  XNOR2_X1  g0836(.A(new_n1035), .B(new_n1036), .ZN(new_n1037));
  AOI21_X1  g0837(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1037), .A2(new_n711), .A3(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1034), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n705), .A2(new_n206), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1001), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n774), .A2(G294), .B1(new_n790), .B2(G283), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(G311), .A2(new_n802), .B1(new_n797), .B2(G317), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n1044), .B1(new_n846), .B2(new_n784), .C1(new_n793), .C2(new_n787), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT48), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1043), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT113), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1048), .B1(new_n1046), .B2(new_n1045), .ZN(new_n1049));
  OR2_X1    g0849(.A1(new_n1049), .A2(KEYINPUT49), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n1049), .A2(KEYINPUT49), .B1(G116), .B2(new_n776), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n780), .A2(G326), .ZN(new_n1052));
  NAND4_X1  g0852(.A1(new_n1050), .A2(new_n1051), .A3(new_n299), .A4(new_n1052), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n284), .A2(new_n769), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(G77), .A2(new_n774), .B1(new_n780), .B2(G150), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n1055), .B1(new_n219), .B2(new_n784), .C1(new_n205), .C2(new_n775), .ZN(new_n1056));
  AOI211_X1 g0856(.A(new_n1054), .B(new_n1056), .C1(G159), .C2(new_n788), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n790), .A2(new_n408), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1057), .B(new_n1058), .C1(new_n202), .C2(new_n794), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1053), .B1(new_n299), .B2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1042), .B1(new_n1060), .B2(new_n763), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n1061), .B(new_n748), .C1(new_n694), .C2(new_n754), .ZN(new_n1062));
  OAI211_X1 g0862(.A(new_n1032), .B(new_n1062), .C1(new_n746), .C2(new_n1030), .ZN(G393));
  XNOR2_X1  g0863(.A(new_n984), .B(new_n695), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1064), .A2(new_n993), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n998), .A2(new_n709), .A3(new_n1065), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n1064), .A2(new_n746), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n748), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n975), .A2(new_n753), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n764), .B1(new_n205), .B2(new_n224), .C1(new_n248), .C2(new_n1002), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n773), .A2(new_n851), .B1(new_n775), .B2(new_n206), .ZN(new_n1072));
  AOI211_X1 g0872(.A(new_n297), .B(new_n1072), .C1(G322), .C2(new_n780), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n802), .A2(G303), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n787), .A2(new_n1007), .B1(new_n794), .B2(new_n1012), .ZN(new_n1075));
  XOR2_X1   g0875(.A(KEYINPUT114), .B(KEYINPUT52), .Z(new_n1076));
  XNOR2_X1  g0876(.A(new_n1075), .B(new_n1076), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(G294), .A2(new_n785), .B1(new_n790), .B2(G116), .ZN(new_n1078));
  NAND4_X1  g0878(.A1(new_n1073), .A2(new_n1074), .A3(new_n1077), .A4(new_n1078), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n787), .A2(new_n362), .B1(new_n794), .B2(new_n805), .ZN(new_n1080));
  XOR2_X1   g0880(.A(new_n1080), .B(KEYINPUT51), .Z(new_n1081));
  AOI211_X1 g0881(.A(new_n299), .B(new_n1081), .C1(G143), .C2(new_n780), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n789), .A2(new_n432), .ZN(new_n1083));
  AOI211_X1 g0883(.A(new_n1083), .B(new_n848), .C1(G68), .C2(new_n774), .ZN(new_n1084));
  OAI211_X1 g0884(.A(new_n1082), .B(new_n1084), .C1(new_n284), .C2(new_n784), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n769), .A2(new_n202), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1079), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  AOI211_X1 g0887(.A(new_n1068), .B(new_n1071), .C1(new_n763), .C2(new_n1087), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n1067), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1066), .A2(new_n1089), .ZN(G390));
  OAI21_X1  g0890(.A(new_n299), .B1(new_n773), .B2(new_n211), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(new_n1091), .B(KEYINPUT115), .ZN(new_n1092));
  AOI211_X1 g0892(.A(new_n1083), .B(new_n1092), .C1(G294), .C2(new_n780), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n785), .A2(G97), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(G107), .A2(new_n802), .B1(new_n797), .B2(G116), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n839), .B1(G283), .B2(new_n788), .ZN(new_n1096));
  NAND4_X1  g0896(.A1(new_n1093), .A2(new_n1094), .A3(new_n1095), .A4(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(G128), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n787), .A2(new_n1098), .B1(new_n794), .B2(new_n840), .ZN(new_n1099));
  INV_X1    g0899(.A(KEYINPUT53), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1100), .B1(new_n774), .B2(G150), .ZN(new_n1101));
  AOI211_X1 g0901(.A(new_n1099), .B(new_n1101), .C1(G50), .C2(new_n776), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n297), .B1(new_n769), .B2(new_n831), .ZN(new_n1103));
  XOR2_X1   g0903(.A(KEYINPUT54), .B(G143), .Z(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n1105), .A2(new_n784), .ZN(new_n1106));
  AOI211_X1 g0906(.A(new_n1103), .B(new_n1106), .C1(G125), .C2(new_n780), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n790), .A2(G159), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n774), .A2(new_n1100), .A3(G150), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n1102), .A2(new_n1107), .A3(new_n1108), .A4(new_n1109), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1027), .B1(new_n1097), .B2(new_n1110), .ZN(new_n1111));
  AOI211_X1 g0911(.A(new_n1068), .B(new_n1111), .C1(new_n284), .C2(new_n856), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1112), .B1(new_n928), .B2(new_n752), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n823), .B1(new_n915), .B2(new_n916), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n1114), .A2(new_n742), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n917), .ZN(new_n1116));
  AOI211_X1 g0916(.A(new_n918), .B(new_n815), .C1(new_n714), .C2(new_n823), .ZN(new_n1117));
  AOI21_X1  g0917(.A(KEYINPUT101), .B1(new_n824), .B2(new_n816), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1116), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n929), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n928), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n908), .A2(new_n896), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(new_n1120), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n817), .A2(new_n818), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n816), .B1(new_n727), .B2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1123), .B1(new_n1125), .B2(new_n1116), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1115), .B1(new_n1121), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1125), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n1122), .B(new_n1120), .C1(new_n1128), .C2(new_n917), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n828), .A2(new_n866), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n922), .A2(new_n929), .ZN(new_n1131));
  OAI211_X1 g0931(.A(new_n1129), .B(new_n1130), .C1(new_n1131), .C2(new_n928), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1127), .A2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1113), .B1(new_n1133), .B2(new_n746), .ZN(new_n1134));
  NAND4_X1  g0934(.A1(new_n453), .A2(G330), .A3(new_n740), .A4(new_n741), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n932), .A2(new_n1135), .A3(new_n397), .A4(new_n647), .ZN(new_n1136));
  NAND4_X1  g0936(.A1(new_n740), .A2(G330), .A3(new_n741), .A4(new_n823), .ZN(new_n1137));
  AND2_X1   g0937(.A1(new_n1137), .A2(new_n917), .ZN(new_n1138));
  OAI22_X1  g0938(.A1(new_n1138), .A2(new_n1115), .B1(new_n1118), .B2(new_n1117), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n917), .B1(new_n742), .B2(new_n820), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1130), .A2(new_n1140), .A3(new_n1128), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1136), .B1(new_n1139), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n708), .B1(new_n1133), .B2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1127), .A2(new_n1132), .A3(new_n1142), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1134), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(G378));
  NAND2_X1  g0947(.A1(new_n371), .A2(new_n873), .ZN(new_n1148));
  XNOR2_X1  g0948(.A(new_n398), .B(new_n1148), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(new_n1151));
  OR2_X1    g0951(.A1(new_n1149), .A2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1149), .A2(new_n1151), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1152), .A2(KEYINPUT118), .A3(new_n1153), .ZN(new_n1154));
  AND3_X1   g0954(.A1(new_n924), .A2(new_n930), .A3(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1154), .B1(new_n924), .B2(new_n930), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n910), .B(G330), .C1(new_n1155), .C2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n904), .A2(new_n909), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n903), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n902), .B1(new_n898), .B2(new_n899), .ZN(new_n1160));
  OAI211_X1 g0960(.A(G330), .B(new_n1158), .C1(new_n1159), .C2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1154), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n931), .A2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n924), .A2(new_n930), .A3(new_n1154), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1161), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1157), .A2(new_n1165), .A3(new_n747), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1152), .A2(new_n751), .A3(new_n1153), .ZN(new_n1167));
  OAI22_X1  g0967(.A1(new_n794), .A2(new_n1098), .B1(new_n784), .B2(new_n831), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n1105), .A2(new_n773), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1168), .B1(new_n1170), .B2(KEYINPUT117), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n790), .A2(G150), .ZN(new_n1172));
  INV_X1    g0972(.A(KEYINPUT117), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(new_n1169), .A2(new_n1173), .B1(G132), .B2(new_n802), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n788), .A2(G125), .ZN(new_n1175));
  NAND4_X1  g0975(.A1(new_n1171), .A2(new_n1172), .A3(new_n1174), .A4(new_n1175), .ZN(new_n1176));
  XOR2_X1   g0976(.A(new_n1176), .B(KEYINPUT59), .Z(new_n1177));
  OAI21_X1  g0977(.A(new_n259), .B1(new_n775), .B2(new_n805), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(G124), .B2(new_n780), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1177), .A2(new_n460), .A3(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(G41), .B1(KEYINPUT3), .B2(G33), .ZN(new_n1181));
  OAI21_X1  g0981(.A(KEYINPUT116), .B1(new_n1181), .B2(G50), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n769), .A2(new_n205), .B1(new_n775), .B2(new_n837), .ZN(new_n1183));
  AOI211_X1 g0983(.A(new_n297), .B(new_n1183), .C1(G283), .C2(new_n780), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1184), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n787), .A2(new_n484), .ZN(new_n1186));
  AOI21_X1  g0986(.A(G41), .B1(new_n790), .B2(G68), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(G77), .A2(new_n774), .B1(new_n797), .B2(G107), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1189), .B1(new_n409), .B2(new_n784), .ZN(new_n1190));
  NOR4_X1   g0990(.A1(new_n1185), .A2(new_n1186), .A3(new_n1188), .A4(new_n1190), .ZN(new_n1191));
  OR2_X1    g0991(.A1(new_n1191), .A2(KEYINPUT58), .ZN(new_n1192));
  NOR3_X1   g0992(.A1(new_n1181), .A2(KEYINPUT116), .A3(G50), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(new_n1191), .B2(KEYINPUT58), .ZN(new_n1194));
  NAND4_X1  g0994(.A1(new_n1180), .A2(new_n1182), .A3(new_n1192), .A4(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1195), .A2(new_n763), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n856), .A2(new_n202), .ZN(new_n1197));
  NAND4_X1  g0997(.A1(new_n1167), .A2(new_n748), .A3(new_n1196), .A4(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1166), .A2(new_n1198), .ZN(new_n1199));
  XNOR2_X1  g0999(.A(new_n1136), .B(KEYINPUT119), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1145), .A2(new_n1200), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1201), .A2(new_n1157), .A3(new_n1165), .ZN(new_n1202));
  INV_X1    g1002(.A(KEYINPUT57), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n708), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n1201), .A2(new_n1157), .A3(new_n1165), .A4(KEYINPUT57), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1199), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(G375));
  INV_X1    g1007(.A(new_n974), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1139), .A2(new_n1136), .A3(new_n1141), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1143), .A2(new_n1208), .A3(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n856), .A2(new_n219), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n748), .B(new_n1211), .C1(new_n1116), .C2(new_n752), .ZN(new_n1212));
  OAI221_X1 g1012(.A(new_n1058), .B1(new_n851), .B2(new_n794), .C1(new_n846), .C2(new_n779), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(G107), .B2(new_n785), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1214), .B1(new_n205), .B2(new_n773), .ZN(new_n1215));
  OAI221_X1 g1015(.A(new_n1020), .B1(new_n484), .B2(new_n769), .C1(new_n843), .C2(new_n787), .ZN(new_n1216));
  NOR3_X1   g1016(.A1(new_n1215), .A2(new_n297), .A3(new_n1216), .ZN(new_n1217));
  XOR2_X1   g1017(.A(new_n1217), .B(KEYINPUT120), .Z(new_n1218));
  NOR2_X1   g1018(.A1(new_n773), .A2(new_n805), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(G137), .A2(new_n797), .B1(new_n802), .B2(new_n1104), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1220), .B1(new_n840), .B2(new_n787), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT121), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  OAI22_X1  g1023(.A1(new_n837), .A2(new_n775), .B1(new_n784), .B2(new_n362), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n297), .B1(new_n779), .B2(new_n1098), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1226), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1227));
  OAI211_X1 g1027(.A(new_n1225), .B(new_n1227), .C1(new_n202), .C2(new_n789), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1218), .B1(new_n1219), .B2(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1212), .B1(new_n763), .B2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1230), .B1(new_n1231), .B2(new_n747), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1210), .A2(new_n1232), .ZN(G381));
  NAND2_X1  g1033(.A1(new_n1206), .A2(new_n1146), .ZN(new_n1234));
  INV_X1    g1034(.A(G390), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1235), .A2(new_n1000), .A3(new_n1028), .ZN(new_n1236));
  OR3_X1    g1036(.A1(G393), .A2(G381), .A3(G396), .ZN(new_n1237));
  NOR3_X1   g1037(.A1(new_n1236), .A2(G384), .A3(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT122), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1234), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1240), .B1(new_n1239), .B2(new_n1238), .ZN(G407));
  OAI211_X1 g1041(.A(G407), .B(G213), .C1(G343), .C2(new_n1234), .ZN(G409));
  NAND2_X1  g1042(.A1(G387), .A2(G390), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT124), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1243), .A2(new_n1244), .A3(new_n1236), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1245), .A2(KEYINPUT125), .ZN(new_n1246));
  XNOR2_X1  g1046(.A(G393), .B(G396), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1246), .A2(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT125), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1243), .A2(new_n1250), .A3(new_n1236), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1245), .A2(KEYINPUT125), .A3(new_n1247), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1249), .A2(new_n1251), .A3(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1254), .A2(new_n709), .A3(new_n1205), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1199), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1146), .B1(new_n1255), .B2(new_n1256), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1201), .A2(new_n1157), .A3(new_n1165), .A4(new_n1208), .ZN(new_n1258));
  AND3_X1   g1058(.A1(new_n1256), .A2(new_n1146), .A3(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n682), .A2(G213), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  NOR3_X1   g1061(.A1(new_n1257), .A2(new_n1259), .A3(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(G384), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT60), .ZN(new_n1264));
  OAI211_X1 g1064(.A(new_n1143), .B(new_n709), .C1(new_n1264), .C2(new_n1209), .ZN(new_n1265));
  AND2_X1   g1065(.A1(new_n1209), .A2(new_n1264), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1232), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1263), .A2(new_n1267), .ZN(new_n1268));
  OAI211_X1 g1068(.A(G384), .B(new_n1232), .C1(new_n1265), .C2(new_n1266), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT63), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  AOI21_X1  g1072(.A(KEYINPUT61), .B1(new_n1262), .B2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT123), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1274), .B1(new_n1257), .B2(new_n1259), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1256), .A2(new_n1146), .A3(new_n1258), .ZN(new_n1276));
  OAI211_X1 g1076(.A(KEYINPUT123), .B(new_n1276), .C1(new_n1206), .C2(new_n1146), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1275), .A2(new_n1260), .A3(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1261), .A2(G2897), .ZN(new_n1279));
  XOR2_X1   g1079(.A(new_n1270), .B(new_n1279), .Z(new_n1280));
  INV_X1    g1080(.A(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1271), .B1(new_n1278), .B2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1270), .ZN(new_n1283));
  NAND4_X1  g1083(.A1(new_n1275), .A2(new_n1283), .A3(new_n1260), .A4(new_n1277), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1284), .ZN(new_n1285));
  OAI211_X1 g1085(.A(new_n1253), .B(new_n1273), .C1(new_n1282), .C2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1252), .A2(new_n1251), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1247), .B1(new_n1245), .B2(KEYINPUT125), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1268), .A2(new_n1269), .A3(KEYINPUT62), .ZN(new_n1290));
  NOR4_X1   g1090(.A1(new_n1257), .A2(new_n1259), .A3(new_n1290), .A4(new_n1261), .ZN(new_n1291));
  XNOR2_X1  g1091(.A(KEYINPUT127), .B(KEYINPUT62), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1291), .B1(new_n1284), .B2(new_n1292), .ZN(new_n1293));
  XNOR2_X1  g1093(.A(KEYINPUT126), .B(KEYINPUT61), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1294), .B1(new_n1280), .B2(new_n1262), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1289), .B1(new_n1293), .B2(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1286), .A2(new_n1296), .ZN(G405));
  INV_X1    g1097(.A(new_n1234), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1283), .B1(new_n1298), .B2(new_n1257), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1257), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1300), .A2(new_n1234), .A3(new_n1270), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1299), .A2(new_n1301), .ZN(new_n1302));
  XNOR2_X1  g1102(.A(new_n1253), .B(new_n1302), .ZN(G402));
endmodule


