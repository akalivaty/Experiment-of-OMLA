//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 1 0 1 0 0 1 1 0 0 0 0 1 0 1 0 0 1 1 0 1 1 0 1 1 0 0 0 1 1 0 0 1 0 0 1 0 0 1 0 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:54 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n697, new_n698, new_n699,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n710, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n730, new_n731,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n877,
    new_n878, new_n879, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n903, new_n904, new_n905, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952;
  INV_X1    g000(.A(G137), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G134), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT11), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n187), .A2(KEYINPUT11), .A3(G134), .ZN(new_n191));
  INV_X1    g005(.A(G134), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G137), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n190), .A2(new_n191), .A3(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G131), .ZN(new_n195));
  INV_X1    g009(.A(G131), .ZN(new_n196));
  NAND4_X1  g010(.A1(new_n190), .A2(new_n191), .A3(new_n196), .A4(new_n193), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G146), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G143), .ZN(new_n200));
  INV_X1    g014(.A(G143), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G146), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n200), .A2(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(KEYINPUT0), .A2(G128), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT64), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT0), .ZN(new_n206));
  INV_X1    g020(.A(G128), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n205), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  OAI21_X1  g022(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n209));
  NAND4_X1  g023(.A1(new_n203), .A2(new_n204), .A3(new_n208), .A4(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT65), .ZN(new_n211));
  XNOR2_X1  g025(.A(G143), .B(G146), .ZN(new_n212));
  INV_X1    g026(.A(new_n204), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n210), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(new_n209), .ZN(new_n216));
  NOR3_X1   g030(.A1(KEYINPUT64), .A2(KEYINPUT0), .A3(G128), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n218), .A2(new_n211), .A3(new_n204), .A4(new_n203), .ZN(new_n219));
  AND3_X1   g033(.A1(new_n215), .A2(KEYINPUT70), .A3(new_n219), .ZN(new_n220));
  AOI21_X1  g034(.A(KEYINPUT70), .B1(new_n215), .B2(new_n219), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n198), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT2), .ZN(new_n223));
  INV_X1    g037(.A(G113), .ZN(new_n224));
  OAI21_X1  g038(.A(KEYINPUT68), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT68), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n226), .A2(KEYINPUT2), .A3(G113), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n223), .A2(new_n224), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(G119), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(G116), .ZN(new_n232));
  INV_X1    g046(.A(G116), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(G119), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n230), .A2(new_n235), .ZN(new_n236));
  AOI22_X1  g050(.A1(new_n225), .A2(new_n227), .B1(new_n223), .B2(new_n224), .ZN(new_n237));
  INV_X1    g051(.A(new_n235), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  AND3_X1   g053(.A1(new_n236), .A2(KEYINPUT69), .A3(new_n239), .ZN(new_n240));
  AOI21_X1  g054(.A(KEYINPUT69), .B1(new_n236), .B2(new_n239), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n188), .A2(new_n193), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G131), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(KEYINPUT66), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT66), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n243), .A2(new_n246), .A3(G131), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n245), .A2(new_n197), .A3(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT71), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  XNOR2_X1  g064(.A(KEYINPUT67), .B(G128), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n200), .A2(KEYINPUT1), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(new_n203), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT1), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n212), .A2(new_n255), .A3(G128), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n245), .A2(KEYINPUT71), .A3(new_n247), .A4(new_n197), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n250), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n222), .A2(new_n242), .A3(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT72), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND4_X1  g076(.A1(new_n222), .A2(new_n242), .A3(new_n259), .A4(KEYINPUT72), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(G237), .ZN(new_n265));
  INV_X1    g079(.A(G953), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n265), .A2(new_n266), .A3(G210), .ZN(new_n267));
  INV_X1    g081(.A(G101), .ZN(new_n268));
  XNOR2_X1  g082(.A(new_n267), .B(new_n268), .ZN(new_n269));
  XNOR2_X1  g083(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n270));
  XOR2_X1   g084(.A(new_n269), .B(new_n270), .Z(new_n271));
  INV_X1    g085(.A(new_n242), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT30), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n273), .B1(new_n222), .B2(new_n259), .ZN(new_n274));
  AND2_X1   g088(.A1(new_n215), .A2(new_n219), .ZN(new_n275));
  INV_X1    g089(.A(new_n198), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n257), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n278), .A2(new_n248), .ZN(new_n279));
  NOR3_X1   g093(.A1(new_n277), .A2(new_n279), .A3(KEYINPUT30), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n272), .B1(new_n274), .B2(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n264), .A2(new_n271), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(KEYINPUT73), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT73), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n264), .A2(new_n281), .A3(new_n284), .A4(new_n271), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n283), .A2(KEYINPUT31), .A3(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT31), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n282), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n272), .B1(new_n277), .B2(new_n279), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT28), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n260), .A2(new_n291), .ZN(new_n292));
  OAI211_X1 g106(.A(new_n290), .B(new_n292), .C1(new_n264), .C2(new_n291), .ZN(new_n293));
  INV_X1    g107(.A(new_n271), .ZN(new_n294));
  AND2_X1   g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n289), .A2(new_n296), .ZN(new_n297));
  NOR2_X1   g111(.A1(G472), .A2(G902), .ZN(new_n298));
  XOR2_X1   g112(.A(new_n298), .B(KEYINPUT74), .Z(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n297), .A2(KEYINPUT32), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(KEYINPUT76), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT76), .ZN(new_n303));
  NAND4_X1  g117(.A1(new_n297), .A2(new_n303), .A3(KEYINPUT32), .A4(new_n300), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n264), .A2(new_n281), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n307), .A2(new_n271), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n293), .A2(new_n294), .ZN(new_n309));
  NOR3_X1   g123(.A1(new_n308), .A2(new_n309), .A3(KEYINPUT29), .ZN(new_n310));
  INV_X1    g124(.A(G902), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n222), .A2(new_n259), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(new_n272), .ZN(new_n313));
  OAI211_X1 g127(.A(new_n292), .B(new_n313), .C1(new_n264), .C2(new_n291), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n271), .A2(KEYINPUT29), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n311), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  OAI21_X1  g130(.A(G472), .B1(new_n310), .B2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT32), .ZN(new_n318));
  AOI21_X1  g132(.A(KEYINPUT75), .B1(new_n297), .B2(new_n300), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n295), .B1(new_n286), .B2(new_n288), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT75), .ZN(new_n321));
  NOR3_X1   g135(.A1(new_n320), .A2(new_n321), .A3(new_n299), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n318), .B1(new_n319), .B2(new_n322), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n305), .A2(new_n317), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n231), .A2(G128), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n325), .B1(new_n251), .B2(new_n231), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT77), .ZN(new_n327));
  XNOR2_X1  g141(.A(new_n326), .B(new_n327), .ZN(new_n328));
  XOR2_X1   g142(.A(KEYINPUT24), .B(G110), .Z(new_n329));
  NOR2_X1   g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT23), .ZN(new_n331));
  OR2_X1    g145(.A1(new_n326), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n331), .A2(new_n207), .A3(G119), .ZN(new_n333));
  AOI21_X1  g147(.A(G110), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n330), .A2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT16), .ZN(new_n336));
  INV_X1    g150(.A(G140), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(G125), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n337), .A2(G125), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n338), .B1(new_n339), .B2(KEYINPUT78), .ZN(new_n340));
  INV_X1    g154(.A(G125), .ZN(new_n341));
  OR3_X1    g155(.A1(new_n341), .A2(KEYINPUT78), .A3(G140), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n336), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n341), .A2(G140), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n344), .A2(KEYINPUT16), .ZN(new_n345));
  OAI21_X1  g159(.A(G146), .B1(new_n343), .B2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(new_n346), .ZN(new_n347));
  NOR3_X1   g161(.A1(new_n344), .A2(new_n339), .A3(G146), .ZN(new_n348));
  OR2_X1    g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT79), .ZN(new_n350));
  OR3_X1    g164(.A1(new_n335), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n328), .A2(new_n329), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n332), .A2(G110), .A3(new_n333), .ZN(new_n353));
  NOR3_X1   g167(.A1(new_n343), .A2(G146), .A3(new_n345), .ZN(new_n354));
  OAI211_X1 g168(.A(new_n352), .B(new_n353), .C1(new_n347), .C2(new_n354), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n350), .B1(new_n335), .B2(new_n349), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n351), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  XNOR2_X1  g171(.A(KEYINPUT22), .B(G137), .ZN(new_n358));
  INV_X1    g172(.A(G221), .ZN(new_n359));
  INV_X1    g173(.A(G234), .ZN(new_n360));
  NOR3_X1   g174(.A1(new_n359), .A2(new_n360), .A3(G953), .ZN(new_n361));
  XOR2_X1   g175(.A(new_n358), .B(new_n361), .Z(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n357), .A2(new_n363), .ZN(new_n364));
  NAND4_X1  g178(.A1(new_n351), .A2(new_n355), .A3(new_n356), .A4(new_n362), .ZN(new_n365));
  AND2_X1   g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(G217), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n367), .B1(G234), .B2(new_n311), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n368), .A2(G902), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n366), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n364), .A2(new_n311), .A3(new_n365), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT25), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n364), .A2(KEYINPUT25), .A3(new_n311), .A4(new_n365), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n373), .A2(KEYINPUT80), .A3(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT80), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n371), .A2(new_n377), .A3(new_n372), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(new_n368), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n370), .B1(new_n376), .B2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(new_n380), .ZN(new_n381));
  OAI21_X1  g195(.A(KEYINPUT88), .B1(new_n347), .B2(new_n354), .ZN(new_n382));
  OR3_X1    g196(.A1(new_n343), .A2(G146), .A3(new_n345), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT88), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n383), .A2(new_n384), .A3(new_n346), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n265), .A2(new_n266), .A3(G214), .ZN(new_n386));
  XNOR2_X1  g200(.A(new_n386), .B(G143), .ZN(new_n387));
  OR2_X1    g201(.A1(new_n387), .A2(new_n196), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT17), .ZN(new_n389));
  OR2_X1    g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n382), .A2(new_n385), .A3(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT89), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND4_X1  g207(.A1(new_n382), .A2(KEYINPUT89), .A3(new_n385), .A4(new_n390), .ZN(new_n394));
  XNOR2_X1  g208(.A(new_n387), .B(G131), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(new_n389), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n393), .A2(new_n394), .A3(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT18), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n387), .B1(new_n398), .B2(new_n196), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n199), .B1(new_n340), .B2(new_n342), .ZN(new_n400));
  OAI221_X1 g214(.A(new_n399), .B1(new_n348), .B2(new_n400), .C1(new_n388), .C2(new_n398), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n397), .A2(new_n401), .ZN(new_n402));
  XNOR2_X1  g216(.A(G113), .B(G122), .ZN(new_n403));
  INV_X1    g217(.A(G104), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n403), .B(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n402), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n397), .A2(new_n405), .A3(new_n401), .ZN(new_n408));
  AOI21_X1  g222(.A(G902), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n395), .A2(new_n347), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n344), .A2(new_n339), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n340), .A2(new_n342), .ZN(new_n413));
  MUX2_X1   g227(.A(new_n412), .B(new_n413), .S(KEYINPUT19), .Z(new_n414));
  OAI21_X1  g228(.A(new_n411), .B1(G146), .B2(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n405), .B1(new_n415), .B2(new_n401), .ZN(new_n416));
  INV_X1    g230(.A(new_n401), .ZN(new_n417));
  AOI22_X1  g231(.A1(new_n391), .A2(new_n392), .B1(new_n389), .B2(new_n395), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n417), .B1(new_n418), .B2(new_n394), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n416), .B1(new_n419), .B2(new_n405), .ZN(new_n420));
  NOR2_X1   g234(.A1(G475), .A2(G902), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  OAI21_X1  g236(.A(KEYINPUT20), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n416), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n408), .A2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT20), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n425), .A2(new_n426), .A3(new_n421), .ZN(new_n427));
  AOI22_X1  g241(.A1(new_n410), .A2(G475), .B1(new_n423), .B2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(G952), .ZN(new_n429));
  AOI211_X1 g243(.A(G953), .B(new_n429), .C1(G234), .C2(G237), .ZN(new_n430));
  OAI211_X1 g244(.A(G902), .B(G953), .C1(new_n360), .C2(new_n265), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n431), .B(KEYINPUT93), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  XOR2_X1   g247(.A(KEYINPUT21), .B(G898), .Z(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n430), .B1(new_n433), .B2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n207), .A2(G143), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n439), .B1(new_n251), .B2(new_n201), .ZN(new_n440));
  XNOR2_X1  g254(.A(new_n440), .B(G134), .ZN(new_n441));
  INV_X1    g255(.A(G122), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(G116), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n233), .A2(G122), .ZN(new_n444));
  AND2_X1   g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(G107), .ZN(new_n446));
  AND2_X1   g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  OAI21_X1  g261(.A(KEYINPUT90), .B1(new_n444), .B2(KEYINPUT14), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT90), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT14), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n449), .A2(new_n450), .A3(new_n233), .A4(G122), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n444), .A2(KEYINPUT14), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n448), .A2(new_n443), .A3(new_n451), .A4(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n447), .B1(new_n453), .B2(G107), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n441), .A2(new_n454), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n445), .B(new_n446), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT13), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n192), .B1(new_n438), .B2(new_n457), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n458), .B1(new_n440), .B2(new_n457), .ZN(new_n459));
  OAI211_X1 g273(.A(new_n456), .B(new_n459), .C1(G134), .C2(new_n440), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n455), .A2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT91), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  XOR2_X1   g277(.A(KEYINPUT9), .B(G234), .Z(new_n464));
  NAND3_X1  g278(.A1(new_n464), .A2(G217), .A3(new_n266), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n455), .A2(KEYINPUT91), .A3(new_n460), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n463), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n465), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n461), .A2(new_n462), .A3(new_n468), .ZN(new_n469));
  AND2_X1   g283(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT92), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n470), .A2(new_n471), .A3(new_n311), .ZN(new_n472));
  INV_X1    g286(.A(G478), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n473), .A2(KEYINPUT15), .ZN(new_n474));
  OR2_X1    g288(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n470), .A2(new_n311), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n474), .B1(new_n476), .B2(KEYINPUT92), .ZN(new_n477));
  INV_X1    g291(.A(new_n472), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n475), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n428), .A2(new_n437), .A3(new_n480), .ZN(new_n481));
  OAI21_X1  g295(.A(G214), .B1(G237), .B2(G902), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  XNOR2_X1  g297(.A(G110), .B(G122), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n446), .A2(G104), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT3), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n487), .B1(new_n404), .B2(G107), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n446), .A2(KEYINPUT3), .A3(G104), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n486), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  OR3_X1    g304(.A1(new_n490), .A2(KEYINPUT4), .A3(new_n268), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n268), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(KEYINPUT4), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n490), .A2(new_n268), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n491), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n242), .A2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT85), .ZN(new_n497));
  OAI21_X1  g311(.A(G113), .B1(new_n232), .B2(KEYINPUT5), .ZN(new_n498));
  AND3_X1   g312(.A1(new_n232), .A2(new_n234), .A3(KEYINPUT5), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n239), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n404), .A2(G107), .ZN(new_n501));
  OAI21_X1  g315(.A(G101), .B1(new_n486), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n492), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n497), .B1(new_n500), .B2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n503), .ZN(new_n505));
  INV_X1    g319(.A(new_n499), .ZN(new_n506));
  INV_X1    g320(.A(new_n498), .ZN(new_n507));
  AOI22_X1  g321(.A1(new_n506), .A2(new_n507), .B1(new_n237), .B2(new_n238), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n505), .A2(KEYINPUT85), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n504), .A2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n485), .B1(new_n496), .B2(new_n511), .ZN(new_n512));
  OAI211_X1 g326(.A(new_n510), .B(new_n484), .C1(new_n242), .C2(new_n495), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n512), .A2(new_n513), .A3(KEYINPUT6), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT6), .ZN(new_n515));
  OAI211_X1 g329(.A(new_n515), .B(new_n485), .C1(new_n496), .C2(new_n511), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n275), .A2(G125), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n278), .A2(new_n341), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  XOR2_X1   g333(.A(KEYINPUT86), .B(G224), .Z(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(new_n266), .ZN(new_n521));
  XOR2_X1   g335(.A(new_n519), .B(new_n521), .Z(new_n522));
  NAND3_X1  g336(.A1(new_n514), .A2(new_n516), .A3(new_n522), .ZN(new_n523));
  OAI21_X1  g337(.A(G210), .B1(G237), .B2(G902), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n521), .A2(KEYINPUT7), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n519), .A2(new_n525), .ZN(new_n526));
  XNOR2_X1  g340(.A(new_n484), .B(KEYINPUT8), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n508), .A2(new_n503), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT87), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n498), .B1(new_n506), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n499), .A2(KEYINPUT87), .ZN(new_n531));
  AOI22_X1  g345(.A1(new_n530), .A2(new_n531), .B1(new_n237), .B2(new_n238), .ZN(new_n532));
  OAI211_X1 g346(.A(new_n527), .B(new_n528), .C1(new_n532), .C2(new_n503), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n526), .A2(new_n533), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n519), .A2(new_n525), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(G902), .B1(new_n536), .B2(new_n513), .ZN(new_n537));
  AND3_X1   g351(.A1(new_n523), .A2(new_n524), .A3(new_n537), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n524), .B1(new_n523), .B2(new_n537), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n359), .B1(new_n464), .B2(new_n311), .ZN(new_n541));
  INV_X1    g355(.A(G469), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT82), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n256), .A2(new_n543), .ZN(new_n544));
  NAND4_X1  g358(.A1(new_n212), .A2(KEYINPUT82), .A3(new_n255), .A4(G128), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n252), .A2(G128), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(new_n203), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n544), .A2(new_n545), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n505), .A2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT10), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n550), .B1(new_n254), .B2(new_n256), .ZN(new_n551));
  AOI22_X1  g365(.A1(new_n549), .A2(new_n550), .B1(new_n505), .B2(new_n551), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n220), .A2(new_n221), .ZN(new_n553));
  OAI211_X1 g367(.A(new_n552), .B(new_n276), .C1(new_n553), .C2(new_n495), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT84), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n266), .A2(G227), .ZN(new_n556));
  XNOR2_X1  g370(.A(new_n556), .B(KEYINPUT81), .ZN(new_n557));
  XNOR2_X1  g371(.A(G110), .B(G140), .ZN(new_n558));
  XNOR2_X1  g372(.A(new_n557), .B(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  AND3_X1   g374(.A1(new_n554), .A2(new_n555), .A3(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n555), .B1(new_n554), .B2(new_n560), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n505), .A2(new_n257), .ZN(new_n563));
  AOI22_X1  g377(.A1(new_n256), .A2(new_n543), .B1(new_n546), .B2(new_n203), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n503), .B1(new_n545), .B2(new_n564), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n198), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(KEYINPUT83), .A2(KEYINPUT12), .ZN(new_n567));
  NOR2_X1   g381(.A1(KEYINPUT83), .A2(KEYINPUT12), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n566), .A2(new_n567), .A3(new_n569), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n549), .B1(new_n257), .B2(new_n505), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT83), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT12), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n571), .A2(new_n572), .A3(new_n573), .A4(new_n198), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n570), .A2(new_n574), .ZN(new_n575));
  NOR3_X1   g389(.A1(new_n561), .A2(new_n562), .A3(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n552), .B1(new_n553), .B2(new_n495), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(new_n198), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n560), .B1(new_n578), .B2(new_n554), .ZN(new_n579));
  OAI211_X1 g393(.A(new_n542), .B(new_n311), .C1(new_n576), .C2(new_n579), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n542), .A2(new_n311), .ZN(new_n581));
  AND2_X1   g395(.A1(new_n554), .A2(new_n560), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n554), .A2(new_n570), .A3(new_n574), .ZN(new_n583));
  AOI22_X1  g397(.A1(new_n582), .A2(new_n578), .B1(new_n583), .B2(new_n559), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n581), .B1(new_n584), .B2(G469), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n541), .B1(new_n580), .B2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  NOR4_X1   g401(.A1(new_n481), .A2(new_n483), .A3(new_n540), .A4(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n324), .A2(new_n381), .A3(new_n588), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n589), .B(G101), .ZN(G3));
  NAND2_X1  g404(.A1(new_n297), .A2(new_n311), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(G472), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT94), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n591), .A2(KEYINPUT94), .A3(G472), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n319), .ZN(new_n597));
  INV_X1    g411(.A(new_n322), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n600), .A2(new_n587), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(new_n381), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT95), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n539), .A2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n540), .ZN(new_n605));
  OAI211_X1 g419(.A(new_n482), .B(new_n604), .C1(new_n605), .C2(new_n603), .ZN(new_n606));
  AND2_X1   g420(.A1(new_n465), .A2(KEYINPUT98), .ZN(new_n607));
  OAI21_X1  g421(.A(KEYINPUT33), .B1(new_n461), .B2(new_n607), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n608), .B1(new_n461), .B2(new_n607), .ZN(new_n609));
  XNOR2_X1  g423(.A(KEYINPUT96), .B(KEYINPUT33), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n467), .A2(new_n469), .A3(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT97), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n467), .A2(KEYINPUT97), .A3(new_n469), .A4(new_n610), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n609), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n615), .A2(G478), .A3(new_n311), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n476), .A2(new_n473), .ZN(new_n617));
  AND2_X1   g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n428), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(new_n437), .ZN(new_n620));
  NOR3_X1   g434(.A1(new_n602), .A2(new_n606), .A3(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(KEYINPUT34), .B(G104), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n621), .B(new_n622), .ZN(G6));
  NAND2_X1  g437(.A1(new_n604), .A2(new_n482), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n624), .B1(new_n540), .B2(KEYINPUT95), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n423), .A2(new_n427), .ZN(new_n626));
  INV_X1    g440(.A(G475), .ZN(new_n627));
  OAI211_X1 g441(.A(new_n626), .B(new_n479), .C1(new_n627), .C2(new_n409), .ZN(new_n628));
  NOR3_X1   g442(.A1(new_n380), .A2(new_n436), .A3(new_n628), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n601), .A2(new_n625), .A3(new_n629), .ZN(new_n630));
  XOR2_X1   g444(.A(KEYINPUT35), .B(G107), .Z(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G9));
  AOI22_X1  g446(.A1(new_n594), .A2(new_n595), .B1(new_n597), .B2(new_n598), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n363), .A2(KEYINPUT36), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(KEYINPUT99), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n357), .B(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(new_n369), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n637), .B1(new_n376), .B2(new_n379), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n633), .A2(new_n588), .A3(new_n638), .ZN(new_n639));
  XOR2_X1   g453(.A(KEYINPUT37), .B(G110), .Z(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G12));
  INV_X1    g455(.A(new_n379), .ZN(new_n642));
  AOI22_X1  g456(.A1(new_n642), .A2(new_n375), .B1(new_n369), .B2(new_n636), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n643), .A2(new_n587), .ZN(new_n644));
  XNOR2_X1  g458(.A(KEYINPUT100), .B(G900), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n433), .A2(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n430), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  NOR3_X1   g463(.A1(new_n606), .A2(new_n628), .A3(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n324), .A2(new_n644), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(G128), .ZN(G30));
  XNOR2_X1  g466(.A(new_n540), .B(KEYINPUT38), .ZN(new_n653));
  NOR3_X1   g467(.A1(new_n653), .A2(new_n638), .A3(new_n483), .ZN(new_n654));
  XOR2_X1   g468(.A(new_n648), .B(KEYINPUT39), .Z(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n586), .A2(new_n656), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n654), .B1(KEYINPUT40), .B2(new_n657), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n271), .B1(new_n264), .B2(new_n313), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n659), .B1(new_n283), .B2(new_n285), .ZN(new_n660));
  AND2_X1   g474(.A1(new_n660), .A2(KEYINPUT101), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n311), .B1(new_n660), .B2(KEYINPUT101), .ZN(new_n662));
  OAI21_X1  g476(.A(G472), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n305), .A2(new_n323), .A3(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n657), .A2(KEYINPUT40), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n428), .A2(new_n480), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  OR3_X1    g482(.A1(new_n658), .A2(new_n665), .A3(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(G143), .ZN(G45));
  AOI21_X1  g484(.A(new_n426), .B1(new_n425), .B2(new_n421), .ZN(new_n671));
  AOI211_X1 g485(.A(KEYINPUT20), .B(new_n422), .C1(new_n408), .C2(new_n424), .ZN(new_n672));
  OAI22_X1  g486(.A1(new_n671), .A2(new_n672), .B1(new_n409), .B2(new_n627), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n616), .A2(new_n617), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n673), .A2(new_n674), .A3(new_n648), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n606), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n324), .A2(new_n644), .A3(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G146), .ZN(G48));
  INV_X1    g492(.A(new_n576), .ZN(new_n679));
  INV_X1    g493(.A(new_n579), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n542), .B1(new_n681), .B2(new_n311), .ZN(new_n682));
  INV_X1    g496(.A(new_n580), .ZN(new_n683));
  NOR3_X1   g497(.A1(new_n682), .A2(new_n683), .A3(new_n541), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n685), .A2(new_n606), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n620), .A2(new_n380), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n324), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(KEYINPUT102), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT102), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n324), .A2(new_n690), .A3(new_n686), .A4(new_n687), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(KEYINPUT41), .B(G113), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(G15));
  NAND3_X1  g508(.A1(new_n324), .A2(new_n629), .A3(new_n686), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G116), .ZN(G18));
  NOR2_X1   g510(.A1(new_n643), .A2(new_n481), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n324), .A2(new_n686), .A3(new_n697), .ZN(new_n698));
  XOR2_X1   g512(.A(KEYINPUT103), .B(G119), .Z(new_n699));
  XNOR2_X1  g513(.A(new_n698), .B(new_n699), .ZN(G21));
  NAND2_X1  g514(.A1(new_n667), .A2(new_n625), .ZN(new_n701));
  NOR3_X1   g515(.A1(new_n701), .A2(new_n685), .A3(new_n436), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n314), .A2(new_n294), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n289), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(new_n300), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n592), .A2(new_n705), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n706), .A2(new_n380), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n702), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G122), .ZN(G24));
  NAND3_X1  g523(.A1(new_n638), .A2(new_n592), .A3(new_n705), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n711), .A2(new_n676), .A3(new_n684), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G125), .ZN(G27));
  NOR3_X1   g527(.A1(new_n538), .A2(new_n539), .A3(new_n483), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n586), .A2(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT42), .ZN(new_n716));
  NOR3_X1   g530(.A1(new_n675), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n318), .B1(new_n320), .B2(new_n299), .ZN(new_n718));
  NOR3_X1   g532(.A1(new_n320), .A2(new_n318), .A3(new_n299), .ZN(new_n719));
  OAI211_X1 g533(.A(new_n317), .B(new_n718), .C1(new_n719), .C2(KEYINPUT104), .ZN(new_n720));
  AND2_X1   g534(.A1(new_n719), .A2(KEYINPUT104), .ZN(new_n721));
  OAI211_X1 g535(.A(new_n717), .B(new_n381), .C1(new_n720), .C2(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(KEYINPUT105), .ZN(new_n723));
  INV_X1    g537(.A(new_n675), .ZN(new_n724));
  INV_X1    g538(.A(new_n715), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n324), .A2(new_n381), .A3(new_n724), .A4(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(new_n716), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n723), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G131), .ZN(G33));
  NOR2_X1   g543(.A1(new_n628), .A2(new_n649), .ZN(new_n730));
  AND4_X1   g544(.A1(new_n324), .A2(new_n381), .A3(new_n730), .A4(new_n725), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(new_n192), .ZN(G36));
  NOR3_X1   g546(.A1(new_n618), .A2(new_n673), .A3(KEYINPUT43), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n428), .A2(KEYINPUT107), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT107), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n673), .A2(new_n735), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n734), .A2(new_n674), .A3(new_n736), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n733), .B1(new_n737), .B2(KEYINPUT43), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n600), .A2(new_n638), .A3(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT44), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n600), .A2(KEYINPUT44), .A3(new_n638), .A4(new_n738), .ZN(new_n742));
  INV_X1    g556(.A(new_n541), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT45), .ZN(new_n744));
  AND2_X1   g558(.A1(new_n582), .A2(new_n578), .ZN(new_n745));
  AND2_X1   g559(.A1(new_n583), .A2(new_n559), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n744), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n584), .A2(KEYINPUT45), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n747), .A2(G469), .A3(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(new_n581), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n749), .A2(KEYINPUT46), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(new_n580), .ZN(new_n752));
  AOI21_X1  g566(.A(KEYINPUT46), .B1(new_n749), .B2(new_n750), .ZN(new_n753));
  OAI211_X1 g567(.A(new_n743), .B(new_n656), .C1(new_n752), .C2(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT106), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n754), .B(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(new_n714), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n741), .A2(new_n742), .A3(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G137), .ZN(G39));
  OAI21_X1  g574(.A(new_n743), .B1(new_n752), .B2(new_n753), .ZN(new_n761));
  AND2_X1   g575(.A1(new_n761), .A2(KEYINPUT47), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT47), .ZN(new_n763));
  OAI211_X1 g577(.A(new_n763), .B(new_n743), .C1(new_n752), .C2(new_n753), .ZN(new_n764));
  INV_X1    g578(.A(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n724), .A2(new_n380), .A3(new_n714), .ZN(new_n766));
  OR4_X1    g580(.A1(new_n324), .A2(new_n762), .A3(new_n765), .A4(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G140), .ZN(G42));
  NAND2_X1  g582(.A1(new_n737), .A2(KEYINPUT43), .ZN(new_n769));
  INV_X1    g583(.A(new_n733), .ZN(new_n770));
  AND3_X1   g584(.A1(new_n684), .A2(new_n430), .A3(new_n714), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n769), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n772), .A2(new_n710), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT113), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT51), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n773), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n673), .A2(new_n674), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n665), .A2(new_n381), .A3(new_n771), .A4(new_n777), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n682), .A2(new_n683), .ZN(new_n779));
  OR2_X1    g593(.A1(new_n779), .A2(KEYINPUT112), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(KEYINPUT112), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n780), .A2(new_n541), .A3(new_n781), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n782), .B1(new_n762), .B2(new_n765), .ZN(new_n783));
  NOR3_X1   g597(.A1(new_n706), .A2(new_n380), .A3(new_n647), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n783), .A2(new_n714), .A3(new_n738), .A4(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n776), .A2(new_n778), .A3(new_n785), .ZN(new_n786));
  AND2_X1   g600(.A1(new_n653), .A2(new_n483), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n784), .A2(new_n738), .A3(new_n684), .A4(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(KEYINPUT50), .ZN(new_n789));
  OAI22_X1  g603(.A1(new_n786), .A2(new_n789), .B1(new_n774), .B2(new_n775), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n776), .A2(new_n785), .ZN(new_n791));
  INV_X1    g605(.A(new_n789), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n774), .A2(new_n775), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n791), .A2(new_n792), .A3(new_n793), .A4(new_n778), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n381), .B1(new_n720), .B2(new_n721), .ZN(new_n795));
  OR3_X1    g609(.A1(new_n772), .A2(new_n795), .A3(KEYINPUT48), .ZN(new_n796));
  OAI21_X1  g610(.A(KEYINPUT48), .B1(new_n772), .B2(new_n795), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n665), .A2(new_n381), .A3(new_n619), .A4(new_n771), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n784), .A2(new_n738), .A3(new_n625), .A4(new_n684), .ZN(new_n800));
  AND3_X1   g614(.A1(new_n800), .A2(G952), .A3(new_n266), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n798), .A2(new_n799), .A3(new_n801), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n802), .A2(KEYINPUT114), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n802), .A2(KEYINPUT114), .ZN(new_n804));
  OAI211_X1 g618(.A(new_n790), .B(new_n794), .C1(new_n803), .C2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT115), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n805), .B(new_n806), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n695), .A2(new_n698), .A3(new_n708), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n808), .B1(new_n691), .B2(new_n689), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n731), .B1(new_n723), .B2(new_n727), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n605), .A2(new_n437), .A3(new_n482), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT109), .ZN(new_n812));
  AOI22_X1  g626(.A1(new_n628), .A2(new_n812), .B1(new_n673), .B2(new_n674), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n428), .A2(KEYINPUT109), .A3(new_n479), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n811), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n633), .A2(new_n815), .A3(new_n381), .A4(new_n586), .ZN(new_n816));
  AND3_X1   g630(.A1(new_n816), .A2(new_n589), .A3(new_n639), .ZN(new_n817));
  NOR4_X1   g631(.A1(new_n757), .A2(new_n673), .A3(new_n479), .A4(new_n649), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n324), .A2(new_n644), .A3(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n711), .A2(new_n724), .A3(new_n725), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n809), .A2(new_n810), .A3(new_n817), .A4(new_n821), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n638), .A2(new_n587), .A3(new_n649), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n664), .A2(new_n625), .A3(new_n667), .A4(new_n823), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n824), .A2(new_n651), .A3(new_n677), .A4(new_n712), .ZN(new_n825));
  XNOR2_X1  g639(.A(new_n825), .B(KEYINPUT52), .ZN(new_n826));
  OAI21_X1  g640(.A(KEYINPUT53), .B1(new_n822), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n810), .A2(new_n821), .ZN(new_n828));
  AND3_X1   g642(.A1(new_n695), .A2(new_n698), .A3(new_n708), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n817), .A2(new_n692), .A3(new_n829), .ZN(new_n830));
  OR3_X1    g644(.A1(new_n828), .A2(KEYINPUT53), .A3(new_n830), .ZN(new_n831));
  AND3_X1   g645(.A1(new_n651), .A2(new_n677), .A3(new_n712), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n832), .A2(KEYINPUT52), .A3(new_n824), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT52), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n825), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n833), .A2(KEYINPUT110), .A3(new_n835), .ZN(new_n836));
  OR3_X1    g650(.A1(new_n825), .A2(KEYINPUT110), .A3(new_n834), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  OAI211_X1 g652(.A(new_n827), .B(KEYINPUT54), .C1(new_n831), .C2(new_n838), .ZN(new_n839));
  AND3_X1   g653(.A1(new_n692), .A2(new_n829), .A3(KEYINPUT111), .ZN(new_n840));
  AOI21_X1  g654(.A(KEYINPUT111), .B1(new_n692), .B2(new_n829), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT53), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n731), .A2(new_n843), .ZN(new_n844));
  AND4_X1   g658(.A1(new_n728), .A2(new_n817), .A3(new_n821), .A4(new_n844), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n842), .A2(new_n837), .A3(new_n836), .A4(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT54), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n843), .B1(new_n822), .B2(new_n826), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n846), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n839), .A2(new_n849), .ZN(new_n850));
  OAI22_X1  g664(.A1(new_n807), .A2(new_n850), .B1(G952), .B2(G953), .ZN(new_n851));
  XNOR2_X1  g665(.A(new_n779), .B(KEYINPUT49), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n852), .A2(new_n482), .A3(new_n743), .A4(new_n653), .ZN(new_n853));
  NOR4_X1   g667(.A1(new_n853), .A2(new_n664), .A3(new_n380), .A4(new_n737), .ZN(new_n854));
  XNOR2_X1  g668(.A(new_n854), .B(KEYINPUT108), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n851), .A2(new_n855), .ZN(G75));
  NAND2_X1  g670(.A1(new_n846), .A2(new_n848), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n857), .A2(G210), .A3(G902), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT56), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n514), .A2(new_n516), .ZN(new_n860));
  XNOR2_X1  g674(.A(new_n860), .B(KEYINPUT116), .ZN(new_n861));
  XNOR2_X1  g675(.A(new_n522), .B(KEYINPUT55), .ZN(new_n862));
  XNOR2_X1  g676(.A(new_n861), .B(new_n862), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n858), .A2(new_n859), .A3(new_n863), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n863), .B1(new_n858), .B2(new_n859), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n266), .A2(G952), .ZN(new_n866));
  XOR2_X1   g680(.A(new_n866), .B(KEYINPUT117), .Z(new_n867));
  NOR3_X1   g681(.A1(new_n864), .A2(new_n865), .A3(new_n867), .ZN(G51));
  XNOR2_X1  g682(.A(new_n581), .B(KEYINPUT57), .ZN(new_n869));
  AND3_X1   g683(.A1(new_n846), .A2(new_n847), .A3(new_n848), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n847), .B1(new_n846), .B2(new_n848), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n869), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n872), .A2(new_n681), .ZN(new_n873));
  XNOR2_X1  g687(.A(new_n749), .B(KEYINPUT118), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n857), .A2(G902), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n866), .B1(new_n873), .B2(new_n875), .ZN(G54));
  NAND4_X1  g690(.A1(new_n857), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n877));
  AND2_X1   g691(.A1(new_n877), .A2(new_n420), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n877), .A2(new_n420), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n878), .A2(new_n879), .A3(new_n866), .ZN(G60));
  NAND2_X1  g694(.A1(G478), .A2(G902), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n881), .B(KEYINPUT59), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n615), .B1(new_n850), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n615), .A2(new_n882), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n857), .A2(KEYINPUT54), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n884), .B1(new_n885), .B2(new_n849), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n883), .A2(new_n886), .A3(new_n867), .ZN(G63));
  INV_X1    g701(.A(KEYINPUT61), .ZN(new_n888));
  XNOR2_X1  g702(.A(KEYINPUT119), .B(KEYINPUT60), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n367), .A2(new_n311), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n889), .B(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n857), .A2(new_n636), .A3(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(new_n867), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n366), .B(KEYINPUT120), .ZN(new_n895));
  INV_X1    g709(.A(new_n895), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n896), .B1(new_n857), .B2(new_n891), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n888), .B1(new_n894), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n857), .A2(new_n891), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n899), .A2(new_n895), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n900), .A2(KEYINPUT61), .A3(new_n893), .A4(new_n892), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n898), .A2(new_n901), .ZN(G66));
  AOI21_X1  g716(.A(new_n266), .B1(new_n434), .B2(new_n520), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n903), .B1(new_n830), .B2(new_n266), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n861), .B1(G898), .B2(new_n266), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n904), .B(new_n905), .Z(G69));
  NOR2_X1   g720(.A1(new_n274), .A2(new_n280), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n907), .B(new_n414), .ZN(new_n908));
  NAND2_X1  g722(.A1(G900), .A2(G953), .ZN(new_n909));
  OR3_X1    g723(.A1(new_n756), .A2(new_n701), .A3(new_n795), .ZN(new_n910));
  AND3_X1   g724(.A1(new_n759), .A2(new_n767), .A3(new_n910), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n651), .A2(new_n677), .A3(new_n712), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(KEYINPUT121), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT121), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n832), .A2(new_n914), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n911), .A2(new_n810), .A3(new_n913), .A4(new_n915), .ZN(new_n916));
  OAI211_X1 g730(.A(new_n908), .B(new_n909), .C1(new_n916), .C2(G953), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n915), .A2(new_n669), .A3(new_n913), .ZN(new_n918));
  NAND2_X1  g732(.A1(KEYINPUT122), .A2(KEYINPUT62), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n918), .B(new_n919), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n767), .B1(KEYINPUT122), .B2(KEYINPUT62), .ZN(new_n921));
  AND2_X1   g735(.A1(new_n324), .A2(new_n381), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n655), .B1(new_n813), .B2(new_n814), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n922), .A2(new_n725), .A3(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT123), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND4_X1  g740(.A1(new_n922), .A2(KEYINPUT123), .A3(new_n725), .A4(new_n923), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n759), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(KEYINPUT124), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT124), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n759), .A2(new_n926), .A3(new_n930), .A4(new_n927), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n921), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  AOI21_X1  g746(.A(G953), .B1(new_n920), .B2(new_n932), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n917), .B1(new_n933), .B2(new_n908), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n266), .B1(G227), .B2(G900), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n935), .B1(new_n917), .B2(KEYINPUT125), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  OAI221_X1 g751(.A(new_n917), .B1(KEYINPUT125), .B2(new_n935), .C1(new_n933), .C2(new_n908), .ZN(new_n938));
  AND2_X1   g752(.A1(new_n937), .A2(new_n938), .ZN(G72));
  NAND2_X1  g753(.A1(G472), .A2(G902), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n940), .B(KEYINPUT63), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n941), .B(KEYINPUT126), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n942), .B1(new_n916), .B2(new_n830), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n306), .A2(new_n271), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n866), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n308), .B1(new_n283), .B2(new_n285), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n946), .A2(new_n941), .ZN(new_n947));
  OAI211_X1 g761(.A(new_n827), .B(new_n947), .C1(new_n831), .C2(new_n838), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n945), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n920), .A2(new_n932), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n942), .B1(new_n950), .B2(new_n830), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n307), .A2(new_n294), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n949), .B1(new_n951), .B2(new_n952), .ZN(G57));
endmodule


