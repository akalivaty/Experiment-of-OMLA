//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 1 0 0 1 0 1 1 0 1 0 0 1 0 1 0 1 0 0 0 0 1 1 1 1 1 0 1 0 0 1 0 0 1 0 0 0 0 0 1 1 1 1 0 0 1 1 1 0 1 1 0 0 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:47 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n438, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n578, new_n579, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n594, new_n595,
    new_n597, new_n598, new_n599, new_n600, new_n601, new_n602, new_n603,
    new_n605, new_n606, new_n607, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n640, new_n642, new_n643, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n856, new_n857,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1225;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  OR2_X1    g011(.A1(new_n436), .A2(KEYINPUT64), .ZN(new_n437));
  NAND2_X1  g012(.A1(new_n436), .A2(KEYINPUT64), .ZN(new_n438));
  NAND2_X1  g013(.A1(new_n437), .A2(new_n438), .ZN(G220));
  XOR2_X1   g014(.A(KEYINPUT65), .B(G96), .Z(G221));
  XNOR2_X1  g015(.A(KEYINPUT66), .B(G69), .ZN(G235));
  INV_X1    g016(.A(G120), .ZN(G236));
  INV_X1    g017(.A(G57), .ZN(G237));
  INV_X1    g018(.A(G108), .ZN(G238));
  NAND4_X1  g019(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT67), .Z(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR3_X1   g030(.A1(G221), .A2(G218), .A3(G219), .ZN(new_n456));
  NAND3_X1  g031(.A1(new_n456), .A2(new_n438), .A3(new_n437), .ZN(new_n457));
  XNOR2_X1  g032(.A(new_n457), .B(KEYINPUT2), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n455), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  NAND2_X1  g035(.A1(new_n455), .A2(G567), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n458), .A2(G2106), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT68), .ZN(new_n463));
  OAI21_X1  g038(.A(new_n461), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n464), .B1(new_n463), .B2(new_n462), .ZN(new_n465));
  XNOR2_X1  g040(.A(new_n465), .B(KEYINPUT69), .ZN(G319));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT72), .ZN(new_n469));
  AND3_X1   g044(.A1(new_n468), .A2(new_n469), .A3(G101), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n469), .B1(new_n468), .B2(G101), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n472), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(G137), .ZN(new_n477));
  OAI22_X1  g052(.A1(new_n470), .A2(new_n471), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  OAI21_X1  g053(.A(KEYINPUT70), .B1(new_n474), .B2(new_n475), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT3), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(new_n467), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT70), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n481), .A2(new_n482), .A3(new_n473), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n479), .A2(G125), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(KEYINPUT71), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT71), .ZN(new_n486));
  NAND4_X1  g061(.A1(new_n479), .A2(new_n483), .A3(new_n486), .A4(G125), .ZN(new_n487));
  NAND2_X1  g062(.A1(G113), .A2(G2104), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n485), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n478), .B1(new_n489), .B2(G2105), .ZN(G160));
  INV_X1    g065(.A(new_n476), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G136), .ZN(new_n492));
  XOR2_X1   g067(.A(new_n492), .B(KEYINPUT73), .Z(new_n493));
  OAI21_X1  g068(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(G112), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n494), .B1(new_n495), .B2(G2105), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n472), .B1(new_n481), .B2(new_n473), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n496), .B1(new_n497), .B2(G124), .ZN(new_n498));
  AND2_X1   g073(.A1(new_n493), .A2(new_n498), .ZN(G162));
  INV_X1    g074(.A(KEYINPUT74), .ZN(new_n500));
  OAI21_X1  g075(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n501));
  INV_X1    g076(.A(G114), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n501), .B1(new_n502), .B2(G2105), .ZN(new_n503));
  NAND2_X1  g078(.A1(G126), .A2(G2105), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n504), .B1(new_n481), .B2(new_n473), .ZN(new_n505));
  OAI21_X1  g080(.A(new_n500), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  OAI211_X1 g081(.A(G126), .B(G2105), .C1(new_n474), .C2(new_n475), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n502), .A2(G2105), .ZN(new_n508));
  OAI211_X1 g083(.A(new_n508), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n507), .A2(new_n509), .A3(KEYINPUT74), .ZN(new_n510));
  INV_X1    g085(.A(G138), .ZN(new_n511));
  OAI21_X1  g086(.A(KEYINPUT4), .B1(new_n476), .B2(new_n511), .ZN(new_n512));
  NOR3_X1   g087(.A1(new_n511), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n479), .A2(new_n483), .A3(new_n513), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n506), .A2(new_n510), .B1(new_n512), .B2(new_n514), .ZN(G164));
  XNOR2_X1  g090(.A(KEYINPUT6), .B(G651), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT5), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G543), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT75), .ZN(new_n519));
  INV_X1    g094(.A(G543), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n519), .B1(KEYINPUT5), .B2(new_n520), .ZN(new_n521));
  NOR3_X1   g096(.A1(new_n517), .A2(KEYINPUT75), .A3(G543), .ZN(new_n522));
  OAI211_X1 g097(.A(new_n516), .B(new_n518), .C1(new_n521), .C2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT76), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  OAI21_X1  g100(.A(KEYINPUT75), .B1(new_n517), .B2(G543), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n519), .A2(new_n520), .A3(KEYINPUT5), .ZN(new_n527));
  AOI22_X1  g102(.A1(new_n526), .A2(new_n527), .B1(new_n517), .B2(G543), .ZN(new_n528));
  AOI21_X1  g103(.A(KEYINPUT76), .B1(new_n528), .B2(new_n516), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n525), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(G88), .ZN(new_n531));
  NAND2_X1  g106(.A1(G75), .A2(G543), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n518), .B1(new_n521), .B2(new_n522), .ZN(new_n533));
  INV_X1    g108(.A(G62), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  AND2_X1   g110(.A1(KEYINPUT6), .A2(G651), .ZN(new_n536));
  NOR2_X1   g111(.A1(KEYINPUT6), .A2(G651), .ZN(new_n537));
  OAI21_X1  g112(.A(G543), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(new_n538), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n535), .A2(G651), .B1(G50), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n531), .A2(new_n540), .ZN(G303));
  INV_X1    g116(.A(G303), .ZN(G166));
  NAND2_X1  g117(.A1(new_n523), .A2(new_n524), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n528), .A2(KEYINPUT76), .A3(new_n516), .ZN(new_n544));
  AND3_X1   g119(.A1(new_n543), .A2(G89), .A3(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(KEYINPUT77), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n538), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n516), .A2(KEYINPUT77), .A3(G543), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G51), .ZN(new_n550));
  AND2_X1   g125(.A1(G63), .A2(G651), .ZN(new_n551));
  OAI211_X1 g126(.A(new_n518), .B(new_n551), .C1(new_n521), .C2(new_n522), .ZN(new_n552));
  NAND3_X1  g127(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT7), .ZN(new_n554));
  AND2_X1   g129(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n550), .A2(new_n555), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n545), .A2(new_n556), .ZN(G168));
  AOI22_X1  g132(.A1(new_n528), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n558));
  INV_X1    g133(.A(G651), .ZN(new_n559));
  OR2_X1    g134(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n543), .A2(G90), .A3(new_n544), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT79), .ZN(new_n562));
  XOR2_X1   g137(.A(KEYINPUT78), .B(G52), .Z(new_n563));
  NAND2_X1  g138(.A1(new_n549), .A2(new_n563), .ZN(new_n564));
  AND3_X1   g139(.A1(new_n561), .A2(new_n562), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n562), .B1(new_n561), .B2(new_n564), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n560), .B1(new_n565), .B2(new_n566), .ZN(G301));
  INV_X1    g142(.A(G301), .ZN(G171));
  NAND2_X1  g143(.A1(G68), .A2(G543), .ZN(new_n569));
  INV_X1    g144(.A(G56), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n569), .B1(new_n533), .B2(new_n570), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n571), .A2(G651), .B1(new_n549), .B2(G43), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n543), .A2(G81), .A3(new_n544), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(G860), .ZN(G153));
  NAND4_X1  g151(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g152(.A1(G1), .A2(G3), .ZN(new_n578));
  XNOR2_X1  g153(.A(new_n578), .B(KEYINPUT8), .ZN(new_n579));
  NAND4_X1  g154(.A1(G319), .A2(G483), .A3(G661), .A4(new_n579), .ZN(G188));
  NAND3_X1  g155(.A1(new_n516), .A2(G53), .A3(G543), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT9), .ZN(new_n582));
  XNOR2_X1  g157(.A(new_n581), .B(new_n582), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n528), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT81), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n559), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(G78), .A2(G543), .ZN(new_n587));
  INV_X1    g162(.A(G65), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n533), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n589), .A2(KEYINPUT81), .ZN(new_n590));
  AOI21_X1  g165(.A(new_n583), .B1(new_n586), .B2(new_n590), .ZN(new_n591));
  OAI21_X1  g166(.A(KEYINPUT80), .B1(new_n525), .B2(new_n529), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT80), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n543), .A2(new_n593), .A3(new_n544), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n592), .A2(G91), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n591), .A2(new_n595), .ZN(G299));
  INV_X1    g171(.A(G51), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n597), .B1(new_n547), .B2(new_n548), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n552), .A2(new_n554), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n543), .A2(G89), .A3(new_n544), .ZN(new_n601));
  AND3_X1   g176(.A1(new_n600), .A2(new_n601), .A3(KEYINPUT82), .ZN(new_n602));
  AOI21_X1  g177(.A(KEYINPUT82), .B1(new_n600), .B2(new_n601), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n602), .A2(new_n603), .ZN(G286));
  NAND3_X1  g179(.A1(new_n592), .A2(G87), .A3(new_n594), .ZN(new_n605));
  OR2_X1    g180(.A1(new_n528), .A2(G74), .ZN(new_n606));
  AOI22_X1  g181(.A1(new_n606), .A2(G651), .B1(G49), .B2(new_n539), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n605), .A2(new_n607), .ZN(G288));
  NAND3_X1  g183(.A1(new_n592), .A2(G86), .A3(new_n594), .ZN(new_n609));
  NAND2_X1  g184(.A1(G73), .A2(G543), .ZN(new_n610));
  INV_X1    g185(.A(G61), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n533), .B2(new_n611), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n612), .A2(G651), .B1(G48), .B2(new_n539), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n609), .A2(new_n613), .ZN(G305));
  AOI22_X1  g189(.A1(new_n530), .A2(G85), .B1(G47), .B2(new_n549), .ZN(new_n615));
  AND2_X1   g190(.A1(G72), .A2(G543), .ZN(new_n616));
  AOI21_X1  g191(.A(new_n616), .B1(new_n528), .B2(G60), .ZN(new_n617));
  INV_X1    g192(.A(KEYINPUT83), .ZN(new_n618));
  AND2_X1   g193(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  OAI21_X1  g194(.A(G651), .B1(new_n617), .B2(new_n618), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n615), .B1(new_n619), .B2(new_n620), .ZN(G290));
  NAND2_X1  g196(.A1(G301), .A2(G868), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n549), .A2(G54), .ZN(new_n623));
  NAND2_X1  g198(.A1(G79), .A2(G543), .ZN(new_n624));
  INV_X1    g199(.A(G66), .ZN(new_n625));
  OAI211_X1 g200(.A(KEYINPUT84), .B(new_n624), .C1(new_n533), .C2(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n626), .A2(G651), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n528), .A2(G66), .ZN(new_n628));
  AOI21_X1  g203(.A(KEYINPUT84), .B1(new_n628), .B2(new_n624), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n623), .B1(new_n627), .B2(new_n629), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n592), .A2(G92), .A3(new_n594), .ZN(new_n631));
  INV_X1    g206(.A(KEYINPUT10), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND4_X1  g208(.A1(new_n592), .A2(KEYINPUT10), .A3(G92), .A4(new_n594), .ZN(new_n634));
  AOI21_X1  g209(.A(new_n630), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n622), .B1(new_n635), .B2(G868), .ZN(G284));
  OAI21_X1  g211(.A(new_n622), .B1(new_n635), .B2(G868), .ZN(G321));
  MUX2_X1   g212(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g213(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g214(.A(G559), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n635), .B1(new_n640), .B2(G860), .ZN(G148));
  NAND2_X1  g216(.A1(new_n635), .A2(new_n640), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n642), .A2(G868), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n643), .B1(G868), .B2(new_n575), .ZN(G323));
  XNOR2_X1  g219(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g220(.A1(new_n479), .A2(new_n483), .A3(new_n468), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT12), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT13), .ZN(new_n648));
  INV_X1    g223(.A(G2100), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n648), .A2(new_n649), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n497), .A2(G123), .ZN(new_n652));
  INV_X1    g227(.A(G135), .ZN(new_n653));
  NOR2_X1   g228(.A1(new_n472), .A2(G111), .ZN(new_n654));
  OAI21_X1  g229(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n655));
  OAI221_X1 g230(.A(new_n652), .B1(new_n653), .B2(new_n476), .C1(new_n654), .C2(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n656), .B(G2096), .Z(new_n657));
  NAND3_X1  g232(.A1(new_n650), .A2(new_n651), .A3(new_n657), .ZN(G156));
  XNOR2_X1  g233(.A(KEYINPUT15), .B(G2435), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(G2438), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2427), .B(G2430), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n662), .A2(KEYINPUT14), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT86), .ZN(new_n664));
  OAI21_X1  g239(.A(new_n664), .B1(new_n660), .B2(new_n661), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1341), .B(G1348), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n665), .B(new_n666), .Z(new_n667));
  XOR2_X1   g242(.A(G2451), .B(G2454), .Z(new_n668));
  XNOR2_X1  g243(.A(KEYINPUT85), .B(KEYINPUT16), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  OR2_X1    g245(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n667), .A2(new_n670), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G2443), .B(G2446), .ZN(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n671), .A2(new_n674), .A3(new_n672), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n676), .A2(new_n677), .A3(G14), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT87), .ZN(G401));
  XOR2_X1   g254(.A(G2072), .B(G2078), .Z(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(G2084), .B(G2090), .Z(new_n682));
  XNOR2_X1  g257(.A(G2067), .B(G2678), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n681), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(new_n684), .B(KEYINPUT18), .Z(new_n685));
  XOR2_X1   g260(.A(KEYINPUT89), .B(KEYINPUT17), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n680), .B(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(new_n682), .ZN(new_n688));
  OR3_X1    g263(.A1(new_n687), .A2(new_n688), .A3(new_n683), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n687), .A2(new_n683), .ZN(new_n690));
  INV_X1    g265(.A(KEYINPUT88), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n688), .B1(new_n681), .B2(new_n683), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n690), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(new_n692), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n694), .A2(KEYINPUT88), .ZN(new_n695));
  OAI211_X1 g270(.A(new_n685), .B(new_n689), .C1(new_n693), .C2(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(G2096), .B(G2100), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(G227));
  XNOR2_X1  g274(.A(G1971), .B(G1976), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT19), .ZN(new_n701));
  XNOR2_X1  g276(.A(G1956), .B(G2474), .ZN(new_n702));
  XNOR2_X1  g277(.A(G1961), .B(G1966), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n701), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n702), .A2(new_n703), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n701), .A2(KEYINPUT92), .ZN(new_n708));
  XOR2_X1   g283(.A(new_n707), .B(new_n708), .Z(new_n709));
  NOR3_X1   g284(.A1(new_n701), .A2(new_n702), .A3(new_n703), .ZN(new_n710));
  XOR2_X1   g285(.A(KEYINPUT90), .B(KEYINPUT20), .Z(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT91), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n710), .B(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n709), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  XOR2_X1   g291(.A(G1991), .B(G1996), .Z(new_n717));
  INV_X1    g292(.A(new_n717), .ZN(new_n718));
  OR2_X1    g293(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n716), .A2(new_n718), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g296(.A(G1981), .B(G1986), .ZN(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g299(.A1(new_n719), .A2(new_n722), .A3(new_n720), .ZN(new_n725));
  AND2_X1   g300(.A1(new_n724), .A2(new_n725), .ZN(G229));
  INV_X1    g301(.A(G16), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n727), .A2(G5), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(G171), .B2(new_n727), .ZN(new_n729));
  INV_X1    g304(.A(KEYINPUT100), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n729), .B(new_n730), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n731), .A2(G1961), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n731), .A2(G1961), .ZN(new_n733));
  INV_X1    g308(.A(G29), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(G33), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n472), .A2(G103), .A3(G2104), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(KEYINPUT25), .Z(new_n737));
  INV_X1    g312(.A(KEYINPUT98), .ZN(new_n738));
  AND3_X1   g313(.A1(new_n491), .A2(new_n738), .A3(G139), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n738), .B1(new_n491), .B2(G139), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n737), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n479), .A2(G127), .A3(new_n483), .ZN(new_n742));
  INV_X1    g317(.A(G115), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n742), .B1(new_n743), .B2(new_n467), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n741), .B1(G2105), .B2(new_n744), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n735), .B1(new_n745), .B2(new_n734), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(G2072), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n727), .A2(G21), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G168), .B2(new_n727), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(G1966), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n734), .A2(G27), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT101), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(G164), .B2(new_n734), .ZN(new_n753));
  INV_X1    g328(.A(G2078), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT30), .B(G28), .ZN(new_n756));
  OR2_X1    g331(.A1(KEYINPUT31), .A2(G11), .ZN(new_n757));
  NAND2_X1  g332(.A1(KEYINPUT31), .A2(G11), .ZN(new_n758));
  AOI22_X1  g333(.A1(new_n756), .A2(new_n734), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(new_n656), .B2(new_n734), .ZN(new_n760));
  AND2_X1   g335(.A1(new_n734), .A2(G32), .ZN(new_n761));
  NAND3_X1  g336(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT26), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(new_n497), .B2(G129), .ZN(new_n764));
  AOI22_X1  g339(.A1(new_n491), .A2(G141), .B1(G105), .B2(new_n468), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n761), .B1(new_n766), .B2(G29), .ZN(new_n767));
  XNOR2_X1  g342(.A(KEYINPUT27), .B(G1996), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n760), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  OAI211_X1 g344(.A(new_n755), .B(new_n769), .C1(new_n767), .C2(new_n768), .ZN(new_n770));
  XNOR2_X1  g345(.A(KEYINPUT99), .B(KEYINPUT24), .ZN(new_n771));
  INV_X1    g346(.A(new_n771), .ZN(new_n772));
  AOI21_X1  g347(.A(G29), .B1(new_n772), .B2(G34), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G34), .B2(new_n772), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(G160), .B2(new_n734), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(G2084), .ZN(new_n776));
  NOR4_X1   g351(.A1(new_n747), .A2(new_n750), .A3(new_n770), .A4(new_n776), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n732), .A2(new_n733), .A3(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(KEYINPUT102), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND4_X1  g355(.A1(new_n732), .A2(new_n777), .A3(KEYINPUT102), .A4(new_n733), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n727), .A2(G4), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(new_n635), .B2(new_n727), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n783), .A2(G1348), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n734), .A2(G35), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(G162), .B2(new_n734), .ZN(new_n786));
  XNOR2_X1  g361(.A(KEYINPUT29), .B(G2090), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  XOR2_X1   g363(.A(KEYINPUT95), .B(G16), .Z(new_n789));
  INV_X1    g364(.A(new_n789), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n790), .A2(G19), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(new_n575), .B2(new_n790), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(G1341), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n497), .A2(G128), .ZN(new_n794));
  INV_X1    g369(.A(G140), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n472), .A2(G116), .ZN(new_n796));
  OAI21_X1  g371(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n797));
  OAI221_X1 g372(.A(new_n794), .B1(new_n795), .B2(new_n476), .C1(new_n796), .C2(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n798), .A2(G29), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n734), .A2(G26), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT28), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(G2067), .ZN(new_n803));
  NOR3_X1   g378(.A1(new_n788), .A2(new_n793), .A3(new_n803), .ZN(new_n804));
  OR2_X1    g379(.A1(new_n783), .A2(G1348), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n789), .A2(G20), .ZN(new_n806));
  XNOR2_X1  g381(.A(KEYINPUT103), .B(KEYINPUT23), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n808), .B1(G299), .B2(G16), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(G1956), .ZN(new_n810));
  AND4_X1   g385(.A1(new_n784), .A2(new_n804), .A3(new_n805), .A4(new_n810), .ZN(new_n811));
  NAND3_X1  g386(.A1(new_n780), .A2(new_n781), .A3(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n812), .A2(KEYINPUT104), .ZN(new_n813));
  INV_X1    g388(.A(KEYINPUT104), .ZN(new_n814));
  NAND4_X1  g389(.A1(new_n780), .A2(new_n814), .A3(new_n781), .A4(new_n811), .ZN(new_n815));
  MUX2_X1   g390(.A(G6), .B(G305), .S(G16), .Z(new_n816));
  XOR2_X1   g391(.A(KEYINPUT32), .B(G1981), .Z(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  AND2_X1   g393(.A1(new_n605), .A2(new_n607), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n819), .A2(new_n727), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n820), .B1(new_n727), .B2(G23), .ZN(new_n821));
  XNOR2_X1  g396(.A(KEYINPUT33), .B(G1976), .ZN(new_n822));
  OR2_X1    g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n821), .A2(new_n822), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n790), .A2(G22), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n825), .B1(G166), .B2(new_n790), .ZN(new_n826));
  XNOR2_X1  g401(.A(KEYINPUT97), .B(G1971), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n826), .B(new_n827), .ZN(new_n828));
  AND4_X1   g403(.A1(new_n818), .A2(new_n823), .A3(new_n824), .A4(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(KEYINPUT96), .B(KEYINPUT34), .ZN(new_n830));
  OR2_X1    g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n829), .A2(new_n830), .ZN(new_n832));
  MUX2_X1   g407(.A(G24), .B(G290), .S(new_n790), .Z(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(G1986), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n734), .A2(G25), .ZN(new_n835));
  OAI21_X1  g410(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n836));
  INV_X1    g411(.A(new_n836), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n837), .B1(G107), .B2(new_n472), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT93), .ZN(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n497), .A2(G119), .ZN(new_n841));
  INV_X1    g416(.A(G131), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n841), .B1(new_n842), .B2(new_n476), .ZN(new_n843));
  OR2_X1    g418(.A1(new_n840), .A2(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(new_n844), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n835), .B1(new_n845), .B2(new_n734), .ZN(new_n846));
  XNOR2_X1  g421(.A(KEYINPUT35), .B(G1991), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT94), .ZN(new_n848));
  XOR2_X1   g423(.A(new_n846), .B(new_n848), .Z(new_n849));
  NOR2_X1   g424(.A1(new_n834), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n831), .A2(new_n832), .A3(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n851), .A2(KEYINPUT36), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT36), .ZN(new_n853));
  NAND4_X1  g428(.A1(new_n831), .A2(new_n853), .A3(new_n832), .A4(new_n850), .ZN(new_n854));
  AOI22_X1  g429(.A1(new_n813), .A2(new_n815), .B1(new_n852), .B2(new_n854), .ZN(G311));
  NAND2_X1  g430(.A1(new_n813), .A2(new_n815), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n852), .A2(new_n854), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(new_n857), .ZN(G150));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n859));
  INV_X1    g434(.A(new_n630), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n861), .A2(new_n640), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT105), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n862), .B(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n864), .A2(KEYINPUT38), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n862), .B(KEYINPUT105), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT38), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(G80), .A2(G543), .ZN(new_n869));
  INV_X1    g444(.A(G67), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n869), .B1(new_n533), .B2(new_n870), .ZN(new_n871));
  AOI22_X1  g446(.A1(new_n871), .A2(G651), .B1(new_n549), .B2(G55), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n543), .A2(G93), .A3(new_n544), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n574), .A2(new_n874), .ZN(new_n875));
  AOI22_X1  g450(.A1(new_n573), .A2(new_n572), .B1(new_n872), .B2(new_n873), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  AND3_X1   g452(.A1(new_n865), .A2(new_n868), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n877), .B1(new_n865), .B2(new_n868), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT39), .ZN(new_n881));
  AOI21_X1  g456(.A(G860), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  OR2_X1    g457(.A1(new_n875), .A2(new_n876), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n866), .A2(new_n867), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n864), .A2(KEYINPUT38), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n883), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n865), .A2(new_n868), .A3(new_n877), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g463(.A(KEYINPUT106), .B1(new_n888), .B2(KEYINPUT39), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT106), .ZN(new_n890));
  AOI211_X1 g465(.A(new_n890), .B(new_n881), .C1(new_n886), .C2(new_n887), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n882), .B1(new_n889), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n874), .A2(G860), .ZN(new_n893));
  XOR2_X1   g468(.A(new_n893), .B(KEYINPUT37), .Z(new_n894));
  NAND2_X1  g469(.A1(new_n892), .A2(new_n894), .ZN(G145));
  XNOR2_X1  g470(.A(new_n844), .B(new_n647), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n491), .A2(G142), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT107), .ZN(new_n898));
  OR3_X1    g473(.A1(new_n898), .A2(new_n472), .A3(G118), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n898), .B1(new_n472), .B2(G118), .ZN(new_n900));
  OR2_X1    g475(.A1(G106), .A2(G2105), .ZN(new_n901));
  NAND4_X1  g476(.A1(new_n899), .A2(G2104), .A3(new_n900), .A4(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n497), .A2(G130), .ZN(new_n903));
  AND3_X1   g478(.A1(new_n897), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  XOR2_X1   g479(.A(new_n896), .B(new_n904), .Z(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n766), .B(new_n798), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n507), .A2(new_n509), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n908), .B1(new_n512), .B2(new_n514), .ZN(new_n909));
  XOR2_X1   g484(.A(new_n907), .B(new_n909), .Z(new_n910));
  OR2_X1    g485(.A1(new_n910), .A2(new_n745), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n745), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT108), .ZN(new_n914));
  NOR3_X1   g489(.A1(new_n906), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  XNOR2_X1  g490(.A(G160), .B(new_n656), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n916), .B(G162), .ZN(new_n917));
  AND2_X1   g492(.A1(new_n917), .A2(KEYINPUT109), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n917), .A2(KEYINPUT109), .ZN(new_n919));
  AOI22_X1  g494(.A1(new_n905), .A2(KEYINPUT108), .B1(new_n911), .B2(new_n912), .ZN(new_n920));
  NOR4_X1   g495(.A1(new_n915), .A2(new_n918), .A3(new_n919), .A4(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n906), .A2(new_n912), .A3(new_n911), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n913), .A2(new_n905), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n922), .A2(new_n917), .A3(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(G37), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n921), .A2(new_n926), .ZN(new_n927));
  XOR2_X1   g502(.A(KEYINPUT110), .B(KEYINPUT40), .Z(new_n928));
  XNOR2_X1  g503(.A(new_n927), .B(new_n928), .ZN(G395));
  XNOR2_X1  g504(.A(G290), .B(G288), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT112), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n930), .B(new_n931), .ZN(new_n932));
  XNOR2_X1  g507(.A(G305), .B(G303), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  AND2_X1   g509(.A1(new_n930), .A2(new_n931), .ZN(new_n935));
  OR2_X1    g510(.A1(new_n935), .A2(new_n933), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(KEYINPUT42), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n935), .A2(new_n933), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n939), .B1(new_n932), .B2(new_n933), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT42), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n630), .B1(new_n591), .B2(new_n595), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n859), .A2(new_n943), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n944), .B1(G299), .B2(new_n635), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT41), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n946), .B1(new_n859), .B2(new_n943), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n947), .B1(G299), .B2(new_n635), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(KEYINPUT111), .ZN(new_n949));
  INV_X1    g524(.A(G299), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n861), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT111), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n951), .A2(new_n952), .A3(new_n947), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n945), .A2(new_n946), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n949), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n642), .B(new_n877), .ZN(new_n956));
  MUX2_X1   g531(.A(new_n945), .B(new_n955), .S(new_n956), .Z(new_n957));
  AND3_X1   g532(.A1(new_n938), .A2(new_n942), .A3(new_n957), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n957), .B1(new_n938), .B2(new_n942), .ZN(new_n959));
  OAI21_X1  g534(.A(G868), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(new_n874), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n960), .B1(G868), .B2(new_n961), .ZN(G295));
  OAI21_X1  g537(.A(new_n960), .B1(G868), .B2(new_n961), .ZN(G331));
  INV_X1    g538(.A(KEYINPUT82), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n964), .B1(new_n545), .B2(new_n556), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n600), .A2(KEYINPUT82), .A3(new_n601), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n561), .A2(new_n564), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(KEYINPUT79), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n561), .A2(new_n562), .A3(new_n564), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n967), .A2(new_n971), .A3(new_n560), .ZN(new_n972));
  INV_X1    g547(.A(G168), .ZN(new_n973));
  NAND2_X1  g548(.A1(G301), .A2(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n972), .A2(new_n974), .A3(new_n877), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(KEYINPUT113), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT113), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n972), .A2(new_n974), .A3(new_n877), .A4(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n972), .A2(new_n974), .ZN(new_n980));
  AOI22_X1  g555(.A1(new_n951), .A2(new_n944), .B1(new_n980), .B2(new_n883), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n979), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(KEYINPUT116), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n954), .A2(new_n948), .ZN(new_n984));
  NOR2_X1   g559(.A1(G301), .A2(G286), .ZN(new_n985));
  AOI21_X1  g560(.A(G168), .B1(new_n971), .B2(new_n560), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n883), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(new_n975), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n984), .A2(KEYINPUT115), .A3(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT115), .ZN(new_n990));
  AOI22_X1  g565(.A1(new_n945), .A2(new_n946), .B1(new_n951), .B2(new_n947), .ZN(new_n991));
  AND3_X1   g566(.A1(new_n972), .A2(new_n974), .A3(new_n877), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n877), .B1(new_n972), .B2(new_n974), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n990), .B1(new_n991), .B2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT116), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n979), .A2(new_n981), .A3(new_n996), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n983), .A2(new_n989), .A3(new_n995), .A4(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(new_n940), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n979), .A2(new_n987), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n987), .A2(new_n945), .A3(new_n975), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(KEYINPUT114), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT114), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n987), .A2(new_n945), .A3(new_n1003), .A4(new_n975), .ZN(new_n1004));
  AOI22_X1  g579(.A1(new_n955), .A2(new_n1000), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(G37), .B1(new_n1005), .B2(new_n937), .ZN(new_n1006));
  AND3_X1   g581(.A1(new_n999), .A2(KEYINPUT43), .A3(new_n1006), .ZN(new_n1007));
  OR2_X1    g582(.A1(new_n1005), .A2(new_n937), .ZN(new_n1008));
  AOI21_X1  g583(.A(KEYINPUT43), .B1(new_n1008), .B2(new_n1006), .ZN(new_n1009));
  OAI21_X1  g584(.A(KEYINPUT44), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT44), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT43), .ZN(new_n1012));
  AND3_X1   g587(.A1(new_n999), .A2(new_n1012), .A3(new_n1006), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1012), .B1(new_n1008), .B2(new_n1006), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1011), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1010), .A2(new_n1015), .ZN(G397));
  AND2_X1   g591(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1017));
  NOR2_X1   g592(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n506), .A2(new_n510), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n512), .A2(new_n514), .ZN(new_n1021));
  AOI21_X1  g596(.A(G1384), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g597(.A(KEYINPUT117), .B1(new_n1022), .B2(KEYINPUT45), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT117), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT45), .ZN(new_n1025));
  OAI211_X1 g600(.A(new_n1024), .B(new_n1025), .C1(G164), .C2(G1384), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1023), .A2(new_n1026), .ZN(new_n1027));
  AOI22_X1  g602(.A1(new_n484), .A2(KEYINPUT71), .B1(G113), .B2(G2104), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n472), .B1(new_n1028), .B2(new_n487), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1025), .A2(G1384), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(new_n908), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1031), .B1(new_n1021), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(G40), .ZN(new_n1034));
  NOR4_X1   g609(.A1(new_n1029), .A2(new_n1033), .A3(new_n1034), .A4(new_n478), .ZN(new_n1035));
  AND2_X1   g610(.A1(new_n1027), .A2(new_n1035), .ZN(new_n1036));
  XNOR2_X1  g611(.A(KEYINPUT56), .B(G2072), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NOR3_X1   g613(.A1(new_n1029), .A2(new_n1034), .A3(new_n478), .ZN(new_n1039));
  XOR2_X1   g614(.A(KEYINPUT118), .B(KEYINPUT50), .Z(new_n1040));
  INV_X1    g615(.A(new_n1040), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1041), .B1(new_n909), .B2(G1384), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT50), .ZN(new_n1043));
  AND3_X1   g618(.A1(new_n1022), .A2(KEYINPUT122), .A3(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(KEYINPUT122), .B1(new_n1022), .B2(new_n1043), .ZN(new_n1045));
  OAI211_X1 g620(.A(new_n1039), .B(new_n1042), .C1(new_n1044), .C2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(G1956), .ZN(new_n1047));
  AND3_X1   g622(.A1(new_n1046), .A2(KEYINPUT126), .A3(new_n1047), .ZN(new_n1048));
  AOI21_X1  g623(.A(KEYINPUT126), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1049));
  OAI211_X1 g624(.A(new_n1019), .B(new_n1038), .C1(new_n1048), .C2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT126), .ZN(new_n1051));
  NAND3_X1  g626(.A1(G160), .A2(G40), .A3(new_n1042), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1045), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1022), .A2(KEYINPUT122), .A3(new_n1043), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1052), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1051), .B1(new_n1055), .B2(G1956), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1046), .A2(KEYINPUT126), .A3(new_n1047), .ZN(new_n1057));
  AOI22_X1  g632(.A1(new_n1056), .A2(new_n1057), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1058), .A2(new_n1019), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n909), .A2(G1384), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1039), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(G2067), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1060), .A2(new_n1040), .ZN(new_n1064));
  OAI21_X1  g639(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1039), .A2(new_n1064), .A3(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(G1348), .ZN(new_n1067));
  AOI22_X1  g642(.A1(new_n1062), .A2(new_n1063), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1068), .A2(new_n861), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1050), .B1(new_n1059), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(G1996), .ZN(new_n1071));
  AND3_X1   g646(.A1(new_n1027), .A2(new_n1035), .A3(new_n1071), .ZN(new_n1072));
  XOR2_X1   g647(.A(KEYINPUT58), .B(G1341), .Z(new_n1073));
  INV_X1    g648(.A(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1074), .B1(new_n1039), .B2(new_n1060), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n575), .B1(new_n1072), .B2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(KEYINPUT59), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT59), .ZN(new_n1078));
  OAI211_X1 g653(.A(new_n1078), .B(new_n575), .C1(new_n1072), .C2(new_n1075), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n635), .A2(KEYINPUT60), .ZN(new_n1080));
  AND3_X1   g655(.A1(new_n1039), .A2(new_n1064), .A3(new_n1065), .ZN(new_n1081));
  OAI22_X1  g656(.A1(new_n1081), .A2(G1348), .B1(G2067), .B2(new_n1061), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n635), .A2(KEYINPUT60), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1080), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1068), .A2(KEYINPUT60), .A3(new_n635), .ZN(new_n1085));
  AOI22_X1  g660(.A1(new_n1077), .A2(new_n1079), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  OAI211_X1 g661(.A(new_n1050), .B(KEYINPUT61), .C1(new_n1058), .C2(new_n1019), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1038), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1089), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1090));
  AOI21_X1  g665(.A(KEYINPUT61), .B1(new_n1090), .B2(new_n1050), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1070), .B1(new_n1088), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT52), .ZN(new_n1093));
  OAI211_X1 g668(.A(KEYINPUT120), .B(new_n1093), .C1(new_n819), .C2(G1976), .ZN(new_n1094));
  XNOR2_X1  g669(.A(KEYINPUT119), .B(G8), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1095), .B1(new_n1039), .B2(new_n1060), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT120), .ZN(new_n1097));
  AOI21_X1  g672(.A(G1976), .B1(new_n605), .B2(new_n607), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1097), .B1(new_n1098), .B2(KEYINPUT52), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n819), .A2(G1976), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1094), .A2(new_n1096), .A3(new_n1099), .A4(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1096), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(KEYINPUT52), .ZN(new_n1103));
  INV_X1    g678(.A(G1981), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n609), .A2(new_n1104), .A3(new_n613), .ZN(new_n1105));
  INV_X1    g680(.A(G86), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n543), .A2(new_n544), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n613), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(G1981), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1105), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT49), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1105), .A2(new_n1109), .A3(KEYINPUT49), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1112), .A2(new_n1096), .A3(new_n1113), .ZN(new_n1114));
  AND3_X1   g689(.A1(new_n1101), .A2(new_n1103), .A3(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(G303), .A2(G8), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT55), .ZN(new_n1117));
  XNOR2_X1  g692(.A(new_n1116), .B(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(G1971), .B1(new_n1027), .B2(new_n1035), .ZN(new_n1120));
  INV_X1    g695(.A(G2090), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1120), .B1(new_n1121), .B2(new_n1055), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1119), .B1(new_n1122), .B2(new_n1095), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1066), .A2(G2090), .ZN(new_n1124));
  OAI211_X1 g699(.A(new_n1118), .B(G8), .C1(new_n1124), .C2(new_n1120), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1115), .A2(new_n1123), .A3(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(G1966), .ZN(new_n1127));
  OAI21_X1  g702(.A(KEYINPUT123), .B1(G164), .B2(new_n1031), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT123), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1129), .A2(new_n1130), .A3(new_n1030), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1025), .B1(new_n909), .B2(G1384), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1128), .A2(new_n1131), .A3(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(G160), .A2(G40), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1127), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(G2084), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1039), .A2(new_n1136), .A3(new_n1064), .A4(new_n1065), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1095), .B1(new_n1135), .B2(new_n1137), .ZN(new_n1138));
  NOR2_X1   g713(.A1(G168), .A2(new_n1095), .ZN(new_n1139));
  OR2_X1    g714(.A1(new_n1139), .A2(KEYINPUT51), .ZN(new_n1140));
  OR2_X1    g715(.A1(new_n1138), .A2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1138), .A2(new_n973), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(G8), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1144), .B1(new_n1135), .B2(new_n1137), .ZN(new_n1145));
  OAI21_X1  g720(.A(KEYINPUT51), .B1(new_n1145), .B2(new_n1139), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1141), .B1(new_n1143), .B2(new_n1146), .ZN(new_n1147));
  XOR2_X1   g722(.A(G301), .B(KEYINPUT54), .Z(new_n1148));
  NAND3_X1  g723(.A1(new_n1027), .A2(new_n1035), .A3(new_n754), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT53), .ZN(new_n1150));
  INV_X1    g725(.A(G1961), .ZN(new_n1151));
  AOI22_X1  g726(.A1(new_n1149), .A2(new_n1150), .B1(new_n1151), .B2(new_n1066), .ZN(new_n1152));
  NOR3_X1   g727(.A1(new_n1033), .A2(new_n1150), .A3(G2078), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1039), .A2(new_n1132), .A3(new_n1153), .ZN(new_n1154));
  AND3_X1   g729(.A1(new_n1148), .A2(new_n1152), .A3(new_n1154), .ZN(new_n1155));
  OR4_X1    g730(.A1(new_n1150), .A2(new_n1133), .A3(new_n1134), .A4(G2078), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1148), .B1(new_n1152), .B2(new_n1156), .ZN(new_n1157));
  NOR4_X1   g732(.A1(new_n1126), .A2(new_n1147), .A3(new_n1155), .A4(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1092), .A2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g734(.A(G301), .B1(new_n1152), .B2(new_n1156), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1115), .A2(new_n1123), .A3(new_n1125), .A4(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT62), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1147), .A2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1162), .A2(new_n1164), .A3(KEYINPUT127), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT127), .ZN(new_n1166));
  OAI211_X1 g741(.A(new_n1142), .B(KEYINPUT51), .C1(new_n1139), .C2(new_n1145), .ZN(new_n1167));
  AOI21_X1  g742(.A(KEYINPUT62), .B1(new_n1167), .B2(new_n1141), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1166), .B1(new_n1168), .B2(new_n1161), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1167), .A2(KEYINPUT62), .A3(new_n1141), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1165), .A2(new_n1169), .A3(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(new_n1105), .ZN(new_n1172));
  NOR2_X1   g747(.A1(G288), .A2(G1976), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1172), .B1(new_n1114), .B2(new_n1173), .ZN(new_n1174));
  AND2_X1   g749(.A1(new_n1174), .A2(KEYINPUT121), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1096), .B1(new_n1174), .B2(KEYINPUT121), .ZN(new_n1176));
  INV_X1    g751(.A(new_n1115), .ZN(new_n1177));
  OAI22_X1  g752(.A1(new_n1175), .A2(new_n1176), .B1(new_n1177), .B2(new_n1125), .ZN(new_n1178));
  INV_X1    g753(.A(new_n1138), .ZN(new_n1179));
  NOR3_X1   g754(.A1(new_n1179), .A2(KEYINPUT124), .A3(G286), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT124), .ZN(new_n1181));
  AOI21_X1  g756(.A(new_n1181), .B1(new_n1138), .B2(new_n967), .ZN(new_n1182));
  OR2_X1    g757(.A1(new_n1180), .A2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1125), .A2(KEYINPUT63), .ZN(new_n1184));
  OAI21_X1  g759(.A(G8), .B1(new_n1124), .B2(new_n1120), .ZN(new_n1185));
  AOI21_X1  g760(.A(new_n1184), .B1(new_n1119), .B2(new_n1185), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n1183), .A2(new_n1186), .A3(new_n1115), .ZN(new_n1187));
  XOR2_X1   g762(.A(KEYINPUT125), .B(KEYINPUT63), .Z(new_n1188));
  NOR2_X1   g763(.A1(new_n1180), .A2(new_n1182), .ZN(new_n1189));
  OAI21_X1  g764(.A(new_n1188), .B1(new_n1189), .B2(new_n1126), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n1178), .B1(new_n1187), .B2(new_n1190), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1159), .A2(new_n1171), .A3(new_n1191), .ZN(new_n1192));
  NOR2_X1   g767(.A1(new_n1134), .A2(new_n1132), .ZN(new_n1193));
  OR2_X1    g768(.A1(new_n845), .A2(new_n848), .ZN(new_n1194));
  XNOR2_X1  g769(.A(new_n798), .B(new_n1063), .ZN(new_n1195));
  XNOR2_X1  g770(.A(new_n766), .B(new_n1071), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n845), .A2(new_n848), .ZN(new_n1197));
  NAND4_X1  g772(.A1(new_n1194), .A2(new_n1195), .A3(new_n1196), .A4(new_n1197), .ZN(new_n1198));
  NOR2_X1   g773(.A1(G290), .A2(G1986), .ZN(new_n1199));
  OR2_X1    g774(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  AND2_X1   g775(.A1(G290), .A2(G1986), .ZN(new_n1201));
  OAI21_X1  g776(.A(new_n1193), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1192), .A2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1199), .A2(new_n1193), .ZN(new_n1204));
  INV_X1    g779(.A(new_n1204), .ZN(new_n1205));
  NOR2_X1   g780(.A1(new_n1205), .A2(KEYINPUT48), .ZN(new_n1206));
  AND2_X1   g781(.A1(new_n1205), .A2(KEYINPUT48), .ZN(new_n1207));
  AOI211_X1 g782(.A(new_n1206), .B(new_n1207), .C1(new_n1193), .C2(new_n1198), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1193), .A2(new_n1071), .ZN(new_n1209));
  XNOR2_X1  g784(.A(new_n1209), .B(KEYINPUT46), .ZN(new_n1210));
  INV_X1    g785(.A(new_n1195), .ZN(new_n1211));
  OAI21_X1  g786(.A(new_n1193), .B1(new_n1211), .B2(new_n766), .ZN(new_n1212));
  NAND2_X1  g787(.A1(new_n1210), .A2(new_n1212), .ZN(new_n1213));
  XOR2_X1   g788(.A(new_n1213), .B(KEYINPUT47), .Z(new_n1214));
  NAND2_X1  g789(.A1(new_n1196), .A2(new_n1195), .ZN(new_n1215));
  OAI22_X1  g790(.A1(new_n1197), .A2(new_n1215), .B1(G2067), .B2(new_n798), .ZN(new_n1216));
  AOI211_X1 g791(.A(new_n1208), .B(new_n1214), .C1(new_n1193), .C2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g792(.A1(new_n1203), .A2(new_n1217), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g793(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1220));
  NAND2_X1  g794(.A1(G319), .A2(new_n698), .ZN(new_n1221));
  AOI21_X1  g795(.A(new_n1221), .B1(new_n724), .B2(new_n725), .ZN(new_n1222));
  OAI211_X1 g796(.A(new_n1222), .B(new_n678), .C1(new_n921), .C2(new_n926), .ZN(new_n1223));
  NOR2_X1   g797(.A1(new_n1220), .A2(new_n1223), .ZN(G308));
  AND2_X1   g798(.A1(new_n678), .A2(new_n1222), .ZN(new_n1225));
  OAI221_X1 g799(.A(new_n1225), .B1(new_n921), .B2(new_n926), .C1(new_n1013), .C2(new_n1014), .ZN(G225));
endmodule


