

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
         n1047, n1048, n1049, n1050;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XOR2_X1 U562 ( .A(KEYINPUT65), .B(n534), .Z(n531) );
  OR2_X1 U563 ( .A1(n642), .A2(n968), .ZN(n643) );
  BUF_X1 U564 ( .A(n642), .Z(n668) );
  INV_X1 U565 ( .A(KEYINPUT29), .ZN(n662) );
  OR2_X1 U566 ( .A1(n684), .A2(n683), .ZN(n697) );
  NAND2_X1 U567 ( .A1(n607), .A2(n712), .ZN(n642) );
  INV_X1 U568 ( .A(KEYINPUT17), .ZN(n532) );
  INV_X1 U569 ( .A(KEYINPUT100), .ZN(n709) );
  NAND2_X1 U570 ( .A1(n900), .A2(G138), .ZN(n554) );
  NOR2_X1 U571 ( .A1(G651), .A2(n586), .ZN(n806) );
  XNOR2_X1 U572 ( .A(n556), .B(KEYINPUT89), .ZN(n558) );
  NOR2_X1 U573 ( .A1(G2104), .A2(G2105), .ZN(n533) );
  XNOR2_X2 U574 ( .A(n533), .B(n532), .ZN(n900) );
  NAND2_X1 U575 ( .A1(n900), .A2(G137), .ZN(n537) );
  AND2_X1 U576 ( .A1(G2104), .A2(G2105), .ZN(n905) );
  NAND2_X1 U577 ( .A1(G113), .A2(n905), .ZN(n534) );
  INV_X1 U578 ( .A(G2105), .ZN(n538) );
  NOR2_X2 U579 ( .A1(G2104), .A2(n538), .ZN(n903) );
  NAND2_X1 U580 ( .A1(G125), .A2(n903), .ZN(n535) );
  AND2_X1 U581 ( .A1(n531), .A2(n535), .ZN(n536) );
  AND2_X1 U582 ( .A1(n537), .A2(n536), .ZN(n541) );
  AND2_X1 U583 ( .A1(n538), .A2(G2104), .ZN(n899) );
  NAND2_X1 U584 ( .A1(G101), .A2(n899), .ZN(n539) );
  XOR2_X1 U585 ( .A(KEYINPUT23), .B(n539), .Z(n540) );
  NAND2_X1 U586 ( .A1(n541), .A2(n540), .ZN(n542) );
  XOR2_X2 U587 ( .A(KEYINPUT64), .B(n542), .Z(G160) );
  INV_X1 U588 ( .A(G651), .ZN(n547) );
  NOR2_X1 U589 ( .A1(G543), .A2(n547), .ZN(n543) );
  XOR2_X1 U590 ( .A(KEYINPUT1), .B(n543), .Z(n544) );
  XNOR2_X1 U591 ( .A(KEYINPUT66), .B(n544), .ZN(n807) );
  NAND2_X1 U592 ( .A1(n807), .A2(G64), .ZN(n546) );
  XOR2_X1 U593 ( .A(KEYINPUT0), .B(G543), .Z(n586) );
  NAND2_X1 U594 ( .A1(n806), .A2(G52), .ZN(n545) );
  AND2_X1 U595 ( .A1(n546), .A2(n545), .ZN(n553) );
  XNOR2_X1 U596 ( .A(KEYINPUT9), .B(KEYINPUT68), .ZN(n551) );
  NOR2_X1 U597 ( .A1(G651), .A2(G543), .ZN(n802) );
  NAND2_X1 U598 ( .A1(G90), .A2(n802), .ZN(n549) );
  NOR2_X1 U599 ( .A1(n586), .A2(n547), .ZN(n803) );
  NAND2_X1 U600 ( .A1(G77), .A2(n803), .ZN(n548) );
  NAND2_X1 U601 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U602 ( .A(n551), .B(n550), .ZN(n552) );
  NAND2_X1 U603 ( .A1(n553), .A2(n552), .ZN(G301) );
  INV_X1 U604 ( .A(G301), .ZN(G171) );
  NAND2_X1 U605 ( .A1(G102), .A2(n899), .ZN(n555) );
  NAND2_X1 U606 ( .A1(n555), .A2(n554), .ZN(n556) );
  NAND2_X1 U607 ( .A1(G126), .A2(n903), .ZN(n557) );
  NAND2_X1 U608 ( .A1(n558), .A2(n557), .ZN(n561) );
  NAND2_X1 U609 ( .A1(G114), .A2(n905), .ZN(n559) );
  XOR2_X1 U610 ( .A(KEYINPUT88), .B(n559), .Z(n560) );
  NOR2_X1 U611 ( .A1(n561), .A2(n560), .ZN(G164) );
  NAND2_X1 U612 ( .A1(n802), .A2(G89), .ZN(n562) );
  XNOR2_X1 U613 ( .A(n562), .B(KEYINPUT4), .ZN(n564) );
  NAND2_X1 U614 ( .A1(G76), .A2(n803), .ZN(n563) );
  NAND2_X1 U615 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U616 ( .A(n565), .B(KEYINPUT5), .ZN(n570) );
  NAND2_X1 U617 ( .A1(n806), .A2(G51), .ZN(n567) );
  NAND2_X1 U618 ( .A1(G63), .A2(n807), .ZN(n566) );
  NAND2_X1 U619 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U620 ( .A(KEYINPUT6), .B(n568), .Z(n569) );
  NAND2_X1 U621 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U622 ( .A(n571), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U623 ( .A1(G91), .A2(n802), .ZN(n573) );
  NAND2_X1 U624 ( .A1(G78), .A2(n803), .ZN(n572) );
  NAND2_X1 U625 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U626 ( .A(KEYINPUT69), .B(n574), .ZN(n578) );
  NAND2_X1 U627 ( .A1(n807), .A2(G65), .ZN(n576) );
  NAND2_X1 U628 ( .A1(n806), .A2(G53), .ZN(n575) );
  AND2_X1 U629 ( .A1(n576), .A2(n575), .ZN(n577) );
  NAND2_X1 U630 ( .A1(n578), .A2(n577), .ZN(G299) );
  XOR2_X1 U631 ( .A(G168), .B(KEYINPUT8), .Z(n579) );
  XNOR2_X1 U632 ( .A(KEYINPUT76), .B(n579), .ZN(G286) );
  NAND2_X1 U633 ( .A1(G88), .A2(n802), .ZN(n581) );
  NAND2_X1 U634 ( .A1(G75), .A2(n803), .ZN(n580) );
  NAND2_X1 U635 ( .A1(n581), .A2(n580), .ZN(n585) );
  NAND2_X1 U636 ( .A1(n806), .A2(G50), .ZN(n583) );
  NAND2_X1 U637 ( .A1(G62), .A2(n807), .ZN(n582) );
  NAND2_X1 U638 ( .A1(n583), .A2(n582), .ZN(n584) );
  NOR2_X1 U639 ( .A1(n585), .A2(n584), .ZN(G166) );
  NAND2_X1 U640 ( .A1(G87), .A2(n586), .ZN(n588) );
  NAND2_X1 U641 ( .A1(G74), .A2(G651), .ZN(n587) );
  NAND2_X1 U642 ( .A1(n588), .A2(n587), .ZN(n589) );
  NOR2_X1 U643 ( .A1(n807), .A2(n589), .ZN(n591) );
  NAND2_X1 U644 ( .A1(n806), .A2(G49), .ZN(n590) );
  NAND2_X1 U645 ( .A1(n591), .A2(n590), .ZN(G288) );
  INV_X1 U646 ( .A(G166), .ZN(G303) );
  NAND2_X1 U647 ( .A1(G48), .A2(n806), .ZN(n598) );
  NAND2_X1 U648 ( .A1(G86), .A2(n802), .ZN(n593) );
  NAND2_X1 U649 ( .A1(G61), .A2(n807), .ZN(n592) );
  NAND2_X1 U650 ( .A1(n593), .A2(n592), .ZN(n596) );
  NAND2_X1 U651 ( .A1(n803), .A2(G73), .ZN(n594) );
  XOR2_X1 U652 ( .A(KEYINPUT2), .B(n594), .Z(n595) );
  NOR2_X1 U653 ( .A1(n596), .A2(n595), .ZN(n597) );
  NAND2_X1 U654 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U655 ( .A(n599), .B(KEYINPUT84), .ZN(G305) );
  NAND2_X1 U656 ( .A1(G85), .A2(n802), .ZN(n601) );
  NAND2_X1 U657 ( .A1(G60), .A2(n807), .ZN(n600) );
  NAND2_X1 U658 ( .A1(n601), .A2(n600), .ZN(n605) );
  NAND2_X1 U659 ( .A1(G72), .A2(n803), .ZN(n603) );
  NAND2_X1 U660 ( .A1(G47), .A2(n806), .ZN(n602) );
  NAND2_X1 U661 ( .A1(n603), .A2(n602), .ZN(n604) );
  NOR2_X1 U662 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X1 U663 ( .A(KEYINPUT67), .B(n606), .ZN(G290) );
  INV_X1 U664 ( .A(KEYINPUT32), .ZN(n677) );
  NAND2_X1 U665 ( .A1(G40), .A2(G160), .ZN(n711) );
  INV_X1 U666 ( .A(n711), .ZN(n607) );
  NOR2_X1 U667 ( .A1(G164), .A2(G1384), .ZN(n712) );
  XNOR2_X1 U668 ( .A(KEYINPUT97), .B(n642), .ZN(n619) );
  BUF_X1 U669 ( .A(n619), .Z(n648) );
  XNOR2_X1 U670 ( .A(KEYINPUT25), .B(G2078), .ZN(n967) );
  NAND2_X1 U671 ( .A1(n648), .A2(n967), .ZN(n609) );
  INV_X1 U672 ( .A(G1961), .ZN(n1033) );
  NAND2_X1 U673 ( .A1(n668), .A2(n1033), .ZN(n608) );
  NAND2_X1 U674 ( .A1(n609), .A2(n608), .ZN(n618) );
  NOR2_X1 U675 ( .A1(G171), .A2(n618), .ZN(n615) );
  NAND2_X2 U676 ( .A1(G8), .A2(n642), .ZN(n706) );
  NOR2_X1 U677 ( .A1(G1966), .A2(n706), .ZN(n681) );
  NOR2_X1 U678 ( .A1(G2084), .A2(n642), .ZN(n680) );
  INV_X1 U679 ( .A(n680), .ZN(n610) );
  NAND2_X1 U680 ( .A1(G8), .A2(n610), .ZN(n611) );
  OR2_X1 U681 ( .A1(n681), .A2(n611), .ZN(n612) );
  XNOR2_X1 U682 ( .A(n612), .B(KEYINPUT30), .ZN(n613) );
  NOR2_X1 U683 ( .A1(G168), .A2(n613), .ZN(n614) );
  NOR2_X1 U684 ( .A1(n615), .A2(n614), .ZN(n616) );
  XOR2_X1 U685 ( .A(n616), .B(KEYINPUT31), .Z(n617) );
  XNOR2_X1 U686 ( .A(KEYINPUT98), .B(n617), .ZN(n678) );
  NAND2_X1 U687 ( .A1(n618), .A2(G171), .ZN(n665) );
  INV_X1 U688 ( .A(G299), .ZN(n813) );
  NAND2_X1 U689 ( .A1(n619), .A2(G2072), .ZN(n620) );
  XNOR2_X1 U690 ( .A(n620), .B(KEYINPUT27), .ZN(n622) );
  INV_X1 U691 ( .A(G1956), .ZN(n1028) );
  NOR2_X1 U692 ( .A1(n1028), .A2(n648), .ZN(n621) );
  NOR2_X1 U693 ( .A1(n622), .A2(n621), .ZN(n657) );
  NAND2_X1 U694 ( .A1(n813), .A2(n657), .ZN(n656) );
  NAND2_X1 U695 ( .A1(G92), .A2(n802), .ZN(n624) );
  NAND2_X1 U696 ( .A1(G79), .A2(n803), .ZN(n623) );
  NAND2_X1 U697 ( .A1(n624), .A2(n623), .ZN(n628) );
  NAND2_X1 U698 ( .A1(n806), .A2(G54), .ZN(n626) );
  NAND2_X1 U699 ( .A1(G66), .A2(n807), .ZN(n625) );
  NAND2_X1 U700 ( .A1(n626), .A2(n625), .ZN(n627) );
  NOR2_X1 U701 ( .A1(n628), .A2(n627), .ZN(n629) );
  XOR2_X1 U702 ( .A(KEYINPUT15), .B(n629), .Z(n630) );
  XNOR2_X1 U703 ( .A(KEYINPUT74), .B(n630), .ZN(n916) );
  NAND2_X1 U704 ( .A1(n802), .A2(G81), .ZN(n631) );
  XNOR2_X1 U705 ( .A(n631), .B(KEYINPUT12), .ZN(n633) );
  NAND2_X1 U706 ( .A1(G68), .A2(n803), .ZN(n632) );
  NAND2_X1 U707 ( .A1(n633), .A2(n632), .ZN(n634) );
  XNOR2_X1 U708 ( .A(n634), .B(KEYINPUT13), .ZN(n638) );
  NAND2_X1 U709 ( .A1(n807), .A2(G56), .ZN(n635) );
  XNOR2_X1 U710 ( .A(n635), .B(KEYINPUT70), .ZN(n636) );
  XNOR2_X1 U711 ( .A(KEYINPUT14), .B(n636), .ZN(n637) );
  NAND2_X1 U712 ( .A1(n638), .A2(n637), .ZN(n639) );
  XNOR2_X1 U713 ( .A(n639), .B(KEYINPUT71), .ZN(n641) );
  NAND2_X1 U714 ( .A1(G43), .A2(n806), .ZN(n640) );
  NAND2_X1 U715 ( .A1(n641), .A2(n640), .ZN(n1011) );
  INV_X1 U716 ( .A(G1996), .ZN(n968) );
  XNOR2_X1 U717 ( .A(n643), .B(KEYINPUT26), .ZN(n645) );
  NAND2_X1 U718 ( .A1(n668), .A2(G1341), .ZN(n644) );
  NAND2_X1 U719 ( .A1(n645), .A2(n644), .ZN(n646) );
  NOR2_X1 U720 ( .A1(n1011), .A2(n646), .ZN(n647) );
  OR2_X1 U721 ( .A1(n916), .A2(n647), .ZN(n654) );
  NAND2_X1 U722 ( .A1(n647), .A2(n916), .ZN(n652) );
  NAND2_X1 U723 ( .A1(n648), .A2(G2067), .ZN(n650) );
  NAND2_X1 U724 ( .A1(G1348), .A2(n668), .ZN(n649) );
  NAND2_X1 U725 ( .A1(n650), .A2(n649), .ZN(n651) );
  NAND2_X1 U726 ( .A1(n652), .A2(n651), .ZN(n653) );
  NAND2_X1 U727 ( .A1(n654), .A2(n653), .ZN(n655) );
  NAND2_X1 U728 ( .A1(n656), .A2(n655), .ZN(n661) );
  NOR2_X1 U729 ( .A1(n813), .A2(n657), .ZN(n659) );
  INV_X1 U730 ( .A(KEYINPUT28), .ZN(n658) );
  XNOR2_X1 U731 ( .A(n659), .B(n658), .ZN(n660) );
  NAND2_X1 U732 ( .A1(n661), .A2(n660), .ZN(n663) );
  XNOR2_X1 U733 ( .A(n663), .B(n662), .ZN(n664) );
  NAND2_X1 U734 ( .A1(n665), .A2(n664), .ZN(n679) );
  NAND2_X1 U735 ( .A1(n678), .A2(n679), .ZN(n666) );
  NAND2_X1 U736 ( .A1(n666), .A2(G286), .ZN(n675) );
  INV_X1 U737 ( .A(G8), .ZN(n673) );
  NOR2_X1 U738 ( .A1(G1971), .A2(n706), .ZN(n667) );
  XNOR2_X1 U739 ( .A(KEYINPUT99), .B(n667), .ZN(n671) );
  NOR2_X1 U740 ( .A1(G2090), .A2(n668), .ZN(n669) );
  NOR2_X1 U741 ( .A1(G166), .A2(n669), .ZN(n670) );
  NAND2_X1 U742 ( .A1(n671), .A2(n670), .ZN(n672) );
  OR2_X1 U743 ( .A1(n673), .A2(n672), .ZN(n674) );
  NAND2_X1 U744 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U745 ( .A(n677), .B(n676), .ZN(n696) );
  AND2_X1 U746 ( .A1(n679), .A2(n678), .ZN(n684) );
  AND2_X1 U747 ( .A1(G8), .A2(n680), .ZN(n682) );
  OR2_X1 U748 ( .A1(n682), .A2(n681), .ZN(n683) );
  NAND2_X1 U749 ( .A1(G1976), .A2(G288), .ZN(n686) );
  AND2_X1 U750 ( .A1(n697), .A2(n686), .ZN(n685) );
  NAND2_X1 U751 ( .A1(n696), .A2(n685), .ZN(n689) );
  INV_X1 U752 ( .A(n686), .ZN(n999) );
  NOR2_X1 U753 ( .A1(G1976), .A2(G288), .ZN(n1000) );
  NOR2_X1 U754 ( .A1(G1971), .A2(G303), .ZN(n998) );
  NOR2_X1 U755 ( .A1(n1000), .A2(n998), .ZN(n687) );
  OR2_X1 U756 ( .A1(n999), .A2(n687), .ZN(n688) );
  AND2_X1 U757 ( .A1(n689), .A2(n688), .ZN(n690) );
  NOR2_X1 U758 ( .A1(n690), .A2(n706), .ZN(n691) );
  NOR2_X1 U759 ( .A1(KEYINPUT33), .A2(n691), .ZN(n694) );
  NAND2_X1 U760 ( .A1(n1000), .A2(KEYINPUT33), .ZN(n692) );
  NOR2_X1 U761 ( .A1(n692), .A2(n706), .ZN(n693) );
  NOR2_X1 U762 ( .A1(n694), .A2(n693), .ZN(n695) );
  XOR2_X1 U763 ( .A(G1981), .B(G305), .Z(n991) );
  NAND2_X1 U764 ( .A1(n695), .A2(n991), .ZN(n703) );
  NAND2_X1 U765 ( .A1(n697), .A2(n696), .ZN(n700) );
  NOR2_X1 U766 ( .A1(G2090), .A2(G303), .ZN(n698) );
  NAND2_X1 U767 ( .A1(G8), .A2(n698), .ZN(n699) );
  NAND2_X1 U768 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U769 ( .A1(n701), .A2(n706), .ZN(n702) );
  NAND2_X1 U770 ( .A1(n703), .A2(n702), .ZN(n708) );
  NOR2_X1 U771 ( .A1(G1981), .A2(G305), .ZN(n704) );
  XOR2_X1 U772 ( .A(n704), .B(KEYINPUT24), .Z(n705) );
  NOR2_X1 U773 ( .A1(n706), .A2(n705), .ZN(n707) );
  NOR2_X1 U774 ( .A1(n708), .A2(n707), .ZN(n710) );
  XNOR2_X1 U775 ( .A(n710), .B(n709), .ZN(n748) );
  XNOR2_X1 U776 ( .A(G1986), .B(G290), .ZN(n1008) );
  NOR2_X1 U777 ( .A1(n712), .A2(n711), .ZN(n760) );
  NAND2_X1 U778 ( .A1(n1008), .A2(n760), .ZN(n746) );
  XNOR2_X1 U779 ( .A(G2067), .B(KEYINPUT37), .ZN(n757) );
  NAND2_X1 U780 ( .A1(G104), .A2(n899), .ZN(n714) );
  NAND2_X1 U781 ( .A1(G140), .A2(n900), .ZN(n713) );
  NAND2_X1 U782 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U783 ( .A(KEYINPUT34), .B(n715), .ZN(n722) );
  NAND2_X1 U784 ( .A1(n905), .A2(G116), .ZN(n716) );
  XNOR2_X1 U785 ( .A(n716), .B(KEYINPUT90), .ZN(n718) );
  NAND2_X1 U786 ( .A1(G128), .A2(n903), .ZN(n717) );
  NAND2_X1 U787 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U788 ( .A(KEYINPUT35), .B(n719), .ZN(n720) );
  XNOR2_X1 U789 ( .A(KEYINPUT91), .B(n720), .ZN(n721) );
  NOR2_X1 U790 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U791 ( .A(KEYINPUT36), .B(n723), .ZN(n895) );
  NOR2_X1 U792 ( .A1(n757), .A2(n895), .ZN(n940) );
  NAND2_X1 U793 ( .A1(n760), .A2(n940), .ZN(n755) );
  INV_X1 U794 ( .A(n755), .ZN(n744) );
  XOR2_X1 U795 ( .A(n760), .B(KEYINPUT95), .Z(n742) );
  NAND2_X1 U796 ( .A1(G119), .A2(n903), .ZN(n724) );
  XOR2_X1 U797 ( .A(KEYINPUT92), .B(n724), .Z(n729) );
  NAND2_X1 U798 ( .A1(G95), .A2(n899), .ZN(n726) );
  NAND2_X1 U799 ( .A1(G131), .A2(n900), .ZN(n725) );
  NAND2_X1 U800 ( .A1(n726), .A2(n725), .ZN(n727) );
  XOR2_X1 U801 ( .A(KEYINPUT93), .B(n727), .Z(n728) );
  NOR2_X1 U802 ( .A1(n729), .A2(n728), .ZN(n731) );
  NAND2_X1 U803 ( .A1(n905), .A2(G107), .ZN(n730) );
  NAND2_X1 U804 ( .A1(n731), .A2(n730), .ZN(n885) );
  NAND2_X1 U805 ( .A1(G1991), .A2(n885), .ZN(n741) );
  XOR2_X1 U806 ( .A(KEYINPUT94), .B(KEYINPUT38), .Z(n733) );
  NAND2_X1 U807 ( .A1(G105), .A2(n899), .ZN(n732) );
  XNOR2_X1 U808 ( .A(n733), .B(n732), .ZN(n737) );
  NAND2_X1 U809 ( .A1(G141), .A2(n900), .ZN(n735) );
  NAND2_X1 U810 ( .A1(G117), .A2(n905), .ZN(n734) );
  NAND2_X1 U811 ( .A1(n735), .A2(n734), .ZN(n736) );
  NOR2_X1 U812 ( .A1(n737), .A2(n736), .ZN(n739) );
  NAND2_X1 U813 ( .A1(n903), .A2(G129), .ZN(n738) );
  NAND2_X1 U814 ( .A1(n739), .A2(n738), .ZN(n887) );
  NAND2_X1 U815 ( .A1(G1996), .A2(n887), .ZN(n740) );
  NAND2_X1 U816 ( .A1(n741), .A2(n740), .ZN(n948) );
  NAND2_X1 U817 ( .A1(n742), .A2(n948), .ZN(n743) );
  XOR2_X1 U818 ( .A(KEYINPUT96), .B(n743), .Z(n752) );
  NOR2_X1 U819 ( .A1(n744), .A2(n752), .ZN(n745) );
  AND2_X1 U820 ( .A1(n746), .A2(n745), .ZN(n747) );
  NAND2_X1 U821 ( .A1(n748), .A2(n747), .ZN(n763) );
  NOR2_X1 U822 ( .A1(G1996), .A2(n887), .ZN(n749) );
  XOR2_X1 U823 ( .A(KEYINPUT101), .B(n749), .Z(n944) );
  NOR2_X1 U824 ( .A1(G1986), .A2(G290), .ZN(n750) );
  NOR2_X1 U825 ( .A1(G1991), .A2(n885), .ZN(n939) );
  NOR2_X1 U826 ( .A1(n750), .A2(n939), .ZN(n751) );
  NOR2_X1 U827 ( .A1(n752), .A2(n751), .ZN(n753) );
  NOR2_X1 U828 ( .A1(n944), .A2(n753), .ZN(n754) );
  XNOR2_X1 U829 ( .A(n754), .B(KEYINPUT39), .ZN(n756) );
  NAND2_X1 U830 ( .A1(n756), .A2(n755), .ZN(n758) );
  NAND2_X1 U831 ( .A1(n757), .A2(n895), .ZN(n953) );
  NAND2_X1 U832 ( .A1(n758), .A2(n953), .ZN(n759) );
  XNOR2_X1 U833 ( .A(KEYINPUT102), .B(n759), .ZN(n761) );
  NAND2_X1 U834 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U835 ( .A1(n763), .A2(n762), .ZN(n764) );
  XNOR2_X1 U836 ( .A(n764), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U837 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U838 ( .A(G132), .ZN(G219) );
  INV_X1 U839 ( .A(G82), .ZN(G220) );
  INV_X1 U840 ( .A(G57), .ZN(G237) );
  INV_X1 U841 ( .A(G120), .ZN(G236) );
  NAND2_X1 U842 ( .A1(G7), .A2(G661), .ZN(n765) );
  XNOR2_X1 U843 ( .A(n765), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U844 ( .A(G223), .ZN(n840) );
  NAND2_X1 U845 ( .A1(n840), .A2(G567), .ZN(n766) );
  XOR2_X1 U846 ( .A(KEYINPUT11), .B(n766), .Z(G234) );
  INV_X1 U847 ( .A(G860), .ZN(n801) );
  NOR2_X1 U848 ( .A1(n1011), .A2(n801), .ZN(n767) );
  XOR2_X1 U849 ( .A(KEYINPUT72), .B(n767), .Z(G153) );
  INV_X1 U850 ( .A(G868), .ZN(n822) );
  NOR2_X1 U851 ( .A1(KEYINPUT73), .A2(G171), .ZN(n768) );
  NOR2_X1 U852 ( .A1(KEYINPUT75), .A2(n768), .ZN(n769) );
  NOR2_X1 U853 ( .A1(n822), .A2(n769), .ZN(n775) );
  NAND2_X1 U854 ( .A1(G301), .A2(G868), .ZN(n770) );
  NAND2_X1 U855 ( .A1(n770), .A2(KEYINPUT73), .ZN(n773) );
  NOR2_X1 U856 ( .A1(KEYINPUT75), .A2(n916), .ZN(n771) );
  NAND2_X1 U857 ( .A1(n822), .A2(n771), .ZN(n772) );
  NAND2_X1 U858 ( .A1(n773), .A2(n772), .ZN(n774) );
  NOR2_X1 U859 ( .A1(n775), .A2(n774), .ZN(n777) );
  NAND2_X1 U860 ( .A1(KEYINPUT75), .A2(n916), .ZN(n776) );
  NAND2_X1 U861 ( .A1(n777), .A2(n776), .ZN(G284) );
  XNOR2_X1 U862 ( .A(KEYINPUT77), .B(G868), .ZN(n778) );
  NOR2_X1 U863 ( .A1(G286), .A2(n778), .ZN(n780) );
  NOR2_X1 U864 ( .A1(G868), .A2(G299), .ZN(n779) );
  NOR2_X1 U865 ( .A1(n780), .A2(n779), .ZN(G297) );
  NAND2_X1 U866 ( .A1(n801), .A2(G559), .ZN(n781) );
  NAND2_X1 U867 ( .A1(n781), .A2(n916), .ZN(n782) );
  XNOR2_X1 U868 ( .A(n782), .B(KEYINPUT78), .ZN(n783) );
  XNOR2_X1 U869 ( .A(KEYINPUT16), .B(n783), .ZN(G148) );
  INV_X1 U870 ( .A(n916), .ZN(n994) );
  NOR2_X1 U871 ( .A1(n994), .A2(n822), .ZN(n784) );
  XNOR2_X1 U872 ( .A(n784), .B(KEYINPUT79), .ZN(n785) );
  NOR2_X1 U873 ( .A1(G559), .A2(n785), .ZN(n787) );
  NOR2_X1 U874 ( .A1(G868), .A2(n1011), .ZN(n786) );
  NOR2_X1 U875 ( .A1(n787), .A2(n786), .ZN(G282) );
  XOR2_X1 U876 ( .A(G2100), .B(KEYINPUT82), .Z(n798) );
  NAND2_X1 U877 ( .A1(G123), .A2(n903), .ZN(n788) );
  XOR2_X1 U878 ( .A(KEYINPUT18), .B(n788), .Z(n794) );
  NAND2_X1 U879 ( .A1(n905), .A2(G111), .ZN(n789) );
  XNOR2_X1 U880 ( .A(n789), .B(KEYINPUT80), .ZN(n791) );
  NAND2_X1 U881 ( .A1(G99), .A2(n899), .ZN(n790) );
  NAND2_X1 U882 ( .A1(n791), .A2(n790), .ZN(n792) );
  XOR2_X1 U883 ( .A(KEYINPUT81), .B(n792), .Z(n793) );
  NOR2_X1 U884 ( .A1(n794), .A2(n793), .ZN(n796) );
  NAND2_X1 U885 ( .A1(n900), .A2(G135), .ZN(n795) );
  NAND2_X1 U886 ( .A1(n796), .A2(n795), .ZN(n941) );
  XOR2_X1 U887 ( .A(G2096), .B(n941), .Z(n797) );
  NAND2_X1 U888 ( .A1(n798), .A2(n797), .ZN(G156) );
  XNOR2_X1 U889 ( .A(n1011), .B(KEYINPUT83), .ZN(n800) );
  NAND2_X1 U890 ( .A1(n916), .A2(G559), .ZN(n799) );
  XNOR2_X1 U891 ( .A(n800), .B(n799), .ZN(n819) );
  NAND2_X1 U892 ( .A1(n801), .A2(n819), .ZN(n812) );
  NAND2_X1 U893 ( .A1(G93), .A2(n802), .ZN(n805) );
  NAND2_X1 U894 ( .A1(G80), .A2(n803), .ZN(n804) );
  NAND2_X1 U895 ( .A1(n805), .A2(n804), .ZN(n811) );
  NAND2_X1 U896 ( .A1(n806), .A2(G55), .ZN(n809) );
  NAND2_X1 U897 ( .A1(G67), .A2(n807), .ZN(n808) );
  NAND2_X1 U898 ( .A1(n809), .A2(n808), .ZN(n810) );
  NOR2_X1 U899 ( .A1(n811), .A2(n810), .ZN(n821) );
  XOR2_X1 U900 ( .A(n812), .B(n821), .Z(G145) );
  XNOR2_X1 U901 ( .A(G288), .B(KEYINPUT19), .ZN(n815) );
  XNOR2_X1 U902 ( .A(n813), .B(G305), .ZN(n814) );
  XNOR2_X1 U903 ( .A(n815), .B(n814), .ZN(n816) );
  XNOR2_X1 U904 ( .A(n821), .B(n816), .ZN(n818) );
  XNOR2_X1 U905 ( .A(G290), .B(G166), .ZN(n817) );
  XNOR2_X1 U906 ( .A(n818), .B(n817), .ZN(n914) );
  XOR2_X1 U907 ( .A(n914), .B(n819), .Z(n820) );
  NOR2_X1 U908 ( .A1(n822), .A2(n820), .ZN(n824) );
  AND2_X1 U909 ( .A1(n822), .A2(n821), .ZN(n823) );
  NOR2_X1 U910 ( .A1(n824), .A2(n823), .ZN(G295) );
  NAND2_X1 U911 ( .A1(G2078), .A2(G2084), .ZN(n825) );
  XNOR2_X1 U912 ( .A(n825), .B(KEYINPUT85), .ZN(n826) );
  XNOR2_X1 U913 ( .A(KEYINPUT20), .B(n826), .ZN(n827) );
  NAND2_X1 U914 ( .A1(n827), .A2(G2090), .ZN(n828) );
  XNOR2_X1 U915 ( .A(KEYINPUT21), .B(n828), .ZN(n829) );
  NAND2_X1 U916 ( .A1(n829), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U917 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U918 ( .A1(G236), .A2(G237), .ZN(n830) );
  NAND2_X1 U919 ( .A1(G69), .A2(n830), .ZN(n831) );
  XNOR2_X1 U920 ( .A(KEYINPUT87), .B(n831), .ZN(n832) );
  NAND2_X1 U921 ( .A1(n832), .A2(G108), .ZN(n845) );
  NAND2_X1 U922 ( .A1(n845), .A2(G567), .ZN(n838) );
  NOR2_X1 U923 ( .A1(G220), .A2(G219), .ZN(n833) );
  XOR2_X1 U924 ( .A(KEYINPUT22), .B(n833), .Z(n834) );
  NOR2_X1 U925 ( .A1(G218), .A2(n834), .ZN(n835) );
  NAND2_X1 U926 ( .A1(G96), .A2(n835), .ZN(n846) );
  NAND2_X1 U927 ( .A1(G2106), .A2(n846), .ZN(n836) );
  XNOR2_X1 U928 ( .A(KEYINPUT86), .B(n836), .ZN(n837) );
  NAND2_X1 U929 ( .A1(n838), .A2(n837), .ZN(n848) );
  NAND2_X1 U930 ( .A1(G483), .A2(G661), .ZN(n839) );
  NOR2_X1 U931 ( .A1(n848), .A2(n839), .ZN(n844) );
  NAND2_X1 U932 ( .A1(n844), .A2(G36), .ZN(G176) );
  NAND2_X1 U933 ( .A1(G2106), .A2(n840), .ZN(G217) );
  AND2_X1 U934 ( .A1(G15), .A2(G2), .ZN(n841) );
  NAND2_X1 U935 ( .A1(G661), .A2(n841), .ZN(G259) );
  NAND2_X1 U936 ( .A1(G3), .A2(G1), .ZN(n842) );
  XOR2_X1 U937 ( .A(KEYINPUT105), .B(n842), .Z(n843) );
  NAND2_X1 U938 ( .A1(n844), .A2(n843), .ZN(G188) );
  INV_X1 U940 ( .A(G108), .ZN(G238) );
  INV_X1 U941 ( .A(G96), .ZN(G221) );
  NOR2_X1 U942 ( .A1(n846), .A2(n845), .ZN(n847) );
  XNOR2_X1 U943 ( .A(n847), .B(KEYINPUT106), .ZN(G325) );
  INV_X1 U944 ( .A(G325), .ZN(G261) );
  INV_X1 U945 ( .A(n848), .ZN(G319) );
  XOR2_X1 U946 ( .A(KEYINPUT42), .B(G2072), .Z(n850) );
  XNOR2_X1 U947 ( .A(G2067), .B(G2084), .ZN(n849) );
  XNOR2_X1 U948 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U949 ( .A(n851), .B(G2096), .Z(n853) );
  XNOR2_X1 U950 ( .A(G2078), .B(G2090), .ZN(n852) );
  XNOR2_X1 U951 ( .A(n853), .B(n852), .ZN(n857) );
  XOR2_X1 U952 ( .A(G2100), .B(KEYINPUT43), .Z(n855) );
  XNOR2_X1 U953 ( .A(G2678), .B(KEYINPUT107), .ZN(n854) );
  XNOR2_X1 U954 ( .A(n855), .B(n854), .ZN(n856) );
  XOR2_X1 U955 ( .A(n857), .B(n856), .Z(G227) );
  XOR2_X1 U956 ( .A(G2474), .B(G1956), .Z(n859) );
  XNOR2_X1 U957 ( .A(G1986), .B(G1961), .ZN(n858) );
  XNOR2_X1 U958 ( .A(n859), .B(n858), .ZN(n860) );
  XOR2_X1 U959 ( .A(n860), .B(KEYINPUT108), .Z(n862) );
  XNOR2_X1 U960 ( .A(G1996), .B(G1991), .ZN(n861) );
  XNOR2_X1 U961 ( .A(n862), .B(n861), .ZN(n866) );
  XOR2_X1 U962 ( .A(G1976), .B(G1981), .Z(n864) );
  XNOR2_X1 U963 ( .A(G1966), .B(G1971), .ZN(n863) );
  XNOR2_X1 U964 ( .A(n864), .B(n863), .ZN(n865) );
  XOR2_X1 U965 ( .A(n866), .B(n865), .Z(n868) );
  XNOR2_X1 U966 ( .A(KEYINPUT41), .B(KEYINPUT109), .ZN(n867) );
  XNOR2_X1 U967 ( .A(n868), .B(n867), .ZN(G229) );
  NAND2_X1 U968 ( .A1(G124), .A2(n903), .ZN(n869) );
  XNOR2_X1 U969 ( .A(n869), .B(KEYINPUT44), .ZN(n872) );
  NAND2_X1 U970 ( .A1(G112), .A2(n905), .ZN(n870) );
  XOR2_X1 U971 ( .A(KEYINPUT111), .B(n870), .Z(n871) );
  NAND2_X1 U972 ( .A1(n872), .A2(n871), .ZN(n877) );
  NAND2_X1 U973 ( .A1(G136), .A2(n900), .ZN(n873) );
  XNOR2_X1 U974 ( .A(n873), .B(KEYINPUT110), .ZN(n875) );
  NAND2_X1 U975 ( .A1(n899), .A2(G100), .ZN(n874) );
  NAND2_X1 U976 ( .A1(n875), .A2(n874), .ZN(n876) );
  NOR2_X1 U977 ( .A1(n877), .A2(n876), .ZN(G162) );
  NAND2_X1 U978 ( .A1(G118), .A2(n905), .ZN(n879) );
  NAND2_X1 U979 ( .A1(G130), .A2(n903), .ZN(n878) );
  NAND2_X1 U980 ( .A1(n879), .A2(n878), .ZN(n884) );
  NAND2_X1 U981 ( .A1(G106), .A2(n899), .ZN(n881) );
  NAND2_X1 U982 ( .A1(G142), .A2(n900), .ZN(n880) );
  NAND2_X1 U983 ( .A1(n881), .A2(n880), .ZN(n882) );
  XOR2_X1 U984 ( .A(n882), .B(KEYINPUT45), .Z(n883) );
  NOR2_X1 U985 ( .A1(n884), .A2(n883), .ZN(n886) );
  XNOR2_X1 U986 ( .A(n886), .B(n885), .ZN(n894) );
  XNOR2_X1 U987 ( .A(KEYINPUT115), .B(KEYINPUT46), .ZN(n889) );
  XNOR2_X1 U988 ( .A(n887), .B(KEYINPUT48), .ZN(n888) );
  XNOR2_X1 U989 ( .A(n889), .B(n888), .ZN(n890) );
  XOR2_X1 U990 ( .A(n890), .B(KEYINPUT114), .Z(n892) );
  XNOR2_X1 U991 ( .A(G164), .B(KEYINPUT112), .ZN(n891) );
  XNOR2_X1 U992 ( .A(n892), .B(n891), .ZN(n893) );
  XNOR2_X1 U993 ( .A(n894), .B(n893), .ZN(n898) );
  XNOR2_X1 U994 ( .A(G162), .B(G160), .ZN(n896) );
  XNOR2_X1 U995 ( .A(n896), .B(n895), .ZN(n897) );
  XNOR2_X1 U996 ( .A(n898), .B(n897), .ZN(n912) );
  NAND2_X1 U997 ( .A1(G103), .A2(n899), .ZN(n902) );
  NAND2_X1 U998 ( .A1(G139), .A2(n900), .ZN(n901) );
  NAND2_X1 U999 ( .A1(n902), .A2(n901), .ZN(n910) );
  NAND2_X1 U1000 ( .A1(n903), .A2(G127), .ZN(n904) );
  XOR2_X1 U1001 ( .A(KEYINPUT113), .B(n904), .Z(n907) );
  NAND2_X1 U1002 ( .A1(n905), .A2(G115), .ZN(n906) );
  NAND2_X1 U1003 ( .A1(n907), .A2(n906), .ZN(n908) );
  XOR2_X1 U1004 ( .A(KEYINPUT47), .B(n908), .Z(n909) );
  NOR2_X1 U1005 ( .A1(n910), .A2(n909), .ZN(n957) );
  XOR2_X1 U1006 ( .A(n941), .B(n957), .Z(n911) );
  XNOR2_X1 U1007 ( .A(n912), .B(n911), .ZN(n913) );
  NOR2_X1 U1008 ( .A1(G37), .A2(n913), .ZN(G395) );
  XNOR2_X1 U1009 ( .A(n914), .B(n1011), .ZN(n915) );
  XNOR2_X1 U1010 ( .A(n915), .B(G286), .ZN(n918) );
  XOR2_X1 U1011 ( .A(n916), .B(G171), .Z(n917) );
  XNOR2_X1 U1012 ( .A(n918), .B(n917), .ZN(n919) );
  NOR2_X1 U1013 ( .A1(G37), .A2(n919), .ZN(G397) );
  XNOR2_X1 U1014 ( .A(G2451), .B(G2427), .ZN(n929) );
  XOR2_X1 U1015 ( .A(G2430), .B(G2443), .Z(n921) );
  XNOR2_X1 U1016 ( .A(KEYINPUT103), .B(G2438), .ZN(n920) );
  XNOR2_X1 U1017 ( .A(n921), .B(n920), .ZN(n925) );
  XOR2_X1 U1018 ( .A(G2435), .B(G2454), .Z(n923) );
  XNOR2_X1 U1019 ( .A(G1341), .B(G1348), .ZN(n922) );
  XNOR2_X1 U1020 ( .A(n923), .B(n922), .ZN(n924) );
  XOR2_X1 U1021 ( .A(n925), .B(n924), .Z(n927) );
  XNOR2_X1 U1022 ( .A(G2446), .B(KEYINPUT104), .ZN(n926) );
  XNOR2_X1 U1023 ( .A(n927), .B(n926), .ZN(n928) );
  XNOR2_X1 U1024 ( .A(n929), .B(n928), .ZN(n930) );
  NAND2_X1 U1025 ( .A1(n930), .A2(G14), .ZN(n938) );
  NAND2_X1 U1026 ( .A1(G319), .A2(n938), .ZN(n935) );
  XNOR2_X1 U1027 ( .A(KEYINPUT49), .B(KEYINPUT117), .ZN(n932) );
  NOR2_X1 U1028 ( .A1(G227), .A2(G229), .ZN(n931) );
  XNOR2_X1 U1029 ( .A(n932), .B(n931), .ZN(n933) );
  XOR2_X1 U1030 ( .A(KEYINPUT116), .B(n933), .Z(n934) );
  NOR2_X1 U1031 ( .A1(n935), .A2(n934), .ZN(n937) );
  NOR2_X1 U1032 ( .A1(G395), .A2(G397), .ZN(n936) );
  NAND2_X1 U1033 ( .A1(n937), .A2(n936), .ZN(G225) );
  INV_X1 U1034 ( .A(G225), .ZN(G308) );
  INV_X1 U1035 ( .A(G69), .ZN(G235) );
  INV_X1 U1036 ( .A(n938), .ZN(G401) );
  NOR2_X1 U1037 ( .A1(n940), .A2(n939), .ZN(n942) );
  NAND2_X1 U1038 ( .A1(n942), .A2(n941), .ZN(n952) );
  XOR2_X1 U1039 ( .A(G2090), .B(G162), .Z(n943) );
  NOR2_X1 U1040 ( .A1(n944), .A2(n943), .ZN(n945) );
  XOR2_X1 U1041 ( .A(KEYINPUT118), .B(n945), .Z(n946) );
  XNOR2_X1 U1042 ( .A(KEYINPUT51), .B(n946), .ZN(n950) );
  XOR2_X1 U1043 ( .A(G2084), .B(G160), .Z(n947) );
  NOR2_X1 U1044 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1045 ( .A1(n950), .A2(n949), .ZN(n951) );
  NOR2_X1 U1046 ( .A1(n952), .A2(n951), .ZN(n954) );
  NAND2_X1 U1047 ( .A1(n954), .A2(n953), .ZN(n955) );
  XOR2_X1 U1048 ( .A(KEYINPUT119), .B(n955), .Z(n962) );
  XOR2_X1 U1049 ( .A(G164), .B(G2078), .Z(n956) );
  XNOR2_X1 U1050 ( .A(KEYINPUT120), .B(n956), .ZN(n959) );
  XOR2_X1 U1051 ( .A(G2072), .B(n957), .Z(n958) );
  NOR2_X1 U1052 ( .A1(n959), .A2(n958), .ZN(n960) );
  XOR2_X1 U1053 ( .A(KEYINPUT50), .B(n960), .Z(n961) );
  NOR2_X1 U1054 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1055 ( .A(KEYINPUT52), .B(n963), .ZN(n964) );
  INV_X1 U1056 ( .A(KEYINPUT55), .ZN(n987) );
  NAND2_X1 U1057 ( .A1(n964), .A2(n987), .ZN(n965) );
  NAND2_X1 U1058 ( .A1(n965), .A2(G29), .ZN(n1049) );
  XNOR2_X1 U1059 ( .A(G2090), .B(G35), .ZN(n980) );
  XOR2_X1 U1060 ( .A(G2072), .B(G33), .Z(n966) );
  NAND2_X1 U1061 ( .A1(n966), .A2(G28), .ZN(n977) );
  XNOR2_X1 U1062 ( .A(n967), .B(G27), .ZN(n970) );
  XNOR2_X1 U1063 ( .A(n968), .B(G32), .ZN(n969) );
  NAND2_X1 U1064 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1065 ( .A(KEYINPUT121), .B(n971), .ZN(n975) );
  XNOR2_X1 U1066 ( .A(G2067), .B(G26), .ZN(n973) );
  XNOR2_X1 U1067 ( .A(G1991), .B(G25), .ZN(n972) );
  NOR2_X1 U1068 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1069 ( .A1(n975), .A2(n974), .ZN(n976) );
  NOR2_X1 U1070 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1071 ( .A(KEYINPUT53), .B(n978), .ZN(n979) );
  NOR2_X1 U1072 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1073 ( .A(KEYINPUT122), .B(n981), .ZN(n985) );
  XNOR2_X1 U1074 ( .A(KEYINPUT54), .B(KEYINPUT123), .ZN(n982) );
  XNOR2_X1 U1075 ( .A(n982), .B(G34), .ZN(n983) );
  XNOR2_X1 U1076 ( .A(G2084), .B(n983), .ZN(n984) );
  NAND2_X1 U1077 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1078 ( .A(n987), .B(n986), .ZN(n989) );
  INV_X1 U1079 ( .A(G29), .ZN(n988) );
  NAND2_X1 U1080 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1081 ( .A1(G11), .A2(n990), .ZN(n1047) );
  XNOR2_X1 U1082 ( .A(G16), .B(KEYINPUT56), .ZN(n1017) );
  XNOR2_X1 U1083 ( .A(G1966), .B(G168), .ZN(n992) );
  NAND2_X1 U1084 ( .A1(n992), .A2(n991), .ZN(n993) );
  XNOR2_X1 U1085 ( .A(n993), .B(KEYINPUT57), .ZN(n1015) );
  XNOR2_X1 U1086 ( .A(G301), .B(G1961), .ZN(n996) );
  XNOR2_X1 U1087 ( .A(n994), .B(G1348), .ZN(n995) );
  NOR2_X1 U1088 ( .A1(n996), .A2(n995), .ZN(n997) );
  XNOR2_X1 U1089 ( .A(KEYINPUT124), .B(n997), .ZN(n1010) );
  NOR2_X1 U1090 ( .A1(n999), .A2(n998), .ZN(n1006) );
  XNOR2_X1 U1091 ( .A(KEYINPUT125), .B(n1000), .ZN(n1002) );
  NAND2_X1 U1092 ( .A1(G1971), .A2(G303), .ZN(n1001) );
  NAND2_X1 U1093 ( .A1(n1002), .A2(n1001), .ZN(n1004) );
  XNOR2_X1 U1094 ( .A(G1956), .B(G299), .ZN(n1003) );
  NOR2_X1 U1095 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1096 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NOR2_X1 U1097 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1098 ( .A1(n1010), .A2(n1009), .ZN(n1013) );
  XNOR2_X1 U1099 ( .A(G1341), .B(n1011), .ZN(n1012) );
  NOR2_X1 U1100 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1101 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1102 ( .A1(n1017), .A2(n1016), .ZN(n1045) );
  INV_X1 U1103 ( .A(G16), .ZN(n1043) );
  XOR2_X1 U1104 ( .A(G1976), .B(G23), .Z(n1019) );
  XOR2_X1 U1105 ( .A(G1971), .B(G22), .Z(n1018) );
  NAND2_X1 U1106 ( .A1(n1019), .A2(n1018), .ZN(n1021) );
  XNOR2_X1 U1107 ( .A(G24), .B(G1986), .ZN(n1020) );
  NOR2_X1 U1108 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XOR2_X1 U1109 ( .A(KEYINPUT58), .B(n1022), .Z(n1040) );
  XNOR2_X1 U1110 ( .A(G1348), .B(KEYINPUT59), .ZN(n1023) );
  XNOR2_X1 U1111 ( .A(n1023), .B(G4), .ZN(n1027) );
  XNOR2_X1 U1112 ( .A(G1341), .B(G19), .ZN(n1025) );
  XNOR2_X1 U1113 ( .A(G6), .B(G1981), .ZN(n1024) );
  NOR2_X1 U1114 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NAND2_X1 U1115 ( .A1(n1027), .A2(n1026), .ZN(n1031) );
  XOR2_X1 U1116 ( .A(KEYINPUT126), .B(n1028), .Z(n1029) );
  XNOR2_X1 U1117 ( .A(G20), .B(n1029), .ZN(n1030) );
  NOR2_X1 U1118 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  XNOR2_X1 U1119 ( .A(KEYINPUT60), .B(n1032), .ZN(n1035) );
  XNOR2_X1 U1120 ( .A(n1033), .B(G5), .ZN(n1034) );
  NAND2_X1 U1121 ( .A1(n1035), .A2(n1034), .ZN(n1037) );
  XNOR2_X1 U1122 ( .A(G21), .B(G1966), .ZN(n1036) );
  NOR2_X1 U1123 ( .A1(n1037), .A2(n1036), .ZN(n1038) );
  XNOR2_X1 U1124 ( .A(KEYINPUT127), .B(n1038), .ZN(n1039) );
  NOR2_X1 U1125 ( .A1(n1040), .A2(n1039), .ZN(n1041) );
  XNOR2_X1 U1126 ( .A(KEYINPUT61), .B(n1041), .ZN(n1042) );
  NAND2_X1 U1127 ( .A1(n1043), .A2(n1042), .ZN(n1044) );
  NAND2_X1 U1128 ( .A1(n1045), .A2(n1044), .ZN(n1046) );
  NOR2_X1 U1129 ( .A1(n1047), .A2(n1046), .ZN(n1048) );
  NAND2_X1 U1130 ( .A1(n1049), .A2(n1048), .ZN(n1050) );
  XOR2_X1 U1131 ( .A(KEYINPUT62), .B(n1050), .Z(G311) );
  INV_X1 U1132 ( .A(G311), .ZN(G150) );
endmodule

