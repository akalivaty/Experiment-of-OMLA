//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 1 0 0 0 0 0 1 1 0 0 0 0 1 0 0 0 1 1 1 1 1 0 0 0 1 0 0 1 1 0 1 0 0 1 0 1 0 0 0 0 1 1 0 1 1 0 0 0 0 0 1 0 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n696,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n735, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n829, new_n830, new_n831, new_n832, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n905, new_n906, new_n908, new_n909, new_n910,
    new_n911, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n930, new_n931, new_n932, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n962, new_n963;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  INV_X1    g002(.A(G169gat), .ZN(new_n204));
  INV_X1    g003(.A(G176gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NOR2_X1   g005(.A1(G169gat), .A2(G176gat), .ZN(new_n207));
  NOR3_X1   g006(.A1(new_n206), .A2(KEYINPUT26), .A3(new_n207), .ZN(new_n208));
  AOI211_X1 g007(.A(new_n203), .B(new_n208), .C1(KEYINPUT26), .C2(new_n207), .ZN(new_n209));
  XNOR2_X1  g008(.A(KEYINPUT27), .B(G183gat), .ZN(new_n210));
  INV_X1    g009(.A(G190gat), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT64), .ZN(new_n212));
  AOI22_X1  g011(.A1(new_n210), .A2(new_n211), .B1(new_n212), .B2(KEYINPUT28), .ZN(new_n213));
  OR3_X1    g012(.A1(new_n213), .A2(new_n212), .A3(KEYINPUT28), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n213), .B1(new_n212), .B2(KEYINPUT28), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n209), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n207), .A2(KEYINPUT23), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n217), .A2(new_n206), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT24), .ZN(new_n219));
  AOI22_X1  g018(.A1(new_n203), .A2(new_n219), .B1(new_n207), .B2(KEYINPUT23), .ZN(new_n220));
  INV_X1    g019(.A(G183gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(new_n211), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n222), .A2(KEYINPUT24), .A3(new_n202), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n218), .A2(new_n220), .A3(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT25), .ZN(new_n225));
  XNOR2_X1  g024(.A(new_n224), .B(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n216), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(G226gat), .ZN(new_n228));
  INV_X1    g027(.A(G233gat), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n227), .A2(new_n230), .ZN(new_n231));
  AOI21_X1  g030(.A(KEYINPUT29), .B1(new_n216), .B2(new_n226), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n231), .B1(new_n230), .B2(new_n232), .ZN(new_n233));
  XNOR2_X1  g032(.A(KEYINPUT72), .B(G197gat), .ZN(new_n234));
  INV_X1    g033(.A(G204gat), .ZN(new_n235));
  AND2_X1   g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n234), .A2(new_n235), .ZN(new_n237));
  INV_X1    g036(.A(G211gat), .ZN(new_n238));
  INV_X1    g037(.A(G218gat), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  OAI22_X1  g039(.A1(new_n236), .A2(new_n237), .B1(KEYINPUT22), .B2(new_n240), .ZN(new_n241));
  XOR2_X1   g040(.A(G211gat), .B(G218gat), .Z(new_n242));
  AND2_X1   g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NOR2_X1   g042(.A1(new_n241), .A2(new_n242), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(KEYINPUT73), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n241), .B(new_n242), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT73), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n246), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n233), .A2(new_n250), .ZN(new_n251));
  XNOR2_X1  g050(.A(G8gat), .B(G36gat), .ZN(new_n252));
  XNOR2_X1  g051(.A(G64gat), .B(G92gat), .ZN(new_n253));
  XOR2_X1   g052(.A(new_n252), .B(new_n253), .Z(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  OAI211_X1 g054(.A(new_n231), .B(new_n245), .C1(new_n230), .C2(new_n232), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n251), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(KEYINPUT30), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n255), .B1(new_n251), .B2(new_n256), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  AOI211_X1 g059(.A(KEYINPUT30), .B(new_n255), .C1(new_n251), .C2(new_n256), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT39), .ZN(new_n263));
  INV_X1    g062(.A(G155gat), .ZN(new_n264));
  INV_X1    g063(.A(G162gat), .ZN(new_n265));
  OAI21_X1  g064(.A(KEYINPUT2), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n266), .B(KEYINPUT75), .ZN(new_n267));
  XNOR2_X1  g066(.A(G155gat), .B(G162gat), .ZN(new_n268));
  XNOR2_X1  g067(.A(G141gat), .B(G148gat), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT74), .ZN(new_n270));
  OR2_X1    g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n269), .A2(new_n270), .ZN(new_n272));
  NAND4_X1  g071(.A1(new_n267), .A2(new_n268), .A3(new_n271), .A4(new_n272), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n269), .A2(KEYINPUT2), .ZN(new_n274));
  OR2_X1    g073(.A1(new_n274), .A2(new_n268), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(G113gat), .ZN(new_n277));
  INV_X1    g076(.A(G120gat), .ZN(new_n278));
  AOI21_X1  g077(.A(KEYINPUT1), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n279), .B1(new_n277), .B2(new_n278), .ZN(new_n280));
  XOR2_X1   g079(.A(G127gat), .B(G134gat), .Z(new_n281));
  OR2_X1    g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n280), .A2(new_n281), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n276), .B(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(G225gat), .A2(G233gat), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT80), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n263), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n276), .A2(KEYINPUT3), .ZN(new_n291));
  XOR2_X1   g090(.A(KEYINPUT76), .B(KEYINPUT3), .Z(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  OAI211_X1 g092(.A(new_n291), .B(new_n284), .C1(new_n276), .C2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT4), .ZN(new_n295));
  OR3_X1    g094(.A1(new_n276), .A2(new_n295), .A3(new_n284), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT65), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n284), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n282), .A2(KEYINPUT65), .A3(new_n283), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n295), .B1(new_n300), .B2(new_n276), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n294), .A2(new_n296), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(new_n287), .ZN(new_n303));
  OAI211_X1 g102(.A(new_n290), .B(new_n303), .C1(new_n289), .C2(new_n288), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n302), .A2(new_n263), .A3(new_n287), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT79), .ZN(new_n306));
  XNOR2_X1  g105(.A(G1gat), .B(G29gat), .ZN(new_n307));
  XNOR2_X1  g106(.A(new_n307), .B(KEYINPUT0), .ZN(new_n308));
  XNOR2_X1  g107(.A(G57gat), .B(G85gat), .ZN(new_n309));
  XOR2_X1   g108(.A(new_n308), .B(new_n309), .Z(new_n310));
  AND3_X1   g109(.A1(new_n305), .A2(new_n306), .A3(new_n310), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n306), .B1(new_n305), .B2(new_n310), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n304), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT40), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(new_n276), .ZN(new_n316));
  NAND4_X1  g115(.A1(new_n316), .A2(KEYINPUT4), .A3(new_n298), .A4(new_n299), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n295), .B1(new_n276), .B2(new_n284), .ZN(new_n318));
  NAND4_X1  g117(.A1(new_n294), .A2(new_n317), .A3(new_n318), .A4(new_n286), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT5), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n320), .B1(new_n285), .B2(new_n287), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n287), .A2(KEYINPUT5), .ZN(new_n323));
  NAND4_X1  g122(.A1(new_n294), .A2(new_n301), .A3(new_n296), .A4(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT81), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n310), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n322), .A2(KEYINPUT81), .A3(new_n324), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  OAI211_X1 g128(.A(KEYINPUT40), .B(new_n304), .C1(new_n311), .C2(new_n312), .ZN(new_n330));
  NAND4_X1  g129(.A1(new_n262), .A2(new_n315), .A3(new_n329), .A4(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT82), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n261), .ZN(new_n334));
  INV_X1    g133(.A(new_n259), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n335), .A2(KEYINPUT30), .A3(new_n257), .ZN(new_n336));
  AND3_X1   g135(.A1(new_n329), .A2(new_n334), .A3(new_n336), .ZN(new_n337));
  NAND4_X1  g136(.A1(new_n337), .A2(KEYINPUT82), .A3(new_n330), .A4(new_n315), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n333), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT29), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n340), .B1(new_n243), .B2(new_n244), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n291), .B1(new_n341), .B2(new_n316), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT77), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  OAI211_X1 g143(.A(KEYINPUT77), .B(new_n291), .C1(new_n341), .C2(new_n316), .ZN(new_n345));
  INV_X1    g144(.A(G228gat), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n346), .A2(new_n229), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n340), .B1(new_n276), .B2(new_n293), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n246), .A2(new_n249), .A3(new_n348), .ZN(new_n349));
  NAND4_X1  g148(.A1(new_n344), .A2(new_n345), .A3(new_n347), .A4(new_n349), .ZN(new_n350));
  AND2_X1   g149(.A1(new_n348), .A2(new_n245), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n316), .B1(new_n341), .B2(new_n292), .ZN(new_n352));
  OAI22_X1  g151(.A1(new_n351), .A2(new_n352), .B1(new_n346), .B2(new_n229), .ZN(new_n353));
  INV_X1    g152(.A(G22gat), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n350), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(KEYINPUT78), .ZN(new_n356));
  XNOR2_X1  g155(.A(G78gat), .B(G106gat), .ZN(new_n357));
  XNOR2_X1  g156(.A(KEYINPUT31), .B(G50gat), .ZN(new_n358));
  XNOR2_X1  g157(.A(new_n357), .B(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n356), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n350), .A2(new_n353), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(G22gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(new_n355), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n360), .A2(new_n363), .ZN(new_n364));
  NAND4_X1  g163(.A1(new_n356), .A2(new_n362), .A3(new_n355), .A4(new_n359), .ZN(new_n365));
  AND2_X1   g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  OR2_X1    g165(.A1(new_n254), .A2(KEYINPUT38), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT37), .ZN(new_n368));
  INV_X1    g167(.A(new_n233), .ZN(new_n369));
  INV_X1    g168(.A(new_n250), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n368), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n233), .A2(new_n247), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n367), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n251), .A2(new_n256), .ZN(new_n374));
  AOI21_X1  g173(.A(KEYINPUT83), .B1(new_n374), .B2(new_n368), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT83), .ZN(new_n376));
  AOI211_X1 g175(.A(new_n376), .B(KEYINPUT37), .C1(new_n251), .C2(new_n256), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n373), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(new_n335), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n310), .B1(new_n322), .B2(new_n324), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(KEYINPUT6), .ZN(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n322), .A2(new_n310), .A3(new_n324), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT6), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n385), .B1(new_n327), .B2(new_n328), .ZN(new_n386));
  NOR3_X1   g185(.A1(new_n379), .A2(new_n382), .A3(new_n386), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n255), .B1(new_n374), .B2(new_n368), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT84), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n390), .B1(new_n375), .B2(new_n377), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n388), .A2(new_n389), .ZN(new_n392));
  OAI21_X1  g191(.A(KEYINPUT38), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n366), .B1(new_n387), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n339), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT36), .ZN(new_n396));
  XOR2_X1   g195(.A(G15gat), .B(G43gat), .Z(new_n397));
  XNOR2_X1  g196(.A(new_n397), .B(KEYINPUT68), .ZN(new_n398));
  XOR2_X1   g197(.A(G71gat), .B(G99gat), .Z(new_n399));
  XNOR2_X1  g198(.A(new_n398), .B(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(G227gat), .A2(G233gat), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  NAND4_X1  g201(.A1(new_n216), .A2(new_n226), .A3(new_n298), .A4(new_n299), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  AOI22_X1  g203(.A1(new_n216), .A2(new_n226), .B1(new_n298), .B2(new_n299), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n402), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  XNOR2_X1  g205(.A(KEYINPUT66), .B(KEYINPUT33), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n400), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT67), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n227), .A2(new_n300), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n401), .B1(new_n410), .B2(new_n403), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT32), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n409), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n406), .A2(KEYINPUT67), .A3(KEYINPUT32), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n408), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n410), .A2(new_n401), .A3(new_n403), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT70), .ZN(new_n417));
  AND3_X1   g216(.A1(new_n416), .A2(new_n417), .A3(KEYINPUT34), .ZN(new_n418));
  AOI21_X1  g217(.A(KEYINPUT34), .B1(new_n416), .B2(new_n417), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  AND2_X1   g219(.A1(new_n400), .A2(KEYINPUT69), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n400), .A2(KEYINPUT69), .ZN(new_n422));
  OR3_X1    g221(.A1(new_n421), .A2(new_n422), .A3(new_n407), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n423), .A2(KEYINPUT32), .A3(new_n406), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n415), .A2(new_n420), .A3(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT71), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n420), .B1(new_n415), .B2(new_n424), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  AOI211_X1 g228(.A(new_n426), .B(new_n420), .C1(new_n424), .C2(new_n415), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n396), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n425), .ZN(new_n432));
  OAI21_X1  g231(.A(KEYINPUT36), .B1(new_n432), .B2(new_n428), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n381), .B1(new_n385), .B2(new_n380), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  OAI211_X1 g234(.A(new_n365), .B(new_n364), .C1(new_n435), .C2(new_n262), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n431), .A2(new_n433), .A3(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n364), .A2(new_n365), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n336), .A2(new_n334), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n432), .A2(new_n428), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n439), .A2(new_n434), .A3(new_n440), .A4(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(KEYINPUT35), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n440), .B1(new_n386), .B2(new_n382), .ZN(new_n444));
  AOI21_X1  g243(.A(KEYINPUT35), .B1(new_n444), .B2(KEYINPUT85), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n415), .A2(new_n424), .ZN(new_n446));
  INV_X1    g245(.A(new_n420), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n448), .A2(new_n426), .A3(new_n425), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n427), .A2(new_n428), .ZN(new_n450));
  AOI22_X1  g249(.A1(new_n449), .A2(new_n450), .B1(new_n365), .B2(new_n364), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT85), .ZN(new_n452));
  OAI211_X1 g251(.A(new_n440), .B(new_n452), .C1(new_n386), .C2(new_n382), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n445), .A2(new_n451), .A3(new_n453), .ZN(new_n454));
  AOI22_X1  g253(.A1(new_n395), .A2(new_n438), .B1(new_n443), .B2(new_n454), .ZN(new_n455));
  XNOR2_X1  g254(.A(G113gat), .B(G141gat), .ZN(new_n456));
  XNOR2_X1  g255(.A(new_n456), .B(G197gat), .ZN(new_n457));
  XOR2_X1   g256(.A(KEYINPUT11), .B(G169gat), .Z(new_n458));
  XNOR2_X1  g257(.A(new_n457), .B(new_n458), .ZN(new_n459));
  XNOR2_X1  g258(.A(new_n459), .B(KEYINPUT12), .ZN(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(G229gat), .A2(G233gat), .ZN(new_n462));
  XNOR2_X1  g261(.A(G43gat), .B(G50gat), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(KEYINPUT15), .ZN(new_n464));
  XNOR2_X1  g263(.A(KEYINPUT86), .B(G43gat), .ZN(new_n465));
  INV_X1    g264(.A(G50gat), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  XNOR2_X1  g266(.A(KEYINPUT87), .B(G50gat), .ZN(new_n468));
  INV_X1    g267(.A(G43gat), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(KEYINPUT15), .B1(new_n467), .B2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT14), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n472), .A2(G29gat), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(G36gat), .ZN(new_n474));
  INV_X1    g273(.A(G36gat), .ZN(new_n475));
  INV_X1    g274(.A(G29gat), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n475), .B1(new_n476), .B2(KEYINPUT14), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n474), .B1(new_n477), .B2(new_n473), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n464), .B1(new_n471), .B2(new_n479), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n478), .A2(KEYINPUT15), .A3(new_n463), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n354), .A2(G15gat), .ZN(new_n484));
  INV_X1    g283(.A(G15gat), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(G22gat), .ZN(new_n486));
  INV_X1    g285(.A(G1gat), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(KEYINPUT16), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n484), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(new_n489), .ZN(new_n490));
  AOI21_X1  g289(.A(G1gat), .B1(new_n484), .B2(new_n486), .ZN(new_n491));
  XOR2_X1   g290(.A(KEYINPUT90), .B(G8gat), .Z(new_n492));
  NOR3_X1   g291(.A1(new_n490), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(G8gat), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT88), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n495), .B1(new_n491), .B2(new_n496), .ZN(new_n497));
  XNOR2_X1  g296(.A(G15gat), .B(G22gat), .ZN(new_n498));
  OAI211_X1 g297(.A(new_n489), .B(KEYINPUT88), .C1(G1gat), .C2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT89), .ZN(new_n500));
  AND3_X1   g299(.A1(new_n497), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n500), .B1(new_n497), .B2(new_n499), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n494), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT91), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT17), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n483), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n480), .A2(new_n506), .A3(new_n481), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n503), .B1(new_n504), .B2(new_n508), .ZN(new_n509));
  OAI211_X1 g308(.A(KEYINPUT18), .B(new_n462), .C1(new_n507), .C2(new_n509), .ZN(new_n510));
  XOR2_X1   g309(.A(new_n462), .B(KEYINPUT13), .Z(new_n511));
  NOR2_X1   g310(.A1(new_n483), .A2(new_n503), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n497), .A2(new_n499), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(KEYINPUT89), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n497), .A2(new_n499), .A3(new_n500), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n493), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n516), .A2(new_n482), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n511), .B1(new_n512), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n510), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g318(.A(KEYINPUT17), .B1(new_n503), .B2(new_n504), .ZN(new_n520));
  AND2_X1   g319(.A1(new_n508), .A2(new_n504), .ZN(new_n521));
  OAI22_X1  g320(.A1(new_n483), .A2(new_n520), .B1(new_n521), .B2(new_n503), .ZN(new_n522));
  AOI21_X1  g321(.A(KEYINPUT18), .B1(new_n522), .B2(new_n462), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n461), .B1(new_n519), .B2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT92), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT18), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n506), .B1(new_n516), .B2(KEYINPUT91), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n509), .B1(new_n482), .B2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(new_n462), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n526), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND4_X1  g329(.A1(new_n530), .A2(new_n460), .A3(new_n510), .A4(new_n518), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n524), .A2(new_n525), .A3(new_n531), .ZN(new_n532));
  OAI211_X1 g331(.A(KEYINPUT92), .B(new_n461), .C1(new_n519), .C2(new_n523), .ZN(new_n533));
  AND3_X1   g332(.A1(new_n532), .A2(KEYINPUT93), .A3(new_n533), .ZN(new_n534));
  AOI21_X1  g333(.A(KEYINPUT93), .B1(new_n532), .B2(new_n533), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n455), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(G99gat), .A2(G106gat), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT96), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(KEYINPUT96), .A2(G99gat), .A3(G106gat), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n540), .A2(KEYINPUT8), .A3(new_n541), .ZN(new_n542));
  OR2_X1    g341(.A1(KEYINPUT97), .A2(G85gat), .ZN(new_n543));
  INV_X1    g342(.A(G92gat), .ZN(new_n544));
  NAND2_X1  g343(.A1(KEYINPUT97), .A2(G85gat), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(G85gat), .A2(G92gat), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(KEYINPUT7), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT7), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n549), .A2(G85gat), .A3(G92gat), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n542), .A2(new_n546), .A3(new_n551), .ZN(new_n552));
  XOR2_X1   g351(.A(G99gat), .B(G106gat), .Z(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(KEYINPUT98), .ZN(new_n555));
  OAI21_X1  g354(.A(KEYINPUT94), .B1(G71gat), .B2(G78gat), .ZN(new_n556));
  XNOR2_X1  g355(.A(G57gat), .B(G64gat), .ZN(new_n557));
  AOI21_X1  g356(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(G71gat), .B(G78gat), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  OAI211_X1 g361(.A(new_n560), .B(new_n556), .C1(new_n557), .C2(new_n558), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AND3_X1   g363(.A1(new_n542), .A2(new_n546), .A3(new_n551), .ZN(new_n565));
  INV_X1    g364(.A(new_n553), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT98), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n552), .A2(new_n568), .A3(new_n553), .ZN(new_n569));
  NAND4_X1  g368(.A1(new_n555), .A2(new_n564), .A3(new_n567), .A4(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT99), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT10), .ZN(new_n573));
  AOI22_X1  g372(.A1(new_n562), .A2(new_n563), .B1(new_n565), .B2(new_n566), .ZN(new_n574));
  NAND4_X1  g373(.A1(new_n574), .A2(KEYINPUT99), .A3(new_n569), .A4(new_n555), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n567), .A2(new_n554), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n576), .A2(new_n562), .A3(new_n563), .ZN(new_n577));
  NAND4_X1  g376(.A1(new_n572), .A2(new_n573), .A3(new_n575), .A4(new_n577), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n564), .A2(new_n567), .A3(KEYINPUT10), .A4(new_n554), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(G230gat), .A2(G233gat), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  AND2_X1   g381(.A1(new_n575), .A2(new_n577), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n583), .A2(new_n572), .ZN(new_n584));
  INV_X1    g383(.A(new_n581), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(G120gat), .B(G148gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(G176gat), .B(G204gat), .ZN(new_n588));
  XOR2_X1   g387(.A(new_n587), .B(new_n588), .Z(new_n589));
  NAND3_X1  g388(.A1(new_n582), .A2(new_n586), .A3(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT100), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND4_X1  g391(.A1(new_n582), .A2(KEYINPUT100), .A3(new_n586), .A4(new_n589), .ZN(new_n593));
  INV_X1    g392(.A(new_n589), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n585), .B1(new_n578), .B2(new_n579), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n581), .B1(new_n583), .B2(new_n572), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n594), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT101), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  OAI211_X1 g398(.A(KEYINPUT101), .B(new_n594), .C1(new_n595), .C2(new_n596), .ZN(new_n600));
  AOI22_X1  g399(.A1(new_n592), .A2(new_n593), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(new_n264), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT95), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n564), .A2(KEYINPUT21), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n605), .B1(new_n516), .B2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n516), .A2(new_n605), .A3(new_n606), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n604), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n609), .ZN(new_n611));
  NOR3_X1   g410(.A1(new_n611), .A2(new_n607), .A3(new_n603), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(G183gat), .B(G211gat), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n564), .A2(KEYINPUT21), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(G231gat), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n617), .A2(new_n229), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n618), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n615), .A2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(G127gat), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n619), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n622), .B1(new_n619), .B2(new_n621), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n614), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n625), .ZN(new_n627));
  INV_X1    g426(.A(new_n614), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n627), .A2(new_n628), .A3(new_n623), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n613), .A2(new_n626), .A3(new_n629), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n628), .B1(new_n627), .B2(new_n623), .ZN(new_n631));
  NOR3_X1   g430(.A1(new_n624), .A2(new_n625), .A3(new_n614), .ZN(new_n632));
  OAI22_X1  g431(.A1(new_n631), .A2(new_n632), .B1(new_n612), .B2(new_n610), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n576), .A2(new_n506), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n483), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n482), .A2(new_n506), .A3(new_n576), .ZN(new_n636));
  AND2_X1   g435(.A1(G232gat), .A2(G233gat), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n637), .A2(KEYINPUT41), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n635), .A2(new_n636), .A3(new_n638), .ZN(new_n639));
  XOR2_X1   g438(.A(G190gat), .B(G218gat), .Z(new_n640));
  NOR2_X1   g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n637), .A2(KEYINPUT41), .ZN(new_n643));
  XNOR2_X1  g442(.A(G134gat), .B(G162gat), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n643), .B(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n639), .A2(new_n640), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n642), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n645), .ZN(new_n648));
  INV_X1    g447(.A(new_n646), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n648), .B1(new_n649), .B2(new_n641), .ZN(new_n650));
  AOI22_X1  g449(.A1(new_n630), .A2(new_n633), .B1(new_n647), .B2(new_n650), .ZN(new_n651));
  AND2_X1   g450(.A1(new_n601), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n537), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n653), .A2(new_n434), .ZN(new_n654));
  XOR2_X1   g453(.A(KEYINPUT102), .B(G1gat), .Z(new_n655));
  XNOR2_X1  g454(.A(new_n654), .B(new_n655), .ZN(G1324gat));
  OR3_X1    g455(.A1(new_n653), .A2(KEYINPUT103), .A3(new_n440), .ZN(new_n657));
  OAI21_X1  g456(.A(KEYINPUT103), .B1(new_n653), .B2(new_n440), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n657), .A2(G8gat), .A3(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n653), .ZN(new_n660));
  XOR2_X1   g459(.A(KEYINPUT16), .B(G8gat), .Z(new_n661));
  NAND4_X1  g460(.A1(new_n660), .A2(KEYINPUT42), .A3(new_n262), .A4(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n661), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n663), .B1(new_n657), .B2(new_n658), .ZN(new_n664));
  OAI211_X1 g463(.A(new_n659), .B(new_n662), .C1(new_n664), .C2(KEYINPUT42), .ZN(G1325gat));
  NAND2_X1  g464(.A1(new_n431), .A2(new_n433), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  OAI21_X1  g466(.A(G15gat), .B1(new_n653), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n449), .A2(new_n450), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n669), .A2(new_n485), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n668), .B1(new_n653), .B2(new_n670), .ZN(G1326gat));
  NAND2_X1  g470(.A1(new_n660), .A2(new_n366), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(KEYINPUT104), .ZN(new_n673));
  XNOR2_X1  g472(.A(KEYINPUT43), .B(G22gat), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n673), .B(new_n674), .ZN(G1327gat));
  NAND2_X1  g474(.A1(new_n630), .A2(new_n633), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n650), .A2(new_n647), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  AND3_X1   g477(.A1(new_n537), .A2(new_n601), .A3(new_n678), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n679), .A2(new_n476), .A3(new_n435), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n680), .B(KEYINPUT45), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT44), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n682), .B1(new_n455), .B2(new_n677), .ZN(new_n683));
  INV_X1    g482(.A(new_n677), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n437), .B1(new_n339), .B2(new_n394), .ZN(new_n685));
  AND3_X1   g484(.A1(new_n669), .A2(new_n439), .A3(new_n453), .ZN(new_n686));
  AOI22_X1  g485(.A1(new_n686), .A2(new_n445), .B1(new_n442), .B2(KEYINPUT35), .ZN(new_n687));
  OAI211_X1 g486(.A(KEYINPUT44), .B(new_n684), .C1(new_n685), .C2(new_n687), .ZN(new_n688));
  AND2_X1   g487(.A1(new_n683), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n532), .A2(new_n533), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n676), .ZN(new_n692));
  NAND4_X1  g491(.A1(new_n689), .A2(new_n691), .A3(new_n692), .A4(new_n601), .ZN(new_n693));
  OAI21_X1  g492(.A(G29gat), .B1(new_n693), .B2(new_n434), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n681), .A2(new_n694), .ZN(G1328gat));
  NAND3_X1  g494(.A1(new_n679), .A2(new_n475), .A3(new_n262), .ZN(new_n696));
  XOR2_X1   g495(.A(new_n696), .B(KEYINPUT46), .Z(new_n697));
  OAI21_X1  g496(.A(G36gat), .B1(new_n693), .B2(new_n440), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(G1329gat));
  OAI21_X1  g498(.A(new_n465), .B1(new_n693), .B2(new_n667), .ZN(new_n700));
  INV_X1    g499(.A(new_n669), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n701), .A2(new_n465), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT47), .ZN(new_n703));
  AOI22_X1  g502(.A1(new_n679), .A2(new_n702), .B1(KEYINPUT105), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n700), .A2(new_n704), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n703), .A2(KEYINPUT105), .ZN(new_n706));
  XOR2_X1   g505(.A(new_n705), .B(new_n706), .Z(G1330gat));
  OAI21_X1  g506(.A(new_n468), .B1(new_n693), .B2(new_n439), .ZN(new_n708));
  AOI21_X1  g507(.A(KEYINPUT48), .B1(new_n708), .B2(KEYINPUT106), .ZN(new_n709));
  INV_X1    g508(.A(new_n468), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n679), .A2(new_n366), .A3(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n708), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n709), .B(new_n712), .ZN(G1331gat));
  NOR2_X1   g512(.A1(new_n455), .A2(new_n691), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n592), .A2(new_n593), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n599), .A2(new_n600), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  AND2_X1   g516(.A1(new_n717), .A2(new_n651), .ZN(new_n718));
  AND2_X1   g517(.A1(new_n714), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(new_n435), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(G57gat), .ZN(G1332gat));
  INV_X1    g520(.A(new_n719), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n722), .A2(new_n440), .ZN(new_n723));
  NOR2_X1   g522(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n724));
  AND2_X1   g523(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n723), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n726), .B1(new_n723), .B2(new_n724), .ZN(G1333gat));
  NAND3_X1  g526(.A1(new_n719), .A2(G71gat), .A3(new_n666), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT107), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n728), .B(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(G71gat), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n731), .B1(new_n722), .B2(new_n701), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g533(.A1(new_n719), .A2(new_n366), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g535(.A1(new_n543), .A2(new_n545), .ZN(new_n737));
  NOR3_X1   g536(.A1(new_n691), .A2(new_n676), .A3(new_n601), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n689), .A2(new_n738), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n737), .B1(new_n739), .B2(new_n434), .ZN(new_n740));
  OAI211_X1 g539(.A(new_n690), .B(new_n678), .C1(new_n685), .C2(new_n687), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT51), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n741), .B(new_n742), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n601), .B1(new_n743), .B2(KEYINPUT108), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n744), .B1(KEYINPUT108), .B2(new_n743), .ZN(new_n745));
  OR2_X1    g544(.A1(new_n434), .A2(new_n737), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n740), .B1(new_n745), .B2(new_n746), .ZN(G1336gat));
  NOR3_X1   g546(.A1(new_n440), .A2(new_n601), .A3(G92gat), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n743), .A2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT52), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n683), .A2(new_n262), .A3(new_n688), .A4(new_n738), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(G92gat), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n749), .A2(new_n750), .A3(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT110), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n741), .A2(KEYINPUT109), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(new_n742), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n741), .A2(KEYINPUT109), .A3(KEYINPUT51), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n756), .A2(new_n757), .A3(new_n748), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(new_n752), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n754), .B1(new_n759), .B2(KEYINPUT52), .ZN(new_n760));
  AOI211_X1 g559(.A(KEYINPUT110), .B(new_n750), .C1(new_n758), .C2(new_n752), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n753), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT111), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  OAI211_X1 g563(.A(new_n753), .B(KEYINPUT111), .C1(new_n760), .C2(new_n761), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(G1337gat));
  OAI21_X1  g565(.A(G99gat), .B1(new_n739), .B2(new_n667), .ZN(new_n767));
  OR2_X1    g566(.A1(new_n701), .A2(G99gat), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n767), .B1(new_n745), .B2(new_n768), .ZN(G1338gat));
  NAND3_X1  g568(.A1(new_n689), .A2(new_n366), .A3(new_n738), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(G106gat), .ZN(new_n771));
  NOR3_X1   g570(.A1(new_n439), .A2(G106gat), .A3(new_n601), .ZN(new_n772));
  AOI21_X1  g571(.A(KEYINPUT53), .B1(new_n743), .B2(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n771), .A2(new_n773), .ZN(new_n774));
  AND2_X1   g573(.A1(new_n756), .A2(new_n757), .ZN(new_n775));
  AOI22_X1  g574(.A1(new_n775), .A2(new_n772), .B1(new_n770), .B2(G106gat), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT53), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n774), .B1(new_n776), .B2(new_n777), .ZN(G1339gat));
  NAND2_X1  g577(.A1(new_n652), .A2(new_n690), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT55), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n578), .A2(new_n585), .A3(new_n579), .ZN(new_n781));
  NAND4_X1  g580(.A1(new_n582), .A2(KEYINPUT112), .A3(KEYINPUT54), .A4(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT54), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n589), .B1(new_n595), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n595), .A2(new_n783), .ZN(new_n786));
  AOI21_X1  g585(.A(KEYINPUT112), .B1(new_n786), .B2(new_n781), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n780), .B1(new_n785), .B2(new_n787), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n582), .A2(KEYINPUT54), .A3(new_n781), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT112), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n791), .A2(KEYINPUT55), .A3(new_n782), .A4(new_n784), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n788), .A2(new_n715), .A3(new_n792), .ZN(new_n793));
  OR2_X1    g592(.A1(new_n512), .A2(new_n517), .ZN(new_n794));
  OAI22_X1  g593(.A1(new_n462), .A2(new_n522), .B1(new_n794), .B2(new_n511), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(new_n459), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n531), .A2(new_n796), .ZN(new_n797));
  NOR3_X1   g596(.A1(new_n793), .A2(new_n677), .A3(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT113), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n799), .B1(new_n601), .B2(new_n797), .ZN(new_n800));
  INV_X1    g599(.A(new_n797), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n717), .A2(KEYINPUT113), .A3(new_n801), .ZN(new_n802));
  OAI211_X1 g601(.A(new_n800), .B(new_n802), .C1(new_n793), .C2(new_n690), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n798), .B1(new_n803), .B2(new_n677), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n779), .B1(new_n804), .B2(new_n676), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(KEYINPUT114), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT114), .ZN(new_n807));
  OAI211_X1 g606(.A(new_n807), .B(new_n779), .C1(new_n804), .C2(new_n676), .ZN(new_n808));
  AND2_X1   g607(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n809), .A2(new_n435), .A3(new_n439), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT115), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n669), .A2(new_n440), .ZN(new_n812));
  OR3_X1    g611(.A1(new_n810), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(new_n536), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n811), .B1(new_n810), .B2(new_n812), .ZN(new_n815));
  AND4_X1   g614(.A1(G113gat), .A2(new_n813), .A3(new_n814), .A4(new_n815), .ZN(new_n816));
  AND2_X1   g615(.A1(new_n809), .A2(new_n435), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n817), .A2(new_n439), .A3(new_n441), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n818), .A2(new_n262), .ZN(new_n819));
  AOI21_X1  g618(.A(G113gat), .B1(new_n819), .B2(new_n691), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n816), .A2(new_n820), .ZN(G1340gat));
  NAND4_X1  g620(.A1(new_n813), .A2(G120gat), .A3(new_n717), .A4(new_n815), .ZN(new_n822));
  NOR3_X1   g621(.A1(new_n818), .A2(new_n262), .A3(new_n601), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n822), .B1(G120gat), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(KEYINPUT116), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT116), .ZN(new_n826));
  OAI211_X1 g625(.A(new_n822), .B(new_n826), .C1(G120gat), .C2(new_n823), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n825), .A2(new_n827), .ZN(G1341gat));
  NAND4_X1  g627(.A1(new_n813), .A2(G127gat), .A3(new_n676), .A4(new_n815), .ZN(new_n829));
  AND2_X1   g628(.A1(new_n829), .A2(KEYINPUT117), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n829), .A2(KEYINPUT117), .ZN(new_n831));
  AOI21_X1  g630(.A(G127gat), .B1(new_n819), .B2(new_n676), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n830), .A2(new_n831), .A3(new_n832), .ZN(G1342gat));
  OR3_X1    g632(.A1(new_n262), .A2(G134gat), .A3(new_n677), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT118), .ZN(new_n835));
  OAI22_X1  g634(.A1(new_n818), .A2(new_n834), .B1(new_n835), .B2(KEYINPUT56), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT56), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n836), .B1(KEYINPUT118), .B2(new_n837), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n813), .A2(new_n684), .A3(new_n815), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(G134gat), .ZN(new_n840));
  OAI211_X1 g639(.A(new_n835), .B(KEYINPUT56), .C1(new_n818), .C2(new_n834), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n838), .A2(new_n840), .A3(new_n841), .ZN(G1343gat));
  NAND2_X1  g641(.A1(new_n667), .A2(new_n366), .ZN(new_n843));
  XNOR2_X1  g642(.A(new_n843), .B(KEYINPUT120), .ZN(new_n844));
  AND3_X1   g643(.A1(new_n817), .A2(new_n440), .A3(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(G141gat), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n845), .A2(new_n846), .A3(new_n814), .ZN(new_n847));
  NOR3_X1   g646(.A1(new_n666), .A2(new_n434), .A3(new_n262), .ZN(new_n848));
  INV_X1    g647(.A(new_n848), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n806), .A2(new_n366), .A3(new_n808), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT57), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT93), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n690), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n532), .A2(KEYINPUT93), .A3(new_n533), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n793), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n601), .A2(new_n797), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n677), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT119), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n798), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  AND3_X1   g659(.A1(new_n788), .A2(new_n715), .A3(new_n792), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n861), .B1(new_n534), .B2(new_n535), .ZN(new_n862));
  INV_X1    g661(.A(new_n857), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n684), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(KEYINPUT119), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n676), .B1(new_n860), .B2(new_n865), .ZN(new_n866));
  INV_X1    g665(.A(new_n779), .ZN(new_n867));
  OAI211_X1 g666(.A(KEYINPUT57), .B(new_n366), .C1(new_n866), .C2(new_n867), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n849), .B1(new_n852), .B2(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(new_n869), .ZN(new_n870));
  OAI21_X1  g669(.A(G141gat), .B1(new_n870), .B2(new_n536), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT58), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n847), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  OAI21_X1  g672(.A(G141gat), .B1(new_n870), .B2(new_n690), .ZN(new_n874));
  AND2_X1   g673(.A1(new_n847), .A2(new_n874), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n873), .B1(new_n875), .B2(new_n872), .ZN(G1344gat));
  INV_X1    g675(.A(G148gat), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n845), .A2(new_n877), .A3(new_n717), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT59), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT121), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n880), .B1(new_n536), .B2(new_n652), .ZN(new_n881));
  AND4_X1   g680(.A1(new_n880), .A2(new_n854), .A3(new_n652), .A4(new_n855), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(new_n798), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n858), .A2(new_n884), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n883), .B1(new_n885), .B2(new_n692), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT122), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n439), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n692), .B1(new_n864), .B2(new_n798), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n854), .A2(new_n652), .A3(new_n855), .ZN(new_n890));
  XNOR2_X1  g689(.A(new_n890), .B(KEYINPUT121), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n887), .B1(new_n889), .B2(new_n891), .ZN(new_n892));
  INV_X1    g691(.A(new_n892), .ZN(new_n893));
  AOI21_X1  g692(.A(KEYINPUT57), .B1(new_n888), .B2(new_n893), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n806), .A2(KEYINPUT57), .A3(new_n366), .A4(new_n808), .ZN(new_n895));
  INV_X1    g694(.A(new_n895), .ZN(new_n896));
  OAI211_X1 g695(.A(new_n717), .B(new_n848), .C1(new_n894), .C2(new_n896), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n879), .B1(new_n897), .B2(G148gat), .ZN(new_n898));
  AOI211_X1 g697(.A(KEYINPUT59), .B(new_n877), .C1(new_n869), .C2(new_n717), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n878), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(KEYINPUT123), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT123), .ZN(new_n902));
  OAI211_X1 g701(.A(new_n878), .B(new_n902), .C1(new_n898), .C2(new_n899), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n901), .A2(new_n903), .ZN(G1345gat));
  NAND3_X1  g703(.A1(new_n845), .A2(new_n264), .A3(new_n676), .ZN(new_n905));
  OAI21_X1  g704(.A(G155gat), .B1(new_n870), .B2(new_n692), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(new_n906), .ZN(G1346gat));
  NOR3_X1   g706(.A1(new_n262), .A2(G162gat), .A3(new_n677), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n817), .A2(new_n844), .A3(new_n908), .ZN(new_n909));
  XNOR2_X1  g708(.A(new_n909), .B(KEYINPUT124), .ZN(new_n910));
  OAI21_X1  g709(.A(G162gat), .B1(new_n870), .B2(new_n677), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(G1347gat));
  NOR2_X1   g711(.A1(new_n435), .A2(new_n440), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n809), .A2(new_n451), .A3(new_n913), .ZN(new_n914));
  NOR3_X1   g713(.A1(new_n914), .A2(new_n204), .A3(new_n536), .ZN(new_n915));
  AND4_X1   g714(.A1(new_n439), .A2(new_n809), .A3(new_n441), .A4(new_n913), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(new_n691), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n915), .B1(new_n917), .B2(new_n204), .ZN(G1348gat));
  NAND3_X1  g717(.A1(new_n916), .A2(new_n205), .A3(new_n717), .ZN(new_n919));
  OAI21_X1  g718(.A(G176gat), .B1(new_n914), .B2(new_n601), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  XOR2_X1   g720(.A(new_n921), .B(KEYINPUT125), .Z(G1349gat));
  AND2_X1   g721(.A1(new_n676), .A2(new_n210), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT126), .ZN(new_n924));
  AOI22_X1  g723(.A1(new_n916), .A2(new_n923), .B1(new_n924), .B2(KEYINPUT60), .ZN(new_n925));
  OAI21_X1  g724(.A(G183gat), .B1(new_n914), .B2(new_n692), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n924), .A2(KEYINPUT60), .ZN(new_n928));
  XOR2_X1   g727(.A(new_n927), .B(new_n928), .Z(G1350gat));
  OAI21_X1  g728(.A(G190gat), .B1(new_n914), .B2(new_n677), .ZN(new_n930));
  XNOR2_X1  g729(.A(new_n930), .B(KEYINPUT61), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n916), .A2(new_n211), .A3(new_n684), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(G1351gat));
  NAND2_X1  g732(.A1(new_n667), .A2(new_n913), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n850), .A2(new_n934), .ZN(new_n935));
  AOI21_X1  g734(.A(G197gat), .B1(new_n935), .B2(new_n691), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n862), .A2(new_n863), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n798), .B1(new_n937), .B2(new_n677), .ZN(new_n938));
  OAI211_X1 g737(.A(new_n887), .B(new_n891), .C1(new_n938), .C2(new_n676), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n939), .A2(new_n366), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n851), .B1(new_n940), .B2(new_n892), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n934), .B1(new_n941), .B2(new_n895), .ZN(new_n942));
  AND2_X1   g741(.A1(new_n814), .A2(G197gat), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n936), .B1(new_n942), .B2(new_n943), .ZN(G1352gat));
  INV_X1    g743(.A(new_n935), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n717), .A2(new_n235), .ZN(new_n946));
  OR3_X1    g745(.A1(new_n945), .A2(KEYINPUT62), .A3(new_n946), .ZN(new_n947));
  OAI21_X1  g746(.A(KEYINPUT62), .B1(new_n945), .B2(new_n946), .ZN(new_n948));
  AOI211_X1 g747(.A(new_n601), .B(new_n934), .C1(new_n941), .C2(new_n895), .ZN(new_n949));
  OAI211_X1 g748(.A(new_n947), .B(new_n948), .C1(new_n235), .C2(new_n949), .ZN(G1353gat));
  NAND3_X1  g749(.A1(new_n935), .A2(new_n238), .A3(new_n676), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT63), .ZN(new_n952));
  AOI211_X1 g751(.A(new_n952), .B(new_n238), .C1(new_n942), .C2(new_n676), .ZN(new_n953));
  INV_X1    g752(.A(new_n934), .ZN(new_n954));
  OAI211_X1 g753(.A(new_n676), .B(new_n954), .C1(new_n894), .C2(new_n896), .ZN(new_n955));
  AOI21_X1  g754(.A(KEYINPUT63), .B1(new_n955), .B2(G211gat), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n951), .B1(new_n953), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n957), .A2(KEYINPUT127), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT127), .ZN(new_n959));
  OAI211_X1 g758(.A(new_n959), .B(new_n951), .C1(new_n953), .C2(new_n956), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n958), .A2(new_n960), .ZN(G1354gat));
  NAND3_X1  g760(.A1(new_n935), .A2(new_n239), .A3(new_n684), .ZN(new_n962));
  AND2_X1   g761(.A1(new_n942), .A2(new_n684), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n962), .B1(new_n963), .B2(new_n239), .ZN(G1355gat));
endmodule


