//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 0 0 1 1 1 0 0 0 1 0 1 0 1 1 1 0 1 0 0 1 0 1 0 0 0 1 0 0 0 1 0 1 1 1 0 1 1 1 0 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:41 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1248, new_n1249, new_n1250, new_n1251,
    new_n1252, new_n1253, new_n1254, new_n1255;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(new_n202));
  XOR2_X1   g0002(.A(new_n202), .B(KEYINPUT64), .Z(G355));
  NAND2_X1  g0003(.A1(G1), .A2(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G13), .ZN(new_n205));
  OAI211_X1 g0005(.A(new_n205), .B(G250), .C1(G257), .C2(G264), .ZN(new_n206));
  XOR2_X1   g0006(.A(new_n206), .B(KEYINPUT0), .Z(new_n207));
  INV_X1    g0007(.A(G50), .ZN(new_n208));
  INV_X1    g0008(.A(G226), .ZN(new_n209));
  INV_X1    g0009(.A(G68), .ZN(new_n210));
  INV_X1    g0010(.A(G238), .ZN(new_n211));
  OAI22_X1  g0011(.A1(new_n208), .A2(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT65), .ZN(new_n214));
  AOI211_X1 g0014(.A(new_n212), .B(new_n214), .C1(G77), .C2(G244), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G116), .A2(G270), .ZN(new_n216));
  INV_X1    g0016(.A(G58), .ZN(new_n217));
  INV_X1    g0017(.A(G232), .ZN(new_n218));
  OAI211_X1 g0018(.A(new_n215), .B(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(G107), .ZN(new_n220));
  INV_X1    g0020(.A(G264), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n204), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT1), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  INV_X1    g0025(.A(G20), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n217), .A2(new_n210), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n228), .A2(G50), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  AOI211_X1 g0030(.A(new_n207), .B(new_n224), .C1(new_n227), .C2(new_n230), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G226), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(new_n221), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G270), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n236), .B(new_n239), .Z(G358));
  XOR2_X1   g0040(.A(G68), .B(G77), .Z(new_n241));
  XNOR2_X1  g0041(.A(G50), .B(G58), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G107), .B(G116), .Z(new_n244));
  XNOR2_X1  g0044(.A(G87), .B(G97), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  INV_X1    g0047(.A(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n226), .A2(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(new_n249), .ZN(new_n250));
  NAND3_X1  g0050(.A1(new_n208), .A2(new_n217), .A3(new_n210), .ZN(new_n251));
  AOI22_X1  g0051(.A1(new_n250), .A2(G150), .B1(new_n251), .B2(G20), .ZN(new_n252));
  XNOR2_X1  g0052(.A(KEYINPUT8), .B(G58), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT69), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  OR3_X1    g0055(.A1(new_n254), .A2(new_n217), .A3(KEYINPUT8), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n226), .A2(G33), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n252), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  OAI21_X1  g0059(.A(KEYINPUT68), .B1(new_n204), .B2(new_n248), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT68), .ZN(new_n261));
  NAND4_X1  g0061(.A1(new_n261), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n260), .A2(new_n225), .A3(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G1), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G20), .ZN(new_n265));
  NAND4_X1  g0065(.A1(new_n260), .A2(new_n225), .A3(new_n265), .A4(new_n262), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  AOI22_X1  g0067(.A1(new_n259), .A2(new_n263), .B1(G50), .B2(new_n267), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n226), .A2(G1), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G13), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(new_n208), .ZN(new_n272));
  AND2_X1   g0072(.A1(new_n268), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT9), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n268), .A2(new_n272), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(KEYINPUT9), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n225), .B1(G33), .B2(G41), .ZN(new_n279));
  INV_X1    g0079(.A(G41), .ZN(new_n280));
  INV_X1    g0080(.A(G45), .ZN(new_n281));
  AOI21_X1  g0081(.A(G1), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(KEYINPUT67), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT67), .ZN(new_n284));
  NOR2_X1   g0084(.A1(G41), .A2(G45), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n284), .B1(new_n285), .B2(G1), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n279), .B1(new_n283), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(G226), .ZN(new_n288));
  XNOR2_X1  g0088(.A(KEYINPUT3), .B(G33), .ZN(new_n289));
  INV_X1    g0089(.A(G1698), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(G222), .ZN(new_n291));
  NAND2_X1  g0091(.A1(G223), .A2(G1698), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n289), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  OAI211_X1 g0093(.A(new_n293), .B(new_n279), .C1(G77), .C2(new_n289), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n282), .A2(G274), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n288), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(G200), .ZN(new_n297));
  INV_X1    g0097(.A(new_n296), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(G190), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n278), .A2(new_n297), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(KEYINPUT71), .A2(KEYINPUT10), .ZN(new_n301));
  OR2_X1    g0101(.A1(KEYINPUT71), .A2(KEYINPUT10), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n300), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  AOI22_X1  g0103(.A1(new_n275), .A2(new_n277), .B1(G190), .B2(new_n298), .ZN(new_n304));
  NAND4_X1  g0104(.A1(new_n304), .A2(KEYINPUT71), .A3(KEYINPUT10), .A4(new_n297), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n276), .B1(new_n298), .B2(G169), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT70), .ZN(new_n307));
  OR2_X1    g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n306), .A2(new_n307), .ZN(new_n309));
  OAI211_X1 g0109(.A(new_n308), .B(new_n309), .C1(G179), .C2(new_n296), .ZN(new_n310));
  NAND2_X1  g0110(.A1(G20), .A2(G77), .ZN(new_n311));
  XNOR2_X1  g0111(.A(KEYINPUT15), .B(G87), .ZN(new_n312));
  OAI221_X1 g0112(.A(new_n311), .B1(new_n253), .B2(new_n249), .C1(new_n258), .C2(new_n312), .ZN(new_n313));
  AOI22_X1  g0113(.A1(new_n313), .A2(new_n263), .B1(new_n267), .B2(G77), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n314), .B1(G77), .B2(new_n270), .ZN(new_n315));
  NAND2_X1  g0115(.A1(G238), .A2(G1698), .ZN(new_n316));
  OAI211_X1 g0116(.A(new_n289), .B(new_n316), .C1(new_n218), .C2(G1698), .ZN(new_n317));
  OAI211_X1 g0117(.A(new_n317), .B(new_n279), .C1(G107), .C2(new_n289), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n287), .A2(G244), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n318), .A2(new_n295), .A3(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n315), .B1(new_n321), .B2(G190), .ZN(new_n322));
  INV_X1    g0122(.A(G200), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n322), .B1(new_n323), .B2(new_n321), .ZN(new_n324));
  NAND4_X1  g0124(.A1(new_n303), .A2(new_n305), .A3(new_n310), .A4(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT75), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n326), .B1(new_n248), .B2(KEYINPUT3), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT3), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n328), .A2(KEYINPUT75), .A3(G33), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n248), .A2(KEYINPUT3), .ZN(new_n331));
  NAND4_X1  g0131(.A1(new_n330), .A2(G223), .A3(new_n290), .A4(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(KEYINPUT79), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n328), .A2(G33), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n334), .B1(new_n327), .B2(new_n329), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n209), .A2(new_n290), .ZN(new_n336));
  AOI22_X1  g0136(.A1(new_n335), .A2(new_n336), .B1(G33), .B2(G87), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT79), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n335), .A2(new_n338), .A3(G223), .A4(new_n290), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n333), .A2(new_n337), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(new_n279), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n287), .A2(G232), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(new_n295), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n341), .A2(G179), .A3(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(G169), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n343), .B1(new_n340), .B2(new_n279), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n345), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  AND3_X1   g0148(.A1(new_n328), .A2(KEYINPUT75), .A3(G33), .ZN(new_n349));
  AOI21_X1  g0149(.A(KEYINPUT75), .B1(new_n328), .B2(G33), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n331), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NOR2_X1   g0151(.A1(KEYINPUT76), .A2(KEYINPUT7), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n351), .A2(new_n226), .A3(new_n352), .ZN(new_n353));
  XOR2_X1   g0153(.A(KEYINPUT76), .B(KEYINPUT7), .Z(new_n354));
  OAI21_X1  g0154(.A(new_n354), .B1(new_n335), .B2(G20), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n353), .A2(new_n355), .A3(G68), .ZN(new_n356));
  NAND2_X1  g0156(.A1(G58), .A2(G68), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n226), .B1(new_n228), .B2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT77), .ZN(new_n360));
  INV_X1    g0160(.A(G159), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n249), .A2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n359), .A2(new_n360), .A3(new_n363), .ZN(new_n364));
  OAI21_X1  g0164(.A(KEYINPUT77), .B1(new_n358), .B2(new_n362), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n356), .A2(KEYINPUT16), .A3(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT16), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT7), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n369), .B1(new_n289), .B2(G20), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n328), .A2(G33), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(new_n331), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n372), .A2(KEYINPUT7), .A3(new_n226), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n210), .B1(new_n370), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n359), .A2(new_n363), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n368), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n367), .A2(new_n263), .A3(new_n376), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n255), .A2(new_n265), .A3(new_n256), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT78), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n270), .A2(new_n225), .A3(new_n260), .A4(new_n262), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n255), .A2(KEYINPUT78), .A3(new_n265), .A4(new_n256), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n380), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n257), .A2(new_n271), .ZN(new_n385));
  AND2_X1   g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n377), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n348), .A2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT18), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n348), .A2(KEYINPUT18), .A3(new_n387), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n390), .A2(KEYINPUT80), .A3(new_n391), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n347), .A2(new_n323), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n387), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT82), .ZN(new_n395));
  INV_X1    g0195(.A(G190), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(KEYINPUT81), .ZN(new_n397));
  OR2_X1    g0197(.A1(new_n396), .A2(KEYINPUT81), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n341), .A2(new_n397), .A3(new_n398), .A4(new_n344), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n394), .A2(new_n395), .A3(KEYINPUT17), .A4(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT17), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n341), .A2(new_n344), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(G200), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n403), .A2(new_n399), .A3(new_n377), .A4(new_n386), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n401), .B1(new_n404), .B2(KEYINPUT82), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT80), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n388), .A2(new_n406), .A3(new_n389), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n392), .A2(new_n400), .A3(new_n405), .A4(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(G97), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n248), .A2(new_n409), .ZN(new_n410));
  NOR2_X1   g0210(.A1(G226), .A2(G1698), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n411), .B1(new_n218), .B2(G1698), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n410), .B1(new_n412), .B2(new_n289), .ZN(new_n413));
  INV_X1    g0213(.A(new_n279), .ZN(new_n414));
  OR2_X1    g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT13), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n287), .A2(G238), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n415), .A2(new_n416), .A3(new_n417), .A4(new_n295), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n295), .B1(new_n413), .B2(new_n414), .ZN(new_n419));
  AOI211_X1 g0219(.A(new_n211), .B(new_n279), .C1(new_n283), .C2(new_n286), .ZN(new_n420));
  OAI21_X1  g0220(.A(KEYINPUT13), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n418), .A2(new_n421), .ZN(new_n422));
  OAI21_X1  g0222(.A(KEYINPUT72), .B1(new_n422), .B2(new_n396), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n226), .A2(G33), .A3(G77), .ZN(new_n424));
  OAI221_X1 g0224(.A(new_n424), .B1(new_n226), .B2(G68), .C1(new_n249), .C2(new_n208), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(new_n263), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(KEYINPUT73), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT73), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n425), .A2(new_n428), .A3(new_n263), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT11), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n271), .A2(KEYINPUT12), .A3(new_n210), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT12), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n434), .B1(new_n270), .B2(G68), .ZN(new_n435));
  OAI211_X1 g0235(.A(new_n433), .B(new_n435), .C1(new_n210), .C2(new_n266), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n427), .A2(KEYINPUT11), .A3(new_n429), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n432), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n422), .A2(G200), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT72), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n418), .A2(new_n421), .A3(new_n442), .A4(G190), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n423), .A2(new_n440), .A3(new_n441), .A4(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT74), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n439), .B1(G200), .B2(new_n422), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n447), .A2(KEYINPUT74), .A3(new_n423), .A4(new_n443), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n422), .A2(G169), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(KEYINPUT14), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT14), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n422), .A2(new_n452), .A3(G169), .ZN(new_n453));
  INV_X1    g0253(.A(G179), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n451), .B(new_n453), .C1(new_n454), .C2(new_n422), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(new_n439), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n449), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n321), .A2(new_n454), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n320), .A2(new_n346), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n458), .A2(new_n315), .A3(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  NOR4_X1   g0261(.A1(new_n325), .A2(new_n408), .A3(new_n457), .A4(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(G250), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(new_n290), .ZN(new_n464));
  INV_X1    g0264(.A(G257), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(G1698), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n330), .A2(new_n331), .A3(new_n464), .A4(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(G33), .A2(G294), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(new_n279), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT86), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT5), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT84), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n473), .B1(new_n474), .B2(G41), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n280), .A2(KEYINPUT84), .A3(KEYINPUT5), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n281), .A2(G1), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n475), .A2(new_n476), .A3(new_n477), .A4(G274), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n475), .A2(new_n477), .A3(new_n476), .ZN(new_n480));
  AND2_X1   g0280(.A1(new_n414), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n479), .B1(new_n481), .B2(G264), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n469), .A2(KEYINPUT86), .A3(new_n279), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n472), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT87), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n472), .A2(KEYINPUT87), .A3(new_n482), .A4(new_n483), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n486), .A2(new_n396), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(KEYINPUT88), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT88), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n486), .A2(new_n490), .A3(new_n396), .A4(new_n487), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n470), .A2(new_n482), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(new_n323), .ZN(new_n493));
  XOR2_X1   g0293(.A(new_n493), .B(KEYINPUT89), .Z(new_n494));
  NAND3_X1  g0294(.A1(new_n489), .A2(new_n491), .A3(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n335), .A2(KEYINPUT22), .A3(G87), .ZN(new_n496));
  NAND2_X1  g0296(.A1(G33), .A2(G116), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(new_n226), .ZN(new_n499));
  INV_X1    g0299(.A(G87), .ZN(new_n500));
  NOR3_X1   g0300(.A1(new_n372), .A2(G20), .A3(new_n500), .ZN(new_n501));
  OR2_X1    g0301(.A1(new_n501), .A2(KEYINPUT22), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n226), .A2(G107), .ZN(new_n503));
  XNOR2_X1  g0303(.A(new_n503), .B(KEYINPUT23), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n499), .A2(new_n502), .A3(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT24), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n499), .A2(KEYINPUT24), .A3(new_n502), .A4(new_n504), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n507), .A2(new_n263), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n271), .A2(new_n220), .ZN(new_n510));
  XNOR2_X1  g0310(.A(new_n510), .B(KEYINPUT25), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n248), .A2(G1), .ZN(new_n513));
  INV_X1    g0313(.A(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n382), .A2(KEYINPUT83), .A3(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT83), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n516), .B1(new_n381), .B2(new_n513), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n515), .A2(G107), .A3(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n509), .A2(new_n512), .A3(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n495), .A2(new_n520), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n346), .B1(new_n486), .B2(new_n487), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n492), .A2(new_n454), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n519), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  AND2_X1   g0324(.A1(new_n521), .A2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(new_n263), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT6), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n409), .A2(new_n220), .ZN(new_n528));
  NOR2_X1   g0328(.A1(G97), .A2(G107), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n220), .A2(KEYINPUT6), .A3(G97), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n226), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n370), .A2(new_n373), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n532), .B1(new_n533), .B2(G107), .ZN(new_n534));
  INV_X1    g0334(.A(G77), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n249), .A2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n526), .B1(new_n534), .B2(new_n537), .ZN(new_n538));
  AND3_X1   g0338(.A1(new_n515), .A2(G97), .A3(new_n517), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n270), .A2(G97), .ZN(new_n540));
  NOR3_X1   g0340(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  AND2_X1   g0341(.A1(new_n481), .A2(G257), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT4), .ZN(new_n543));
  INV_X1    g0343(.A(G244), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n543), .B1(new_n351), .B2(new_n544), .ZN(new_n545));
  OAI21_X1  g0345(.A(KEYINPUT4), .B1(new_n372), .B2(new_n463), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(G1698), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n289), .A2(KEYINPUT4), .A3(G244), .A4(new_n290), .ZN(new_n548));
  NAND2_X1  g0348(.A1(G33), .A2(G283), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n545), .A2(new_n547), .A3(new_n548), .A4(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n542), .B1(new_n550), .B2(new_n279), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n551), .A2(G190), .A3(new_n478), .ZN(new_n552));
  AOI211_X1 g0352(.A(new_n479), .B(new_n542), .C1(new_n279), .C2(new_n550), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n541), .B(new_n552), .C1(new_n323), .C2(new_n553), .ZN(new_n554));
  NOR2_X1   g0354(.A1(G238), .A2(G1698), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n555), .B1(new_n544), .B2(G1698), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n335), .A2(new_n556), .B1(G33), .B2(G116), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n477), .A2(G250), .ZN(new_n558));
  INV_X1    g0358(.A(G274), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n477), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n414), .A2(new_n560), .ZN(new_n561));
  OAI22_X1  g0361(.A1(new_n557), .A2(new_n414), .B1(new_n558), .B2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(G190), .ZN(new_n564));
  INV_X1    g0364(.A(new_n312), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n565), .A2(new_n270), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n335), .A2(new_n226), .A3(G68), .ZN(new_n567));
  NOR3_X1   g0367(.A1(new_n248), .A2(new_n409), .A3(G20), .ZN(new_n568));
  OR2_X1    g0368(.A1(new_n568), .A2(KEYINPUT19), .ZN(new_n569));
  AOI21_X1  g0369(.A(G20), .B1(new_n410), .B2(KEYINPUT19), .ZN(new_n570));
  NOR3_X1   g0370(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n567), .B(new_n569), .C1(new_n570), .C2(new_n571), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n566), .B1(new_n572), .B2(new_n263), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n562), .A2(G200), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n515), .A2(G87), .A3(new_n517), .ZN(new_n575));
  AND3_X1   g0375(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n515), .A2(new_n565), .A3(new_n517), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n573), .A2(new_n577), .B1(new_n346), .B2(new_n562), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n563), .A2(new_n454), .ZN(new_n579));
  AOI22_X1  g0379(.A1(new_n564), .A2(new_n576), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(new_n540), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n515), .A2(G97), .A3(new_n517), .ZN(new_n582));
  AOI211_X1 g0382(.A(new_n536), .B(new_n532), .C1(G107), .C2(new_n533), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n581), .B(new_n582), .C1(new_n583), .C2(new_n526), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n551), .A2(new_n454), .A3(new_n478), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n584), .B(new_n585), .C1(new_n553), .C2(G169), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n554), .A2(new_n580), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n465), .A2(new_n290), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n221), .A2(G1698), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n335), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n372), .A2(G303), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n279), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n414), .A2(new_n480), .A3(G270), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n478), .ZN(new_n595));
  INV_X1    g0395(.A(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  NOR2_X1   g0397(.A1(KEYINPUT85), .A2(KEYINPUT20), .ZN(new_n598));
  INV_X1    g0398(.A(G116), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(G20), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n549), .B(new_n226), .C1(G33), .C2(new_n409), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n263), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n602), .A2(KEYINPUT85), .A3(KEYINPUT20), .ZN(new_n603));
  NAND2_X1  g0403(.A1(KEYINPUT85), .A2(KEYINPUT20), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n263), .A2(new_n604), .A3(new_n600), .A4(new_n601), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n598), .B1(new_n603), .B2(new_n605), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n271), .A2(G116), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n382), .A2(new_n514), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n607), .B1(new_n608), .B2(G116), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n597), .B(G169), .C1(new_n606), .C2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT21), .ZN(new_n611));
  OR2_X1    g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n610), .A2(new_n611), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n414), .B1(new_n590), .B2(new_n591), .ZN(new_n614));
  NOR3_X1   g0414(.A1(new_n614), .A2(new_n595), .A3(new_n454), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n615), .B1(new_n606), .B2(new_n609), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n606), .A2(new_n609), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n597), .A2(G200), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n398), .A2(new_n397), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n617), .B(new_n618), .C1(new_n619), .C2(new_n597), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n612), .A2(new_n613), .A3(new_n616), .A4(new_n620), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n587), .A2(new_n621), .ZN(new_n622));
  AND3_X1   g0422(.A1(new_n462), .A2(new_n525), .A3(new_n622), .ZN(G372));
  INV_X1    g0423(.A(new_n310), .ZN(new_n624));
  AND3_X1   g0424(.A1(new_n348), .A2(KEYINPUT18), .A3(new_n387), .ZN(new_n625));
  AOI21_X1  g0425(.A(KEYINPUT18), .B1(new_n348), .B2(new_n387), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  AOI22_X1  g0428(.A1(new_n449), .A2(new_n461), .B1(new_n439), .B2(new_n455), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n405), .A2(new_n400), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n628), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  XNOR2_X1  g0431(.A(new_n631), .B(KEYINPUT90), .ZN(new_n632));
  AND2_X1   g0432(.A1(new_n303), .A2(new_n305), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n624), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n587), .ZN(new_n635));
  AND3_X1   g0435(.A1(new_n612), .A2(new_n613), .A3(new_n616), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(new_n524), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n521), .A2(new_n635), .A3(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n586), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n639), .A2(KEYINPUT26), .A3(new_n580), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT26), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n576), .A2(new_n564), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n578), .A2(new_n579), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n641), .B1(new_n644), .B2(new_n586), .ZN(new_n645));
  AOI22_X1  g0445(.A1(new_n640), .A2(new_n645), .B1(new_n579), .B2(new_n578), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n638), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n462), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n634), .A2(new_n648), .ZN(G369));
  INV_X1    g0449(.A(G330), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n636), .A2(KEYINPUT92), .A3(new_n620), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT92), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n621), .A2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(G13), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n654), .A2(G20), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(new_n225), .ZN(new_n656));
  OR3_X1    g0456(.A1(new_n656), .A2(KEYINPUT91), .A3(KEYINPUT27), .ZN(new_n657));
  INV_X1    g0457(.A(G213), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n658), .B1(new_n656), .B2(KEYINPUT27), .ZN(new_n659));
  OAI21_X1  g0459(.A(KEYINPUT91), .B1(new_n656), .B2(KEYINPUT27), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n657), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(G343), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  OAI211_X1 g0464(.A(new_n651), .B(new_n653), .C1(new_n617), .C2(new_n664), .ZN(new_n665));
  OAI211_X1 g0465(.A(new_n636), .B(new_n663), .C1(new_n609), .C2(new_n606), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(KEYINPUT93), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT93), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n665), .A2(new_n669), .A3(new_n666), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n650), .B1(new_n668), .B2(new_n670), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n525), .B1(new_n520), .B2(new_n664), .ZN(new_n672));
  OR2_X1    g0472(.A1(new_n524), .A2(new_n664), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  AND2_X1   g0475(.A1(new_n521), .A2(new_n637), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(new_n664), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n675), .A2(new_n677), .ZN(G399));
  INV_X1    g0478(.A(new_n205), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n679), .A2(G41), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(G1), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n571), .A2(new_n599), .ZN(new_n683));
  OAI22_X1  g0483(.A1(new_n682), .A2(new_n683), .B1(new_n229), .B2(new_n681), .ZN(new_n684));
  XNOR2_X1  g0484(.A(new_n684), .B(KEYINPUT28), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n663), .B1(new_n638), .B2(new_n646), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n687), .A2(KEYINPUT29), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n554), .A2(new_n586), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT96), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n554), .A2(KEYINPUT96), .A3(new_n586), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n693), .A2(new_n521), .A3(new_n642), .A4(new_n637), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n663), .B1(new_n694), .B2(new_n646), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT29), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  AND2_X1   g0497(.A1(new_n470), .A2(new_n482), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n551), .A2(new_n698), .A3(new_n563), .A4(new_n615), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(KEYINPUT94), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(KEYINPUT30), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n698), .B1(new_n551), .B2(new_n478), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n454), .B1(new_n614), .B2(new_n595), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  AOI21_X1  g0504(.A(KEYINPUT95), .B1(new_n704), .B2(new_n562), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT95), .ZN(new_n706));
  NOR3_X1   g0506(.A1(new_n703), .A2(new_n563), .A3(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n702), .B1(new_n705), .B2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT30), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n699), .A2(KEYINPUT94), .A3(new_n709), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n701), .A2(new_n708), .A3(new_n710), .ZN(new_n711));
  AND3_X1   g0511(.A1(new_n711), .A2(KEYINPUT31), .A3(new_n663), .ZN(new_n712));
  AOI21_X1  g0512(.A(KEYINPUT31), .B1(new_n711), .B2(new_n663), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n521), .A2(new_n622), .A3(new_n524), .A4(new_n664), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n650), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NOR3_X1   g0516(.A1(new_n688), .A2(new_n697), .A3(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n685), .B1(new_n717), .B2(G1), .ZN(G364));
  NAND3_X1  g0518(.A1(new_n668), .A2(new_n650), .A3(new_n670), .ZN(new_n719));
  XOR2_X1   g0519(.A(new_n719), .B(KEYINPUT97), .Z(new_n720));
  INV_X1    g0520(.A(new_n671), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n682), .B1(G45), .B2(new_n655), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n720), .A2(new_n721), .A3(new_n723), .ZN(new_n724));
  XOR2_X1   g0524(.A(new_n722), .B(KEYINPUT98), .Z(new_n725));
  NOR2_X1   g0525(.A1(new_n226), .A2(new_n454), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(G200), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n619), .A2(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n226), .A2(G179), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n729), .A2(new_n396), .A3(G200), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  AOI22_X1  g0531(.A1(new_n728), .A2(G50), .B1(G107), .B2(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n727), .A2(G190), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n454), .A2(new_n323), .ZN(new_n735));
  XNOR2_X1  g0535(.A(new_n735), .B(KEYINPUT100), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n736), .A2(G20), .A3(new_n396), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  AOI21_X1  g0538(.A(KEYINPUT32), .B1(new_n738), .B2(G159), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT32), .ZN(new_n740));
  NOR3_X1   g0540(.A1(new_n737), .A2(new_n740), .A3(new_n361), .ZN(new_n741));
  OAI221_X1 g0541(.A(new_n732), .B1(new_n210), .B2(new_n734), .C1(new_n739), .C2(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n736), .A2(G190), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(G20), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(G97), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n726), .A2(new_n323), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n619), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n746), .A2(G190), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  OAI221_X1 g0550(.A(new_n745), .B1(new_n217), .B2(new_n748), .C1(new_n535), .C2(new_n750), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n729), .A2(G190), .A3(G200), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(new_n500), .ZN(new_n753));
  NOR4_X1   g0553(.A1(new_n742), .A2(new_n751), .A3(new_n372), .A4(new_n753), .ZN(new_n754));
  XOR2_X1   g0554(.A(new_n754), .B(KEYINPUT101), .Z(new_n755));
  AOI21_X1  g0555(.A(new_n289), .B1(new_n738), .B2(G329), .ZN(new_n756));
  INV_X1    g0556(.A(G283), .ZN(new_n757));
  XOR2_X1   g0557(.A(KEYINPUT33), .B(G317), .Z(new_n758));
  OAI221_X1 g0558(.A(new_n756), .B1(new_n757), .B2(new_n730), .C1(new_n734), .C2(new_n758), .ZN(new_n759));
  AOI22_X1  g0559(.A1(new_n744), .A2(G294), .B1(G326), .B2(new_n728), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n759), .B1(KEYINPUT102), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n749), .A2(G311), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n747), .A2(G322), .ZN(new_n763));
  OR2_X1    g0563(.A1(new_n760), .A2(KEYINPUT102), .ZN(new_n764));
  NAND4_X1  g0564(.A1(new_n761), .A2(new_n762), .A3(new_n763), .A4(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n752), .ZN(new_n766));
  AND2_X1   g0566(.A1(new_n766), .A2(G303), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n755), .B1(new_n765), .B2(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n225), .B1(G20), .B2(new_n346), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n725), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  OR3_X1    g0570(.A1(KEYINPUT99), .A2(G13), .A3(G33), .ZN(new_n771));
  OAI21_X1  g0571(.A(KEYINPUT99), .B1(G13), .B2(G33), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(G20), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n667), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n679), .A2(new_n372), .ZN(new_n777));
  NAND2_X1  g0577(.A1(G355), .A2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n243), .A2(new_n281), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n335), .A2(new_n679), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n780), .B1(G45), .B2(new_n229), .ZN(new_n781));
  OAI221_X1 g0581(.A(new_n778), .B1(G116), .B2(new_n205), .C1(new_n779), .C2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n775), .A2(new_n769), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n770), .A2(new_n776), .A3(new_n784), .ZN(new_n785));
  XNOR2_X1  g0585(.A(new_n785), .B(KEYINPUT103), .ZN(new_n786));
  AND2_X1   g0586(.A1(new_n724), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(G396));
  NAND2_X1  g0588(.A1(new_n315), .A2(new_n663), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n324), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(new_n460), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n461), .A2(new_n664), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  XNOR2_X1  g0594(.A(new_n686), .B(new_n794), .ZN(new_n795));
  XOR2_X1   g0595(.A(new_n795), .B(new_n716), .Z(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(new_n722), .ZN(new_n797));
  INV_X1    g0597(.A(new_n769), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n728), .A2(G303), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n799), .B1(new_n220), .B2(new_n752), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n289), .B1(new_n731), .B2(G87), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n747), .A2(G294), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n745), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  AOI211_X1 g0603(.A(new_n800), .B(new_n803), .C1(G311), .C2(new_n738), .ZN(new_n804));
  OAI221_X1 g0604(.A(new_n804), .B1(new_n599), .B2(new_n750), .C1(new_n757), .C2(new_n734), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n730), .A2(new_n210), .ZN(new_n806));
  AOI211_X1 g0606(.A(new_n351), .B(new_n806), .C1(G50), .C2(new_n766), .ZN(new_n807));
  INV_X1    g0607(.A(G132), .ZN(new_n808));
  INV_X1    g0608(.A(new_n744), .ZN(new_n809));
  OAI221_X1 g0609(.A(new_n807), .B1(new_n808), .B2(new_n737), .C1(new_n809), .C2(new_n217), .ZN(new_n810));
  XNOR2_X1  g0610(.A(new_n810), .B(KEYINPUT105), .ZN(new_n811));
  AOI22_X1  g0611(.A1(new_n747), .A2(G143), .B1(new_n749), .B2(G159), .ZN(new_n812));
  INV_X1    g0612(.A(G137), .ZN(new_n813));
  INV_X1    g0613(.A(new_n728), .ZN(new_n814));
  INV_X1    g0614(.A(G150), .ZN(new_n815));
  OAI221_X1 g0615(.A(new_n812), .B1(new_n813), .B2(new_n814), .C1(new_n815), .C2(new_n734), .ZN(new_n816));
  XNOR2_X1  g0616(.A(new_n816), .B(KEYINPUT34), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n811), .A2(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n798), .B1(new_n805), .B2(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n773), .A2(new_n769), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n725), .B1(new_n535), .B2(new_n820), .ZN(new_n821));
  XOR2_X1   g0621(.A(new_n821), .B(KEYINPUT104), .Z(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  AOI211_X1 g0623(.A(new_n819), .B(new_n823), .C1(new_n773), .C2(new_n793), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n797), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(G384));
  OAI21_X1  g0626(.A(new_n462), .B1(new_n688), .B2(new_n697), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n634), .A2(new_n827), .ZN(new_n828));
  XNOR2_X1  g0628(.A(new_n828), .B(KEYINPUT111), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT110), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n367), .A2(new_n263), .ZN(new_n831));
  AOI21_X1  g0631(.A(KEYINPUT16), .B1(new_n356), .B2(new_n366), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n386), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n661), .ZN(new_n834));
  AND3_X1   g0634(.A1(new_n833), .A2(KEYINPUT107), .A3(new_n834), .ZN(new_n835));
  AOI21_X1  g0635(.A(KEYINPUT107), .B1(new_n833), .B2(new_n834), .ZN(new_n836));
  OR2_X1    g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n405), .A2(new_n400), .A3(new_n407), .ZN(new_n838));
  NOR3_X1   g0638(.A1(new_n625), .A2(new_n626), .A3(new_n406), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n837), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n387), .B1(new_n348), .B2(new_n834), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT37), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n841), .A2(new_n842), .A3(new_n404), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n348), .A2(new_n833), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(new_n404), .ZN(new_n845));
  NOR3_X1   g0645(.A1(new_n845), .A2(new_n835), .A3(new_n836), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n843), .B1(new_n846), .B2(new_n842), .ZN(new_n847));
  AND3_X1   g0647(.A1(new_n840), .A2(new_n847), .A3(KEYINPUT38), .ZN(new_n848));
  AOI21_X1  g0648(.A(KEYINPUT38), .B1(new_n840), .B2(new_n847), .ZN(new_n849));
  OAI21_X1  g0649(.A(KEYINPUT39), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n387), .A2(new_n834), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n852), .B1(new_n630), .B2(new_n627), .ZN(new_n853));
  AND4_X1   g0653(.A1(new_n842), .A2(new_n388), .A3(new_n404), .A4(new_n851), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n842), .B1(new_n841), .B2(new_n404), .ZN(new_n855));
  OAI21_X1  g0655(.A(KEYINPUT109), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n388), .A2(new_n404), .A3(new_n851), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(KEYINPUT37), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT109), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n858), .A2(new_n859), .A3(new_n843), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n853), .A2(new_n856), .A3(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT38), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT39), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n840), .A2(new_n847), .A3(KEYINPUT38), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n830), .B1(new_n850), .B2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n455), .A2(new_n439), .A3(new_n664), .ZN(new_n869));
  XNOR2_X1  g0669(.A(new_n869), .B(KEYINPUT108), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n850), .A2(new_n866), .A3(new_n830), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n868), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n439), .A2(new_n663), .ZN(new_n873));
  AND3_X1   g0673(.A1(new_n449), .A2(new_n456), .A3(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n873), .B1(new_n449), .B2(new_n456), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n647), .A2(new_n664), .A3(new_n794), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n876), .B1(new_n877), .B2(new_n792), .ZN(new_n878));
  INV_X1    g0678(.A(new_n849), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(new_n865), .ZN(new_n880));
  AOI22_X1  g0680(.A1(new_n878), .A2(new_n880), .B1(new_n627), .B2(new_n661), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n872), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g0682(.A(new_n829), .B(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT40), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n714), .A2(new_n715), .ZN(new_n885));
  INV_X1    g0685(.A(new_n875), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n449), .A2(new_n456), .A3(new_n873), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n793), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  OAI211_X1 g0688(.A(new_n885), .B(new_n888), .C1(new_n848), .C2(new_n849), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n884), .B1(new_n863), .B2(new_n865), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n794), .B1(new_n874), .B2(new_n875), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n891), .B1(new_n715), .B2(new_n714), .ZN(new_n892));
  AOI22_X1  g0692(.A1(new_n884), .A2(new_n889), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n462), .A2(new_n885), .ZN(new_n894));
  XOR2_X1   g0694(.A(new_n893), .B(new_n894), .Z(new_n895));
  NOR2_X1   g0695(.A1(new_n895), .A2(new_n650), .ZN(new_n896));
  XNOR2_X1  g0696(.A(new_n883), .B(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n897), .B1(new_n264), .B2(new_n655), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n530), .A2(new_n531), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n599), .B1(new_n899), .B2(KEYINPUT35), .ZN(new_n900));
  OAI211_X1 g0700(.A(new_n900), .B(new_n227), .C1(KEYINPUT35), .C2(new_n899), .ZN(new_n901));
  XNOR2_X1  g0701(.A(new_n901), .B(KEYINPUT36), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n230), .A2(G77), .A3(new_n357), .ZN(new_n903));
  XOR2_X1   g0703(.A(new_n903), .B(KEYINPUT106), .Z(new_n904));
  OAI21_X1  g0704(.A(new_n904), .B1(G50), .B2(new_n210), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n905), .A2(G1), .A3(new_n654), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n898), .A2(new_n902), .A3(new_n906), .ZN(G367));
  NOR2_X1   g0707(.A1(new_n636), .A2(new_n663), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n525), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n584), .A2(new_n663), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n693), .A2(new_n910), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n912), .B(KEYINPUT42), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n586), .B1(new_n911), .B2(new_n524), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(new_n664), .ZN(new_n915));
  AND2_X1   g0715(.A1(new_n573), .A2(new_n575), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n580), .B1(new_n916), .B2(new_n664), .ZN(new_n917));
  OR3_X1    g0717(.A1(new_n643), .A2(new_n916), .A3(new_n664), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  AOI22_X1  g0719(.A1(new_n913), .A2(new_n915), .B1(KEYINPUT43), .B2(new_n919), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n919), .A2(KEYINPUT43), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n920), .B(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(new_n675), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n911), .B1(new_n586), .B2(new_n664), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n922), .B(new_n925), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n680), .B(KEYINPUT41), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT112), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n924), .A2(new_n677), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT45), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n930), .B(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n676), .A2(new_n911), .A3(new_n664), .ZN(new_n933));
  XOR2_X1   g0733(.A(new_n933), .B(KEYINPUT44), .Z(new_n934));
  NAND2_X1  g0734(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(new_n923), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n932), .A2(new_n675), .A3(new_n934), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n909), .B1(new_n674), .B2(new_n908), .ZN(new_n939));
  OR2_X1    g0739(.A1(new_n939), .A2(new_n671), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n671), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(new_n717), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n929), .B1(new_n938), .B2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(new_n717), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n945), .B1(new_n940), .B2(new_n941), .ZN(new_n946));
  NAND4_X1  g0746(.A1(new_n946), .A2(KEYINPUT112), .A3(new_n937), .A4(new_n936), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n944), .A2(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n928), .B1(new_n948), .B2(new_n717), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n264), .B1(new_n655), .B2(G45), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n926), .B1(new_n949), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n744), .A2(G68), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n953), .B1(new_n815), .B2(new_n748), .ZN(new_n954));
  XOR2_X1   g0754(.A(new_n954), .B(KEYINPUT116), .Z(new_n955));
  AND2_X1   g0755(.A1(new_n728), .A2(G143), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n730), .A2(new_n535), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n957), .B1(G58), .B2(new_n766), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n958), .B1(new_n208), .B2(new_n750), .ZN(new_n959));
  NOR4_X1   g0759(.A1(new_n955), .A2(new_n372), .A3(new_n956), .A4(new_n959), .ZN(new_n960));
  OAI221_X1 g0760(.A(new_n960), .B1(new_n813), .B2(new_n737), .C1(new_n361), .C2(new_n734), .ZN(new_n961));
  AOI22_X1  g0761(.A1(new_n744), .A2(G107), .B1(G283), .B2(new_n749), .ZN(new_n962));
  XOR2_X1   g0762(.A(new_n962), .B(KEYINPUT113), .Z(new_n963));
  AOI22_X1  g0763(.A1(G303), .A2(new_n747), .B1(new_n728), .B2(G311), .ZN(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  AND2_X1   g0765(.A1(new_n965), .A2(KEYINPUT114), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n965), .A2(KEYINPUT114), .ZN(new_n967));
  NOR4_X1   g0767(.A1(new_n963), .A2(new_n335), .A3(new_n966), .A4(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n731), .A2(G97), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n733), .A2(G294), .ZN(new_n970));
  AOI21_X1  g0770(.A(KEYINPUT46), .B1(new_n766), .B2(G116), .ZN(new_n971));
  AND3_X1   g0771(.A1(new_n766), .A2(KEYINPUT46), .A3(G116), .ZN(new_n972));
  XNOR2_X1  g0772(.A(KEYINPUT115), .B(G317), .ZN(new_n973));
  AOI211_X1 g0773(.A(new_n971), .B(new_n972), .C1(new_n738), .C2(new_n973), .ZN(new_n974));
  NAND4_X1  g0774(.A1(new_n968), .A2(new_n969), .A3(new_n970), .A4(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n961), .A2(new_n975), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(KEYINPUT47), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n977), .A2(new_n769), .ZN(new_n978));
  INV_X1    g0778(.A(new_n725), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n917), .A2(new_n918), .A3(new_n775), .ZN(new_n980));
  INV_X1    g0780(.A(new_n780), .ZN(new_n981));
  OAI221_X1 g0781(.A(new_n783), .B1(new_n205), .B2(new_n312), .C1(new_n239), .C2(new_n981), .ZN(new_n982));
  NAND4_X1  g0782(.A1(new_n978), .A2(new_n979), .A3(new_n980), .A4(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n952), .A2(new_n983), .ZN(G387));
  NAND3_X1  g0784(.A1(new_n945), .A2(new_n941), .A3(new_n940), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n943), .A2(new_n680), .A3(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n942), .A2(new_n951), .ZN(new_n987));
  AOI22_X1  g0787(.A1(G303), .A2(new_n749), .B1(new_n733), .B2(G311), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n747), .A2(new_n973), .ZN(new_n989));
  INV_X1    g0789(.A(G322), .ZN(new_n990));
  OAI211_X1 g0790(.A(new_n988), .B(new_n989), .C1(new_n990), .C2(new_n814), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(KEYINPUT48), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n766), .A2(G294), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n992), .B(new_n993), .C1(new_n757), .C2(new_n809), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n994), .B(KEYINPUT49), .Z(new_n995));
  AOI21_X1  g0795(.A(new_n335), .B1(new_n738), .B2(G326), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n996), .B1(new_n599), .B2(new_n730), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(KEYINPUT117), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n995), .A2(new_n998), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n335), .B1(new_n734), .B2(new_n257), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(new_n744), .A2(new_n565), .B1(G68), .B2(new_n749), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n752), .A2(new_n535), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n1002), .B1(new_n738), .B2(G150), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n728), .A2(G159), .ZN(new_n1004));
  NAND4_X1  g0804(.A1(new_n1001), .A2(new_n1003), .A3(new_n969), .A4(new_n1004), .ZN(new_n1005));
  AOI211_X1 g0805(.A(new_n1000), .B(new_n1005), .C1(G50), .C2(new_n747), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n769), .B1(new_n999), .B2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n981), .B1(new_n236), .B2(G45), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1008), .B1(new_n683), .B2(new_n777), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n253), .A2(G50), .ZN(new_n1010));
  XOR2_X1   g0810(.A(new_n1010), .B(KEYINPUT50), .Z(new_n1011));
  NOR2_X1   g0811(.A1(new_n210), .A2(new_n535), .ZN(new_n1012));
  NOR4_X1   g0812(.A1(new_n1011), .A2(G45), .A3(new_n1012), .A4(new_n683), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n1009), .A2(new_n1013), .B1(G107), .B2(new_n205), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n725), .B1(new_n1014), .B2(new_n783), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n775), .ZN(new_n1016));
  OAI211_X1 g0816(.A(new_n1007), .B(new_n1015), .C1(new_n674), .C2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n986), .A2(new_n987), .A3(new_n1017), .ZN(G393));
  NAND3_X1  g0818(.A1(new_n936), .A2(new_n951), .A3(new_n937), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n783), .B1(new_n246), .B2(new_n981), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1020), .B1(G97), .B2(new_n679), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n809), .A2(new_n535), .ZN(new_n1022));
  AOI211_X1 g0822(.A(new_n351), .B(new_n1022), .C1(G143), .C2(new_n738), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n766), .A2(G68), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(G150), .A2(new_n728), .B1(new_n747), .B2(G159), .ZN(new_n1025));
  XOR2_X1   g0825(.A(new_n1025), .B(KEYINPUT51), .Z(new_n1026));
  OAI22_X1  g0826(.A1(new_n734), .A2(new_n208), .B1(new_n750), .B2(new_n253), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1027), .B1(G87), .B2(new_n731), .ZN(new_n1028));
  NAND4_X1  g0828(.A1(new_n1023), .A2(new_n1024), .A3(new_n1026), .A4(new_n1028), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n737), .A2(new_n990), .B1(new_n757), .B2(new_n752), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT118), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1031), .B1(G107), .B2(new_n731), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n744), .A2(G116), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n749), .A2(G294), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n289), .B1(new_n733), .B2(G303), .ZN(new_n1035));
  NAND4_X1  g0835(.A1(new_n1032), .A2(new_n1033), .A3(new_n1034), .A4(new_n1035), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(G311), .A2(new_n747), .B1(new_n728), .B2(G317), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(KEYINPUT52), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1029), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1039));
  AOI211_X1 g0839(.A(new_n725), .B(new_n1021), .C1(new_n1039), .C2(new_n769), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1040), .B1(new_n924), .B2(new_n1016), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1019), .A2(new_n1041), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n944), .A2(new_n947), .B1(new_n938), .B2(new_n943), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1042), .B1(new_n1043), .B2(new_n680), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1044), .ZN(G390));
  NOR3_X1   g0845(.A1(new_n408), .A2(new_n457), .A3(new_n461), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n325), .ZN(new_n1047));
  NAND4_X1  g0847(.A1(new_n885), .A2(G330), .A3(new_n1046), .A4(new_n1047), .ZN(new_n1048));
  INV_X1    g0848(.A(KEYINPUT120), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  NAND4_X1  g0850(.A1(new_n462), .A2(KEYINPUT120), .A3(G330), .A4(new_n885), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  AND3_X1   g0852(.A1(new_n634), .A2(new_n827), .A3(new_n1052), .ZN(new_n1053));
  AND2_X1   g0853(.A1(new_n794), .A2(KEYINPUT121), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n885), .A2(G330), .A3(new_n794), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1055), .A2(new_n876), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n876), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n716), .A2(new_n1057), .A3(new_n794), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1054), .B1(new_n1056), .B2(new_n1058), .ZN(new_n1059));
  AND3_X1   g0859(.A1(new_n716), .A2(KEYINPUT121), .A3(new_n794), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n695), .A2(new_n791), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1061), .A2(new_n792), .ZN(new_n1062));
  NOR3_X1   g0862(.A1(new_n1059), .A2(new_n1060), .A3(new_n1062), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n792), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1064), .B1(new_n686), .B2(new_n794), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1065), .B1(new_n1056), .B2(new_n1058), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1053), .B1(new_n1063), .B2(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT119), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1068), .B1(new_n878), .B2(new_n870), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n870), .ZN(new_n1070));
  OAI211_X1 g0870(.A(KEYINPUT119), .B(new_n1070), .C1(new_n1065), .C2(new_n876), .ZN(new_n1071));
  AND3_X1   g0871(.A1(new_n850), .A2(new_n830), .A3(new_n866), .ZN(new_n1072));
  OAI211_X1 g0872(.A(new_n1069), .B(new_n1071), .C1(new_n1072), .C2(new_n867), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1062), .A2(new_n1057), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n863), .A2(new_n865), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1074), .A2(new_n1075), .A3(new_n1070), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1073), .A2(new_n1058), .A3(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1058), .B1(new_n1073), .B2(new_n1076), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1067), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n1072), .A2(new_n867), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1076), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1058), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1063), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1066), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND4_X1  g0888(.A1(new_n1085), .A2(new_n1088), .A3(new_n1053), .A4(new_n1077), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1080), .A2(new_n1089), .A3(new_n680), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1085), .A2(new_n951), .A3(new_n1077), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n734), .A2(new_n220), .B1(new_n210), .B2(new_n730), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1022), .B1(G116), .B2(new_n747), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n1093), .B(KEYINPUT122), .ZN(new_n1094));
  AOI211_X1 g0894(.A(new_n1092), .B(new_n1094), .C1(G97), .C2(new_n749), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n738), .A2(G294), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n728), .A2(G283), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n753), .A2(new_n289), .ZN(new_n1098));
  NAND4_X1  g0898(.A1(new_n1095), .A2(new_n1096), .A3(new_n1097), .A4(new_n1098), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n752), .A2(new_n815), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(new_n1100), .B(KEYINPUT53), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(new_n728), .A2(G128), .B1(G50), .B2(new_n731), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  XOR2_X1   g0903(.A(KEYINPUT54), .B(G143), .Z(new_n1104));
  AOI21_X1  g0904(.A(new_n372), .B1(new_n749), .B2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1105), .B1(new_n809), .B2(new_n361), .ZN(new_n1106));
  AOI211_X1 g0906(.A(new_n1103), .B(new_n1106), .C1(G125), .C2(new_n738), .ZN(new_n1107));
  OAI221_X1 g0907(.A(new_n1107), .B1(new_n808), .B2(new_n748), .C1(new_n813), .C2(new_n734), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n798), .B1(new_n1099), .B2(new_n1108), .ZN(new_n1109));
  AOI211_X1 g0909(.A(new_n725), .B(new_n1109), .C1(new_n257), .C2(new_n820), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1110), .B1(new_n1081), .B2(new_n774), .ZN(new_n1111));
  AND3_X1   g0911(.A1(new_n1091), .A2(KEYINPUT123), .A3(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(KEYINPUT123), .B1(new_n1091), .B2(new_n1111), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1090), .B1(new_n1112), .B2(new_n1113), .ZN(G378));
  INV_X1    g0914(.A(KEYINPUT125), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n889), .A2(new_n884), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n890), .A2(new_n892), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1116), .A2(new_n1117), .A3(G330), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n303), .A2(new_n305), .A3(new_n310), .ZN(new_n1119));
  XOR2_X1   g0919(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1120));
  XNOR2_X1  g0920(.A(new_n1119), .B(new_n1120), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n273), .A2(new_n661), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(new_n1121), .B(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1118), .A2(new_n1123), .ZN(new_n1124));
  XOR2_X1   g0924(.A(new_n1121), .B(new_n1122), .Z(new_n1125));
  NAND3_X1  g0925(.A1(new_n893), .A2(G330), .A3(new_n1125), .ZN(new_n1126));
  AND4_X1   g0926(.A1(new_n872), .A2(new_n1124), .A3(new_n881), .A4(new_n1126), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(new_n1126), .A2(new_n1124), .B1(new_n872), .B2(new_n881), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1115), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1118), .A2(new_n1123), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1125), .B1(new_n893), .B2(G330), .ZN(new_n1131));
  NOR3_X1   g0931(.A1(new_n1072), .A2(new_n867), .A3(new_n1070), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n881), .ZN(new_n1133));
  OAI22_X1  g0933(.A1(new_n1130), .A2(new_n1131), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  NAND4_X1  g0934(.A1(new_n872), .A2(new_n1124), .A3(new_n1126), .A4(new_n881), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1134), .A2(KEYINPUT125), .A3(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1129), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1089), .A2(new_n1053), .ZN(new_n1138));
  AOI21_X1  g0938(.A(KEYINPUT57), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  AND3_X1   g0939(.A1(new_n1134), .A2(KEYINPUT57), .A3(new_n1135), .ZN(new_n1140));
  NOR3_X1   g0940(.A1(new_n1078), .A2(new_n1079), .A3(new_n1067), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n634), .A2(new_n827), .A3(new_n1052), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1140), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(new_n680), .ZN(new_n1144));
  OR2_X1    g0944(.A1(new_n1139), .A2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1125), .A2(new_n773), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n738), .A2(G283), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n728), .A2(G116), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n730), .A2(new_n217), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  NAND4_X1  g0950(.A1(new_n1147), .A2(new_n953), .A3(new_n1148), .A4(new_n1150), .ZN(new_n1151));
  OAI221_X1 g0951(.A(new_n351), .B1(new_n734), .B2(new_n409), .C1(new_n748), .C2(new_n220), .ZN(new_n1152));
  NOR4_X1   g0952(.A1(new_n1151), .A2(new_n1152), .A3(G41), .A4(new_n1002), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1153), .B1(new_n312), .B2(new_n750), .ZN(new_n1154));
  XOR2_X1   g0954(.A(new_n1154), .B(KEYINPUT124), .Z(new_n1155));
  XNOR2_X1  g0955(.A(new_n1155), .B(KEYINPUT58), .ZN(new_n1156));
  INV_X1    g0956(.A(G124), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n280), .B1(new_n737), .B2(new_n1157), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(new_n744), .A2(G150), .B1(G128), .B2(new_n747), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n728), .A2(G125), .B1(new_n749), .B2(G137), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n1159), .B(new_n1160), .C1(new_n808), .C2(new_n734), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1161), .B1(new_n766), .B2(new_n1104), .ZN(new_n1162));
  INV_X1    g0962(.A(KEYINPUT59), .ZN(new_n1163));
  AOI211_X1 g0963(.A(G33), .B(new_n1158), .C1(new_n1162), .C2(new_n1163), .ZN(new_n1164));
  OAI221_X1 g0964(.A(new_n1164), .B1(new_n1163), .B2(new_n1162), .C1(new_n361), .C2(new_n730), .ZN(new_n1165));
  AOI21_X1  g0965(.A(G41), .B1(new_n330), .B2(G33), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1165), .B1(G50), .B2(new_n1166), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n769), .B1(new_n1156), .B2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n820), .A2(new_n208), .ZN(new_n1169));
  NAND4_X1  g0969(.A1(new_n1146), .A2(new_n722), .A3(new_n1168), .A4(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1171), .B1(new_n1137), .B2(new_n951), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1145), .A2(new_n1172), .ZN(G375));
  NAND2_X1  g0973(.A1(new_n876), .A2(new_n773), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n744), .A2(G50), .B1(G150), .B2(new_n749), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(new_n1175), .B(KEYINPUT126), .ZN(new_n1176));
  AOI211_X1 g0976(.A(new_n351), .B(new_n1176), .C1(G128), .C2(new_n738), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n748), .A2(new_n813), .ZN(new_n1178));
  AOI211_X1 g0978(.A(new_n1149), .B(new_n1178), .C1(new_n733), .C2(new_n1104), .ZN(new_n1179));
  AND2_X1   g0979(.A1(new_n1177), .A2(new_n1179), .ZN(new_n1180));
  OAI221_X1 g0980(.A(new_n1180), .B1(new_n808), .B2(new_n814), .C1(new_n361), .C2(new_n752), .ZN(new_n1181));
  OAI22_X1  g0981(.A1(new_n809), .A2(new_n312), .B1(new_n757), .B2(new_n748), .ZN(new_n1182));
  AOI211_X1 g0982(.A(new_n957), .B(new_n1182), .C1(G303), .C2(new_n738), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n752), .A2(new_n409), .ZN(new_n1184));
  AOI211_X1 g0984(.A(new_n289), .B(new_n1184), .C1(G294), .C2(new_n728), .ZN(new_n1185));
  AND2_X1   g0985(.A1(new_n1183), .A2(new_n1185), .ZN(new_n1186));
  OAI221_X1 g0986(.A(new_n1186), .B1(new_n220), .B2(new_n750), .C1(new_n599), .C2(new_n734), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n798), .B1(new_n1181), .B2(new_n1187), .ZN(new_n1188));
  AOI211_X1 g0988(.A(new_n725), .B(new_n1188), .C1(new_n210), .C2(new_n820), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(new_n1088), .A2(new_n951), .B1(new_n1174), .B2(new_n1189), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1086), .A2(new_n1087), .A3(new_n1142), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1191), .A2(new_n927), .A3(new_n1067), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1190), .A2(new_n1192), .ZN(G381));
  INV_X1    g0993(.A(G375), .ZN(new_n1194));
  AND3_X1   g0994(.A1(new_n1090), .A2(new_n1091), .A3(new_n1111), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n952), .A2(new_n983), .A3(new_n1044), .ZN(new_n1197));
  OR3_X1    g0997(.A1(new_n1196), .A2(G381), .A3(new_n1197), .ZN(new_n1198));
  NOR3_X1   g0998(.A1(G396), .A2(G393), .A3(G384), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1199), .ZN(new_n1200));
  OR2_X1    g1000(.A1(new_n1198), .A2(new_n1200), .ZN(G407));
  OAI221_X1 g1001(.A(G213), .B1(new_n1196), .B2(G343), .C1(new_n1198), .C2(new_n1200), .ZN(G409));
  XNOR2_X1  g1002(.A(G393), .B(new_n787), .ZN(new_n1203));
  AND3_X1   g1003(.A1(new_n952), .A2(new_n983), .A3(new_n1044), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1044), .B1(new_n952), .B2(new_n983), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1203), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(G387), .A2(G390), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1203), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1207), .A2(new_n1197), .A3(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1206), .A2(new_n1209), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n658), .A2(G343), .ZN(new_n1211));
  OAI211_X1 g1011(.A(G378), .B(new_n1172), .C1(new_n1139), .C2(new_n1144), .ZN(new_n1212));
  AND3_X1   g1012(.A1(new_n1137), .A2(new_n927), .A3(new_n1138), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1134), .A2(new_n951), .A3(new_n1135), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1214), .A2(new_n1170), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1195), .B1(new_n1213), .B2(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1211), .B1(new_n1212), .B2(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT60), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n681), .B1(new_n1191), .B2(new_n1218), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n1219), .B(new_n1067), .C1(new_n1218), .C2(new_n1191), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1220), .A2(G384), .A3(new_n1190), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(G384), .B1(new_n1220), .B2(new_n1190), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1217), .A2(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1225), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1210), .B1(new_n1226), .B2(KEYINPUT63), .ZN(new_n1227));
  OAI211_X1 g1027(.A(G2897), .B(new_n1211), .C1(new_n1222), .C2(new_n1223), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1223), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1211), .A2(G2897), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1229), .A2(new_n1221), .A3(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1228), .A2(new_n1231), .ZN(new_n1232));
  OAI21_X1  g1032(.A(KEYINPUT63), .B1(new_n1232), .B2(new_n1217), .ZN(new_n1233));
  AOI21_X1  g1033(.A(KEYINPUT61), .B1(new_n1233), .B2(new_n1225), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1227), .A2(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT61), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1236), .B1(new_n1232), .B2(new_n1217), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1211), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1212), .A2(new_n1216), .ZN(new_n1239));
  OR2_X1    g1039(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n1240));
  AND4_X1   g1040(.A1(new_n1238), .A2(new_n1239), .A3(new_n1224), .A4(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1240), .B1(new_n1217), .B2(new_n1224), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1237), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1245));
  AND2_X1   g1045(.A1(new_n1206), .A2(new_n1209), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1235), .B1(new_n1245), .B2(new_n1246), .ZN(G405));
  NAND2_X1  g1047(.A1(G375), .A2(new_n1195), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1248), .A2(new_n1212), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1246), .A2(new_n1249), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1210), .A2(new_n1212), .A3(new_n1248), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1224), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1250), .A2(new_n1251), .A3(new_n1224), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1254), .A2(new_n1255), .ZN(G402));
endmodule


