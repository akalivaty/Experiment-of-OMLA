//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 0 0 0 1 0 0 0 1 1 0 1 1 1 1 0 1 1 0 1 1 1 1 0 1 1 1 0 0 0 0 1 0 0 0 0 1 0 0 0 1 1 0 0 1 0 0 1 1 0 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:32 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n677, new_n678, new_n679, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n695, new_n696, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n707, new_n708,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n778, new_n779, new_n780, new_n781, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  OAI21_X1  g001(.A(G210), .B1(G237), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(KEYINPUT83), .ZN(new_n190));
  INV_X1    g004(.A(G113), .ZN(new_n191));
  INV_X1    g005(.A(G116), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n192), .A2(G119), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT5), .ZN(new_n194));
  AOI21_X1  g008(.A(new_n191), .B1(new_n193), .B2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G119), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G116), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n192), .A2(G119), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n197), .A2(new_n198), .A3(KEYINPUT5), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n195), .A2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(KEYINPUT78), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n197), .A2(new_n198), .ZN(new_n202));
  XNOR2_X1  g016(.A(KEYINPUT2), .B(G113), .ZN(new_n203));
  OR2_X1    g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G104), .ZN(new_n205));
  OAI21_X1  g019(.A(KEYINPUT3), .B1(new_n205), .B2(G107), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT3), .ZN(new_n207));
  INV_X1    g021(.A(G107), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n207), .A2(new_n208), .A3(G104), .ZN(new_n209));
  INV_X1    g023(.A(G101), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n205), .A2(G107), .ZN(new_n211));
  NAND4_X1  g025(.A1(new_n206), .A2(new_n209), .A3(new_n210), .A4(new_n211), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n208), .A2(G104), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n205), .A2(G107), .ZN(new_n214));
  OAI21_X1  g028(.A(G101), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n212), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT78), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n195), .A2(new_n217), .A3(new_n199), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n201), .A2(new_n204), .A3(new_n216), .A4(new_n218), .ZN(new_n219));
  XNOR2_X1  g033(.A(G110), .B(G122), .ZN(new_n220));
  XNOR2_X1  g034(.A(new_n220), .B(KEYINPUT8), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT79), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n199), .A2(new_n222), .ZN(new_n223));
  NAND4_X1  g037(.A1(new_n197), .A2(new_n198), .A3(KEYINPUT79), .A4(KEYINPUT5), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n223), .A2(new_n195), .A3(new_n224), .ZN(new_n225));
  AND2_X1   g039(.A1(new_n225), .A2(new_n204), .ZN(new_n226));
  OAI211_X1 g040(.A(new_n219), .B(new_n221), .C1(new_n226), .C2(new_n216), .ZN(new_n227));
  INV_X1    g041(.A(G146), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(G143), .ZN(new_n229));
  INV_X1    g043(.A(G143), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G146), .ZN(new_n231));
  NAND2_X1  g045(.A1(KEYINPUT0), .A2(G128), .ZN(new_n232));
  AND3_X1   g046(.A1(new_n229), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(new_n233), .ZN(new_n234));
  OR2_X1    g048(.A1(KEYINPUT0), .A2(G128), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(new_n232), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n229), .A2(new_n231), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n234), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G125), .ZN(new_n240));
  INV_X1    g054(.A(G224), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n241), .A2(G953), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT1), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n229), .A2(new_n231), .A3(new_n243), .A4(G128), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  OAI21_X1  g059(.A(KEYINPUT1), .B1(new_n230), .B2(G146), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT67), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  OAI211_X1 g062(.A(KEYINPUT67), .B(KEYINPUT1), .C1(new_n230), .C2(G146), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n248), .A2(G128), .A3(new_n249), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n245), .B1(new_n250), .B2(new_n237), .ZN(new_n251));
  OAI211_X1 g065(.A(new_n240), .B(new_n242), .C1(G125), .C2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT7), .ZN(new_n253));
  OAI211_X1 g067(.A(new_n240), .B(new_n253), .C1(G125), .C2(new_n251), .ZN(new_n254));
  AND3_X1   g068(.A1(new_n227), .A2(new_n252), .A3(new_n254), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n240), .B1(new_n251), .B2(G125), .ZN(new_n256));
  OR2_X1    g070(.A1(new_n242), .A2(KEYINPUT80), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n253), .B1(new_n242), .B2(KEYINPUT80), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n256), .A2(KEYINPUT81), .A3(new_n257), .A4(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n249), .A2(G128), .ZN(new_n260));
  AOI21_X1  g074(.A(KEYINPUT67), .B1(new_n229), .B2(KEYINPUT1), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n237), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  AOI21_X1  g076(.A(G125), .B1(new_n262), .B2(new_n244), .ZN(new_n263));
  INV_X1    g077(.A(G125), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n264), .B1(new_n234), .B2(new_n238), .ZN(new_n265));
  OAI211_X1 g079(.A(new_n257), .B(new_n258), .C1(new_n263), .C2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT81), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n259), .A2(new_n268), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n206), .A2(new_n209), .A3(new_n211), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(G101), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n271), .A2(KEYINPUT4), .A3(new_n212), .ZN(new_n272));
  XNOR2_X1  g086(.A(new_n202), .B(new_n203), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT4), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n270), .A2(new_n274), .A3(G101), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n272), .A2(new_n273), .A3(new_n275), .ZN(new_n276));
  AND2_X1   g090(.A1(new_n212), .A2(new_n215), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n201), .A2(new_n277), .A3(new_n204), .A4(new_n218), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n276), .A2(new_n278), .A3(new_n220), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n255), .A2(new_n269), .A3(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT82), .ZN(new_n281));
  INV_X1    g095(.A(G902), .ZN(new_n282));
  AND3_X1   g096(.A1(new_n280), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n281), .B1(new_n280), .B2(new_n282), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n279), .A2(KEYINPUT6), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n276), .A2(new_n278), .ZN(new_n287));
  INV_X1    g101(.A(new_n220), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  XNOR2_X1  g103(.A(new_n286), .B(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n256), .B1(new_n241), .B2(G953), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(new_n252), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n190), .B1(new_n285), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n280), .A2(new_n282), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(KEYINPUT82), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n280), .A2(new_n281), .A3(new_n282), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n296), .A2(new_n190), .A3(new_n293), .A4(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n187), .B1(new_n294), .B2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT84), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n296), .A2(new_n293), .A3(new_n297), .ZN(new_n303));
  INV_X1    g117(.A(new_n190), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(new_n298), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n306), .A2(KEYINPUT84), .A3(new_n187), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n302), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(G234), .A2(G237), .ZN(new_n309));
  INV_X1    g123(.A(G953), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n309), .A2(G952), .A3(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  XOR2_X1   g126(.A(KEYINPUT21), .B(G898), .Z(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n309), .A2(G902), .A3(G953), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n312), .B1(new_n314), .B2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(G140), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(G125), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n264), .A2(G140), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(KEYINPUT19), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT19), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n320), .A2(new_n321), .A3(new_n324), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n323), .A2(new_n228), .A3(new_n325), .ZN(new_n326));
  OAI21_X1  g140(.A(KEYINPUT74), .B1(new_n320), .B2(KEYINPUT16), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n320), .A2(new_n321), .A3(KEYINPUT16), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT74), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT16), .ZN(new_n330));
  NAND4_X1  g144(.A1(new_n329), .A2(new_n330), .A3(new_n319), .A4(G125), .ZN(new_n331));
  NAND4_X1  g145(.A1(new_n327), .A2(new_n328), .A3(G146), .A4(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n326), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(KEYINPUT87), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT87), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n326), .A2(new_n335), .A3(new_n332), .ZN(new_n336));
  INV_X1    g150(.A(G237), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(KEYINPUT69), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT69), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(G237), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  AND2_X1   g155(.A1(KEYINPUT85), .A2(G143), .ZN(new_n342));
  NOR2_X1   g156(.A1(KEYINPUT85), .A2(G143), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  AND4_X1   g158(.A1(G214), .A2(new_n341), .A3(new_n344), .A4(new_n310), .ZN(new_n345));
  INV_X1    g159(.A(new_n342), .ZN(new_n346));
  AOI21_X1  g160(.A(G953), .B1(new_n338), .B2(new_n340), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n346), .B1(new_n347), .B2(G214), .ZN(new_n348));
  INV_X1    g162(.A(G131), .ZN(new_n349));
  NOR3_X1   g163(.A1(new_n345), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n341), .A2(G214), .A3(new_n310), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(new_n342), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n347), .A2(G214), .A3(new_n344), .ZN(new_n353));
  AOI21_X1  g167(.A(G131), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  OAI211_X1 g168(.A(new_n334), .B(new_n336), .C1(new_n350), .C2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT18), .ZN(new_n356));
  OAI21_X1  g170(.A(KEYINPUT86), .B1(new_n356), .B2(new_n349), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n352), .A2(new_n357), .A3(new_n353), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n356), .A2(new_n349), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT86), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n358), .A2(new_n361), .ZN(new_n362));
  XNOR2_X1  g176(.A(new_n322), .B(G146), .ZN(new_n363));
  NAND4_X1  g177(.A1(new_n352), .A2(new_n360), .A3(new_n359), .A4(new_n353), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n362), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n355), .A2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT88), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  XNOR2_X1  g182(.A(G113), .B(G122), .ZN(new_n369));
  XNOR2_X1  g183(.A(new_n369), .B(new_n205), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n355), .A2(new_n365), .A3(KEYINPUT88), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n368), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n349), .B1(new_n345), .B2(new_n348), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT17), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n352), .A2(G131), .A3(new_n353), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n374), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n345), .A2(new_n348), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT89), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n378), .A2(new_n379), .A3(KEYINPUT17), .A4(G131), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n327), .A2(new_n328), .A3(new_n331), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(new_n228), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(new_n332), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n352), .A2(KEYINPUT17), .A3(G131), .A4(new_n353), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(KEYINPUT89), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n377), .A2(new_n380), .A3(new_n384), .A4(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n387), .A2(new_n370), .A3(new_n365), .ZN(new_n388));
  AOI21_X1  g202(.A(G475), .B1(new_n373), .B2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT20), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n389), .A2(new_n390), .A3(new_n282), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n390), .B1(new_n389), .B2(new_n282), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT90), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n391), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND4_X1  g208(.A1(new_n389), .A2(KEYINPUT90), .A3(new_n390), .A4(new_n282), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  XNOR2_X1  g210(.A(KEYINPUT9), .B(G234), .ZN(new_n397));
  XOR2_X1   g211(.A(new_n397), .B(KEYINPUT75), .Z(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  XOR2_X1   g213(.A(KEYINPUT73), .B(G217), .Z(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  NOR3_X1   g215(.A1(new_n399), .A2(G953), .A3(new_n401), .ZN(new_n402));
  XNOR2_X1  g216(.A(G128), .B(G143), .ZN(new_n403));
  INV_X1    g217(.A(G134), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n403), .B(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n192), .A2(KEYINPUT14), .A3(G122), .ZN(new_n406));
  XNOR2_X1  g220(.A(G116), .B(G122), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  OAI211_X1 g222(.A(G107), .B(new_n406), .C1(new_n408), .C2(KEYINPUT14), .ZN(new_n409));
  OAI211_X1 g223(.A(new_n405), .B(new_n409), .C1(G107), .C2(new_n408), .ZN(new_n410));
  AOI21_X1  g224(.A(KEYINPUT13), .B1(new_n230), .B2(G128), .ZN(new_n411));
  XOR2_X1   g225(.A(new_n411), .B(KEYINPUT94), .Z(new_n412));
  NAND3_X1  g226(.A1(new_n230), .A2(KEYINPUT13), .A3(G128), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n413), .B1(G128), .B2(new_n230), .ZN(new_n414));
  OAI21_X1  g228(.A(G134), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n407), .B(new_n208), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n403), .A2(new_n404), .ZN(new_n417));
  XNOR2_X1  g231(.A(new_n417), .B(KEYINPUT95), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n415), .A2(new_n416), .A3(new_n418), .ZN(new_n419));
  AND3_X1   g233(.A1(new_n402), .A2(new_n410), .A3(new_n419), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n402), .B1(new_n419), .B2(new_n410), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(G478), .ZN(new_n424));
  OR2_X1    g238(.A1(new_n424), .A2(KEYINPUT15), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n423), .A2(new_n282), .A3(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n425), .B1(new_n423), .B2(new_n282), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT93), .ZN(new_n430));
  INV_X1    g244(.A(new_n388), .ZN(new_n431));
  AND3_X1   g245(.A1(new_n362), .A2(new_n363), .A3(new_n364), .ZN(new_n432));
  AND2_X1   g246(.A1(new_n377), .A2(new_n384), .ZN(new_n433));
  XNOR2_X1  g247(.A(new_n385), .B(new_n379), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n432), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  OAI21_X1  g249(.A(KEYINPUT92), .B1(new_n435), .B2(new_n370), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n387), .A2(new_n365), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT92), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n437), .A2(new_n438), .A3(new_n371), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n431), .B1(new_n436), .B2(new_n439), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n430), .B1(new_n440), .B2(G902), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n438), .B1(new_n437), .B2(new_n371), .ZN(new_n442));
  AOI211_X1 g256(.A(KEYINPUT92), .B(new_n370), .C1(new_n387), .C2(new_n365), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n388), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n444), .A2(KEYINPUT93), .A3(new_n282), .ZN(new_n445));
  XOR2_X1   g259(.A(KEYINPUT91), .B(G475), .Z(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n441), .A2(new_n445), .A3(new_n447), .ZN(new_n448));
  AND4_X1   g262(.A1(new_n318), .A2(new_n396), .A3(new_n429), .A4(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT23), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n450), .B1(new_n196), .B2(G128), .ZN(new_n451));
  INV_X1    g265(.A(G128), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n452), .A2(KEYINPUT23), .A3(G119), .ZN(new_n453));
  OAI211_X1 g267(.A(new_n451), .B(new_n453), .C1(G119), .C2(new_n452), .ZN(new_n454));
  XNOR2_X1  g268(.A(G119), .B(G128), .ZN(new_n455));
  XOR2_X1   g269(.A(KEYINPUT24), .B(G110), .Z(new_n456));
  AOI22_X1  g270(.A1(new_n454), .A2(G110), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n383), .A2(new_n457), .ZN(new_n458));
  OAI22_X1  g272(.A1(new_n454), .A2(G110), .B1(new_n455), .B2(new_n456), .ZN(new_n459));
  OAI211_X1 g273(.A(new_n459), .B(new_n332), .C1(G146), .C2(new_n322), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n310), .A2(G221), .A3(G234), .ZN(new_n462));
  XNOR2_X1  g276(.A(new_n462), .B(KEYINPUT22), .ZN(new_n463));
  INV_X1    g277(.A(G137), .ZN(new_n464));
  XNOR2_X1  g278(.A(new_n463), .B(new_n464), .ZN(new_n465));
  OR2_X1    g279(.A1(new_n461), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n461), .A2(new_n465), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n466), .A2(new_n282), .A3(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT25), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n468), .B(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n401), .B1(G234), .B2(new_n282), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n472), .B1(new_n471), .B2(new_n468), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT68), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n464), .A2(KEYINPUT11), .A3(G134), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n404), .A2(G137), .ZN(new_n476));
  AND2_X1   g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT11), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n478), .B1(new_n404), .B2(G137), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(KEYINPUT65), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n464), .A2(G134), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT65), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n481), .A2(new_n482), .A3(new_n478), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n477), .A2(new_n349), .A3(new_n480), .A4(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT66), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n481), .A2(new_n476), .A3(new_n485), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n486), .B(G131), .C1(new_n485), .C2(new_n481), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n474), .B1(new_n488), .B2(new_n251), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n482), .B1(new_n481), .B2(new_n478), .ZN(new_n490));
  AOI211_X1 g304(.A(KEYINPUT65), .B(KEYINPUT11), .C1(new_n464), .C2(G134), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n349), .B1(new_n492), .B2(new_n477), .ZN(new_n493));
  INV_X1    g307(.A(new_n484), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n239), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n262), .A2(new_n244), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n496), .A2(KEYINPUT68), .A3(new_n484), .A4(new_n487), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n489), .A2(new_n495), .A3(new_n497), .A4(KEYINPUT30), .ZN(new_n498));
  XOR2_X1   g312(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n499));
  NOR2_X1   g313(.A1(new_n488), .A2(new_n251), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n233), .B1(new_n237), .B2(new_n236), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n477), .A2(new_n480), .A3(new_n483), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(G131), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n501), .B1(new_n503), .B2(new_n484), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n499), .B1(new_n500), .B2(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n498), .A2(new_n505), .A3(new_n273), .ZN(new_n506));
  INV_X1    g320(.A(new_n273), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n489), .A2(new_n495), .A3(new_n497), .A4(new_n507), .ZN(new_n508));
  AND2_X1   g322(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT70), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT31), .ZN(new_n511));
  XNOR2_X1  g325(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n512), .B(G101), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n347), .A2(G210), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n513), .B(new_n514), .ZN(new_n515));
  NAND4_X1  g329(.A1(new_n509), .A2(new_n510), .A3(new_n511), .A4(new_n515), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n273), .B1(new_n500), .B2(new_n504), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n508), .A2(new_n517), .ZN(new_n518));
  XNOR2_X1  g332(.A(KEYINPUT71), .B(KEYINPUT28), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n500), .A2(new_n504), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(new_n507), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT28), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n520), .A2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n515), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND4_X1  g341(.A1(new_n506), .A2(new_n510), .A3(new_n508), .A4(new_n515), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(KEYINPUT31), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n516), .A2(new_n527), .A3(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(G472), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n530), .A2(new_n531), .A3(new_n282), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(KEYINPUT32), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT32), .ZN(new_n534));
  NAND4_X1  g348(.A1(new_n530), .A2(new_n534), .A3(new_n531), .A4(new_n282), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT29), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n520), .A2(new_n537), .A3(new_n524), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n489), .A2(new_n495), .A3(new_n497), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(new_n273), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n523), .B1(new_n540), .B2(new_n508), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT72), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n542), .B1(new_n522), .B2(new_n523), .ZN(new_n543));
  AOI211_X1 g357(.A(KEYINPUT72), .B(KEYINPUT28), .C1(new_n521), .C2(new_n507), .ZN(new_n544));
  NOR3_X1   g358(.A1(new_n541), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  OAI211_X1 g359(.A(new_n515), .B(new_n538), .C1(new_n545), .C2(new_n537), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n515), .A2(KEYINPUT29), .ZN(new_n547));
  AOI21_X1  g361(.A(G902), .B1(new_n509), .B2(new_n547), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n531), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n473), .B1(new_n536), .B2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(G469), .ZN(new_n552));
  AOI22_X1  g366(.A1(new_n246), .A2(G128), .B1(new_n229), .B2(new_n231), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n277), .B1(new_n245), .B2(new_n553), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n554), .B1(new_n496), .B2(new_n277), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n493), .A2(new_n494), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(KEYINPUT12), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n496), .A2(KEYINPUT10), .A3(new_n277), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n272), .A2(new_n239), .A3(new_n275), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT10), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n245), .A2(new_n553), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n562), .B1(new_n563), .B2(new_n216), .ZN(new_n564));
  NAND4_X1  g378(.A1(new_n560), .A2(new_n556), .A3(new_n561), .A4(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT12), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n555), .A2(new_n557), .A3(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n559), .A2(new_n565), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n310), .A2(G227), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n569), .B(new_n319), .ZN(new_n570));
  XNOR2_X1  g384(.A(new_n570), .B(KEYINPUT76), .ZN(new_n571));
  XOR2_X1   g385(.A(new_n571), .B(G110), .Z(new_n572));
  NOR2_X1   g386(.A1(new_n568), .A2(new_n572), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n571), .B(G110), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n560), .A2(new_n561), .A3(new_n564), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(new_n557), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n574), .B1(new_n565), .B2(new_n576), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n552), .B(new_n282), .C1(new_n573), .C2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(G469), .A2(G902), .ZN(new_n579));
  AND2_X1   g393(.A1(new_n574), .A2(KEYINPUT77), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n574), .A2(KEYINPUT77), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n568), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n576), .A2(new_n574), .A3(new_n565), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n582), .A2(G469), .A3(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n578), .A2(new_n579), .A3(new_n584), .ZN(new_n585));
  OAI21_X1  g399(.A(G221), .B1(new_n399), .B2(G902), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n308), .A2(new_n449), .A3(new_n551), .A4(new_n588), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n589), .B(G101), .ZN(G3));
  AOI21_X1  g404(.A(new_n531), .B1(new_n530), .B2(new_n282), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  AND2_X1   g406(.A1(new_n592), .A2(new_n532), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  NOR3_X1   g408(.A1(new_n594), .A2(new_n473), .A3(new_n587), .ZN(new_n595));
  AOI21_X1  g409(.A(G478), .B1(new_n423), .B2(new_n282), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT33), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(KEYINPUT96), .ZN(new_n598));
  OR2_X1    g412(.A1(new_n597), .A2(KEYINPUT96), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n423), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n422), .A2(KEYINPUT96), .A3(new_n597), .ZN(new_n601));
  AOI21_X1  g415(.A(G902), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n596), .B1(new_n602), .B2(G478), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n603), .B1(new_n396), .B2(new_n448), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n285), .A2(new_n189), .A3(new_n293), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n303), .A2(new_n188), .ZN(new_n606));
  AND3_X1   g420(.A1(new_n605), .A2(new_n606), .A3(new_n187), .ZN(new_n607));
  AND3_X1   g421(.A1(new_n604), .A2(new_n318), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n595), .A2(new_n608), .ZN(new_n609));
  XOR2_X1   g423(.A(KEYINPUT34), .B(G104), .Z(new_n610));
  XNOR2_X1  g424(.A(new_n609), .B(new_n610), .ZN(G6));
  INV_X1    g425(.A(KEYINPUT100), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT98), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n441), .A2(new_n613), .A3(new_n445), .A4(new_n447), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT97), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n392), .A2(new_n615), .ZN(new_n616));
  AND2_X1   g430(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n429), .ZN(new_n618));
  INV_X1    g432(.A(new_n392), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n619), .A2(KEYINPUT97), .A3(new_n391), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n445), .A2(new_n447), .ZN(new_n621));
  AOI21_X1  g435(.A(KEYINPUT93), .B1(new_n444), .B2(new_n282), .ZN(new_n622));
  OAI21_X1  g436(.A(KEYINPUT98), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n617), .A2(new_n618), .A3(new_n620), .A4(new_n623), .ZN(new_n624));
  XOR2_X1   g438(.A(new_n317), .B(KEYINPUT99), .Z(new_n625));
  OAI21_X1  g439(.A(new_n612), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n623), .A2(new_n620), .A3(new_n614), .A4(new_n616), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n625), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n628), .A2(KEYINPUT100), .A3(new_n618), .A4(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n626), .A2(new_n607), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(KEYINPUT101), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT101), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n626), .A2(new_n633), .A3(new_n607), .A4(new_n630), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(new_n595), .ZN(new_n636));
  XOR2_X1   g450(.A(KEYINPUT35), .B(G107), .Z(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(G9));
  NOR2_X1   g452(.A1(new_n465), .A2(KEYINPUT36), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n461), .B(new_n639), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n471), .A2(G902), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n472), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n449), .A2(new_n643), .ZN(new_n644));
  AOI21_X1  g458(.A(KEYINPUT84), .B1(new_n306), .B2(new_n187), .ZN(new_n645));
  INV_X1    g459(.A(new_n187), .ZN(new_n646));
  AOI211_X1 g460(.A(new_n301), .B(new_n646), .C1(new_n305), .C2(new_n298), .ZN(new_n647));
  OAI211_X1 g461(.A(new_n588), .B(new_n593), .C1(new_n645), .C2(new_n647), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n644), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(KEYINPUT37), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(G110), .ZN(G12));
  AOI21_X1  g465(.A(new_n549), .B1(new_n533), .B2(new_n535), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n605), .A2(new_n643), .A3(new_n606), .A4(new_n187), .ZN(new_n653));
  NOR3_X1   g467(.A1(new_n652), .A2(new_n587), .A3(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n627), .A2(new_n429), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n311), .B1(new_n315), .B2(G900), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n654), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(G128), .ZN(G30));
  XOR2_X1   g472(.A(new_n656), .B(KEYINPUT39), .Z(new_n659));
  NOR2_X1   g473(.A1(new_n587), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(KEYINPUT102), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT40), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n663), .A2(new_n646), .ZN(new_n664));
  INV_X1    g478(.A(new_n509), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n665), .A2(new_n526), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n515), .B1(new_n540), .B2(new_n508), .ZN(new_n667));
  OAI21_X1  g481(.A(new_n282), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(G472), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n643), .B1(new_n536), .B2(new_n669), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n429), .B1(new_n396), .B2(new_n448), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT38), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n306), .B(new_n672), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n673), .B1(new_n661), .B2(new_n662), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n664), .A2(new_n670), .A3(new_n671), .A4(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G143), .ZN(G45));
  INV_X1    g490(.A(new_n656), .ZN(new_n677));
  AOI211_X1 g491(.A(new_n603), .B(new_n677), .C1(new_n396), .C2(new_n448), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n654), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G146), .ZN(G48));
  INV_X1    g494(.A(new_n551), .ZN(new_n681));
  OAI21_X1  g495(.A(new_n282), .B1(new_n573), .B2(new_n577), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n552), .A2(KEYINPUT103), .ZN(new_n683));
  OR2_X1    g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n682), .A2(new_n683), .ZN(new_n685));
  AND3_X1   g499(.A1(new_n684), .A2(new_n586), .A3(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n681), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(new_n608), .ZN(new_n689));
  XNOR2_X1  g503(.A(KEYINPUT41), .B(G113), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n689), .B(new_n690), .ZN(G15));
  INV_X1    g505(.A(new_n688), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n692), .B1(new_n632), .B2(new_n634), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(new_n192), .ZN(G18));
  NAND2_X1  g508(.A1(new_n607), .A2(new_n686), .ZN(new_n695));
  NOR3_X1   g509(.A1(new_n644), .A2(new_n652), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(new_n196), .ZN(G21));
  NAND2_X1  g511(.A1(new_n671), .A2(new_n607), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n531), .A2(new_n282), .ZN(new_n699));
  OR2_X1    g513(.A1(new_n541), .A2(new_n543), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n526), .B1(new_n700), .B2(new_n544), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n528), .B(new_n511), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n699), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  OR3_X1    g517(.A1(new_n473), .A2(new_n591), .A3(new_n703), .ZN(new_n704));
  OR4_X1    g518(.A1(new_n625), .A2(new_n698), .A3(new_n687), .A4(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G122), .ZN(G24));
  INV_X1    g520(.A(new_n695), .ZN(new_n707));
  AOI22_X1  g521(.A1(new_n470), .A2(new_n471), .B1(new_n640), .B2(new_n641), .ZN(new_n708));
  NOR3_X1   g522(.A1(new_n591), .A2(new_n703), .A3(new_n708), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n678), .A2(new_n707), .A3(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G125), .ZN(G27));
  INV_X1    g525(.A(KEYINPUT42), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT105), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n583), .A2(new_n713), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n576), .A2(new_n574), .A3(KEYINPUT105), .A4(new_n565), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n716), .A2(new_n582), .A3(G469), .ZN(new_n717));
  XOR2_X1   g531(.A(new_n579), .B(KEYINPUT104), .Z(new_n718));
  NAND3_X1  g532(.A1(new_n578), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(new_n586), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT106), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n305), .A2(new_n187), .A3(new_n298), .ZN(new_n723));
  AOI21_X1  g537(.A(KEYINPUT106), .B1(new_n719), .B2(new_n586), .ZN(new_n724));
  NOR3_X1   g538(.A1(new_n722), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n551), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n604), .A2(new_n656), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n712), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n678), .A2(new_n551), .A3(new_n725), .A4(KEYINPUT42), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G131), .ZN(G33));
  NAND4_X1  g545(.A1(new_n655), .A2(new_n551), .A3(new_n656), .A4(new_n725), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G134), .ZN(G36));
  NAND2_X1  g547(.A1(new_n396), .A2(new_n448), .ZN(new_n734));
  INV_X1    g548(.A(new_n603), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT43), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  OR2_X1    g551(.A1(new_n734), .A2(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT108), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n396), .A2(new_n740), .A3(new_n448), .ZN(new_n741));
  INV_X1    g555(.A(new_n741), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n740), .B1(new_n396), .B2(new_n448), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n735), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n739), .B1(KEYINPUT43), .B2(new_n744), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n593), .B1(new_n745), .B2(KEYINPUT109), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n734), .A2(KEYINPUT108), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n603), .B1(new_n747), .B2(new_n741), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n738), .B1(new_n748), .B2(new_n736), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT109), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n746), .A2(KEYINPUT44), .A3(new_n643), .A4(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT44), .ZN(new_n753));
  OAI211_X1 g567(.A(KEYINPUT109), .B(new_n738), .C1(new_n748), .C2(new_n736), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n754), .A2(new_n594), .A3(new_n643), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n744), .A2(KEYINPUT43), .ZN(new_n756));
  AOI21_X1  g570(.A(KEYINPUT109), .B1(new_n756), .B2(new_n738), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n753), .B1(new_n755), .B2(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(new_n723), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n582), .A2(new_n583), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT45), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n716), .A2(new_n582), .A3(KEYINPUT45), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n762), .A2(G469), .A3(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n764), .A2(KEYINPUT46), .A3(new_n718), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT107), .ZN(new_n766));
  OR2_X1    g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  AOI21_X1  g581(.A(KEYINPUT46), .B1(new_n764), .B2(new_n718), .ZN(new_n768));
  INV_X1    g582(.A(new_n578), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n765), .A2(new_n766), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n767), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(new_n659), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n772), .A2(new_n586), .A3(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(new_n774), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n752), .A2(new_n758), .A3(new_n759), .A4(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G137), .ZN(G39));
  NAND2_X1  g591(.A1(new_n772), .A2(new_n586), .ZN(new_n778));
  XOR2_X1   g592(.A(new_n778), .B(KEYINPUT47), .Z(new_n779));
  AND2_X1   g593(.A1(new_n652), .A2(new_n473), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n779), .A2(new_n678), .A3(new_n759), .A4(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G140), .ZN(G42));
  NOR2_X1   g596(.A1(new_n687), .A2(new_n723), .ZN(new_n783));
  AND2_X1   g597(.A1(new_n536), .A2(new_n669), .ZN(new_n784));
  INV_X1    g598(.A(new_n473), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n783), .A2(new_n784), .A3(new_n785), .A4(new_n312), .ZN(new_n786));
  INV_X1    g600(.A(new_n604), .ZN(new_n787));
  OAI211_X1 g601(.A(G952), .B(new_n310), .C1(new_n786), .C2(new_n787), .ZN(new_n788));
  NOR3_X1   g602(.A1(new_n749), .A2(new_n311), .A3(new_n704), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n788), .B1(new_n789), .B2(new_n707), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT48), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n749), .A2(new_n311), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n792), .A2(new_n783), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT115), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n792), .A2(KEYINPUT115), .A3(new_n783), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n791), .B1(new_n797), .B2(new_n551), .ZN(new_n798));
  AOI211_X1 g612(.A(KEYINPUT48), .B(new_n681), .C1(new_n795), .C2(new_n796), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n790), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(KEYINPUT117), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n705), .A2(new_n689), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n802), .B1(new_n635), .B2(new_n688), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n396), .A2(new_n618), .A3(new_n448), .ZN(new_n804));
  INV_X1    g618(.A(new_n804), .ZN(new_n805));
  AND4_X1   g619(.A1(new_n532), .A2(new_n785), .A3(new_n592), .A4(new_n629), .ZN(new_n806));
  AND4_X1   g620(.A1(new_n308), .A2(new_n588), .A3(new_n805), .A4(new_n806), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n649), .A2(new_n807), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n308), .A2(new_n588), .A3(new_n604), .A4(new_n806), .ZN(new_n809));
  AND3_X1   g623(.A1(new_n589), .A2(new_n809), .A3(KEYINPUT111), .ZN(new_n810));
  AOI21_X1  g624(.A(KEYINPUT111), .B1(new_n589), .B2(new_n809), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n808), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n734), .A2(new_n709), .A3(new_n735), .A4(new_n656), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n723), .A2(new_n724), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n814), .B1(new_n721), .B2(new_n720), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n643), .A2(new_n429), .A3(new_n656), .ZN(new_n817));
  NOR4_X1   g631(.A1(new_n652), .A2(new_n587), .A3(new_n723), .A4(new_n817), .ZN(new_n818));
  AOI22_X1  g632(.A1(new_n816), .A2(KEYINPUT112), .B1(new_n818), .B2(new_n628), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT112), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n820), .B1(new_n813), .B2(new_n815), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n730), .A2(new_n819), .A3(new_n732), .A4(new_n821), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n812), .A2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(new_n696), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n720), .A2(new_n677), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n670), .A2(new_n607), .A3(new_n671), .A4(new_n825), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n657), .A2(new_n679), .A3(new_n710), .A4(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT52), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  OAI211_X1 g643(.A(new_n654), .B(new_n656), .C1(new_n655), .C2(new_n604), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n830), .A2(KEYINPUT52), .A3(new_n710), .A4(new_n826), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n803), .A2(new_n823), .A3(new_n824), .A4(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n833), .A2(KEYINPUT53), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT113), .ZN(new_n835));
  AND3_X1   g649(.A1(new_n829), .A2(new_n835), .A3(new_n831), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n835), .B1(new_n829), .B2(new_n831), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n693), .A2(new_n696), .A3(new_n802), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT53), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n838), .A2(new_n839), .A3(new_n840), .A4(new_n823), .ZN(new_n841));
  AND2_X1   g655(.A1(new_n834), .A2(new_n841), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n842), .A2(KEYINPUT54), .ZN(new_n843));
  INV_X1    g657(.A(new_n843), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n833), .A2(KEYINPUT53), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n838), .A2(new_n839), .A3(new_n823), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n845), .B1(KEYINPUT53), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(KEYINPUT54), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n801), .A2(new_n844), .A3(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(new_n673), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT114), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n687), .A2(new_n187), .ZN(new_n852));
  INV_X1    g666(.A(new_n852), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n850), .B1(new_n851), .B2(new_n853), .ZN(new_n854));
  OAI211_X1 g668(.A(new_n789), .B(new_n854), .C1(new_n851), .C2(new_n853), .ZN(new_n855));
  XOR2_X1   g669(.A(new_n855), .B(KEYINPUT50), .Z(new_n856));
  INV_X1    g670(.A(new_n709), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n857), .B1(new_n795), .B2(new_n796), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n684), .A2(new_n685), .ZN(new_n859));
  XOR2_X1   g673(.A(new_n859), .B(KEYINPUT110), .Z(new_n860));
  NOR2_X1   g674(.A1(new_n860), .A2(new_n586), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n779), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n789), .A2(new_n759), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n786), .A2(new_n734), .A3(new_n735), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n858), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n856), .A2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT51), .ZN(new_n868));
  INV_X1    g682(.A(new_n864), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n868), .B1(new_n869), .B2(KEYINPUT116), .ZN(new_n870));
  XOR2_X1   g684(.A(new_n867), .B(new_n870), .Z(new_n871));
  OAI22_X1  g685(.A1(new_n849), .A2(new_n871), .B1(G952), .B2(G953), .ZN(new_n872));
  XOR2_X1   g686(.A(new_n860), .B(KEYINPUT49), .Z(new_n873));
  AND4_X1   g687(.A1(new_n187), .A2(new_n873), .A3(new_n586), .A4(new_n748), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n874), .A2(new_n785), .A3(new_n784), .A4(new_n673), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n872), .A2(new_n875), .ZN(G75));
  NAND3_X1  g690(.A1(new_n834), .A2(new_n841), .A3(G902), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n877), .A2(KEYINPUT118), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT118), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n834), .A2(new_n841), .A3(new_n879), .A4(G902), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n878), .A2(new_n189), .A3(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT56), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n290), .B(new_n292), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n883), .B(KEYINPUT55), .ZN(new_n884));
  INV_X1    g698(.A(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n881), .A2(new_n882), .A3(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT119), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n310), .A2(G952), .ZN(new_n889));
  INV_X1    g703(.A(G210), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n882), .B1(new_n877), .B2(new_n890), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n889), .B1(new_n891), .B2(new_n884), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n881), .A2(KEYINPUT119), .A3(new_n882), .A4(new_n885), .ZN(new_n893));
  AND3_X1   g707(.A1(new_n888), .A2(new_n892), .A3(new_n893), .ZN(G51));
  XOR2_X1   g708(.A(new_n718), .B(KEYINPUT57), .Z(new_n895));
  AND2_X1   g709(.A1(new_n842), .A2(KEYINPUT54), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n895), .B1(new_n896), .B2(new_n843), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n897), .B1(new_n577), .B2(new_n573), .ZN(new_n898));
  INV_X1    g712(.A(new_n764), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n878), .A2(new_n899), .A3(new_n880), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n889), .B1(new_n898), .B2(new_n900), .ZN(G54));
  NAND2_X1  g715(.A1(KEYINPUT58), .A2(G475), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(KEYINPUT120), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n878), .A2(new_n880), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n373), .A2(new_n388), .ZN(new_n905));
  INV_X1    g719(.A(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(new_n889), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n878), .A2(new_n905), .A3(new_n880), .A4(new_n903), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n907), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(KEYINPUT121), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT121), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n907), .A2(new_n912), .A3(new_n908), .A4(new_n909), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n911), .A2(new_n913), .ZN(G60));
  NAND2_X1  g728(.A1(new_n600), .A2(new_n601), .ZN(new_n915));
  NAND2_X1  g729(.A1(G478), .A2(G902), .ZN(new_n916));
  XOR2_X1   g730(.A(new_n916), .B(KEYINPUT59), .Z(new_n917));
  INV_X1    g731(.A(new_n917), .ZN(new_n918));
  OAI211_X1 g732(.A(new_n915), .B(new_n918), .C1(new_n896), .C2(new_n843), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n917), .B1(new_n844), .B2(new_n848), .ZN(new_n920));
  OAI211_X1 g734(.A(new_n908), .B(new_n919), .C1(new_n920), .C2(new_n915), .ZN(new_n921));
  INV_X1    g735(.A(new_n921), .ZN(G63));
  NAND2_X1  g736(.A1(G217), .A2(G902), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n923), .B(KEYINPUT60), .Z(new_n924));
  NAND2_X1  g738(.A1(new_n842), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n466), .A2(new_n467), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n889), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n842), .A2(new_n640), .A3(new_n924), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(KEYINPUT122), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT122), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n842), .A2(new_n930), .A3(new_n640), .A4(new_n924), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n927), .A2(new_n929), .A3(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT61), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n927), .A2(new_n929), .A3(KEYINPUT61), .A4(new_n931), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n934), .A2(new_n935), .ZN(G66));
  OR4_X1    g750(.A1(new_n693), .A2(new_n812), .A3(new_n696), .A4(new_n802), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(new_n310), .ZN(new_n938));
  OAI21_X1  g752(.A(G953), .B1(new_n314), .B2(new_n241), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  XOR2_X1   g754(.A(new_n940), .B(KEYINPUT123), .Z(new_n941));
  INV_X1    g755(.A(G898), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n290), .B1(new_n942), .B2(G953), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n941), .B(new_n943), .ZN(G69));
  NAND2_X1  g758(.A1(new_n498), .A2(new_n505), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n323), .A2(new_n325), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n945), .B(new_n946), .Z(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(G900), .A2(G953), .ZN(new_n949));
  AND2_X1   g763(.A1(new_n730), .A2(new_n732), .ZN(new_n950));
  AND2_X1   g764(.A1(new_n830), .A2(new_n710), .ZN(new_n951));
  NAND4_X1  g765(.A1(new_n776), .A2(new_n781), .A3(new_n950), .A4(new_n951), .ZN(new_n952));
  NOR3_X1   g766(.A1(new_n774), .A2(new_n681), .A3(new_n698), .ZN(new_n953));
  XOR2_X1   g767(.A(new_n953), .B(KEYINPUT125), .Z(new_n954));
  OR2_X1    g768(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  OAI211_X1 g769(.A(new_n948), .B(new_n949), .C1(new_n955), .C2(G953), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n675), .A2(new_n951), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n957), .B(KEYINPUT62), .Z(new_n958));
  AOI21_X1  g772(.A(new_n681), .B1(new_n787), .B2(new_n804), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n959), .A2(new_n661), .A3(new_n759), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n958), .A2(new_n776), .A3(new_n781), .A4(new_n960), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(new_n310), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n962), .A2(new_n947), .ZN(new_n963));
  AND2_X1   g777(.A1(new_n956), .A2(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n310), .B1(G227), .B2(G900), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT124), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n965), .B1(new_n956), .B2(new_n966), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n964), .B(new_n967), .ZN(G72));
  NAND2_X1  g782(.A1(G472), .A2(G902), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n969), .B(KEYINPUT63), .Z(new_n970));
  NOR2_X1   g784(.A1(new_n509), .A2(new_n515), .ZN(new_n971));
  OAI211_X1 g785(.A(new_n847), .B(new_n970), .C1(new_n666), .C2(new_n971), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n970), .B1(new_n961), .B2(new_n937), .ZN(new_n973));
  XOR2_X1   g787(.A(new_n509), .B(KEYINPUT126), .Z(new_n974));
  INV_X1    g788(.A(new_n974), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n973), .A2(new_n515), .A3(new_n975), .ZN(new_n976));
  NOR3_X1   g790(.A1(new_n952), .A2(new_n937), .A3(new_n954), .ZN(new_n977));
  INV_X1    g791(.A(new_n970), .ZN(new_n978));
  OAI211_X1 g792(.A(new_n526), .B(new_n974), .C1(new_n977), .C2(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(KEYINPUT127), .ZN(new_n980));
  AND3_X1   g794(.A1(new_n979), .A2(new_n980), .A3(new_n908), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n980), .B1(new_n979), .B2(new_n908), .ZN(new_n982));
  OAI211_X1 g796(.A(new_n972), .B(new_n976), .C1(new_n981), .C2(new_n982), .ZN(new_n983));
  INV_X1    g797(.A(new_n983), .ZN(G57));
endmodule


