//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 1 1 0 1 1 1 0 0 1 0 1 1 1 1 1 0 1 1 1 0 0 1 0 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:02 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n548, new_n549, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n608, new_n609,
    new_n612, new_n614, new_n615, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1152, new_n1153, new_n1154, new_n1155;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT65), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT66), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XNOR2_X1  g017(.A(new_n442), .B(KEYINPUT67), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G219), .A2(G220), .A3(G221), .A4(G218), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  AND2_X1   g030(.A1(new_n452), .A2(G2106), .ZN(new_n456));
  OR2_X1    g031(.A1(new_n456), .A2(KEYINPUT68), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n453), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n456), .A2(KEYINPUT68), .ZN(new_n459));
  NAND3_X1  g034(.A1(new_n457), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  XOR2_X1   g037(.A(new_n462), .B(KEYINPUT69), .Z(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  AND3_X1   g042(.A1(new_n465), .A2(new_n467), .A3(G125), .ZN(new_n468));
  OAI21_X1  g043(.A(G2105), .B1(new_n463), .B2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT71), .ZN(new_n470));
  NOR3_X1   g045(.A1(new_n470), .A2(new_n464), .A3(G2105), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  AOI21_X1  g047(.A(KEYINPUT71), .B1(new_n472), .B2(G2104), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G101), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT70), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n477), .B1(new_n466), .B2(G2104), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n464), .A2(KEYINPUT70), .A3(KEYINPUT3), .ZN(new_n479));
  NAND4_X1  g054(.A1(new_n478), .A2(new_n479), .A3(new_n472), .A4(new_n467), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G137), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n469), .A2(new_n476), .A3(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G160));
  NAND4_X1  g059(.A1(new_n478), .A2(new_n479), .A3(G2105), .A4(new_n467), .ZN(new_n485));
  INV_X1    g060(.A(G124), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n472), .A2(G112), .ZN(new_n487));
  OAI21_X1  g062(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n488));
  OAI22_X1  g063(.A1(new_n485), .A2(new_n486), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n489), .B1(new_n481), .B2(G136), .ZN(G162));
  INV_X1    g065(.A(G126), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n472), .A2(G114), .ZN(new_n492));
  OAI21_X1  g067(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n493));
  OAI22_X1  g068(.A1(new_n485), .A2(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(G138), .ZN(new_n495));
  OAI21_X1  g070(.A(KEYINPUT4), .B1(new_n480), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n465), .A2(new_n467), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(new_n498));
  NOR3_X1   g073(.A1(new_n495), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n494), .B1(new_n496), .B2(new_n500), .ZN(G164));
  INV_X1    g076(.A(KEYINPUT72), .ZN(new_n502));
  INV_X1    g077(.A(G651), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n502), .B1(new_n503), .B2(KEYINPUT6), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT6), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n505), .A2(KEYINPUT72), .A3(G651), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n503), .A2(KEYINPUT6), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n507), .A2(G543), .A3(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G50), .ZN(new_n511));
  XNOR2_X1  g086(.A(KEYINPUT5), .B(G543), .ZN(new_n512));
  AND3_X1   g087(.A1(new_n505), .A2(KEYINPUT72), .A3(G651), .ZN(new_n513));
  AOI21_X1  g088(.A(KEYINPUT72), .B1(new_n505), .B2(G651), .ZN(new_n514));
  OAI211_X1 g089(.A(new_n512), .B(new_n508), .C1(new_n513), .C2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G88), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n512), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n518));
  OR2_X1    g093(.A1(new_n518), .A2(new_n503), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n511), .A2(new_n517), .A3(new_n519), .ZN(G303));
  INV_X1    g095(.A(G303), .ZN(G166));
  NAND2_X1  g096(.A1(new_n516), .A2(G89), .ZN(new_n522));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  XNOR2_X1  g098(.A(new_n523), .B(KEYINPUT7), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n512), .A2(G63), .A3(G651), .ZN(new_n525));
  XNOR2_X1  g100(.A(KEYINPUT73), .B(G51), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n525), .B1(new_n509), .B2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT74), .ZN(new_n528));
  OAI211_X1 g103(.A(new_n522), .B(new_n524), .C1(new_n527), .C2(new_n528), .ZN(new_n529));
  AND2_X1   g104(.A1(new_n527), .A2(new_n528), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n529), .A2(new_n530), .ZN(G168));
  NAND2_X1  g106(.A1(new_n516), .A2(G90), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n512), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n533));
  OR2_X1    g108(.A1(new_n533), .A2(new_n503), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n505), .A2(G651), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n535), .B1(new_n504), .B2(new_n506), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n536), .A2(G52), .A3(G543), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n532), .A2(new_n534), .A3(new_n537), .ZN(G301));
  INV_X1    g113(.A(G301), .ZN(G171));
  NAND2_X1  g114(.A1(new_n510), .A2(G43), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n516), .A2(G81), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n512), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n542));
  OR2_X1    g117(.A1(new_n542), .A2(new_n503), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n540), .A2(new_n541), .A3(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G860), .ZN(G153));
  NAND4_X1  g121(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g122(.A1(G1), .A2(G3), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT8), .ZN(new_n549));
  NAND4_X1  g124(.A1(G319), .A2(G483), .A3(G661), .A4(new_n549), .ZN(G188));
  AND2_X1   g125(.A1(KEYINPUT5), .A2(G543), .ZN(new_n551));
  NOR2_X1   g126(.A1(KEYINPUT5), .A2(G543), .ZN(new_n552));
  OAI21_X1  g127(.A(G65), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(G78), .A2(G543), .ZN(new_n554));
  AOI21_X1  g129(.A(new_n503), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  AND2_X1   g130(.A1(G53), .A2(G543), .ZN(new_n556));
  OAI211_X1 g131(.A(new_n508), .B(new_n556), .C1(new_n513), .C2(new_n514), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(KEYINPUT9), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT9), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n536), .A2(new_n559), .A3(new_n556), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n555), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT75), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n515), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n536), .A2(KEYINPUT75), .A3(new_n512), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n563), .A2(G91), .A3(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT76), .ZN(new_n566));
  AND3_X1   g141(.A1(new_n561), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  AOI21_X1  g142(.A(new_n566), .B1(new_n561), .B2(new_n565), .ZN(new_n568));
  NOR2_X1   g143(.A1(new_n567), .A2(new_n568), .ZN(G299));
  INV_X1    g144(.A(G168), .ZN(G286));
  AND4_X1   g145(.A1(KEYINPUT75), .A2(new_n507), .A3(new_n508), .A4(new_n512), .ZN(new_n571));
  AOI21_X1  g146(.A(KEYINPUT75), .B1(new_n536), .B2(new_n512), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n573), .A2(G87), .ZN(new_n574));
  OR2_X1    g149(.A1(new_n512), .A2(G74), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n510), .A2(G49), .B1(G651), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n574), .A2(new_n576), .ZN(G288));
  NAND2_X1  g152(.A1(new_n573), .A2(G86), .ZN(new_n578));
  NAND2_X1  g153(.A1(G73), .A2(G543), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n551), .A2(new_n552), .ZN(new_n580));
  INV_X1    g155(.A(G61), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n579), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n582), .A2(G651), .ZN(new_n583));
  INV_X1    g158(.A(G48), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n584), .B2(new_n509), .ZN(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n578), .A2(new_n586), .ZN(G305));
  AOI22_X1  g162(.A1(new_n512), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n588), .A2(new_n503), .ZN(new_n589));
  XOR2_X1   g164(.A(new_n589), .B(KEYINPUT77), .Z(new_n590));
  AOI22_X1  g165(.A1(G47), .A2(new_n510), .B1(new_n516), .B2(G85), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(G290));
  NAND2_X1  g167(.A1(G301), .A2(G868), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT78), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n509), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n536), .A2(KEYINPUT78), .A3(G543), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n595), .A2(G54), .A3(new_n596), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n512), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n598));
  OR2_X1    g173(.A1(new_n598), .A2(new_n503), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n573), .A2(KEYINPUT10), .A3(G92), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n563), .A2(G92), .A3(new_n564), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT10), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g179(.A(new_n600), .B1(new_n601), .B2(new_n604), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n593), .B1(new_n605), .B2(G868), .ZN(G284));
  OAI21_X1  g181(.A(new_n593), .B1(new_n605), .B2(G868), .ZN(G321));
  NAND2_X1  g182(.A1(G286), .A2(G868), .ZN(new_n608));
  INV_X1    g183(.A(G299), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n609), .B2(G868), .ZN(G297));
  XNOR2_X1  g185(.A(G297), .B(KEYINPUT79), .ZN(G280));
  INV_X1    g186(.A(G559), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n605), .B1(new_n612), .B2(G860), .ZN(G148));
  NAND2_X1  g188(.A1(new_n605), .A2(new_n612), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(G868), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(G868), .B2(new_n545), .ZN(G323));
  XNOR2_X1  g191(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g192(.A1(new_n475), .A2(new_n498), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT12), .ZN(new_n619));
  XNOR2_X1  g194(.A(KEYINPUT80), .B(G2100), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT13), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n619), .B(new_n621), .ZN(new_n622));
  INV_X1    g197(.A(G123), .ZN(new_n623));
  INV_X1    g198(.A(KEYINPUT81), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n624), .B1(new_n472), .B2(G111), .ZN(new_n625));
  OR2_X1    g200(.A1(G99), .A2(G2105), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n625), .A2(G2104), .A3(new_n626), .ZN(new_n627));
  NOR3_X1   g202(.A1(new_n624), .A2(new_n472), .A3(G111), .ZN(new_n628));
  OAI22_X1  g203(.A1(new_n485), .A2(new_n623), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n629), .B1(new_n481), .B2(G135), .ZN(new_n630));
  INV_X1    g205(.A(G2096), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n630), .A2(new_n631), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n622), .A2(new_n632), .A3(new_n633), .ZN(G156));
  XNOR2_X1  g209(.A(G2427), .B(G2438), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2430), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT15), .B(G2435), .ZN(new_n637));
  OR2_X1    g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n636), .A2(new_n637), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n638), .A2(KEYINPUT14), .A3(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2451), .B(G2454), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT16), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n640), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2443), .B(G2446), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(G1341), .B(G1348), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT82), .ZN(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  INV_X1    g224(.A(KEYINPUT83), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  INV_X1    g226(.A(G14), .ZN(new_n652));
  INV_X1    g227(.A(new_n645), .ZN(new_n653));
  AOI21_X1  g228(.A(new_n652), .B1(new_n653), .B2(new_n647), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(G401));
  INV_X1    g231(.A(KEYINPUT18), .ZN(new_n657));
  XOR2_X1   g232(.A(G2084), .B(G2090), .Z(new_n658));
  XNOR2_X1  g233(.A(G2067), .B(G2678), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n660), .A2(KEYINPUT17), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n658), .A2(new_n659), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n657), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(G2100), .ZN(new_n664));
  XOR2_X1   g239(.A(G2072), .B(G2078), .Z(new_n665));
  AOI21_X1  g240(.A(new_n665), .B1(new_n660), .B2(KEYINPUT18), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(G2096), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n664), .B(new_n667), .ZN(G227));
  XNOR2_X1  g243(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT87), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1961), .B(G1966), .ZN(new_n671));
  AND2_X1   g246(.A1(new_n671), .A2(KEYINPUT84), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n671), .A2(KEYINPUT84), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1956), .B(G2474), .ZN(new_n674));
  OR3_X1    g249(.A1(new_n672), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1971), .B(G1976), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT19), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT20), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n674), .B1(new_n672), .B2(new_n673), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n680), .A2(new_n677), .ZN(new_n681));
  XOR2_X1   g256(.A(new_n681), .B(KEYINPUT85), .Z(new_n682));
  NOR2_X1   g257(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n675), .A2(new_n680), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT86), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n685), .A2(new_n677), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1981), .B(G1986), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n687), .A2(new_n689), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n670), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(new_n692), .ZN(new_n694));
  INV_X1    g269(.A(new_n670), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n694), .A2(new_n695), .A3(new_n690), .ZN(new_n696));
  XNOR2_X1  g271(.A(G1991), .B(G1996), .ZN(new_n697));
  AND3_X1   g272(.A1(new_n693), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n697), .B1(new_n693), .B2(new_n696), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n698), .A2(new_n699), .ZN(G229));
  OAI21_X1  g275(.A(KEYINPUT98), .B1(G16), .B2(G21), .ZN(new_n701));
  NAND2_X1  g276(.A1(G168), .A2(G16), .ZN(new_n702));
  MUX2_X1   g277(.A(KEYINPUT98), .B(new_n701), .S(new_n702), .Z(new_n703));
  INV_X1    g278(.A(G1966), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  XOR2_X1   g280(.A(new_n705), .B(KEYINPUT99), .Z(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT24), .B(G34), .ZN(new_n707));
  INV_X1    g282(.A(G29), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n709), .B(KEYINPUT95), .Z(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(new_n483), .B2(new_n708), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT96), .ZN(new_n712));
  INV_X1    g287(.A(G16), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G5), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(G171), .B2(new_n713), .ZN(new_n715));
  OAI22_X1  g290(.A1(new_n712), .A2(G2084), .B1(G1961), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n708), .A2(G32), .ZN(new_n717));
  NAND3_X1  g292(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT26), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(G129), .ZN(new_n721));
  INV_X1    g296(.A(G105), .ZN(new_n722));
  OAI221_X1 g297(.A(new_n720), .B1(new_n485), .B2(new_n721), .C1(new_n474), .C2(new_n722), .ZN(new_n723));
  AND2_X1   g298(.A1(new_n481), .A2(G141), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  OR2_X1    g300(.A1(new_n725), .A2(KEYINPUT97), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n725), .A2(KEYINPUT97), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(new_n728), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n717), .B1(new_n729), .B2(new_n708), .ZN(new_n730));
  XNOR2_X1  g305(.A(KEYINPUT27), .B(G1996), .ZN(new_n731));
  INV_X1    g306(.A(new_n731), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n716), .B1(new_n730), .B2(new_n732), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT100), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n706), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n713), .A2(G20), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT23), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(new_n609), .B2(new_n713), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT102), .ZN(new_n739));
  INV_X1    g314(.A(G1956), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n730), .A2(new_n732), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n708), .A2(G27), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(G164), .B2(new_n708), .ZN(new_n744));
  XNOR2_X1  g319(.A(KEYINPUT101), .B(G2078), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n744), .B(new_n745), .ZN(new_n746));
  NOR2_X1   g321(.A1(G16), .A2(G19), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(new_n545), .B2(G16), .ZN(new_n748));
  XOR2_X1   g323(.A(KEYINPUT92), .B(G1341), .Z(new_n749));
  AOI22_X1  g324(.A1(new_n748), .A2(new_n749), .B1(new_n715), .B2(G1961), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(new_n748), .B2(new_n749), .ZN(new_n751));
  NOR3_X1   g326(.A1(new_n742), .A2(new_n746), .A3(new_n751), .ZN(new_n752));
  NOR2_X1   g327(.A1(G29), .A2(G35), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(G162), .B2(G29), .ZN(new_n754));
  XNOR2_X1  g329(.A(KEYINPUT29), .B(G2090), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  NOR2_X1   g331(.A1(G29), .A2(G33), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT94), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n481), .A2(G139), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n472), .A2(G103), .A3(G2104), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT25), .Z(new_n761));
  AOI22_X1  g336(.A1(new_n498), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n762));
  OAI211_X1 g337(.A(new_n759), .B(new_n761), .C1(new_n762), .C2(new_n472), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n758), .B1(new_n763), .B2(new_n708), .ZN(new_n764));
  INV_X1    g339(.A(G2072), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n764), .A2(new_n765), .ZN(new_n767));
  INV_X1    g342(.A(KEYINPUT30), .ZN(new_n768));
  AND2_X1   g343(.A1(new_n768), .A2(G28), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n708), .B1(new_n768), .B2(G28), .ZN(new_n770));
  AND2_X1   g345(.A1(KEYINPUT31), .A2(G11), .ZN(new_n771));
  NOR2_X1   g346(.A1(KEYINPUT31), .A2(G11), .ZN(new_n772));
  OAI22_X1  g347(.A1(new_n769), .A2(new_n770), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(new_n630), .B2(G29), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n767), .A2(new_n774), .ZN(new_n775));
  NOR3_X1   g350(.A1(new_n756), .A2(new_n766), .A3(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n708), .A2(G26), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT28), .ZN(new_n778));
  INV_X1    g353(.A(G128), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n472), .A2(G116), .ZN(new_n780));
  OAI21_X1  g355(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n781));
  OAI22_X1  g356(.A1(new_n485), .A2(new_n779), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(new_n481), .B2(G140), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n778), .B1(new_n783), .B2(new_n708), .ZN(new_n784));
  XNOR2_X1  g359(.A(KEYINPUT93), .B(G2067), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(new_n712), .B2(G2084), .ZN(new_n787));
  OAI211_X1 g362(.A(new_n776), .B(new_n787), .C1(new_n703), .C2(new_n704), .ZN(new_n788));
  NOR2_X1   g363(.A1(G4), .A2(G16), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(new_n605), .B2(G16), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(G1348), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n788), .A2(new_n791), .ZN(new_n792));
  NAND4_X1  g367(.A1(new_n735), .A2(new_n741), .A3(new_n752), .A4(new_n792), .ZN(new_n793));
  AND2_X1   g368(.A1(new_n713), .A2(G23), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(G288), .B2(G16), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT90), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT33), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n797), .A2(G1976), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n797), .A2(G1976), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n713), .A2(G22), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(G166), .B2(new_n713), .ZN(new_n801));
  XOR2_X1   g376(.A(new_n801), .B(KEYINPUT91), .Z(new_n802));
  AND2_X1   g377(.A1(new_n802), .A2(G1971), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n802), .A2(G1971), .ZN(new_n804));
  MUX2_X1   g379(.A(G6), .B(G305), .S(G16), .Z(new_n805));
  XNOR2_X1  g380(.A(KEYINPUT32), .B(G1981), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  NOR3_X1   g382(.A1(new_n803), .A2(new_n804), .A3(new_n807), .ZN(new_n808));
  NAND3_X1  g383(.A1(new_n798), .A2(new_n799), .A3(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n809), .A2(KEYINPUT34), .ZN(new_n810));
  INV_X1    g385(.A(KEYINPUT34), .ZN(new_n811));
  NAND4_X1  g386(.A1(new_n798), .A2(new_n811), .A3(new_n799), .A4(new_n808), .ZN(new_n812));
  INV_X1    g387(.A(G131), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n480), .A2(new_n813), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT88), .ZN(new_n815));
  INV_X1    g390(.A(new_n485), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n816), .A2(G119), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n472), .A2(G107), .ZN(new_n818));
  OAI21_X1  g393(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n819));
  OAI211_X1 g394(.A(new_n815), .B(new_n817), .C1(new_n818), .C2(new_n819), .ZN(new_n820));
  MUX2_X1   g395(.A(G25), .B(new_n820), .S(G29), .Z(new_n821));
  XNOR2_X1  g396(.A(KEYINPUT35), .B(G1991), .ZN(new_n822));
  XOR2_X1   g397(.A(new_n821), .B(new_n822), .Z(new_n823));
  MUX2_X1   g398(.A(G24), .B(G290), .S(G16), .Z(new_n824));
  XOR2_X1   g399(.A(KEYINPUT89), .B(G1986), .Z(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  NAND4_X1  g401(.A1(new_n810), .A2(new_n812), .A3(new_n823), .A4(new_n826), .ZN(new_n827));
  OR2_X1    g402(.A1(new_n827), .A2(KEYINPUT36), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n827), .A2(KEYINPUT36), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n793), .B1(new_n828), .B2(new_n829), .ZN(G311));
  INV_X1    g405(.A(G311), .ZN(G150));
  NAND2_X1  g406(.A1(new_n510), .A2(G55), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n516), .A2(G93), .ZN(new_n833));
  AOI22_X1  g408(.A1(new_n512), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n834));
  OR2_X1    g409(.A1(new_n834), .A2(new_n503), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n832), .A2(new_n833), .A3(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT103), .ZN(new_n837));
  OR3_X1    g412(.A1(new_n544), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n836), .A2(new_n837), .ZN(new_n839));
  NAND4_X1  g414(.A1(new_n833), .A2(new_n832), .A3(new_n835), .A4(KEYINPUT103), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n839), .A2(new_n544), .A3(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n838), .A2(new_n841), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n842), .B(KEYINPUT38), .Z(new_n843));
  NAND2_X1  g418(.A1(new_n605), .A2(G559), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n843), .B(new_n844), .ZN(new_n845));
  AND2_X1   g420(.A1(new_n845), .A2(KEYINPUT39), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n845), .A2(KEYINPUT39), .ZN(new_n847));
  NOR3_X1   g422(.A1(new_n846), .A2(new_n847), .A3(G860), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n836), .A2(G860), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(KEYINPUT37), .ZN(new_n850));
  OR2_X1    g425(.A1(new_n848), .A2(new_n850), .ZN(G145));
  XNOR2_X1  g426(.A(new_n728), .B(new_n783), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n481), .A2(G142), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n816), .A2(G130), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n472), .A2(G118), .ZN(new_n855));
  OAI21_X1  g430(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n856));
  OAI211_X1 g431(.A(new_n853), .B(new_n854), .C1(new_n855), .C2(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n852), .B(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n496), .A2(new_n500), .ZN(new_n859));
  INV_X1    g434(.A(new_n494), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n861), .A2(KEYINPUT104), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT104), .ZN(new_n863));
  NAND2_X1  g438(.A1(G164), .A2(new_n863), .ZN(new_n864));
  AND2_X1   g439(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n763), .A2(KEYINPUT105), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n865), .B(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n820), .B(new_n619), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n867), .B(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n858), .B(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n630), .B(new_n483), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(G162), .ZN(new_n872));
  OR2_X1    g447(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g448(.A(G37), .B1(new_n870), .B2(new_n872), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g451(.A(new_n842), .B(new_n614), .ZN(new_n877));
  OAI21_X1  g452(.A(KEYINPUT106), .B1(new_n567), .B2(new_n568), .ZN(new_n878));
  INV_X1    g453(.A(G91), .ZN(new_n879));
  NOR3_X1   g454(.A1(new_n571), .A2(new_n572), .A3(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(new_n555), .ZN(new_n881));
  AND4_X1   g456(.A1(new_n559), .A2(new_n507), .A3(new_n508), .A4(new_n556), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n559), .B1(new_n536), .B2(new_n556), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n881), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  OAI21_X1  g459(.A(KEYINPUT76), .B1(new_n880), .B2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT106), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n561), .A2(new_n565), .A3(new_n566), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n601), .A2(new_n604), .ZN(new_n889));
  INV_X1    g464(.A(new_n600), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n878), .A2(new_n888), .A3(new_n891), .ZN(new_n892));
  OAI211_X1 g467(.A(new_n605), .B(KEYINPUT106), .C1(new_n568), .C2(new_n567), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n877), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(KEYINPUT41), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT107), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT41), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n892), .A2(new_n898), .A3(new_n893), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n896), .A2(new_n897), .A3(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n894), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n901), .A2(KEYINPUT107), .A3(new_n898), .ZN(new_n902));
  AND2_X1   g477(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n895), .B1(new_n903), .B2(new_n877), .ZN(new_n904));
  OR2_X1    g479(.A1(new_n904), .A2(KEYINPUT42), .ZN(new_n905));
  XOR2_X1   g480(.A(G290), .B(G305), .Z(new_n906));
  XNOR2_X1  g481(.A(G288), .B(G166), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n906), .B(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n904), .A2(KEYINPUT42), .ZN(new_n910));
  AND3_X1   g485(.A1(new_n905), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n909), .B1(new_n905), .B2(new_n910), .ZN(new_n912));
  OAI21_X1  g487(.A(G868), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(G868), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n836), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n913), .A2(new_n915), .ZN(G295));
  NAND2_X1  g491(.A1(new_n913), .A2(new_n915), .ZN(G331));
  NAND3_X1  g492(.A1(G168), .A2(KEYINPUT108), .A3(G171), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT108), .ZN(new_n919));
  NAND2_X1  g494(.A1(G301), .A2(new_n919), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n532), .A2(new_n534), .A3(KEYINPUT108), .A4(new_n537), .ZN(new_n921));
  OAI211_X1 g496(.A(new_n920), .B(new_n921), .C1(new_n529), .C2(new_n530), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n918), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n923), .A2(new_n842), .ZN(new_n924));
  NAND4_X1  g499(.A1(new_n918), .A2(new_n922), .A3(new_n838), .A4(new_n841), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n900), .A2(new_n902), .A3(new_n926), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n894), .B1(new_n842), .B2(new_n923), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT109), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n925), .A2(new_n929), .ZN(new_n930));
  OR2_X1    g505(.A1(new_n925), .A2(new_n929), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n928), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n927), .A2(new_n908), .A3(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(G37), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n908), .B1(new_n927), .B2(new_n932), .ZN(new_n936));
  OAI21_X1  g511(.A(KEYINPUT43), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT110), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  OAI211_X1 g514(.A(KEYINPUT110), .B(KEYINPUT43), .C1(new_n935), .C2(new_n936), .ZN(new_n940));
  INV_X1    g515(.A(new_n935), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n931), .A2(new_n924), .A3(new_n930), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT111), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n899), .A2(new_n943), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n892), .A2(new_n893), .A3(KEYINPUT111), .A4(new_n898), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n944), .A2(new_n896), .A3(new_n945), .ZN(new_n946));
  AND2_X1   g521(.A1(new_n942), .A2(new_n946), .ZN(new_n947));
  AND2_X1   g522(.A1(new_n928), .A2(new_n925), .ZN(new_n948));
  OAI211_X1 g523(.A(KEYINPUT112), .B(new_n909), .C1(new_n947), .C2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT43), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT112), .ZN(new_n951));
  AOI22_X1  g526(.A1(new_n942), .A2(new_n946), .B1(new_n925), .B2(new_n928), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n951), .B1(new_n952), .B2(new_n908), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n941), .A2(new_n949), .A3(new_n950), .A4(new_n953), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n939), .A2(new_n940), .A3(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n950), .B1(new_n935), .B2(new_n936), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n941), .A2(new_n949), .A3(new_n953), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n956), .B1(new_n957), .B2(new_n950), .ZN(new_n958));
  MUX2_X1   g533(.A(new_n955), .B(new_n958), .S(KEYINPUT44), .Z(G397));
  XNOR2_X1  g534(.A(KEYINPUT113), .B(G1384), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n865), .A2(new_n960), .ZN(new_n961));
  XOR2_X1   g536(.A(KEYINPUT114), .B(KEYINPUT45), .Z(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND4_X1  g538(.A1(new_n469), .A2(new_n476), .A3(G40), .A4(new_n482), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  OR3_X1    g541(.A1(new_n966), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n967));
  OAI21_X1  g542(.A(KEYINPUT46), .B1(new_n966), .B2(G1996), .ZN(new_n968));
  XNOR2_X1  g543(.A(new_n783), .B(G2067), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n969), .ZN(new_n970));
  AOI22_X1  g545(.A1(new_n967), .A2(new_n968), .B1(new_n965), .B2(new_n970), .ZN(new_n971));
  XOR2_X1   g546(.A(KEYINPUT126), .B(KEYINPUT47), .Z(new_n972));
  XNOR2_X1  g547(.A(new_n971), .B(new_n972), .ZN(new_n973));
  XNOR2_X1  g548(.A(new_n728), .B(G1996), .ZN(new_n974));
  INV_X1    g549(.A(new_n969), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n965), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n820), .A2(new_n822), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(G2067), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n783), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n965), .B1(new_n981), .B2(KEYINPUT125), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n982), .B1(KEYINPUT125), .B2(new_n981), .ZN(new_n983));
  OR3_X1    g558(.A1(new_n966), .A2(G1986), .A3(G290), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT48), .ZN(new_n985));
  AND2_X1   g560(.A1(new_n820), .A2(new_n822), .ZN(new_n986));
  NOR4_X1   g561(.A1(new_n974), .A2(new_n975), .A3(new_n977), .A4(new_n986), .ZN(new_n987));
  OAI22_X1  g562(.A1(new_n984), .A2(new_n985), .B1(new_n966), .B2(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n988), .B1(new_n985), .B2(new_n984), .ZN(new_n989));
  NOR3_X1   g564(.A1(new_n973), .A2(new_n983), .A3(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(G1981), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n578), .A2(new_n991), .A3(new_n586), .ZN(new_n992));
  AND2_X1   g567(.A1(new_n516), .A2(G86), .ZN(new_n993));
  OAI21_X1  g568(.A(G1981), .B1(new_n993), .B2(new_n585), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n992), .A2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT49), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(G1384), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n861), .A2(new_n998), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n999), .A2(new_n964), .ZN(new_n1000));
  XNOR2_X1  g575(.A(KEYINPUT117), .B(G8), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n992), .A2(KEYINPUT49), .A3(new_n994), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n997), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n574), .A2(G1976), .A3(new_n576), .ZN(new_n1005));
  INV_X1    g580(.A(G1976), .ZN(new_n1006));
  AOI21_X1  g581(.A(KEYINPUT52), .B1(G288), .B2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1002), .A2(new_n1005), .A3(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1001), .ZN(new_n1009));
  OAI211_X1 g584(.A(new_n1005), .B(new_n1009), .C1(new_n964), .C2(new_n999), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(KEYINPUT52), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1004), .A2(new_n1008), .A3(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(G303), .A2(G8), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT116), .ZN(new_n1014));
  AND2_X1   g589(.A1(new_n1014), .A2(KEYINPUT55), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1014), .A2(KEYINPUT55), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1013), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1017), .B1(new_n1013), .B2(new_n1016), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n999), .A2(KEYINPUT50), .ZN(new_n1019));
  INV_X1    g594(.A(new_n964), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT115), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT50), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(new_n998), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1021), .B1(G164), .B2(new_n1023), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n861), .A2(KEYINPUT115), .A3(new_n1022), .A4(new_n998), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n1019), .A2(new_n1020), .A3(new_n1024), .A4(new_n1025), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1026), .A2(G2090), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n862), .A2(new_n864), .A3(KEYINPUT45), .A4(new_n960), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n964), .B1(new_n999), .B2(new_n962), .ZN(new_n1029));
  AOI21_X1  g604(.A(G1971), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  OAI211_X1 g605(.A(G8), .B(new_n1018), .C1(new_n1027), .C2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(new_n992), .ZN(new_n1032));
  NOR2_X1   g607(.A1(G288), .A2(G1976), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1032), .B1(new_n1004), .B2(new_n1033), .ZN(new_n1034));
  XNOR2_X1  g609(.A(new_n1002), .B(KEYINPUT118), .ZN(new_n1035));
  OAI22_X1  g610(.A1(new_n1012), .A2(new_n1031), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT61), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n561), .A2(new_n565), .ZN(new_n1038));
  XOR2_X1   g613(.A(new_n1038), .B(KEYINPUT57), .Z(new_n1039));
  NOR2_X1   g614(.A1(G164), .A2(new_n1023), .ZN(new_n1040));
  AOI21_X1  g615(.A(G1384), .B1(new_n859), .B2(new_n860), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1020), .B1(new_n1022), .B2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1040), .B1(new_n1042), .B2(KEYINPUT119), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT119), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1019), .A2(new_n1044), .A3(new_n1020), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1043), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(new_n740), .ZN(new_n1047));
  XNOR2_X1  g622(.A(KEYINPUT56), .B(G2072), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1028), .A2(new_n1029), .A3(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1039), .B1(new_n1047), .B2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(G1956), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1039), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1049), .ZN(new_n1053));
  NOR3_X1   g628(.A1(new_n1051), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1037), .B1(new_n1050), .B2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1047), .A2(new_n1039), .A3(new_n1049), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1052), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1056), .A2(new_n1057), .A3(KEYINPUT61), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1059));
  XNOR2_X1  g634(.A(KEYINPUT58), .B(G1341), .ZN(new_n1060));
  OAI22_X1  g635(.A1(new_n1059), .A2(G1996), .B1(new_n1000), .B2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(new_n545), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(KEYINPUT59), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT59), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1061), .A2(new_n1064), .A3(new_n545), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(G1348), .ZN(new_n1067));
  AOI22_X1  g642(.A1(new_n1026), .A2(new_n1067), .B1(new_n979), .B2(new_n1000), .ZN(new_n1068));
  OR2_X1    g643(.A1(new_n1068), .A2(KEYINPUT60), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1026), .A2(new_n1067), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1000), .A2(new_n979), .ZN(new_n1071));
  AND4_X1   g646(.A1(KEYINPUT60), .A2(new_n1070), .A3(new_n891), .A4(new_n1071), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n891), .B1(new_n1068), .B2(KEYINPUT60), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1069), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1055), .A2(new_n1058), .A3(new_n1066), .A4(new_n1074), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1068), .A2(new_n891), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1056), .B1(new_n1050), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1075), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1025), .A2(new_n1024), .ZN(new_n1079));
  OR3_X1    g654(.A1(new_n1079), .A2(new_n1042), .A3(G2084), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT45), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n999), .A2(new_n1081), .ZN(new_n1082));
  OAI211_X1 g657(.A(new_n1082), .B(new_n1020), .C1(new_n962), .C2(new_n999), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(new_n704), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1080), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(new_n1009), .ZN(new_n1086));
  NOR2_X1   g661(.A1(G168), .A2(new_n1001), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1087), .A2(KEYINPUT51), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(G8), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1090), .B1(new_n1080), .B2(new_n1084), .ZN(new_n1091));
  OAI21_X1  g666(.A(KEYINPUT51), .B1(new_n1091), .B2(new_n1087), .ZN(new_n1092));
  AOI211_X1 g667(.A(G168), .B(new_n1001), .C1(new_n1080), .C2(new_n1084), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1089), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT53), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1095), .B1(new_n1059), .B2(G2078), .ZN(new_n1096));
  XNOR2_X1  g671(.A(KEYINPUT122), .B(G1961), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1026), .A2(new_n1097), .ZN(new_n1098));
  AND2_X1   g673(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1099));
  XNOR2_X1  g674(.A(G301), .B(KEYINPUT54), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1100), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1095), .A2(G2078), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n963), .A2(new_n1020), .A3(new_n1028), .A4(new_n1102), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1099), .A2(new_n1101), .A3(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1083), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(new_n1102), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1106), .A2(new_n1096), .A3(new_n1098), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(new_n1100), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1104), .A2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1012), .ZN(new_n1110));
  INV_X1    g685(.A(G2090), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1043), .A2(new_n1111), .A3(new_n1045), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1030), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1001), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  OAI211_X1 g689(.A(new_n1110), .B(new_n1031), .C1(new_n1114), .C2(new_n1018), .ZN(new_n1115));
  NOR3_X1   g690(.A1(new_n1094), .A2(new_n1109), .A3(new_n1115), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1036), .B1(new_n1078), .B2(new_n1116), .ZN(new_n1117));
  XNOR2_X1  g692(.A(KEYINPUT120), .B(KEYINPUT63), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1085), .A2(G168), .A3(new_n1009), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1118), .B1(new_n1115), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT121), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  OAI211_X1 g697(.A(KEYINPUT121), .B(new_n1118), .C1(new_n1115), .C2(new_n1119), .ZN(new_n1123));
  AND2_X1   g698(.A1(new_n1110), .A2(new_n1031), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1119), .ZN(new_n1125));
  OAI21_X1  g700(.A(G8), .B1(new_n1027), .B2(new_n1030), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1018), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1124), .A2(KEYINPUT63), .A3(new_n1125), .A4(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1122), .A2(new_n1123), .A3(new_n1129), .ZN(new_n1130));
  AND3_X1   g705(.A1(new_n1117), .A2(KEYINPUT123), .A3(new_n1130), .ZN(new_n1131));
  AOI21_X1  g706(.A(KEYINPUT123), .B1(new_n1117), .B2(new_n1130), .ZN(new_n1132));
  AOI211_X1 g707(.A(G301), .B(new_n1115), .C1(new_n1106), .C2(new_n1099), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT124), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT62), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1134), .B1(new_n1094), .B2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1094), .A2(new_n1135), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1133), .A2(new_n1136), .A3(new_n1137), .ZN(new_n1138));
  NOR3_X1   g713(.A1(new_n1094), .A2(new_n1134), .A3(new_n1135), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NOR3_X1   g715(.A1(new_n1131), .A2(new_n1132), .A3(new_n1140), .ZN(new_n1141));
  XOR2_X1   g716(.A(G290), .B(G1986), .Z(new_n1142));
  AOI21_X1  g717(.A(new_n966), .B1(new_n987), .B2(new_n1142), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n990), .B1(new_n1141), .B2(new_n1143), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g719(.A1(new_n460), .A2(G227), .ZN(new_n1146));
  OAI211_X1 g720(.A(new_n655), .B(new_n1146), .C1(new_n698), .C2(new_n699), .ZN(new_n1147));
  AOI21_X1  g721(.A(new_n1147), .B1(new_n873), .B2(new_n874), .ZN(new_n1148));
  AND3_X1   g722(.A1(new_n955), .A2(KEYINPUT127), .A3(new_n1148), .ZN(new_n1149));
  AOI21_X1  g723(.A(KEYINPUT127), .B1(new_n955), .B2(new_n1148), .ZN(new_n1150));
  NOR2_X1   g724(.A1(new_n1149), .A2(new_n1150), .ZN(G308));
  NAND2_X1  g725(.A1(new_n955), .A2(new_n1148), .ZN(new_n1152));
  INV_X1    g726(.A(KEYINPUT127), .ZN(new_n1153));
  NAND2_X1  g727(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g728(.A1(new_n955), .A2(KEYINPUT127), .A3(new_n1148), .ZN(new_n1155));
  NAND2_X1  g729(.A1(new_n1154), .A2(new_n1155), .ZN(G225));
endmodule


